module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
 n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
 n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
 n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
 n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
 n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , 
 n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , 
 n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , 
 n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , 
 n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , 
 n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , 
 n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , 
 n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , 
 n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , 
 n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , 
 n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , 
 n381 , n382 , n383 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 ;
output n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , 
 n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , 
 n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , 
 n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , 
 n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , 
 n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , 
 n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , 
 n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , 
 n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , 
 n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , 
 n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , 
 n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , 
 n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , 
 n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , 
 n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , 
 n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , 
 n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , 
 n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , 
 n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , 
 n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , 
 n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , 
 n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , 
 n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , 
 n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , 
 n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , 
 n379 , n380 , n381 , n382 , n383 ;
wire n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , 
 n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , 
 n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , 
 n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , 
 n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , 
 n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , 
 n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , 
 n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , 
 n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , 
 n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , 
 n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , 
 n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , 
 n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , 
 n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , 
 n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , 
 n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , 
 n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , 
 n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , 
 n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , 
 n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , 
 n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , 
 n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , 
 n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , 
 n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , 
 n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , 
 n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , 
 n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , 
 n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , 
 n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , 
 n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , 
 n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , 
 n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , 
 n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , 
 n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , 
 n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , 
 n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , 
 n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , 
 n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , 
 n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , 
 n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , 
 n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , 
 n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , 
 n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , 
 n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , 
 n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , 
 n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , 
 n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , 
 n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , 
 n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , 
 n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , 
 n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , 
 n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , 
 n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , 
 n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , 
 n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , 
 n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , 
 n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , 
 n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , 
 n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , 
 n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , 
 n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , 
 n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , 
 n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , 
 n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , 
 n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , 
 n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , 
 n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , 
 n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , 
 n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , 
 n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , 
 n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , 
 n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , 
 n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , 
 n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , 
 n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , 
 n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , 
 n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , 
 n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , 
 n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , 
 n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , 
 n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , 
 n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , 
 n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , 
 n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , 
 n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , 
 n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , 
 n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , 
 n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , 
 n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , 
 n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , 
 n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , 
 n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , 
 n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , 
 n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , 
 n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , 
 n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , 
 n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , 
 n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , 
 n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , 
 n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , 
 n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , 
 n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , 
 n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , 
 n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , 
 n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , 
 n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , 
 n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , 
 n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , 
 n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , 
 n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , 
 n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , 
 n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , 
 n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , 
 n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , 
 n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , 
 n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , 
 n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , 
 n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , 
 n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , 
 n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , 
 n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , 
 n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , 
 n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , 
 n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , 
 n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , 
 n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , 
 n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , 
 n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , 
 n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , 
 n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , 
 n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , 
 n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , 
 n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , 
 n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , 
 n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , 
 n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , 
 n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , 
 n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , 
 n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , 
 n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , 
 n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , 
 n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , 
 n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , 
 n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , 
 n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , 
 n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , 
 n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , 
 n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , 
 n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , 
 n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , 
 n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , 
 n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , 
 n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , 
 n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , 
 n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , 
 n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , 
 n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , 
 n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , 
 n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , 
 n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , 
 n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , 
 n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , 
 n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , 
 n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , 
 n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , 
 n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , 
 n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , 
 n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , 
 n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , 
 n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , 
 n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , 
 n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , 
 n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , 
 n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , 
 n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , 
 n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , 
 n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , 
 n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , 
 n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , 
 n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , 
 n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , 
 n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , 
 n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , 
 n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , 
 n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , 
 n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , 
 n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , 
 n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , 
 n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , 
 n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , 
 n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , 
 n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , 
 n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , 
 n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , 
 n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , 
 n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , 
 n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , 
 n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , 
 n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , 
 n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , 
 n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , 
 n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , 
 n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , 
 n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , 
 n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , 
 n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , 
 n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , 
 n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , 
 n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , 
 n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , 
 n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , 
 n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , 
 n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , 
 n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , 
 n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , 
 n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , 
 n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , 
 n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , 
 n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , 
 n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , 
 n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , 
 n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , 
 n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , 
 n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , 
 n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , 
 n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , 
 n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , 
 n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , 
 n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , 
 n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , 
 n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , 
 n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , 
 n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , 
 n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , 
 n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , 
 n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , 
 n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , 
 n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , 
 n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , 
 n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , 
 n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , 
 n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , 
 n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , 
 n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , 
 n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , 
 n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , 
 n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , 
 n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , 
 n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , 
 n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , 
 n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , 
 n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , 
 n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , 
 n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , 
 n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , 
 n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , 
 n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , 
 n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , 
 n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , 
 n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , 
 n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , 
 n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , 
 n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , 
 n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , 
 n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , 
 n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , 
 n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , 
 n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , 
 n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , 
 n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , 
 n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , 
 n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , 
 n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , 
 n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , 
 n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , 
 n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , 
 n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , 
 n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , 
 n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , 
 n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , 
 n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , 
 n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , 
 n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , 
 n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , 
 n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , 
 n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , 
 n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , 
 n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , 
 n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , 
 n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , 
 n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , 
 n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , 
 n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , 
 n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , 
 n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , 
 n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , 
 n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , 
 n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , 
 n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , 
 n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , 
 n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , 
 n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , 
 n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , 
 n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , 
 n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , 
 n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , 
 n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , 
 n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , 
 n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , 
 n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , 
 n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , 
 n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , 
 n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , 
 n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , 
 n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , 
 n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , 
 n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , 
 n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , 
 n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , 
 n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , 
 n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , 
 n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , 
 n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , 
 n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , 
 n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , 
 n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , 
 n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , 
 n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , 
 n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , 
 n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , 
 n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , 
 n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , 
 n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , 
 n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , 
 n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , 
 n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , 
 n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , 
 n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , 
 n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , 
 n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , 
 n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , 
 n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , 
 n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , 
 n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , 
 n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , 
 n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , 
 n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , 
 n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , 
 n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , 
 n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , 
 n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , 
 n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , 
 n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , 
 n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , 
 n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , 
 n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , 
 n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , 
 n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , 
 n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , 
 n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , 
 n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , 
 n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , 
 n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , 
 n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , 
 n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , 
 n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , 
 n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , 
 n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , 
 n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , 
 n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , 
 n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , 
 n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , 
 n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , 
 n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , 
 n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , 
 n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , 
 n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , 
 n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , 
 n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , 
 n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , 
 n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , 
 n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , 
 n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , 
 n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , 
 n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , 
 n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , 
 n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , 
 n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , 
 n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , 
 n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , 
 n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , 
 n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , 
 n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , 
 n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , 
 n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , 
 n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , 
 n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , 
 n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , 
 n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , 
 n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , 
 n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , 
 n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , 
 n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , 
 n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , 
 n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , 
 n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , 
 n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , 
 n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , 
 n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , 
 n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , 
 n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , 
 n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , 
 n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , 
 n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , 
 n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , 
 n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , 
 n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , 
 n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , 
 n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , 
 n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , 
 n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , 
 n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , 
 n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , 
 n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , 
 n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , 
 n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , 
 n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , 
 n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , 
 n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , 
 n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , 
 n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , 
 n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , 
 n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , 
 n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , 
 n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , 
 n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , 
 n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , 
 n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , 
 n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , 
 n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , 
 n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , 
 n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , 
 n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , 
 n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , 
 n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , 
 n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , 
 n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , 
 n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , 
 n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , 
 n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , 
 n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , 
 n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , 
 n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , 
 n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , 
 n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , 
 n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , 
 n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , 
 n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , 
 n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , 
 n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , 
 n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , 
 n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , 
 n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , 
 n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , 
 n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , 
 n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , 
 n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , 
 n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , 
 n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , 
 n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , 
 n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , 
 n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , 
 n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , 
 n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , 
 n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , 
 n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , 
 n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , 
 n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , 
 n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , 
 n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , 
 n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , 
 n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , 
 n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , 
 n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , 
 n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , 
 n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , 
 n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , 
 n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , 
 n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , 
 n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , 
 n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , 
 n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , 
 n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , 
 n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , 
 n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , 
 n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , 
 n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , 
 n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , 
 n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , 
 n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , 
 n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , 
 n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , 
 n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , 
 n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , 
 n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , 
 n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , 
 n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , 
 n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , 
 n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , 
 n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , 
 n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , 
 n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , 
 n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , 
 n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , 
 n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , 
 n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , 
 n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , 
 n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , 
 n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , 
 n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , 
 n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , 
 n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , 
 n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , 
 n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , 
 n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , 
 n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , 
 n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , 
 n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , 
 n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , 
 n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , 
 n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , 
 n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , 
 n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , 
 n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , 
 n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , 
 n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , 
 n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , 
 n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , 
 n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , 
 n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , 
 n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , 
 n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , 
 n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , 
 n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , 
 n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , 
 n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , 
 n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , 
 n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , 
 n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , 
 n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , 
 n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , 
 n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , 
 n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , 
 n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , 
 n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , 
 n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , 
 n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , 
 n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , 
 n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , 
 n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , 
 n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , 
 n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , 
 n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , 
 n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , 
 n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , 
 n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , 
 n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , 
 n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , 
 n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , 
 n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , 
 n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , 
 n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , 
 n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , 
 n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , 
 n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , 
 n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , 
 n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , 
 n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , 
 n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , 
 n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , 
 n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , 
 n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , 
 n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , 
 n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , 
 n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , 
 n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , 
 n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , 
 n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , 
 n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , 
 n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , 
 n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , 
 n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , 
 n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , 
 n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , 
 n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , 
 n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , 
 n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , 
 n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , 
 n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , 
 n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , 
 n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , 
 n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , 
 n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , 
 n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , 
 n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , 
 n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , 
 n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , 
 n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , 
 n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , 
 n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , 
 n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , 
 n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , 
 n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , 
 n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , 
 n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , 
 n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , 
 n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , 
 n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , 
 n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , 
 n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , 
 n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , 
 n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , 
 n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , 
 n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , 
 n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , 
 n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , 
 n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , 
 n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , 
 n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , 
 n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , 
 n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , 
 n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , 
 n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , 
 n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , 
 n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , 
 n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , 
 n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , 
 n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , 
 n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , 
 n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , 
 n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , 
 n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , 
 n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , 
 n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , 
 n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , 
 n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , 
 n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , 
 n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , 
 n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , 
 n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , 
 n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , 
 n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , 
 n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , 
 n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , 
 n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , 
 n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , 
 n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , 
 n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , 
 n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , 
 n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , 
 n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , 
 n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , 
 n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , 
 n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , 
 n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , 
 n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , 
 n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , 
 n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , 
 n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , 
 n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , 
 n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , 
 n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , 
 n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , 
 n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , 
 n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , 
 n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , 
 n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , 
 n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , 
 n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , 
 n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , 
 n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , 
 n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , 
 n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , 
 n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , 
 n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , 
 n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , 
 n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , 
 n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , 
 n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , 
 n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , 
 n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , 
 n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , 
 n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , 
 n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , 
 n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , 
 n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , 
 n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , 
 n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , 
 n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , 
 n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , 
 n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , 
 n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , 
 n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , 
 n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , 
 n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , 
 n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , 
 n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , 
 n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , 
 n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , 
 n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , 
 n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , 
 n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , 
 n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , 
 n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , 
 n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , 
 n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , 
 n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , 
 n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , 
 n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , 
 n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , 
 n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , 
 n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , 
 n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , 
 n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , 
 n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , 
 n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , 
 n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , 
 n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , 
 n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , 
 n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , 
 n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , 
 n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , 
 n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , 
 n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , 
 n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , 
 n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , 
 n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , 
 n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , 
 n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , 
 n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , 
 n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , 
 n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , 
 n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , 
 n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , 
 n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , 
 n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , 
 n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , 
 n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , 
 n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , 
 n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , 
 n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , 
 n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , 
 n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , 
 n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , 
 n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , 
 n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , 
 n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , 
 n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , 
 n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , 
 n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , 
 n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , 
 n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , 
 n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , 
 n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , 
 n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , 
 n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , 
 n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , 
 n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , 
 n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , 
 n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , 
 n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , 
 n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , 
 n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , 
 n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , 
 n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , 
 n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , 
 n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , 
 n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , 
 n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , 
 n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , 
 n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , 
 n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , 
 n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , 
 n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , 
 n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , 
 n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , 
 n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , 
 n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , 
 n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , 
 n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , 
 n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , 
 n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , 
 n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , 
 n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , 
 n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , 
 n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , 
 n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , 
 n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , 
 n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , 
 n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , 
 n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , 
 n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , 
 n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , 
 n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , 
 n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , 
 n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , 
 n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , 
 n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , 
 n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , 
 n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , 
 n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , 
 n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , 
 n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , 
 n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , 
 n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , 
 n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , 
 n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , 
 n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , 
 n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , 
 n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , 
 n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , 
 n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , 
 n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , 
 n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , 
 n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , 
 n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , 
 n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , 
 n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , 
 n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , 
 n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , 
 n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , 
 n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , 
 n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , 
 n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , 
 n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , 
 n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , 
 n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , 
 n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , 
 n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , 
 n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , 
 n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , 
 n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , 
 n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , 
 n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , 
 n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , 
 n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , 
 n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , 
 n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , 
 n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , 
 n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , 
 n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , 
 n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , 
 n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , 
 n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , 
 n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , 
 n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , 
 n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , 
 n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , 
 n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , 
 n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , 
 n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , 
 n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , 
 n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , 
 n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , 
 n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , 
 n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , 
 n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , 
 n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , 
 n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , 
 n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , 
 n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , 
 n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , 
 n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , 
 n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , 
 n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , 
 n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , 
 n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , 
 n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , 
 n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , 
 n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , 
 n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , 
 n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , 
 n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , 
 n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , 
 n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , 
 n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , 
 n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , 
 n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , 
 n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , 
 n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , 
 n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , 
 n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , 
 n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , 
 n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , 
 n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , 
 n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , 
 n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , 
 n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , 
 n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , 
 n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , 
 n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , 
 n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , 
 n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , 
 n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , 
 n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , 
 n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , 
 n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , 
 n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , 
 n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , 
 n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , 
 n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , 
 n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , 
 n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , 
 n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , 
 n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , 
 n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , 
 n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , 
 n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , 
 n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , 
 n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , 
 n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , 
 n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , 
 n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , 
 n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , 
 n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , 
 n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , 
 n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , 
 n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , 
 n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , 
 n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , 
 n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , 
 n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , 
 n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , 
 n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , 
 n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , 
 n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , 
 n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , 
 n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , 
 n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , 
 n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , 
 n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , 
 n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , 
 n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , 
 n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , 
 n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , 
 n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , 
 n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , 
 n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , 
 n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , 
 n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , 
 n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , 
 n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , 
 n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , 
 n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , 
 n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , 
 n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , 
 n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , 
 n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , 
 n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , 
 n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , 
 n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , 
 n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , 
 n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , 
 n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , 
 n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , 
 n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , 
 n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , 
 n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , 
 n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , 
 n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , 
 n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , 
 n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , 
 n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , 
 n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , 
 n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , 
 n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , 
 n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , 
 n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , 
 n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , 
 n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , 
 n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , 
 n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , 
 n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , 
 n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , 
 n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , 
 n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , 
 n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , 
 n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , 
 n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , 
 n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , 
 n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , 
 n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , 
 n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , 
 n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , 
 n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , 
 n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , 
 n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , 
 n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , 
 n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , 
 n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , 
 n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , 
 n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , 
 n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , 
 n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , 
 n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , 
 n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , 
 n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , 
 n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , 
 n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , 
 n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , 
 n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , 
 n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , 
 n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , 
 n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , 
 n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , 
 n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , 
 n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , 
 n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , 
 n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , 
 n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , 
 n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , 
 n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , 
 n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , 
 n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , 
 n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , 
 n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , 
 n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , 
 n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , 
 n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , 
 n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , 
 n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , 
 n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , 
 n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , 
 n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , 
 n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , 
 n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , 
 n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , 
 n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , 
 n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , 
 n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , 
 n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , 
 n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , 
 n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , 
 n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , 
 n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , 
 n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , 
 n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , 
 n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , 
 n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , 
 n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , 
 n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , 
 n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , 
 n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , 
 n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , 
 n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , 
 n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , 
 n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , 
 n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , 
 n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , 
 n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , 
 n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , 
 n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , 
 n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , 
 n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , 
 n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , 
 n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , 
 n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , 
 n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , 
 n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , 
 n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , 
 n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , 
 n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , 
 n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , 
 n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , 
 n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , 
 n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , 
 n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , 
 n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , 
 n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , 
 n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , 
 n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , 
 n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , 
 n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , 
 n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , 
 n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , 
 n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , 
 n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , 
 n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , 
 n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , 
 n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , 
 n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , 
 n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , 
 n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , 
 n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , 
 n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , 
 n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , 
 n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , 
 n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , 
 n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , 
 n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , 
 n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , 
 n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , 
 n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , 
 n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , 
 n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , 
 n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , 
 n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , 
 n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , 
 n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , 
 n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , 
 n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , 
 n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , 
 n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , 
 n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , 
 n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , 
 n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , 
 n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , 
 n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , 
 n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , 
 n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , 
 n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , 
 n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , 
 n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , 
 n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , 
 n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , 
 n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , 
 n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , 
 n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , 
 n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , 
 n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , 
 n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , 
 n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , 
 n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , 
 n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , 
 n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , 
 n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , 
 n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , 
 n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , 
 n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , 
 n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , 
 n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , 
 n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , 
 n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , 
 n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , 
 n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , 
 n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , 
 n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , 
 n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , 
 n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , 
 n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , 
 n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , 
 n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , 
 n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , 
 n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , 
 n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , 
 n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , 
 n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , 
 n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , 
 n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , 
 n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , 
 n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , 
 n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , 
 n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , 
 n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , 
 n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , 
 n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , 
 n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , 
 n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , 
 n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , 
 n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , 
 n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , 
 n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , 
 n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , 
 n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , 
 n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , 
 n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , 
 n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , 
 n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , 
 n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , 
 n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , 
 n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , 
 n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , 
 n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , 
 n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , 
 n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , 
 n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , 
 n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , 
 n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , 
 n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , 
 n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , 
 n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , 
 n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , 
 n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , 
 n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , 
 n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , 
 n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , 
 n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , 
 n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , 
 n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , 
 n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , 
 n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , 
 n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , 
 n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , 
 n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , 
 n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , 
 n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , 
 n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , 
 n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , 
 n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , 
 n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , 
 n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , 
 n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , 
 n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , 
 n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , 
 n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , 
 n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , 
 n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , 
 n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , 
 n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , 
 n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , 
 n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , 
 n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , 
 n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , 
 n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , 
 n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , 
 n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , 
 n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , 
 n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , 
 n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , 
 n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , 
 n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , 
 n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , 
 n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , 
 n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , 
 n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , 
 n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , 
 n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , 
 n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , 
 n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , 
 n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , 
 n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , 
 n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , 
 n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , 
 n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , 
 n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , 
 n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , 
 n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , 
 n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , 
 n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , 
 n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , 
 n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , 
 n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , 
 n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , 
 n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , 
 n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , 
 n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , 
 n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , 
 n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , 
 n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , 
 n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , 
 n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , 
 n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , 
 n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , 
 n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , 
 n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , 
 n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , 
 n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , 
 n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , 
 n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , 
 n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , 
 n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , 
 n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , 
 n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , 
 n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , 
 n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , 
 n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , 
 n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , 
 n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , 
 n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , 
 n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , 
 n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , 
 n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , 
 n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , 
 n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , 
 n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , 
 n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , 
 n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , 
 n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , 
 n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , 
 n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , 
 n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , 
 n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , 
 n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , 
 n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , 
 n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , 
 n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , 
 n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , 
 n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , 
 n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , 
 n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , 
 n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , 
 n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , 
 n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , 
 n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , 
 n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , 
 n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , 
 n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , 
 n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , 
 n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , 
 n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , 
 n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , 
 n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , 
 n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , 
 n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , 
 n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , 
 n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , 
 n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , 
 n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , 
 n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , 
 n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , 
 n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , 
 n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , 
 n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , 
 n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , 
 n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , 
 n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , 
 n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , 
 n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , 
 n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , 
 n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , 
 n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , 
 n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , 
 n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , 
 n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , 
 n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , 
 n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , 
 n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , 
 n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , 
 n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , 
 n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , 
 n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , 
 n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , 
 n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , 
 n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , 
 n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , 
 n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , 
 n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , 
 n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , 
 n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , 
 n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , 
 n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , 
 n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , 
 n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , 
 n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , 
 n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , 
 n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , 
 n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , 
 n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , 
 n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , 
 n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , 
 n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , 
 n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , 
 n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , 
 n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , 
 n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , 
 n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , 
 n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , 
 n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , 
 n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , 
 n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , 
 n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , 
 n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , 
 n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , 
 n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , 
 n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , 
 n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , 
 n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , 
 n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , 
 n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , 
 n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , 
 n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , 
 n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , 
 n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , 
 n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , 
 n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , 
 n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , 
 n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , 
 n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , 
 n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , 
 n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , 
 n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , 
 n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , 
 n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , 
 n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , 
 n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , 
 n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , 
 n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , 
 n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , 
 n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , 
 n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , 
 n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , 
 n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , 
 n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , 
 n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , 
 n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , 
 n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , 
 n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , 
 n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , 
 n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , 
 n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , 
 n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , 
 n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , 
 n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , 
 n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , 
 n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , 
 n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , 
 n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , 
 n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , 
 n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , 
 n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , 
 n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , 
 n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , 
 n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , 
 n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , 
 n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , 
 n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , 
 n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , 
 n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , 
 n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , 
 n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , 
 n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , 
 n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , 
 n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , 
 n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , 
 n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , 
 n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , 
 n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , 
 n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , 
 n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , 
 n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , 
 n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , 
 n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , 
 n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , 
 n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , 
 n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , 
 n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , 
 n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , 
 n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , 
 n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , 
 n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , 
 n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , 
 n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , 
 n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , 
 n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , 
 n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , 
 n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , 
 n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , 
 n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , 
 n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , 
 n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , 
 n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , 
 n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , 
 n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , 
 n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , 
 n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , 
 n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , 
 n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , 
 n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , 
 n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , 
 n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , 
 n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , 
 n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , 
 n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , 
 n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , 
 n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , 
 n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , 
 n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , 
 n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , 
 n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , 
 n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , 
 n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , 
 n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , 
 n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , 
 n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , 
 n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , 
 n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , 
 n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , 
 n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , 
 n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , 
 n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , 
 n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , 
 n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , 
 n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , 
 n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , 
 n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , 
 n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , 
 n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , 
 n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , 
 n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , 
 n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , 
 n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , 
 n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , 
 n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , 
 n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , 
 n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , 
 n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , 
 n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , 
 n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , 
 n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , 
 n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , 
 n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , 
 n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , 
 n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , 
 n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , 
 n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , 
 n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , 
 n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , 
 n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , 
 n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , 
 n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , 
 n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , 
 n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , 
 n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , 
 n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , 
 n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , 
 n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , 
 n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , 
 n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , 
 n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , 
 n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , 
 n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , 
 n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , 
 n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , 
 n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , 
 n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , 
 n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , 
 n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , 
 n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , 
 n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , 
 n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , 
 n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , 
 n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , 
 n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , 
 n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , 
 n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , 
 n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , 
 n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , 
 n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , 
 n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , 
 n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , 
 n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , 
 n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , 
 n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , 
 n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , 
 n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , 
 n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , 
 n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , 
 n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , 
 n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , 
 n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , 
 n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , 
 n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , 
 n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , 
 n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , 
 n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , 
 n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , 
 n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , 
 n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , 
 n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , 
 n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , 
 n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , 
 n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , 
 n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , 
 n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , 
 n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , 
 n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , 
 n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , 
 n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , 
 n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , 
 n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , 
 n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , 
 n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , 
 n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , 
 n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , 
 n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , 
 n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , 
 n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , 
 n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , 
 n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , 
 n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , 
 n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , 
 n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , 
 n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , 
 n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , 
 n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , 
 n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , 
 n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , 
 n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , 
 n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , 
 n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , 
 n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , 
 n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , 
 n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , 
 n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , 
 n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , 
 n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , 
 n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , 
 n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , 
 n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , 
 n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , 
 n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , 
 n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , 
 n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , 
 n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , 
 n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , 
 n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , 
 n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , 
 n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , 
 n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , 
 n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , 
 n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , 
 n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , 
 n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , 
 n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , 
 n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , 
 n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , 
 n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , 
 n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , 
 n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , 
 n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , 
 n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , 
 n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , 
 n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , 
 n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , 
 n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , 
 n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , 
 n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , 
 n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , 
 n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , 
 n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , 
 n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , 
 n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , 
 n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , 
 n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , 
 n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , 
 n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , 
 n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , 
 n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , 
 n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , 
 n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , 
 n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , 
 n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , 
 n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , 
 n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , 
 n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , 
 n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , 
 n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , 
 n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , 
 n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , 
 n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , 
 n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , 
 n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , 
 n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , 
 n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , 
 n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , 
 n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , 
 n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , 
 n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , 
 n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , 
 n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , 
 n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , 
 n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , 
 n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , 
 n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , 
 n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , 
 n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , 
 n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , 
 n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , 
 n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , 
 n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , 
 n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , 
 n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , 
 n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , 
 n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , 
 n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , 
 n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , 
 n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , 
 n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , 
 n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , 
 n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , 
 n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , 
 n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , 
 n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , 
 n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , 
 n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , 
 n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , 
 n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , 
 n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , 
 n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , 
 n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , 
 n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , 
 n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , 
 n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , 
 n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , 
 n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , 
 n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , 
 n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , 
 n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , 
 n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , 
 n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , 
 n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , 
 n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , 
 n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , 
 n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , 
 n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , 
 n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , 
 n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , 
 n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , 
 n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , 
 n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , 
 n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , 
 n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , 
 n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , 
 n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , 
 n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , 
 n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , 
 n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , 
 n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , 
 n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , 
 n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , 
 n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , 
 n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , 
 n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , 
 n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , 
 n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , 
 n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , 
 n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , 
 n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , 
 n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , 
 n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , 
 n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , 
 n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , 
 n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , 
 n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , 
 n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , 
 n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , 
 n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , 
 n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , 
 n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , 
 n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , 
 n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , 
 n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , 
 n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , 
 n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , 
 n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , 
 n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , 
 n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , 
 n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , 
 n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , 
 n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , 
 n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , 
 n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , 
 n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , 
 n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , 
 n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , 
 n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , 
 n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , 
 n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , 
 n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , 
 n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , 
 n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , 
 n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , 
 n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , 
 n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , 
 n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , 
 n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , 
 n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , 
 n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , 
 n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , 
 n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , 
 n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , 
 n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , 
 n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , 
 n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , 
 n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , 
 n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , 
 n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , 
 n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , 
 n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , 
 n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , 
 n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , 
 n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , 
 n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , 
 n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , 
 n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , 
 n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , 
 n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , 
 n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , 
 n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , 
 n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , 
 n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , 
 n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , 
 n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , 
 n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , 
 n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , 
 n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , 
 n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , 
 n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , 
 n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , 
 n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , 
 n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , 
 n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , 
 n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , 
 n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , 
 n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , 
 n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , 
 n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , 
 n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , 
 n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , 
 n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , 
 n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , 
 n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , 
 n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , 
 n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , 
 n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , 
 n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , 
 n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , 
 n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , 
 n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , 
 n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , 
 n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , 
 n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , 
 n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , 
 n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , 
 n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , 
 n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , 
 n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , 
 n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , 
 n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , 
 n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , 
 n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , 
 n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , 
 n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , 
 n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , 
 n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , 
 n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , 
 n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , 
 n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , 
 n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , 
 n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , 
 n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , 
 n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , 
 n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , 
 n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , 
 n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , 
 n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , 
 n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , 
 n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , 
 n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , 
 n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , 
 n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , 
 n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , 
 n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , 
 n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , 
 n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , 
 n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , 
 n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , 
 n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , 
 n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , 
 n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , 
 n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , 
 n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , 
 n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , 
 n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , 
 n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , 
 n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , 
 n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , 
 n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , 
 n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , 
 n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , 
 n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , 
 n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , 
 n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , 
 n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , 
 n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , 
 n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , 
 n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , 
 n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , 
 n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , 
 n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , 
 n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , 
 n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , 
 n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , 
 n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , 
 n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , 
 n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , 
 n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , 
 n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , 
 n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , 
 n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , 
 n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , 
 n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , 
 n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , 
 n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , 
 n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , 
 n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , 
 n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , 
 n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , 
 n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , 
 n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , 
 n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , 
 n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , 
 n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , 
 n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , 
 n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , 
 n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , 
 n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , 
 n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , 
 n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , 
 n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , 
 n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , 
 n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , 
 n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , 
 n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , 
 n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , 
 n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , 
 n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , 
 n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , 
 n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , 
 n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , 
 n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , 
 n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , 
 n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , 
 n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , 
 n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , 
 n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , 
 n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , 
 n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , 
 n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , 
 n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , 
 n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , 
 n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , 
 n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , 
 n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , 
 n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , 
 n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , 
 n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , 
 n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , 
 n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , 
 n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , 
 n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , 
 n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , 
 n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , 
 n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , 
 n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , 
 n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , 
 n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , 
 n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , 
 n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , 
 n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , 
 n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , 
 n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , 
 n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , 
 n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , 
 n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , 
 n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , 
 n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , 
 n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , 
 n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , 
 n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , 
 n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , 
 n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , 
 n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , 
 n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , 
 n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , 
 n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , 
 n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , 
 n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , 
 n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , 
 n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , 
 n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , 
 n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , 
 n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , 
 n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , 
 n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , 
 n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , 
 n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , 
 n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , 
 n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , 
 n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , 
 n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , 
 n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , 
 n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , 
 n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , 
 n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , 
 n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , 
 n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , 
 n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , 
 n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , 
 n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , 
 n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , 
 n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , 
 n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , 
 n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , 
 n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , 
 n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , 
 n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , 
 n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , 
 n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , 
 n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , 
 n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , 
 n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , 
 n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , 
 n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , 
 n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , 
 n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , 
 n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , 
 n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , 
 n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , 
 n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , 
 n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , 
 n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , 
 n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , 
 n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , 
 n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , 
 n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , 
 n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , 
 n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , 
 n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , 
 n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , 
 n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , 
 n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , 
 n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , 
 n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , 
 n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , 
 n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , 
 n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , 
 n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , 
 n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , 
 n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , 
 n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , 
 n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , 
 n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , 
 n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , 
 n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , 
 n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , 
 n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , 
 n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , 
 n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , 
 n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , 
 n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , 
 n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , 
 n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , 
 n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , 
 n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , 
 n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , 
 n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , 
 n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , 
 n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , 
 n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , 
 n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , 
 n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , 
 n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , 
 n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , 
 n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , 
 n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , 
 n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , 
 n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , 
 n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , 
 n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , 
 n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , 
 n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , 
 n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , 
 n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , 
 n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , 
 n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , 
 n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , 
 n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , 
 n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , 
 n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , 
 n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , 
 n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , 
 n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , 
 n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , 
 n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , 
 n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , 
 n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , 
 n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , 
 n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , 
 n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , 
 n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , 
 n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , 
 n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , 
 n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , 
 n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , 
 n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , 
 n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , 
 n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , 
 n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , 
 n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , 
 n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , 
 n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , 
 n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , 
 n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , 
 n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , 
 n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , 
 n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , 
 n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , 
 n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , 
 n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , 
 n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , 
 n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , 
 n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , 
 n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , 
 n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , 
 n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , 
 n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , 
 n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , 
 n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , 
 n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , 
 n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , 
 n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , 
 n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , 
 n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , 
 n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , 
 n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , 
 n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , 
 n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , 
 n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , 
 n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , 
 n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , 
 n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , 
 n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , 
 n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , 
 n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , 
 n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , 
 n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , 
 n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , 
 n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , 
 n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , 
 n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , 
 n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , 
 n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , 
 n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , 
 n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , 
 n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , 
 n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , 
 n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , 
 n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , 
 n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , 
 n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , 
 n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , 
 n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , 
 n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , 
 n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , 
 n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , 
 n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , 
 n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , 
 n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , 
 n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , 
 n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , 
 n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , 
 n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , 
 n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , 
 n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , 
 n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , 
 n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , 
 n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , 
 n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , 
 n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , 
 n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , 
 n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , 
 n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , 
 n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , 
 n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , 
 n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , 
 n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , 
 n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , 
 n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , 
 n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , 
 n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , 
 n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , 
 n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , 
 n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , 
 n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , 
 n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , 
 n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , 
 n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , 
 n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , 
 n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , 
 n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , 
 n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , 
 n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , 
 n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , 
 n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , 
 n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , 
 n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , 
 n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , 
 n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , 
 n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , 
 n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , 
 n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , 
 n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , 
 n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , 
 n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , 
 n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , 
 n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , 
 n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , 
 n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , 
 n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , 
 n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , 
 n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , 
 n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , 
 n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , 
 n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , 
 n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , 
 n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , 
 n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , 
 n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , 
 n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , 
 n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , 
 n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , 
 n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , 
 n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , 
 n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , 
 n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , 
 n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , 
 n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , 
 n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , 
 n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , 
 n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , 
 n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , 
 n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , 
 n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , 
 n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , 
 n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , 
 n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , 
 n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , 
 n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , 
 n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , 
 n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , 
 n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , 
 n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , 
 n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , 
 n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , 
 n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , 
 n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , 
 n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , 
 n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , 
 n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , 
 n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , 
 n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , 
 n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , 
 n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , 
 n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , 
 n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , 
 n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , 
 n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , 
 n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , 
 n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , 
 n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , 
 n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , 
 n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , 
 n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , 
 n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , 
 n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , 
 n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , 
 n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , 
 n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , 
 n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , 
 n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , 
 n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , 
 n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , 
 n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , 
 n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , 
 n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , 
 n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , 
 n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , 
 n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , 
 n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , 
 n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , 
 n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , 
 n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , 
 n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , 
 n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , 
 n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , 
 n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , 
 n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , 
 n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , 
 n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , 
 n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , 
 n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , 
 n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , 
 n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , 
 n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , 
 n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , 
 n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , 
 n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , 
 n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , 
 n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , 
 n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , 
 n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , 
 n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , 
 n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , 
 n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , 
 n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , 
 n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , 
 n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , 
 n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , 
 n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , 
 n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , 
 n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , 
 n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , 
 n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , 
 n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , 
 n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , 
 n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , 
 n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , 
 n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , 
 n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , 
 n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , 
 n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , 
 n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , 
 n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , 
 n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , 
 n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , 
 n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , 
 n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , 
 n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , 
 n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , 
 n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , 
 n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , 
 n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , 
 n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , 
 n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , 
 n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , 
 n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , 
 n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , 
 n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , 
 n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , 
 n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , 
 n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , 
 n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , 
 n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , 
 n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , 
 n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , 
 n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , 
 n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , 
 n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , 
 n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , 
 n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , 
 n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , 
 n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , 
 n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , 
 n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , 
 n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , 
 n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , 
 n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , 
 n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , 
 n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , 
 n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , 
 n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , 
 n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , 
 n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , 
 n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , 
 n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , 
 n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , 
 n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , 
 n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , 
 n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , 
 n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , 
 n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , 
 n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , 
 n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , 
 n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , 
 n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , 
 n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , 
 n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , 
 n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , 
 n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , 
 n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , 
 n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , 
 n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , 
 n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , 
 n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , 
 n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , 
 n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , 
 n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , 
 n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , 
 n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , 
 n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , 
 n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , 
 n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , 
 n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , 
 n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , 
 n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , 
 n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , 
 n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , 
 n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , 
 n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , 
 n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , 
 n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , 
 n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , 
 n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , 
 n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , 
 n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , 
 n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , 
 n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , 
 n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , 
 n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , 
 n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , 
 n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , 
 n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , 
 n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , 
 n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , 
 n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , 
 n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , 
 n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , 
 n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , 
 n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , 
 n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , 
 n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , 
 n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , 
 n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , 
 n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , 
 n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , 
 n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , 
 n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , 
 n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , 
 n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , 
 n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , 
 n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , 
 n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , 
 n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , 
 n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , 
 n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , 
 n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , 
 n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , 
 n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , 
 n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , 
 n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , 
 n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , 
 n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , 
 n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , 
 n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , 
 n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , 
 n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , 
 n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , 
 n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , 
 n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , 
 n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , 
 n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , 
 n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , 
 n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , 
 n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , 
 n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , 
 n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , 
 n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , 
 n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , 
 n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , 
 n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , 
 n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , 
 n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , 
 n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , 
 n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , 
 n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , 
 n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , 
 n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , 
 n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , 
 n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , 
 n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , 
 n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , 
 n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , 
 n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , 
 n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , 
 n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , 
 n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , 
 n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , 
 n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , 
 n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , 
 n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , 
 n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , 
 n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , 
 n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , 
 n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , 
 n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , 
 n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , 
 n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , 
 n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , 
 n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , 
 n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , 
 n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , 
 n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , 
 n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , 
 n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , 
 n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , 
 n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , 
 n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , 
 n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , 
 n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , 
 n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , 
 n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , 
 n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , 
 n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , 
 n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , 
 n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , 
 n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , 
 n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , 
 n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , 
 n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , 
 n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , 
 n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , 
 n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , 
 n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , 
 n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , 
 n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , 
 n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , 
 n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , 
 n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , 
 n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , 
 n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , 
 n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , 
 n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , 
 n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , 
 n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , 
 n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , 
 n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , 
 n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , 
 n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , 
 n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , 
 n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , 
 n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , 
 n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , 
 n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , 
 n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , 
 n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , 
 n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , 
 n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , 
 n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , 
 n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , 
 n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , 
 n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , 
 n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , 
 n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , 
 n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , 
 n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , 
 n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , 
 n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , 
 n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , 
 n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , 
 n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , 
 n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , 
 n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , 
 n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , 
 n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , 
 n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , 
 n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , 
 n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , 
 n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , 
 n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , 
 n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , 
 n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , 
 n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , 
 n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , 
 n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , 
 n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , 
 n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , 
 n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , 
 n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , 
 n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , 
 n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , 
 n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , 
 n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , 
 n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , 
 n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , 
 n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , 
 n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , 
 n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , 
 n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , 
 n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , 
 n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , 
 n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , 
 n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , 
 n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , 
 n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , 
 n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , 
 n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , 
 n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , 
 n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , 
 n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , 
 n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , 
 n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , 
 n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , 
 n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , 
 n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , 
 n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , 
 n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , 
 n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , 
 n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , 
 n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , 
 n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , 
 n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , 
 n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , 
 n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , 
 n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , 
 n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , 
 n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , 
 n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , 
 n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , 
 n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , 
 n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , 
 n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , 
 n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , 
 n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , 
 n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , 
 n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , 
 n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , 
 n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , 
 n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , 
 n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , 
 n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , 
 n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , 
 n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , 
 n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , 
 n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , 
 n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , 
 n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , 
 n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , 
 n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , 
 n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , 
 n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , 
 n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , 
 n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , 
 n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , 
 n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , 
 n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , 
 n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , 
 n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , 
 n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , 
 n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , 
 n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , 
 n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , 
 n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , 
 n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , 
 n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , 
 n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , 
 n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , 
 n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , 
 n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , 
 n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , 
 n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , 
 n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , 
 n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , 
 n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , 
 n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , 
 n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , 
 n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , 
 n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , 
 n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , 
 n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , 
 n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , 
 n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , 
 n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , 
 n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , 
 n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , 
 n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , 
 n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , 
 n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , 
 n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , 
 n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , 
 n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , 
 n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , 
 n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , 
 n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , 
 n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , 
 n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , 
 n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , 
 n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , 
 n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , 
 n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , 
 n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , 
 n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , 
 n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , 
 n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , 
 n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , 
 n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , 
 n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , 
 n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , 
 n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , 
 n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , 
 n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , 
 n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , 
 n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , 
 n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , 
 n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , 
 n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , 
 n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , 
 n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , 
 n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , 
 n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , 
 n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , 
 n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , 
 n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , 
 n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , 
 n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , 
 n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , 
 n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , 
 n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , 
 n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , 
 n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , 
 n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , 
 n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , 
 n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , 
 n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , 
 n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , 
 n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , 
 n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , 
 n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , 
 n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , 
 n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , 
 n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , 
 n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , 
 n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , 
 n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , 
 n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , 
 n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , 
 n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , 
 n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , 
 n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , 
 n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , 
 n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , 
 n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , 
 n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , 
 n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , 
 n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , 
 n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , 
 n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , 
 n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , 
 n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , 
 n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , 
 n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , 
 n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , 
 n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , 
 n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , 
 n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , 
 n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , 
 n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , 
 n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , 
 n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , 
 n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , 
 n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , 
 n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , 
 n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , 
 n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , 
 n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , 
 n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , 
 n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , 
 n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , 
 n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , 
 n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , 
 n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , 
 n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , 
 n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , 
 n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , 
 n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , 
 n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , 
 n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , 
 n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , 
 n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , 
 n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , 
 n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , 
 n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , 
 n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , 
 n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , 
 n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , 
 n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , 
 n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , 
 n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , 
 n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , 
 n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , 
 n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , 
 n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , 
 n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , 
 n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , 
 n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , 
 n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , 
 n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , 
 n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , 
 n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , 
 n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , 
 n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , 
 n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , 
 n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , 
 n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , 
 n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , 
 n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , 
 n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , 
 n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , 
 n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , 
 n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , 
 n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , 
 n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , 
 n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , 
 n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , 
 n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , 
 n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , 
 n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , 
 n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , 
 n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , 
 n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , 
 n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , 
 n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , 
 n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , 
 n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , 
 n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , 
 n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , 
 n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , 
 n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , 
 n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , 
 n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , 
 n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , 
 n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , 
 n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , 
 n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , 
 n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , 
 n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , 
 n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , 
 n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , 
 n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , 
 n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , 
 n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , 
 n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , 
 n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , 
 n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , 
 n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , 
 n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , 
 n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , 
 n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , 
 n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , 
 n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , 
 n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , 
 n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , 
 n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , 
 n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , 
 n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , 
 n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , 
 n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , 
 n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , 
 n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , 
 n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , 
 n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , 
 n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , 
 n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , 
 n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , 
 n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , 
 n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , 
 n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , 
 n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , 
 n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , 
 n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , 
 n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , 
 n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , 
 n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , 
 n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , 
 n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , 
 n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , 
 n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , 
 n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , 
 n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , 
 n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , 
 n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , 
 n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , 
 n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , 
 n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , 
 n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , 
 n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , 
 n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , 
 n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , 
 n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , 
 n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , 
 n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , 
 n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , 
 n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , 
 n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , 
 n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , 
 n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , 
 n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , 
 n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , 
 n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , 
 n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , 
 n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , 
 n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , 
 n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , 
 n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , 
 n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , 
 n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , 
 n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , 
 n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , 
 n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , 
 n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , 
 n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , 
 n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , 
 n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , 
 n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , 
 n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , 
 n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , 
 n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , 
 n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , 
 n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , 
 n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , 
 n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , 
 n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , 
 n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , 
 n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , 
 n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , 
 n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , 
 n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , 
 n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , 
 n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , 
 n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , 
 n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , 
 n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , 
 n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , 
 n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , 
 n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , 
 n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , 
 n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , 
 n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , 
 n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , 
 n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , 
 n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , 
 n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , 
 n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , 
 n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , 
 n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , 
 n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , 
 n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , 
 n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , 
 n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , 
 n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , 
 n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , 
 n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , 
 n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , 
 n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , 
 n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , 
 n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , 
 n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , 
 n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , 
 n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , 
 n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , 
 n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , 
 n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , 
 n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , 
 n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , 
 n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , 
 n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , 
 n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , 
 n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , 
 n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , 
 n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , 
 n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , 
 n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , 
 n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , 
 n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , 
 n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , 
 n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , 
 n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , 
 n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , 
 n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , 
 n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , 
 n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , 
 n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , 
 n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , 
 n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , 
 n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , 
 n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , 
 n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , 
 n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , 
 n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , 
 n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , 
 n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , 
 n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , 
 n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , 
 n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , 
 n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , 
 n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , 
 n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , 
 n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , 
 n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , 
 n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , 
 n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , 
 n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , 
 n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , 
 n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , 
 n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , 
 n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , 
 n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , 
 n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , 
 n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , 
 n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , 
 n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , 
 n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , 
 n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , 
 n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , 
 n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , 
 n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , 
 n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , 
 n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , 
 n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , 
 n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , 
 n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , 
 n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , 
 n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , 
 n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , 
 n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , 
 n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , 
 n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , 
 n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , 
 n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , 
 n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , 
 n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , 
 n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , 
 n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , 
 n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , 
 n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , 
 n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , 
 n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , 
 n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , 
 n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , 
 n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , 
 n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , 
 n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , 
 n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , 
 n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , 
 n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , 
 n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , 
 n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , 
 n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , 
 n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , 
 n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , 
 n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , 
 n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , 
 n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , 
 n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , 
 n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , 
 n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , 
 n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , 
 n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , 
 n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , 
 n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , 
 n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , 
 n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , 
 n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , 
 n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , 
 n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , 
 n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , 
 n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , 
 n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , 
 n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , 
 n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , 
 n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , 
 n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , 
 n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , 
 n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , 
 n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , 
 n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , 
 n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , 
 n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , 
 n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , 
 n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , 
 n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , 
 n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , 
 n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , 
 n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , 
 n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , 
 n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , 
 n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , 
 n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , 
 n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , 
 n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , 
 n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , 
 n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , 
 n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , 
 n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , 
 n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , 
 n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , 
 n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , 
 n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , 
 n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , 
 n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , 
 n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , 
 n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , 
 n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , 
 n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , 
 n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , 
 n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , 
 n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , 
 n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , 
 n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , 
 n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , 
 n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , 
 n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , 
 n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , 
 n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , 
 n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , 
 n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , 
 n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , 
 n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , 
 n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , 
 n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , 
 n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , 
 n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , 
 n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , 
 n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , 
 n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , 
 n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , 
 n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , 
 n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , 
 n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , 
 n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , 
 n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , 
 n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , 
 n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , 
 n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , 
 n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , 
 n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , 
 n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , 
 n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , 
 n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , 
 n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , 
 n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , 
 n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , 
 n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , 
 n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , 
 n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , 
 n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , 
 n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , 
 n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , 
 n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , 
 n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , 
 n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , 
 n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , 
 n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , 
 n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , 
 n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , 
 n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , 
 n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , 
 n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , 
 n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , 
 n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , 
 n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , 
 n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , 
 n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , 
 n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , 
 n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , 
 n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , 
 n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , 
 n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , 
 n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , 
 n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , 
 n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , 
 n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , 
 n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , 
 n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , 
 n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , 
 n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , 
 n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , 
 n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , 
 n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , 
 n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , 
 n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , 
 n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , 
 n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , 
 n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , 
 n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , 
 n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , 
 n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , 
 n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , 
 n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , 
 n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , 
 n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , 
 n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , 
 n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , 
 n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , 
 n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , 
 n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , 
 n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , 
 n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , 
 n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , 
 n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , 
 n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , 
 n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , 
 n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , 
 n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , 
 n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , 
 n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , 
 n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , 
 n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , 
 n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , 
 n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , 
 n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , 
 n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , 
 n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , 
 n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , 
 n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , 
 n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , 
 n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , 
 n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , 
 n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , 
 n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , 
 n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , 
 n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , 
 n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , 
 n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , 
 n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , 
 n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , 
 n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , 
 n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , 
 n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , 
 n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , 
 n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , 
 n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , 
 n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , 
 n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , 
 n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , 
 n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , 
 n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , 
 n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , 
 n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , 
 n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , 
 n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , 
 n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , 
 n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , 
 n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , 
 n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , 
 n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , 
 n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , 
 n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , 
 n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , 
 n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , 
 n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , 
 n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , 
 n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , 
 n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , 
 n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , 
 n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , 
 n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , 
 n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , 
 n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , 
 n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , 
 n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , 
 n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , 
 n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , 
 n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , 
 n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , 
 n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , 
 n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , 
 n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , 
 n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , 
 n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , 
 n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , 
 n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , 
 n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , 
 n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , 
 n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , 
 n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , 
 n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , 
 n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , 
 n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , 
 n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , 
 n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , 
 n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , 
 n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , 
 n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , 
 n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , 
 n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , 
 n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , 
 n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , 
 n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , 
 n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , 
 n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , 
 n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , 
 n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , 
 n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , 
 n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , 
 n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , 
 n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , 
 n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , 
 n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , 
 n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , 
 n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , 
 n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , 
 n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , 
 n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , 
 n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , 
 n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , 
 n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , 
 n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , 
 n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , 
 n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , 
 n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , 
 n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , 
 n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , 
 n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , 
 n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , 
 n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , 
 n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , 
 n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , 
 n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , 
 n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , 
 n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , 
 n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , 
 n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , 
 n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , 
 n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , 
 n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , 
 n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , 
 n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , 
 n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , 
 n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , 
 n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , 
 n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , 
 n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , 
 n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , 
 n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , 
 n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , 
 n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , 
 n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , 
 n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , 
 n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , 
 n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , 
 n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , 
 n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , 
 n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , 
 n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , 
 n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , 
 n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , 
 n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , 
 n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , 
 n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , 
 n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , 
 n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , 
 n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , 
 n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , 
 n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , 
 n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , 
 n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , 
 n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , 
 n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , 
 n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , 
 n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , 
 n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , 
 n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , 
 n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , 
 n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , 
 n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , 
 n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , 
 n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , 
 n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , 
 n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , 
 n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , 
 n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , 
 n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , 
 n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , 
 n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , 
 n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , 
 n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , 
 n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , 
 n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , 
 n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , 
 n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , 
 n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , 
 n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , 
 n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , 
 n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , 
 n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , 
 n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , 
 n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , 
 n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , 
 n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , 
 n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , 
 n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , 
 n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , 
 n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , 
 n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , 
 n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , 
 n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , 
 n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , 
 n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , 
 n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , 
 n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , 
 n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , 
 n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , 
 n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , 
 n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , 
 n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , 
 n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , 
 n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , 
 n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , 
 n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , 
 n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , 
 n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , 
 n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , 
 n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , 
 n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , 
 n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , 
 n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , 
 n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , 
 n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , 
 n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , 
 n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , 
 n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , 
 n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , 
 n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , 
 n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , 
 n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , 
 n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , 
 n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , 
 n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , 
 n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , 
 n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , 
 n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , 
 n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , 
 n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , 
 n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , 
 n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , 
 n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , 
 n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , 
 n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , 
 n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , 
 n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , 
 n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , 
 n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , 
 n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , 
 n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , 
 n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , 
 n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , 
 n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , 
 n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , 
 n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , 
 n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , 
 n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , 
 n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , 
 n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , 
 n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , 
 n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , 
 n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , 
 n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , 
 n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , 
 n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , 
 n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , 
 n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , 
 n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , 
 n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , 
 n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , 
 n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , 
 n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , 
 n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , 
 n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , 
 n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , 
 n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , 
 n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , 
 n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , 
 n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , 
 n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , 
 n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , 
 n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , 
 n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , 
 n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , 
 n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , 
 n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , 
 n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , 
 n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , 
 n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , 
 n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , 
 n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , 
 n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , 
 n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , 
 n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , 
 n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , 
 n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , 
 n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , 
 n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , 
 n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , 
 n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , 
 n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , 
 n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , 
 n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , 
 n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , 
 n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , 
 n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , 
 n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , 
 n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , 
 n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , 
 n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , 
 n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , 
 n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , 
 n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , 
 n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , 
 n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , 
 n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , 
 n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , 
 n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , 
 n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , 
 n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , 
 n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , 
 n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , 
 n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , 
 n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , 
 n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , 
 n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , 
 n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , 
 n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , 
 n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , 
 n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , 
 n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , 
 n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , 
 n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , 
 n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , 
 n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , 
 n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , 
 n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , 
 n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , 
 n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , 
 n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , 
 n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , 
 n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , 
 n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , 
 n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , 
 n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , 
 n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , 
 n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , 
 n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , 
 n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , 
 n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , 
 n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , 
 n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , 
 n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , 
 n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , 
 n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , 
 n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , 
 n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , 
 n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , 
 n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , 
 n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , 
 n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , 
 n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , 
 n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , 
 n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , 
 n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , 
 n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , 
 n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , 
 n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , 
 n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , 
 n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , 
 n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , 
 n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , 
 n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , 
 n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , 
 n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , 
 n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , 
 n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , 
 n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , 
 n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , 
 n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , 
 n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , 
 n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , 
 n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , 
 n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , 
 n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , 
 n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , 
 n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , 
 n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , 
 n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , 
 n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , 
 n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , 
 n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , 
 n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , 
 n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , 
 n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , 
 n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , 
 n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , 
 n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , 
 n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , 
 n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , 
 n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , 
 n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , 
 n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , 
 n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , 
 n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , 
 n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , 
 n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , 
 n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , 
 n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , 
 n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , 
 n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , 
 n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , 
 n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , 
 n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , 
 n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , 
 n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , 
 n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , 
 n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , 
 n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , 
 n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , 
 n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , 
 n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , 
 n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , 
 n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , 
 n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , 
 n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , 
 n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , 
 n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , 
 n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , 
 n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , 
 n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , 
 n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , 
 n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , 
 n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , 
 n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , 
 n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , 
 n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , 
 n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , 
 n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , 
 n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , 
 n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , 
 n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , 
 n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , 
 n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , 
 n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , 
 n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , 
 n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , 
 n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , 
 n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , 
 n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , 
 n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , 
 n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , 
 n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , 
 n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , 
 n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , 
 n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , 
 n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , 
 n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , 
 n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , 
 n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , 
 n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , 
 n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , 
 n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , 
 n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , 
 n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , 
 n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , 
 n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , 
 n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , 
 n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , 
 n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , 
 n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , 
 n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , 
 n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , 
 n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , 
 n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , 
 n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , 
 n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , 
 n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , 
 n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , 
 n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , 
 n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , 
 n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , 
 n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , 
 n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , 
 n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , 
 n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , 
 n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , 
 n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , 
 n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , 
 n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , 
 n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , 
 n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , 
 n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , 
 n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , 
 n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , 
 n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , 
 n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , 
 n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , 
 n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , 
 n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , 
 n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , 
 n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , 
 n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , 
 n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , 
 n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , 
 n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , 
 n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , 
 n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , 
 n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , 
 n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , 
 n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , 
 n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , 
 n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , 
 n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , 
 n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , 
 n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , 
 n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , 
 n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , 
 n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , 
 n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , 
 n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , 
 n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , 
 n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , 
 n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , 
 n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , 
 n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , 
 n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , 
 n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , 
 n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , 
 n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , 
 n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , 
 n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , 
 n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , 
 n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , 
 n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , 
 n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , 
 n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , 
 n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , 
 n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , 
 n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , 
 n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , 
 n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , 
 n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , 
 n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , 
 n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , 
 n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , 
 n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , 
 n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , 
 n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , 
 n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , 
 n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , 
 n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , 
 n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , 
 n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , 
 n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , 
 n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , 
 n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , 
 n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , 
 n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , 
 n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , 
 n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , 
 n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , 
 n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , 
 n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , 
 n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , 
 n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , 
 n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , 
 n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , 
 n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , 
 n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , 
 n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , 
 n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , 
 n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , 
 n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , 
 n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , 
 n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , 
 n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , 
 n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , 
 n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , 
 n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , 
 n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , 
 n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , 
 n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , 
 n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , 
 n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , 
 n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , 
 n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , 
 n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , 
 n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , 
 n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , 
 n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , 
 n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , 
 n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , 
 n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , 
 n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , 
 n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , 
 n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , 
 n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , 
 n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , 
 n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , 
 n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , 
 n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , 
 n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , 
 n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , 
 n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , 
 n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , 
 n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , 
 n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , 
 n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , 
 n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , 
 n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , 
 n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , 
 n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , 
 n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , 
 n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , 
 n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , 
 n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , 
 n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , 
 n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , 
 n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , 
 n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , 
 n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , 
 n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , 
 n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , 
 n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , 
 n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , 
 n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , 
 n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , 
 n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , 
 n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , 
 n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , 
 n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , 
 n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , 
 n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , 
 n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , 
 n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , 
 n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , 
 n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , 
 n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , 
 n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , 
 n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , 
 n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , 
 n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , 
 n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , 
 n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , 
 n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , 
 n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , 
 n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , 
 n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , 
 n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , 
 n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , 
 n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , 
 n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , 
 n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , 
 n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , 
 n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , 
 n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , 
 n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , 
 n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , 
 n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , 
 n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , 
 n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , 
 n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , 
 n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , 
 n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , 
 n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , 
 n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , 
 n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , 
 n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , 
 n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , 
 n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , 
 n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , 
 n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , 
 n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , 
 n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , 
 n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , 
 n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , 
 n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , 
 n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , 
 n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , 
 n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , 
 n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , 
 n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , 
 n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , 
 n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , 
 n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , 
 n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , 
 n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , 
 n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , 
 n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , 
 n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , 
 n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , 
 n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , 
 n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , 
 n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , 
 n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , 
 n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , 
 n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , 
 n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , 
 n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , 
 n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , 
 n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , 
 n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , 
 n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , 
 n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , 
 n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , 
 n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , 
 n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , 
 n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , 
 n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , 
 n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , 
 n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , 
 n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , 
 n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , 
 n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , 
 n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , 
 n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , 
 n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , 
 n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , 
 n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , 
 n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , 
 n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , 
 n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , 
 n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , 
 n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , 
 n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , 
 n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , 
 n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , 
 n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , 
 n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , 
 n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , 
 n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , 
 n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , 
 n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , 
 n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , 
 n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , 
 n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , 
 n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , 
 n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , 
 n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , 
 n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , 
 n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , 
 n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , 
 n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , 
 n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , 
 n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , 
 n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , 
 n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , 
 n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , 
 n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , 
 n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , 
 n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , 
 n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , 
 n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , 
 n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , 
 n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , 
 n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , 
 n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , 
 n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , 
 n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , 
 n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , 
 n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , 
 n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , 
 n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , 
 n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , 
 n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , 
 n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , 
 n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , 
 n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , 
 n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , 
 n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , 
 n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , 
 n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , 
 n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , 
 n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , 
 n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , 
 n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , 
 n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , 
 n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , 
 n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , 
 n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , 
 n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , 
 n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , 
 n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , 
 n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , 
 n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , 
 n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , 
 n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , 
 n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , 
 n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , 
 n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , 
 n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , 
 n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , 
 n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , 
 n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , 
 n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , 
 n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , 
 n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , 
 n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , 
 n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , 
 n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , 
 n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , 
 n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , 
 n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , 
 n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , 
 n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , 
 n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , 
 n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , 
 n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , 
 n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , 
 n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , 
 n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , 
 n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , 
 n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , 
 n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , 
 n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , 
 n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , 
 n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , 
 n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , 
 n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , 
 n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , 
 n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , 
 n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , 
 n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , 
 n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , 
 n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , 
 n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , 
 n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , 
 n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , 
 n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , 
 n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , 
 n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , 
 n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , 
 n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , 
 n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , 
 n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , 
 n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , 
 n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , 
 n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , 
 n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , 
 n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , 
 n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , 
 n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , 
 n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , 
 n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , 
 n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , 
 n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , 
 n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , 
 n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , 
 n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , 
 n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , 
 n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , 
 n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , 
 n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , 
 n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , 
 n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , 
 n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , 
 n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , 
 n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , 
 n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , 
 n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , 
 n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , 
 n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , 
 n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , 
 n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , 
 n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , 
 n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , 
 n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , 
 n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , 
 n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , 
 n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , 
 n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , 
 n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , 
 n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , 
 n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , 
 n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , 
 n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , 
 n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , 
 n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , 
 n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , 
 n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , 
 n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , 
 n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , 
 n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , 
 n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , 
 n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , 
 n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , 
 n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , 
 n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , 
 n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , 
 n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , 
 n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , 
 n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , 
 n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , 
 n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , 
 n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , 
 n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , 
 n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , 
 n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , 
 n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , 
 n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , 
 n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , 
 n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , 
 n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , 
 n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , 
 n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , 
 n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , 
 n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , 
 n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , 
 n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , 
 n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , 
 n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , 
 n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , 
 n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , 
 n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , 
 n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , 
 n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , 
 n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , 
 n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , 
 n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , 
 n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , 
 n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , 
 n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , 
 n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , 
 n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , 
 n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , 
 n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , 
 n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , 
 n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , 
 n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , 
 n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , 
 n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , 
 n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , 
 n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , 
 n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , 
 n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , 
 n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , 
 n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , 
 n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , 
 n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , 
 n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , 
 n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , 
 n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , 
 n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , 
 n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , 
 n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , 
 n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , 
 n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , 
 n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , 
 n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , 
 n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , 
 n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , 
 n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , 
 n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , 
 n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , 
 n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , 
 n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , 
 n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , 
 n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , 
 n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , 
 n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , 
 n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , 
 n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , 
 n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , 
 n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , 
 n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , 
 n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , 
 n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , 
 n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , 
 n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , 
 n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , 
 n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , 
 n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , 
 n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , 
 n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , 
 n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , 
 n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , 
 n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , 
 n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , 
 n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , 
 n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , 
 n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , 
 n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , 
 n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , 
 n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , 
 n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , 
 n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , 
 n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , 
 n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , 
 n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , 
 n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , 
 n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , 
 n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , 
 n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , 
 n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , 
 n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , 
 n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , 
 n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , 
 n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , 
 n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , 
 n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , 
 n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , 
 n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , 
 n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , 
 n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , 
 n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , 
 n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , 
 n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , 
 n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , 
 n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , 
 n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , 
 n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , 
 n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , 
 n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , 
 n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , 
 n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , 
 n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , 
 n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , 
 n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , 
 n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , 
 n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , 
 n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , 
 n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , 
 n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , 
 n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , 
 n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , 
 n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , 
 n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , 
 n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , 
 n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , 
 n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , 
 n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , 
 n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , 
 n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , 
 n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , 
 n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , 
 n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , 
 n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , 
 n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , 
 n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , 
 n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , 
 n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , 
 n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , 
 n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , 
 n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , 
 n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , 
 n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , 
 n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , 
 n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , 
 n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , 
 n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , 
 n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , 
 n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , 
 n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , 
 n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , 
 n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , 
 n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , 
 n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , 
 n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , 
 n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , 
 n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , 
 n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , 
 n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , 
 n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , 
 n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , 
 n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , 
 n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , 
 n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , 
 n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , 
 n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , 
 n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , 
 n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , 
 n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , 
 n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , 
 n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , 
 n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , 
 n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , 
 n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , 
 n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , 
 n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , 
 n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , 
 n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , 
 n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , 
 n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , 
 n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , 
 n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , 
 n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , 
 n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , 
 n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , 
 n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , 
 n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , 
 n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , 
 n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , 
 n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , 
 n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , 
 n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , 
 n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , 
 n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , 
 n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , 
 n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , 
 n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , 
 n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , 
 n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , 
 n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , 
 n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , 
 n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , 
 n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , 
 n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , 
 n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , 
 n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , 
 n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , 
 n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , 
 n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , 
 n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , 
 n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , 
 n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , 
 n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , 
 n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , 
 n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , 
 n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , 
 n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , 
 n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , 
 n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , 
 n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , 
 n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , 
 n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , 
 n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , 
 n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , 
 n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , 
 n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , 
 n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , 
 n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , 
 n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , 
 n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , 
 n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , 
 n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , 
 n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , 
 n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , 
 n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , 
 n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , 
 n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , 
 n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , 
 n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , 
 n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , 
 n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , 
 n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , 
 n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , 
 n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , 
 n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , 
 n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , 
 n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , 
 n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , 
 n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , 
 n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , 
 n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , 
 n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , 
 n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , 
 n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , 
 n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , 
 n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , 
 n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , 
 n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , 
 n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , 
 n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , 
 n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , 
 n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , 
 n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , 
 n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , 
 n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , 
 n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , 
 n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , 
 n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , 
 n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , 
 n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , 
 n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , 
 n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , 
 n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , 
 n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , 
 n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , 
 n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , 
 n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , 
 n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , 
 n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , 
 n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , 
 n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , 
 n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , 
 n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , 
 n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , 
 n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , 
 n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , 
 n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , 
 n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , 
 n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , 
 n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , 
 n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , 
 n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , 
 n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , 
 n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , 
 n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , 
 n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , 
 n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , 
 n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , 
 n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , 
 n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , 
 n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , 
 n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , 
 n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , 
 n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , 
 n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , 
 n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , 
 n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , 
 n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , 
 n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , 
 n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , 
 n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , 
 n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , 
 n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , 
 n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , 
 n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , 
 n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , 
 n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , 
 n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , 
 n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , 
 n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , 
 n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , 
 n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , 
 n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , 
 n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , 
 n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , 
 n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , 
 n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , 
 n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , 
 n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , 
 n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , 
 n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , 
 n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , 
 n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , 
 n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , 
 n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , 
 n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , 
 n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , 
 n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , 
 n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , 
 n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , 
 n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , 
 n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , 
 n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , 
 n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , 
 n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , 
 n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , 
 n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , 
 n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , 
 n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , 
 n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , 
 n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , 
 n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , 
 n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , 
 n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , 
 n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , 
 n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , 
 n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , 
 n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , 
 n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , 
 n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , 
 n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , 
 n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , 
 n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , 
 n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , 
 n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , 
 n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , 
 n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , 
 n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , 
 n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , 
 n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , 
 n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , 
 n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , 
 n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , 
 n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , 
 n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , 
 n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , 
 n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , 
 n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , 
 n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , 
 n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , 
 n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , 
 n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , 
 n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , 
 n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , 
 n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , 
 n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , 
 n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , 
 n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , 
 n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , 
 n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , 
 n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , 
 n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , 
 n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , 
 n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , 
 n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , 
 n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , 
 n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , 
 n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , 
 n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , 
 n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , 
 n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , 
 n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , 
 n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , 
 n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , 
 n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , 
 n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , 
 n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , 
 n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , 
 n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , 
 n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , 
 n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , 
 n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , 
 n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , 
 n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , 
 n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , 
 n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , 
 n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , 
 n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , 
 n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , 
 n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , 
 n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , 
 n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , 
 n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , 
 n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , 
 n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , 
 n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , 
 n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , 
 n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , 
 n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , 
 n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , 
 n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , 
 n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , 
 n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , 
 n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , 
 n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , 
 n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , 
 n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , 
 n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , 
 n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , 
 n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , 
 n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , 
 n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , 
 n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , 
 n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , 
 n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , 
 n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , 
 n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , 
 n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , 
 n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , 
 n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , 
 n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , 
 n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , 
 n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , 
 n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , 
 n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , 
 n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , 
 n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , 
 n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , 
 n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , 
 n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , 
 n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , 
 n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , 
 n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , 
 n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , 
 n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , 
 n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , 
 n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , 
 n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , 
 n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , 
 n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , 
 n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , 
 n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , 
 n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , 
 n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , 
 n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , 
 n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , 
 n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , 
 n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , 
 n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , 
 n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , 
 n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , 
 n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , 
 n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , 
 n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , 
 n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , 
 n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , 
 n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , 
 n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , 
 n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , 
 n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , 
 n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , 
 n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , 
 n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , 
 n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , 
 n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , 
 n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , 
 n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , 
 n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , 
 n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , 
 n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , 
 n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , 
 n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , 
 n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , 
 n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , 
 n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , 
 n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , 
 n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , 
 n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , 
 n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , 
 n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , 
 n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , 
 n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , 
 n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , 
 n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , 
 n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , 
 n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , 
 n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , 
 n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , 
 n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , 
 n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , 
 n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , 
 n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , 
 n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , 
 n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , 
 n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , 
 n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , 
 n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , 
 n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , 
 n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , 
 n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , 
 n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , 
 n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , 
 n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , 
 n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , 
 n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , 
 n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , 
 n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , 
 n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , 
 n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , 
 n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , 
 n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , 
 n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , 
 n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , 
 n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , 
 n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , 
 n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , 
 n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , 
 n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , 
 n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , 
 n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , 
 n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , 
 n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , 
 n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , 
 n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , 
 n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , 
 n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , 
 n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , 
 n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , 
 n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , 
 n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , 
 n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , 
 n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , 
 n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , 
 n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , 
 n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , 
 n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , 
 n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , 
 n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , 
 n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , 
 n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , 
 n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , 
 n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , 
 n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , 
 n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , 
 n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , 
 n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , 
 n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , 
 n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , 
 n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , 
 n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , 
 n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , 
 n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , 
 n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , 
 n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , 
 n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , 
 n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , 
 n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , 
 n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , 
 n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , 
 n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , 
 n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , 
 n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , 
 n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , 
 n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , 
 n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , 
 n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , 
 n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , 
 n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , 
 n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , 
 n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , 
 n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , 
 n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , 
 n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , 
 n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , 
 n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , 
 n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , 
 n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , 
 n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , 
 n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , 
 n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , 
 n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , 
 n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , 
 n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , 
 n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , 
 n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , 
 n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , 
 n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , 
 n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , 
 n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , 
 n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , 
 n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , 
 n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , 
 n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , 
 n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , 
 n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , 
 n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , 
 n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , 
 n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , 
 n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , 
 n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , 
 n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , 
 n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , 
 n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , 
 n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , 
 n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , 
 n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , 
 n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , 
 n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , 
 n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , 
 n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , 
 n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , 
 n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , 
 n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , 
 n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , 
 n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , 
 n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , 
 n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , 
 n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , 
 n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , 
 n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , 
 n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , 
 n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , 
 n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , 
 n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , 
 n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , 
 n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , 
 n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , 
 n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , 
 n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , 
 n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , 
 n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , 
 n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , 
 n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , 
 n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , 
 n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , 
 n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , 
 n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , 
 n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , 
 n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , 
 n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , 
 n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , 
 n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , 
 n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , 
 n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , 
 n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , 
 n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , 
 n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , 
 n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , 
 n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , 
 n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , 
 n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , 
 n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , 
 n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , 
 n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , 
 n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , 
 n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , 
 n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , 
 n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , 
 n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , 
 n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , 
 n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , 
 n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , 
 n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , 
 n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , 
 n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , 
 n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , 
 n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , 
 n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , 
 n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , 
 n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , 
 n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , 
 n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , 
 n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , 
 n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , 
 n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , 
 n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , 
 n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , 
 n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , 
 n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , 
 n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , 
 n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , 
 n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , 
 n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , 
 n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , 
 n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , 
 n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , 
 n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , 
 n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , 
 n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , 
 n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , 
 n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , 
 n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , 
 n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , 
 n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , 
 n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , 
 n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , 
 n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , 
 n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , 
 n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , 
 n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , 
 n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , 
 n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , 
 n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , 
 n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , 
 n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , 
 n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , 
 n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , 
 n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , 
 n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , 
 n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , 
 n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , 
 n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , 
 n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , 
 n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , 
 n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , 
 n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , 
 n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , 
 n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , 
 n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , 
 n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , 
 n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , 
 n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , 
 n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , 
 n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , 
 n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , 
 n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , 
 n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , 
 n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , 
 n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , 
 n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , 
 n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , 
 n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , 
 n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , 
 n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , 
 n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , 
 n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , 
 n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , 
 n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , 
 n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , 
 n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , 
 n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , 
 n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , 
 n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , 
 n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , 
 n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , 
 n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , 
 n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , 
 n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , 
 n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , 
 n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , 
 n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , 
 n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , 
 n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , 
 n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , 
 n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , 
 n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , 
 n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , 
 n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , 
 n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , 
 n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , 
 n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , 
 n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , 
 n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , 
 n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , 
 n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , 
 n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , 
 n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , 
 n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , 
 n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , 
 n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , 
 n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , 
 n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , 
 n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , 
 n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , 
 n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , 
 n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , 
 n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , 
 n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , 
 n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , 
 n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , 
 n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , 
 n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , 
 n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , 
 n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , 
 n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , 
 n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , 
 n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , 
 n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , 
 n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , 
 n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , 
 n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , 
 n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , 
 n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , 
 n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , 
 n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , 
 n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , 
 n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , 
 n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , 
 n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , 
 n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , 
 n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , 
 n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , 
 n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , 
 n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , 
 n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , 
 n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , 
 n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , 
 n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , 
 n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , 
 n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , 
 n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , 
 n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , 
 n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , 
 n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , 
 n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , 
 n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , 
 n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , 
 n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , 
 n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , 
 n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , 
 n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , 
 n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , 
 n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , 
 n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , 
 n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , 
 n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , 
 n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , 
 n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , 
 n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , 
 n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , 
 n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , 
 n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , 
 n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , 
 n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , 
 n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , 
 n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , 
 n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , 
 n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , 
 n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , 
 n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , 
 n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , 
 n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , 
 n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , 
 n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , 
 n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , 
 n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , 
 n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , 
 n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , 
 n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , 
 n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , 
 n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , 
 n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , 
 n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , 
 n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , 
 n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , 
 n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , 
 n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , n50527 , n50528 , 
 n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , 
 n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , 
 n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , 
 n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , 
 n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , 
 n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , 
 n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , 
 n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , 
 n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , 
 n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , 
 n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , 
 n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , 
 n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , 
 n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , 
 n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , 
 n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , 
 n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , 
 n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , 
 n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , 
 n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , 
 n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , 
 n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , 
 n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , 
 n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , 
 n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , 
 n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , 
 n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , 
 n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , 
 n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , 
 n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , 
 n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , 
 n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , 
 n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , 
 n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , 
 n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , 
 n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , 
 n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , 
 n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , 
 n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , 
 n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , 
 n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , 
 n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , 
 n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , 
 n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , 
 n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , 
 n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , 
 n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , 
 n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , 
 n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , 
 n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , 
 n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , 
 n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , 
 n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , 
 n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , 
 n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , 
 n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , 
 n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , 
 n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , 
 n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , 
 n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , 
 n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , 
 n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , 
 n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , 
 n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , 
 n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , 
 n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , 
 n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , n51197 , n51198 , 
 n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , 
 n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , 
 n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , 
 n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , 
 n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , 
 n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , 
 n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , 
 n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , n51277 , n51278 , 
 n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , n51287 , n51288 , 
 n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , n51297 , n51298 , 
 n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , n51307 , n51308 , 
 n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , n51317 , n51318 , 
 n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , n51327 , n51328 , 
 n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , 
 n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , n51347 , n51348 , 
 n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , n51357 , n51358 , 
 n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , n51367 , n51368 , 
 n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , n51377 , n51378 , 
 n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , n51387 , n51388 , 
 n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , n51397 , n51398 , 
 n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , n51407 , n51408 , 
 n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , n51417 , n51418 , 
 n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , n51427 , n51428 , 
 n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , n51437 , n51438 , 
 n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , n51447 , n51448 , 
 n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , n51457 , n51458 , 
 n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , n51467 , n51468 , 
 n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , n51477 , n51478 , 
 n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , n51487 , n51488 , 
 n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , n51497 , n51498 , 
 n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , n51507 , n51508 , 
 n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , n51517 , n51518 , 
 n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , n51527 , n51528 , 
 n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , n51537 , n51538 , 
 n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , n51547 , n51548 , 
 n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , n51557 , n51558 , 
 n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , n51567 , n51568 , 
 n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , n51577 , n51578 , 
 n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , n51587 , n51588 , 
 n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , n51597 , n51598 , 
 n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , n51607 , n51608 , 
 n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , n51617 , n51618 , 
 n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , n51627 , n51628 , 
 n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , n51637 , n51638 , 
 n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , n51647 , n51648 , 
 n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , n51657 , n51658 , 
 n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , n51667 , n51668 , 
 n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , n51677 , n51678 , 
 n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , n51687 , n51688 , 
 n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , n51697 , n51698 , 
 n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , n51707 , n51708 , 
 n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , n51717 , n51718 , 
 n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , n51727 , n51728 , 
 n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , n51737 , n51738 , 
 n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , n51747 , n51748 , 
 n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , n51757 , n51758 , 
 n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , n51767 , n51768 , 
 n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , n51777 , n51778 , 
 n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , n51787 , n51788 , 
 n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , n51797 , n51798 , 
 n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , n51807 , n51808 , 
 n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , n51817 , n51818 , 
 n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n51827 , n51828 , 
 n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , n51837 , n51838 , 
 n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , n51847 , n51848 , 
 n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , n51857 , n51858 , 
 n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , n51867 , n51868 , 
 n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , n51877 , n51878 , 
 n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , n51887 , n51888 , 
 n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , n51897 , n51898 , 
 n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , n51908 , 
 n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , n51917 , n51918 , 
 n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , n51927 , n51928 , 
 n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , n51937 , n51938 , 
 n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , n51947 , n51948 , 
 n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , n51957 , n51958 , 
 n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , n51967 , n51968 , 
 n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , n51977 , n51978 , 
 n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , n51987 , n51988 , 
 n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , n51997 , n51998 , 
 n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , n52007 , n52008 , 
 n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , n52017 , n52018 , 
 n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , n52027 , n52028 , 
 n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , n52037 , n52038 , 
 n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , n52047 , n52048 , 
 n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , n52057 , n52058 , 
 n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , n52067 , n52068 , 
 n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , n52077 , n52078 , 
 n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , n52087 , n52088 , 
 n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , n52097 , n52098 , 
 n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , n52107 , n52108 , 
 n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , n52117 , n52118 , 
 n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , n52127 , n52128 , 
 n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , n52137 , n52138 , 
 n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , n52147 , n52148 , 
 n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , n52157 , n52158 , 
 n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , n52167 , n52168 , 
 n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , n52177 , n52178 , 
 n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , n52187 , n52188 , 
 n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , n52197 , n52198 , 
 n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , n52207 , n52208 , 
 n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , n52217 , n52218 , 
 n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , n52227 , n52228 , 
 n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , n52237 , n52238 , 
 n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , n52247 , n52248 , 
 n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , n52257 , n52258 , 
 n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , n52267 , n52268 , 
 n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , n52277 , n52278 , 
 n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , n52287 , n52288 , 
 n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , n52297 , n52298 , 
 n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , n52307 , n52308 , 
 n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , n52317 , n52318 , 
 n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , n52327 , n52328 , 
 n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , n52337 , n52338 , 
 n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , n52347 , n52348 , 
 n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , n52357 , n52358 , 
 n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , 
 n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , 
 n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , n52387 , n52388 , 
 n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , n52397 , n52398 , 
 n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , n52407 , n52408 , 
 n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , n52417 , n52418 , 
 n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , n52427 , n52428 , 
 n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , n52437 , n52438 , 
 n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , n52447 , n52448 , 
 n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , n52457 , n52458 , 
 n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , n52467 , n52468 , 
 n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , n52477 , n52478 , 
 n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , n52487 , n52488 , 
 n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , n52497 , n52498 , 
 n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , n52507 , n52508 , 
 n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , n52517 , n52518 , 
 n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , 
 n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , n52537 , n52538 , 
 n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , n52547 , n52548 , 
 n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , n52557 , n52558 , 
 n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , 
 n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , 
 n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , n52587 , n52588 , 
 n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , n52597 , n52598 , 
 n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , n52607 , n52608 , 
 n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , n52617 , n52618 , 
 n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , n52627 , n52628 , 
 n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , n52637 , n52638 , 
 n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , n52647 , n52648 , 
 n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , n52657 , n52658 , 
 n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , n52667 , n52668 , 
 n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , n52677 , n52678 , 
 n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , n52687 , n52688 , 
 n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , n52697 , n52698 , 
 n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , 
 n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , 
 n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , n52727 , n52728 , 
 n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , 
 n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , 
 n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , 
 n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , 
 n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , 
 n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , 
 n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , 
 n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , 
 n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , 
 n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , 
 n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , 
 n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , n52847 , n52848 , 
 n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , n52857 , n52858 , 
 n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , n52867 , n52868 , 
 n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , n52877 , n52878 , 
 n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , n52887 , n52888 , 
 n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , n52897 , n52898 , 
 n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , n52907 , n52908 , 
 n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , n52917 , n52918 , 
 n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , n52927 , n52928 , 
 n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , n52937 , n52938 , 
 n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , n52947 , n52948 , 
 n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , n52957 , n52958 , 
 n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , n52967 , n52968 , 
 n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , n52977 , n52978 , 
 n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , n52987 , n52988 , 
 n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , n52997 , n52998 , 
 n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , n53007 , n53008 , 
 n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , n53017 , n53018 , 
 n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , n53027 , n53028 , 
 n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , n53037 , n53038 , 
 n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , n53047 , n53048 , 
 n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , n53057 , n53058 , 
 n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , n53067 , n53068 , 
 n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , n53077 , n53078 , 
 n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , n53087 , n53088 , 
 n53089 , n53090 , n53091 , n53092 , n53093 , n53094 , n53095 , n53096 , n53097 , n53098 , 
 n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , n53107 , n53108 , 
 n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , n53117 , n53118 , 
 n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , n53127 , n53128 , 
 n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , n53137 , n53138 , 
 n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , n53147 , n53148 , 
 n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , n53157 , n53158 , 
 n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , n53167 , n53168 , 
 n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , n53177 , n53178 , 
 n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , n53187 , n53188 , 
 n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , n53197 , n53198 , 
 n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , n53207 , n53208 , 
 n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , n53217 , n53218 , 
 n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , n53227 , n53228 , 
 n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , n53237 , n53238 , 
 n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , n53247 , n53248 , 
 n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , n53257 , n53258 , 
 n53259 , n53260 , n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , n53267 , n53268 , 
 n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , n53277 , n53278 , 
 n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , n53287 , n53288 , 
 n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , n53297 , n53298 , 
 n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , n53307 , n53308 , 
 n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , n53317 , n53318 , 
 n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , 
 n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , 
 n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , 
 n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , 
 n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , 
 n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , 
 n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , 
 n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , 
 n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , 
 n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , n53417 , n53418 , 
 n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , 
 n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , 
 n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , 
 n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , 
 n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , 
 n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , 
 n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , 
 n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , 
 n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , 
 n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , 
 n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , 
 n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , 
 n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , 
 n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , n53557 , n53558 , 
 n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , 
 n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , 
 n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , 
 n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , 
 n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , 
 n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , 
 n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , 
 n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , 
 n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , 
 n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , 
 n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , 
 n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , 
 n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , n53687 , n53688 , 
 n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , 
 n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , 
 n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , 
 n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , 
 n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , n53737 , n53738 , 
 n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , 
 n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , 
 n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , 
 n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , 
 n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , 
 n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , 
 n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , 
 n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , 
 n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , 
 n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , 
 n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , 
 n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , 
 n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , n53867 , n53868 , 
 n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , n53877 , n53878 , 
 n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , n53887 , n53888 , 
 n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , n53897 , n53898 , 
 n53899 , n53900 , n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , n53907 , n53908 , 
 n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , n53917 , n53918 , 
 n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , n53927 , n53928 , 
 n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , n53937 , n53938 , 
 n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , n53947 , n53948 , 
 n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , n53957 , n53958 , 
 n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , n53967 , n53968 , 
 n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , 
 n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , n53987 , n53988 , 
 n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , n53997 , n53998 , 
 n53999 , n54000 , n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , n54007 , n54008 , 
 n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , n54017 , n54018 , 
 n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , n54027 , n54028 , 
 n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , n54037 , n54038 , 
 n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , n54047 , n54048 , 
 n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , n54057 , n54058 , 
 n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , n54067 , n54068 , 
 n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , n54077 , n54078 , 
 n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , n54087 , n54088 , 
 n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , n54097 , n54098 , 
 n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , n54107 , n54108 , 
 n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , n54117 , n54118 , 
 n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , 
 n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , n54137 , n54138 , 
 n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , n54147 , n54148 , 
 n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , n54157 , n54158 , 
 n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , n54167 , n54168 , 
 n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , n54177 , n54178 , 
 n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , n54187 , n54188 , 
 n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , n54197 , n54198 , 
 n54199 , n54200 , n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , n54207 , n54208 , 
 n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , n54217 , n54218 , 
 n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , n54227 , n54228 , 
 n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , n54237 , n54238 , 
 n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , n54247 , n54248 , 
 n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , n54257 , n54258 , 
 n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , n54267 , n54268 , 
 n54269 , n54270 , n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , n54277 , n54278 , 
 n54279 , n54280 , n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , n54287 , n54288 , 
 n54289 , n54290 , n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , n54297 , n54298 , 
 n54299 , n54300 , n54301 , n54302 , n54303 , n54304 , n54305 , n54306 , n54307 , n54308 , 
 n54309 , n54310 , n54311 , n54312 , n54313 , n54314 , n54315 , n54316 , n54317 , n54318 , 
 n54319 , n54320 , n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , n54327 , n54328 , 
 n54329 , n54330 , n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , n54337 , n54338 , 
 n54339 , n54340 , n54341 , n54342 , n54343 , n54344 , n54345 , n54346 , n54347 , n54348 , 
 n54349 , n54350 , n54351 , n54352 , n54353 , n54354 , n54355 , n54356 , n54357 , n54358 , 
 n54359 , n54360 , n54361 , n54362 , n54363 , n54364 , n54365 , n54366 , n54367 , n54368 , 
 n54369 , n54370 , n54371 , n54372 , n54373 , n54374 , n54375 , n54376 , n54377 , n54378 , 
 n54379 , n54380 , n54381 , n54382 , n54383 , n54384 , n54385 , n54386 , n54387 , n54388 , 
 n54389 , n54390 , n54391 , n54392 , n54393 , n54394 , n54395 , n54396 , n54397 , n54398 , 
 n54399 , n54400 , n54401 , n54402 , n54403 , n54404 , n54405 , n54406 , n54407 , n54408 , 
 n54409 , n54410 , n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , n54417 , n54418 , 
 n54419 , n54420 , n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , n54427 , n54428 , 
 n54429 , n54430 , n54431 , n54432 , n54433 , n54434 , n54435 , n54436 , n54437 , n54438 , 
 n54439 , n54440 , n54441 , n54442 , n54443 , n54444 , n54445 , n54446 , n54447 , n54448 , 
 n54449 , n54450 , n54451 , n54452 , n54453 , n54454 , n54455 , n54456 , n54457 , n54458 , 
 n54459 , n54460 , n54461 , n54462 , n54463 , n54464 , n54465 , n54466 , n54467 , n54468 , 
 n54469 , n54470 , n54471 , n54472 , n54473 , n54474 , n54475 , n54476 , n54477 , n54478 , 
 n54479 , n54480 , n54481 , n54482 , n54483 , n54484 , n54485 , n54486 , n54487 , n54488 , 
 n54489 , n54490 , n54491 , n54492 , n54493 , n54494 , n54495 , n54496 , n54497 , n54498 , 
 n54499 , n54500 , n54501 , n54502 , n54503 , n54504 , n54505 , n54506 , n54507 , n54508 , 
 n54509 , n54510 , n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , n54517 , n54518 , 
 n54519 , n54520 , n54521 , n54522 , n54523 , n54524 , n54525 , n54526 , n54527 , n54528 , 
 n54529 , n54530 , n54531 , n54532 , n54533 , n54534 , n54535 , n54536 , n54537 , n54538 , 
 n54539 , n54540 , n54541 , n54542 , n54543 , n54544 , n54545 , n54546 , n54547 , n54548 , 
 n54549 , n54550 , n54551 , n54552 , n54553 , n54554 , n54555 , n54556 , n54557 , n54558 , 
 n54559 , n54560 , n54561 , n54562 , n54563 , n54564 , n54565 , n54566 , n54567 , n54568 , 
 n54569 , n54570 , n54571 , n54572 , n54573 , n54574 , n54575 , n54576 , n54577 , n54578 , 
 n54579 , n54580 , n54581 , n54582 , n54583 , n54584 , n54585 , n54586 , n54587 , n54588 , 
 n54589 , n54590 , n54591 , n54592 , n54593 , n54594 , n54595 , n54596 , n54597 , n54598 , 
 n54599 , n54600 , n54601 , n54602 , n54603 , n54604 , n54605 , n54606 , n54607 , n54608 , 
 n54609 , n54610 , n54611 , n54612 , n54613 , n54614 , n54615 , n54616 , n54617 , n54618 , 
 n54619 , n54620 , n54621 , n54622 , n54623 , n54624 , n54625 , n54626 , n54627 , n54628 , 
 n54629 , n54630 , n54631 , n54632 , n54633 , n54634 , n54635 , n54636 , n54637 , n54638 , 
 n54639 , n54640 , n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , n54647 , n54648 , 
 n54649 , n54650 , n54651 , n54652 , n54653 , n54654 , n54655 , n54656 , n54657 , n54658 , 
 n54659 , n54660 , n54661 , n54662 , n54663 , n54664 , n54665 , n54666 , n54667 , n54668 , 
 n54669 , n54670 , n54671 , n54672 , n54673 , n54674 , n54675 , n54676 , n54677 , n54678 , 
 n54679 , n54680 , n54681 , n54682 , n54683 , n54684 , n54685 , n54686 , n54687 , n54688 , 
 n54689 , n54690 , n54691 , n54692 , n54693 , n54694 , n54695 , n54696 , n54697 , n54698 , 
 n54699 , n54700 , n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , n54707 , n54708 , 
 n54709 , n54710 , n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , n54717 , n54718 , 
 n54719 , n54720 , n54721 , n54722 , n54723 , n54724 , n54725 , n54726 , n54727 , n54728 , 
 n54729 , n54730 , n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , n54737 , n54738 , 
 n54739 , n54740 , n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , n54747 , n54748 , 
 n54749 , n54750 , n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , n54757 , n54758 , 
 n54759 , n54760 , n54761 , n54762 , n54763 , n54764 , n54765 , n54766 , n54767 , n54768 , 
 n54769 , n54770 , n54771 , n54772 , n54773 , n54774 , n54775 , n54776 , n54777 , n54778 , 
 n54779 , n54780 , n54781 , n54782 , n54783 , n54784 , n54785 , n54786 , n54787 , n54788 , 
 n54789 , n54790 , n54791 , n54792 , n54793 , n54794 , n54795 , n54796 , n54797 , n54798 , 
 n54799 , n54800 , n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , n54807 , n54808 , 
 n54809 , n54810 , n54811 , n54812 , n54813 , n54814 , n54815 , n54816 , n54817 , n54818 , 
 n54819 , n54820 , n54821 , n54822 , n54823 , n54824 , n54825 , n54826 , n54827 , n54828 , 
 n54829 , n54830 , n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , n54837 , n54838 , 
 n54839 , n54840 , n54841 , n54842 , n54843 , n54844 , n54845 , n54846 , n54847 , n54848 , 
 n54849 , n54850 , n54851 , n54852 , n54853 , n54854 , n54855 , n54856 , n54857 , n54858 , 
 n54859 , n54860 , n54861 , n54862 , n54863 , n54864 , n54865 , n54866 , n54867 , n54868 , 
 n54869 , n54870 , n54871 , n54872 , n54873 , n54874 , n54875 , n54876 , n54877 , n54878 , 
 n54879 , n54880 , n54881 , n54882 , n54883 , n54884 , n54885 , n54886 , n54887 , n54888 , 
 n54889 , n54890 , n54891 , n54892 , n54893 , n54894 , n54895 , n54896 , n54897 , n54898 , 
 n54899 , n54900 , n54901 , n54902 , n54903 , n54904 , n54905 , n54906 , n54907 , n54908 , 
 n54909 , n54910 , n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , n54917 , n54918 , 
 n54919 , n54920 , n54921 , n54922 , n54923 , n54924 , n54925 , n54926 , n54927 , n54928 , 
 n54929 , n54930 , n54931 , n54932 , n54933 , n54934 , n54935 , n54936 , n54937 , n54938 , 
 n54939 , n54940 , n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , n54947 , n54948 , 
 n54949 , n54950 , n54951 , n54952 , n54953 , n54954 , n54955 , n54956 , n54957 , n54958 , 
 n54959 , n54960 , n54961 , n54962 , n54963 , n54964 , n54965 , n54966 , n54967 , n54968 , 
 n54969 , n54970 , n54971 , n54972 , n54973 , n54974 , n54975 , n54976 , n54977 , n54978 , 
 n54979 , n54980 , n54981 , n54982 , n54983 , n54984 , n54985 , n54986 , n54987 , n54988 , 
 n54989 , n54990 , n54991 , n54992 , n54993 , n54994 , n54995 , n54996 , n54997 , n54998 , 
 n54999 , n55000 , n55001 , n55002 , n55003 , n55004 , n55005 , n55006 , n55007 , n55008 , 
 n55009 , n55010 , n55011 , n55012 , n55013 , n55014 , n55015 , n55016 , n55017 , n55018 , 
 n55019 , n55020 , n55021 , n55022 , n55023 , n55024 , n55025 , n55026 , n55027 , n55028 , 
 n55029 , n55030 , n55031 , n55032 , n55033 , n55034 , n55035 , n55036 , n55037 , n55038 , 
 n55039 , n55040 , n55041 , n55042 , n55043 , n55044 , n55045 , n55046 , n55047 , n55048 , 
 n55049 , n55050 , n55051 , n55052 , n55053 , n55054 , n55055 , n55056 , n55057 , n55058 , 
 n55059 , n55060 , n55061 , n55062 , n55063 , n55064 , n55065 , n55066 , n55067 , n55068 , 
 n55069 , n55070 , n55071 , n55072 , n55073 , n55074 , n55075 , n55076 , n55077 , n55078 , 
 n55079 , n55080 , n55081 , n55082 , n55083 , n55084 , n55085 , n55086 , n55087 , n55088 , 
 n55089 , n55090 , n55091 , n55092 , n55093 , n55094 , n55095 , n55096 , n55097 , n55098 , 
 n55099 , n55100 , n55101 , n55102 , n55103 , n55104 , n55105 , n55106 , n55107 , n55108 , 
 n55109 , n55110 , n55111 , n55112 , n55113 , n55114 , n55115 , n55116 , n55117 , n55118 , 
 n55119 , n55120 , n55121 , n55122 , n55123 , n55124 , n55125 , n55126 , n55127 , n55128 , 
 n55129 , n55130 , n55131 , n55132 , n55133 , n55134 , n55135 , n55136 , n55137 , n55138 , 
 n55139 , n55140 , n55141 , n55142 , n55143 , n55144 , n55145 , n55146 , n55147 , n55148 , 
 n55149 , n55150 , n55151 , n55152 , n55153 , n55154 , n55155 , n55156 , n55157 , n55158 , 
 n55159 , n55160 , n55161 , n55162 , n55163 , n55164 , n55165 , n55166 , n55167 , n55168 , 
 n55169 , n55170 , n55171 , n55172 , n55173 , n55174 , n55175 , n55176 , n55177 , n55178 , 
 n55179 , n55180 , n55181 , n55182 , n55183 , n55184 , n55185 , n55186 , n55187 , n55188 , 
 n55189 , n55190 , n55191 , n55192 , n55193 , n55194 , n55195 , n55196 , n55197 , n55198 , 
 n55199 , n55200 , n55201 , n55202 , n55203 , n55204 , n55205 , n55206 , n55207 , n55208 , 
 n55209 , n55210 , n55211 , n55212 , n55213 , n55214 , n55215 , n55216 , n55217 , n55218 , 
 n55219 , n55220 , n55221 , n55222 , n55223 , n55224 , n55225 , n55226 , n55227 , n55228 , 
 n55229 , n55230 , n55231 , n55232 , n55233 , n55234 , n55235 , n55236 , n55237 , n55238 , 
 n55239 , n55240 , n55241 , n55242 , n55243 , n55244 , n55245 , n55246 , n55247 , n55248 , 
 n55249 , n55250 , n55251 , n55252 , n55253 , n55254 , n55255 , n55256 , n55257 , n55258 , 
 n55259 , n55260 , n55261 , n55262 , n55263 , n55264 , n55265 , n55266 , n55267 , n55268 , 
 n55269 , n55270 , n55271 , n55272 , n55273 , n55274 , n55275 , n55276 , n55277 , n55278 , 
 n55279 , n55280 , n55281 , n55282 , n55283 , n55284 , n55285 , n55286 , n55287 , n55288 , 
 n55289 , n55290 , n55291 , n55292 , n55293 , n55294 , n55295 , n55296 , n55297 , n55298 , 
 n55299 , n55300 , n55301 , n55302 , n55303 , n55304 , n55305 , n55306 , n55307 , n55308 , 
 n55309 , n55310 , n55311 , n55312 , n55313 , n55314 , n55315 , n55316 , n55317 , n55318 , 
 n55319 , n55320 , n55321 , n55322 , n55323 , n55324 , n55325 , n55326 , n55327 , n55328 , 
 n55329 , n55330 , n55331 , n55332 , n55333 , n55334 , n55335 , n55336 , n55337 , n55338 , 
 n55339 , n55340 , n55341 , n55342 , n55343 , n55344 , n55345 , n55346 , n55347 , n55348 , 
 n55349 , n55350 , n55351 , n55352 , n55353 , n55354 , n55355 , n55356 , n55357 , n55358 , 
 n55359 , n55360 , n55361 , n55362 , n55363 , n55364 , n55365 , n55366 , n55367 , n55368 , 
 n55369 , n55370 , n55371 , n55372 , n55373 , n55374 , n55375 , n55376 , n55377 , n55378 , 
 n55379 , n55380 , n55381 , n55382 , n55383 , n55384 , n55385 , n55386 , n55387 , n55388 , 
 n55389 , n55390 , n55391 , n55392 , n55393 , n55394 , n55395 , n55396 , n55397 , n55398 , 
 n55399 , n55400 , n55401 , n55402 , n55403 , n55404 , n55405 , n55406 , n55407 , n55408 , 
 n55409 , n55410 , n55411 , n55412 , n55413 , n55414 , n55415 , n55416 , n55417 , n55418 , 
 n55419 , n55420 , n55421 , n55422 , n55423 , n55424 , n55425 , n55426 , n55427 , n55428 , 
 n55429 , n55430 , n55431 , n55432 , n55433 , n55434 , n55435 , n55436 , n55437 , n55438 , 
 n55439 , n55440 , n55441 , n55442 , n55443 , n55444 , n55445 , n55446 , n55447 , n55448 , 
 n55449 , n55450 , n55451 , n55452 , n55453 , n55454 , n55455 , n55456 , n55457 , n55458 , 
 n55459 , n55460 , n55461 , n55462 , n55463 , n55464 , n55465 , n55466 , n55467 , n55468 , 
 n55469 , n55470 , n55471 , n55472 , n55473 , n55474 , n55475 , n55476 , n55477 , n55478 , 
 n55479 , n55480 , n55481 , n55482 , n55483 , n55484 , n55485 , n55486 , n55487 , n55488 , 
 n55489 , n55490 , n55491 , n55492 , n55493 , n55494 , n55495 , n55496 , n55497 , n55498 , 
 n55499 , n55500 , n55501 , n55502 , n55503 , n55504 , n55505 , n55506 , n55507 , n55508 , 
 n55509 , n55510 , n55511 , n55512 , n55513 , n55514 , n55515 , n55516 , n55517 , n55518 , 
 n55519 , n55520 , n55521 , n55522 , n55523 , n55524 , n55525 , n55526 , n55527 , n55528 , 
 n55529 , n55530 , n55531 , n55532 , n55533 , n55534 , n55535 , n55536 , n55537 , n55538 , 
 n55539 , n55540 , n55541 , n55542 , n55543 , n55544 , n55545 , n55546 , n55547 , n55548 , 
 n55549 , n55550 , n55551 , n55552 , n55553 , n55554 , n55555 , n55556 , n55557 , n55558 , 
 n55559 , n55560 , n55561 , n55562 , n55563 , n55564 , n55565 , n55566 , n55567 , n55568 , 
 n55569 , n55570 , n55571 , n55572 , n55573 , n55574 , n55575 , n55576 , n55577 , n55578 , 
 n55579 , n55580 , n55581 , n55582 , n55583 , n55584 , n55585 , n55586 , n55587 , n55588 , 
 n55589 , n55590 , n55591 , n55592 , n55593 , n55594 , n55595 , n55596 , n55597 , n55598 , 
 n55599 , n55600 , n55601 , n55602 , n55603 , n55604 , n55605 , n55606 , n55607 , n55608 , 
 n55609 , n55610 , n55611 , n55612 , n55613 , n55614 , n55615 , n55616 , n55617 , n55618 , 
 n55619 , n55620 , n55621 , n55622 , n55623 , n55624 , n55625 , n55626 , n55627 , n55628 , 
 n55629 , n55630 , n55631 , n55632 , n55633 , n55634 , n55635 , n55636 , n55637 , n55638 , 
 n55639 , n55640 , n55641 , n55642 , n55643 , n55644 , n55645 , n55646 , n55647 , n55648 , 
 n55649 , n55650 , n55651 , n55652 , n55653 , n55654 , n55655 , n55656 , n55657 , n55658 , 
 n55659 , n55660 , n55661 , n55662 , n55663 , n55664 , n55665 , n55666 , n55667 , n55668 , 
 n55669 , n55670 , n55671 , n55672 , n55673 , n55674 , n55675 , n55676 , n55677 , n55678 , 
 n55679 , n55680 , n55681 , n55682 , n55683 , n55684 , n55685 , n55686 , n55687 , n55688 , 
 n55689 , n55690 , n55691 , n55692 , n55693 , n55694 , n55695 , n55696 , n55697 , n55698 , 
 n55699 , n55700 , n55701 , n55702 , n55703 , n55704 , n55705 , n55706 , n55707 , n55708 , 
 n55709 , n55710 , n55711 , n55712 , n55713 , n55714 , n55715 , n55716 , n55717 , n55718 , 
 n55719 , n55720 , n55721 , n55722 , n55723 , n55724 , n55725 , n55726 , n55727 , n55728 , 
 n55729 , n55730 , n55731 , n55732 , n55733 , n55734 , n55735 , n55736 , n55737 , n55738 , 
 n55739 , n55740 , n55741 , n55742 , n55743 , n55744 , n55745 , n55746 , n55747 , n55748 , 
 n55749 , n55750 , n55751 , n55752 , n55753 , n55754 , n55755 , n55756 , n55757 , n55758 , 
 n55759 , n55760 , n55761 , n55762 , n55763 , n55764 , n55765 , n55766 , n55767 , n55768 , 
 n55769 , n55770 , n55771 , n55772 , n55773 , n55774 , n55775 , n55776 , n55777 , n55778 , 
 n55779 , n55780 , n55781 , n55782 , n55783 , n55784 , n55785 , n55786 , n55787 , n55788 , 
 n55789 , n55790 , n55791 , n55792 , n55793 , n55794 , n55795 , n55796 , n55797 , n55798 , 
 n55799 , n55800 , n55801 , n55802 , n55803 , n55804 , n55805 , n55806 , n55807 , n55808 , 
 n55809 , n55810 , n55811 , n55812 , n55813 , n55814 , n55815 , n55816 , n55817 , n55818 , 
 n55819 , n55820 , n55821 , n55822 , n55823 , n55824 , n55825 , n55826 , n55827 , n55828 , 
 n55829 , n55830 , n55831 , n55832 , n55833 , n55834 , n55835 , n55836 , n55837 , n55838 , 
 n55839 , n55840 , n55841 , n55842 , n55843 , n55844 , n55845 , n55846 , n55847 , n55848 , 
 n55849 , n55850 , n55851 , n55852 , n55853 , n55854 , n55855 , n55856 , n55857 , n55858 , 
 n55859 , n55860 , n55861 , n55862 , n55863 , n55864 , n55865 , n55866 , n55867 , n55868 , 
 n55869 , n55870 , n55871 , n55872 , n55873 , n55874 , n55875 , n55876 , n55877 , n55878 , 
 n55879 , n55880 , n55881 , n55882 , n55883 , n55884 , n55885 , n55886 , n55887 , n55888 , 
 n55889 , n55890 , n55891 , n55892 , n55893 , n55894 , n55895 , n55896 , n55897 , n55898 , 
 n55899 , n55900 , n55901 , n55902 , n55903 , n55904 , n55905 , n55906 , n55907 , n55908 , 
 n55909 , n55910 , n55911 , n55912 , n55913 , n55914 , n55915 , n55916 , n55917 , n55918 , 
 n55919 , n55920 , n55921 , n55922 , n55923 , n55924 , n55925 , n55926 , n55927 , n55928 , 
 n55929 , n55930 , n55931 , n55932 , n55933 , n55934 , n55935 , n55936 , n55937 , n55938 , 
 n55939 , n55940 , n55941 , n55942 , n55943 , n55944 , n55945 , n55946 , n55947 , n55948 , 
 n55949 , n55950 , n55951 , n55952 , n55953 , n55954 , n55955 , n55956 , n55957 , n55958 , 
 n55959 , n55960 , n55961 , n55962 , n55963 , n55964 , n55965 , n55966 , n55967 , n55968 , 
 n55969 , n55970 , n55971 , n55972 , n55973 , n55974 , n55975 , n55976 , n55977 , n55978 , 
 n55979 , n55980 , n55981 , n55982 , n55983 , n55984 , n55985 , n55986 , n55987 , n55988 , 
 n55989 , n55990 , n55991 , n55992 , n55993 , n55994 , n55995 , n55996 , n55997 , n55998 , 
 n55999 , n56000 , n56001 , n56002 , n56003 , n56004 , n56005 , n56006 , n56007 , n56008 , 
 n56009 , n56010 , n56011 , n56012 , n56013 , n56014 , n56015 , n56016 , n56017 , n56018 , 
 n56019 , n56020 , n56021 , n56022 , n56023 , n56024 , n56025 , n56026 , n56027 , n56028 , 
 n56029 , n56030 , n56031 , n56032 , n56033 , n56034 , n56035 , n56036 , n56037 , n56038 , 
 n56039 , n56040 , n56041 , n56042 , n56043 , n56044 , n56045 , n56046 , n56047 , n56048 , 
 n56049 , n56050 , n56051 , n56052 , n56053 , n56054 , n56055 , n56056 , n56057 , n56058 , 
 n56059 , n56060 , n56061 , n56062 , n56063 , n56064 , n56065 , n56066 , n56067 , n56068 , 
 n56069 , n56070 , n56071 , n56072 , n56073 , n56074 , n56075 , n56076 , n56077 , n56078 , 
 n56079 , n56080 , n56081 , n56082 , n56083 , n56084 , n56085 , n56086 , n56087 , n56088 , 
 n56089 , n56090 , n56091 , n56092 , n56093 , n56094 , n56095 , n56096 , n56097 , n56098 , 
 n56099 , n56100 , n56101 , n56102 , n56103 , n56104 , n56105 , n56106 , n56107 , n56108 , 
 n56109 , n56110 , n56111 , n56112 , n56113 , n56114 , n56115 , n56116 , n56117 , n56118 , 
 n56119 , n56120 , n56121 , n56122 , n56123 , n56124 , n56125 , n56126 , n56127 , n56128 , 
 n56129 , n56130 , n56131 , n56132 , n56133 , n56134 , n56135 , n56136 , n56137 , n56138 , 
 n56139 , n56140 , n56141 , n56142 , n56143 , n56144 , n56145 , n56146 , n56147 , n56148 , 
 n56149 , n56150 , n56151 , n56152 , n56153 , n56154 , n56155 , n56156 , n56157 , n56158 , 
 n56159 , n56160 , n56161 , n56162 , n56163 , n56164 , n56165 , n56166 , n56167 , n56168 , 
 n56169 , n56170 , n56171 , n56172 , n56173 , n56174 , n56175 , n56176 , n56177 , n56178 , 
 n56179 , n56180 , n56181 , n56182 , n56183 , n56184 , n56185 , n56186 , n56187 , n56188 , 
 n56189 , n56190 , n56191 , n56192 , n56193 , n56194 , n56195 , n56196 , n56197 , n56198 , 
 n56199 , n56200 , n56201 , n56202 , n56203 , n56204 , n56205 , n56206 , n56207 , n56208 , 
 n56209 , n56210 , n56211 , n56212 , n56213 , n56214 , n56215 , n56216 , n56217 , n56218 , 
 n56219 , n56220 , n56221 , n56222 , n56223 , n56224 , n56225 , n56226 , n56227 , n56228 , 
 n56229 , n56230 , n56231 , n56232 , n56233 , n56234 , n56235 , n56236 , n56237 , n56238 , 
 n56239 , n56240 , n56241 , n56242 , n56243 , n56244 , n56245 , n56246 , n56247 , n56248 , 
 n56249 , n56250 , n56251 , n56252 , n56253 , n56254 , n56255 , n56256 , n56257 , n56258 , 
 n56259 , n56260 , n56261 , n56262 , n56263 , n56264 , n56265 , n56266 , n56267 , n56268 , 
 n56269 , n56270 , n56271 , n56272 , n56273 , n56274 , n56275 , n56276 , n56277 , n56278 , 
 n56279 , n56280 , n56281 , n56282 , n56283 , n56284 , n56285 , n56286 , n56287 , n56288 , 
 n56289 , n56290 , n56291 , n56292 , n56293 , n56294 , n56295 , n56296 , n56297 , n56298 , 
 n56299 , n56300 , n56301 , n56302 , n56303 , n56304 , n56305 , n56306 , n56307 , n56308 , 
 n56309 , n56310 , n56311 , n56312 , n56313 , n56314 , n56315 , n56316 , n56317 , n56318 , 
 n56319 , n56320 , n56321 , n56322 , n56323 , n56324 , n56325 , n56326 , n56327 , n56328 , 
 n56329 , n56330 , n56331 , n56332 , n56333 , n56334 , n56335 , n56336 , n56337 , n56338 , 
 n56339 , n56340 , n56341 , n56342 , n56343 , n56344 , n56345 , n56346 , n56347 , n56348 , 
 n56349 , n56350 , n56351 , n56352 , n56353 , n56354 , n56355 , n56356 , n56357 , n56358 , 
 n56359 , n56360 , n56361 , n56362 , n56363 , n56364 , n56365 , n56366 , n56367 , n56368 , 
 n56369 , n56370 , n56371 , n56372 , n56373 , n56374 , n56375 , n56376 , n56377 , n56378 , 
 n56379 , n56380 , n56381 , n56382 , n56383 , n56384 , n56385 , n56386 , n56387 , n56388 , 
 n56389 , n56390 , n56391 , n56392 , n56393 , n56394 , n56395 , n56396 , n56397 , n56398 , 
 n56399 , n56400 , n56401 , n56402 , n56403 , n56404 , n56405 , n56406 , n56407 , n56408 , 
 n56409 , n56410 , n56411 , n56412 , n56413 , n56414 , n56415 , n56416 , n56417 , n56418 , 
 n56419 , n56420 , n56421 , n56422 , n56423 , n56424 , n56425 , n56426 , n56427 , n56428 , 
 n56429 , n56430 , n56431 , n56432 , n56433 , n56434 , n56435 , n56436 , n56437 , n56438 , 
 n56439 , n56440 , n56441 , n56442 , n56443 , n56444 , n56445 , n56446 , n56447 , n56448 , 
 n56449 , n56450 , n56451 , n56452 , n56453 , n56454 , n56455 , n56456 , n56457 , n56458 , 
 n56459 , n56460 , n56461 , n56462 , n56463 , n56464 , n56465 , n56466 , n56467 , n56468 , 
 n56469 , n56470 , n56471 , n56472 , n56473 , n56474 , n56475 , n56476 , n56477 , n56478 , 
 n56479 , n56480 , n56481 , n56482 , n56483 , n56484 , n56485 , n56486 , n56487 , n56488 , 
 n56489 , n56490 , n56491 , n56492 , n56493 , n56494 , n56495 , n56496 , n56497 , n56498 , 
 n56499 , n56500 , n56501 , n56502 , n56503 , n56504 , n56505 , n56506 , n56507 , n56508 , 
 n56509 , n56510 , n56511 , n56512 , n56513 , n56514 , n56515 , n56516 , n56517 , n56518 , 
 n56519 , n56520 , n56521 , n56522 , n56523 , n56524 , n56525 , n56526 , n56527 , n56528 , 
 n56529 , n56530 , n56531 , n56532 , n56533 , n56534 , n56535 , n56536 , n56537 , n56538 , 
 n56539 , n56540 , n56541 , n56542 , n56543 , n56544 , n56545 , n56546 , n56547 , n56548 , 
 n56549 , n56550 , n56551 , n56552 , n56553 , n56554 , n56555 , n56556 , n56557 , n56558 , 
 n56559 , n56560 , n56561 , n56562 , n56563 , n56564 , n56565 , n56566 , n56567 , n56568 , 
 n56569 , n56570 , n56571 , n56572 , n56573 , n56574 , n56575 , n56576 , n56577 , n56578 , 
 n56579 , n56580 , n56581 , n56582 , n56583 , n56584 , n56585 , n56586 , n56587 , n56588 , 
 n56589 , n56590 , n56591 , n56592 , n56593 , n56594 , n56595 , n56596 , n56597 , n56598 , 
 n56599 , n56600 , n56601 , n56602 , n56603 , n56604 , n56605 , n56606 , n56607 , n56608 , 
 n56609 , n56610 , n56611 , n56612 , n56613 , n56614 , n56615 , n56616 , n56617 , n56618 , 
 n56619 , n56620 , n56621 , n56622 , n56623 , n56624 , n56625 , n56626 , n56627 , n56628 , 
 n56629 , n56630 , n56631 , n56632 , n56633 , n56634 , n56635 , n56636 , n56637 , n56638 , 
 n56639 , n56640 , n56641 , n56642 , n56643 , n56644 , n56645 , n56646 , n56647 , n56648 , 
 n56649 , n56650 , n56651 , n56652 , n56653 , n56654 , n56655 , n56656 , n56657 , n56658 , 
 n56659 , n56660 , n56661 , n56662 , n56663 , n56664 , n56665 , n56666 , n56667 , n56668 , 
 n56669 , n56670 , n56671 , n56672 , n56673 , n56674 , n56675 , n56676 , n56677 , n56678 , 
 n56679 , n56680 , n56681 , n56682 , n56683 , n56684 , n56685 , n56686 , n56687 , n56688 , 
 n56689 , n56690 , n56691 , n56692 , n56693 , n56694 , n56695 , n56696 , n56697 , n56698 , 
 n56699 , n56700 , n56701 , n56702 , n56703 , n56704 , n56705 , n56706 , n56707 , n56708 , 
 n56709 , n56710 , n56711 , n56712 , n56713 , n56714 , n56715 , n56716 , n56717 , n56718 , 
 n56719 , n56720 , n56721 , n56722 , n56723 , n56724 , n56725 , n56726 , n56727 , n56728 , 
 n56729 , n56730 , n56731 , n56732 , n56733 , n56734 , n56735 , n56736 , n56737 , n56738 , 
 n56739 , n56740 , n56741 , n56742 , n56743 , n56744 , n56745 , n56746 , n56747 , n56748 , 
 n56749 , n56750 , n56751 , n56752 , n56753 , n56754 , n56755 , n56756 , n56757 , n56758 , 
 n56759 , n56760 , n56761 , n56762 , n56763 , n56764 , n56765 , n56766 , n56767 , n56768 , 
 n56769 , n56770 , n56771 , n56772 , n56773 , n56774 , n56775 , n56776 , n56777 , n56778 , 
 n56779 , n56780 , n56781 , n56782 , n56783 , n56784 , n56785 , n56786 , n56787 , n56788 , 
 n56789 , n56790 , n56791 , n56792 , n56793 , n56794 , n56795 , n56796 , n56797 , n56798 , 
 n56799 , n56800 , n56801 , n56802 , n56803 , n56804 , n56805 , n56806 , n56807 , n56808 , 
 n56809 , n56810 , n56811 , n56812 , n56813 , n56814 , n56815 , n56816 , n56817 , n56818 , 
 n56819 , n56820 , n56821 , n56822 , n56823 , n56824 , n56825 , n56826 , n56827 , n56828 , 
 n56829 , n56830 , n56831 , n56832 , n56833 , n56834 , n56835 , n56836 , n56837 , n56838 , 
 n56839 , n56840 , n56841 , n56842 , n56843 , n56844 , n56845 , n56846 , n56847 , n56848 , 
 n56849 , n56850 , n56851 , n56852 , n56853 , n56854 , n56855 , n56856 , n56857 , n56858 , 
 n56859 , n56860 , n56861 , n56862 , n56863 , n56864 , n56865 , n56866 , n56867 , n56868 , 
 n56869 , n56870 , n56871 , n56872 , n56873 , n56874 , n56875 , n56876 , n56877 , n56878 , 
 n56879 , n56880 , n56881 , n56882 , n56883 , n56884 , n56885 , n56886 , n56887 , n56888 , 
 n56889 , n56890 , n56891 , n56892 , n56893 , n56894 , n56895 , n56896 , n56897 , n56898 , 
 n56899 , n56900 , n56901 , n56902 , n56903 , n56904 , n56905 , n56906 , n56907 , n56908 , 
 n56909 , n56910 , n56911 , n56912 , n56913 , n56914 , n56915 , n56916 , n56917 , n56918 , 
 n56919 , n56920 , n56921 , n56922 , n56923 , n56924 , n56925 , n56926 , n56927 , n56928 , 
 n56929 , n56930 , n56931 , n56932 , n56933 , n56934 , n56935 , n56936 , n56937 , n56938 , 
 n56939 , n56940 , n56941 , n56942 , n56943 , n56944 , n56945 , n56946 , n56947 , n56948 , 
 n56949 , n56950 , n56951 , n56952 , n56953 , n56954 , n56955 , n56956 , n56957 , n56958 , 
 n56959 , n56960 , n56961 , n56962 , n56963 , n56964 , n56965 , n56966 , n56967 , n56968 , 
 n56969 , n56970 , n56971 , n56972 , n56973 , n56974 , n56975 , n56976 , n56977 , n56978 , 
 n56979 , n56980 , n56981 , n56982 , n56983 , n56984 , n56985 , n56986 , n56987 , n56988 , 
 n56989 , n56990 , n56991 , n56992 , n56993 , n56994 , n56995 , n56996 , n56997 , n56998 , 
 n56999 , n57000 , n57001 , n57002 , n57003 , n57004 , n57005 , n57006 , n57007 , n57008 , 
 n57009 , n57010 , n57011 , n57012 , n57013 , n57014 , n57015 , n57016 , n57017 , n57018 , 
 n57019 , n57020 , n57021 , n57022 , n57023 , n57024 , n57025 , n57026 , n57027 , n57028 , 
 n57029 , n57030 , n57031 , n57032 , n57033 , n57034 , n57035 , n57036 , n57037 , n57038 , 
 n57039 , n57040 , n57041 , n57042 , n57043 , n57044 , n57045 , n57046 , n57047 , n57048 , 
 n57049 , n57050 , n57051 , n57052 , n57053 , n57054 , n57055 , n57056 , n57057 , n57058 , 
 n57059 , n57060 , n57061 , n57062 , n57063 , n57064 , n57065 , n57066 , n57067 , n57068 , 
 n57069 , n57070 , n57071 , n57072 , n57073 , n57074 , n57075 , n57076 , n57077 , n57078 , 
 n57079 , n57080 , n57081 , n57082 , n57083 , n57084 , n57085 , n57086 , n57087 , n57088 , 
 n57089 , n57090 , n57091 , n57092 , n57093 , n57094 , n57095 , n57096 , n57097 , n57098 , 
 n57099 , n57100 , n57101 , n57102 , n57103 , n57104 , n57105 , n57106 , n57107 , n57108 , 
 n57109 , n57110 , n57111 , n57112 , n57113 , n57114 , n57115 , n57116 , n57117 , n57118 , 
 n57119 , n57120 , n57121 , n57122 , n57123 , n57124 , n57125 , n57126 , n57127 , n57128 , 
 n57129 , n57130 , n57131 , n57132 , n57133 , n57134 , n57135 , n57136 , n57137 , n57138 , 
 n57139 , n57140 , n57141 , n57142 , n57143 , n57144 , n57145 , n57146 , n57147 , n57148 , 
 n57149 , n57150 , n57151 , n57152 , n57153 , n57154 , n57155 , n57156 , n57157 , n57158 , 
 n57159 , n57160 , n57161 , n57162 , n57163 , n57164 , n57165 , n57166 , n57167 , n57168 , 
 n57169 , n57170 , n57171 , n57172 , n57173 , n57174 , n57175 , n57176 , n57177 , n57178 , 
 n57179 , n57180 , n57181 , n57182 , n57183 , n57184 , n57185 , n57186 , n57187 , n57188 , 
 n57189 , n57190 , n57191 , n57192 , n57193 , n57194 , n57195 , n57196 , n57197 , n57198 , 
 n57199 , n57200 , n57201 , n57202 , n57203 , n57204 , n57205 , n57206 , n57207 , n57208 , 
 n57209 , n57210 , n57211 , n57212 , n57213 , n57214 , n57215 , n57216 , n57217 , n57218 , 
 n57219 , n57220 , n57221 , n57222 , n57223 , n57224 , n57225 , n57226 , n57227 , n57228 , 
 n57229 , n57230 , n57231 , n57232 , n57233 , n57234 , n57235 , n57236 , n57237 , n57238 , 
 n57239 , n57240 , n57241 , n57242 , n57243 , n57244 , n57245 , n57246 , n57247 , n57248 , 
 n57249 , n57250 , n57251 , n57252 , n57253 , n57254 , n57255 , n57256 , n57257 , n57258 , 
 n57259 , n57260 , n57261 , n57262 , n57263 , n57264 , n57265 , n57266 , n57267 , n57268 , 
 n57269 , n57270 , n57271 , n57272 , n57273 , n57274 , n57275 , n57276 , n57277 , n57278 , 
 n57279 , n57280 , n57281 , n57282 , n57283 , n57284 , n57285 , n57286 , n57287 , n57288 , 
 n57289 , n57290 , n57291 , n57292 , n57293 , n57294 , n57295 , n57296 , n57297 , n57298 , 
 n57299 , n57300 , n57301 , n57302 , n57303 , n57304 , n57305 , n57306 , n57307 , n57308 , 
 n57309 , n57310 , n57311 , n57312 , n57313 , n57314 , n57315 , n57316 , n57317 , n57318 , 
 n57319 , n57320 , n57321 , n57322 , n57323 , n57324 , n57325 , n57326 , n57327 , n57328 , 
 n57329 , n57330 , n57331 , n57332 , n57333 , n57334 , n57335 , n57336 , n57337 , n57338 , 
 n57339 , n57340 , n57341 , n57342 , n57343 , n57344 , n57345 , n57346 , n57347 , n57348 , 
 n57349 , n57350 , n57351 , n57352 , n57353 , n57354 , n57355 , n57356 , n57357 , n57358 , 
 n57359 , n57360 , n57361 , n57362 , n57363 , n57364 , n57365 , n57366 , n57367 , n57368 , 
 n57369 , n57370 , n57371 , n57372 , n57373 , n57374 , n57375 , n57376 , n57377 , n57378 , 
 n57379 , n57380 , n57381 , n57382 , n57383 , n57384 , n57385 , n57386 , n57387 , n57388 , 
 n57389 , n57390 , n57391 , n57392 , n57393 , n57394 , n57395 , n57396 , n57397 , n57398 , 
 n57399 , n57400 , n57401 , n57402 , n57403 , n57404 , n57405 , n57406 , n57407 , n57408 , 
 n57409 , n57410 , n57411 , n57412 , n57413 , n57414 , n57415 , n57416 , n57417 , n57418 , 
 n57419 , n57420 , n57421 , n57422 , n57423 , n57424 , n57425 , n57426 , n57427 , n57428 , 
 n57429 , n57430 , n57431 , n57432 , n57433 , n57434 , n57435 , n57436 , n57437 , n57438 , 
 n57439 , n57440 , n57441 , n57442 , n57443 , n57444 , n57445 , n57446 , n57447 , n57448 , 
 n57449 , n57450 , n57451 , n57452 , n57453 , n57454 , n57455 , n57456 , n57457 , n57458 , 
 n57459 , n57460 , n57461 , n57462 , n57463 , n57464 , n57465 , n57466 , n57467 , n57468 , 
 n57469 , n57470 , n57471 , n57472 , n57473 , n57474 , n57475 , n57476 , n57477 , n57478 , 
 n57479 , n57480 , n57481 , n57482 , n57483 , n57484 , n57485 , n57486 , n57487 , n57488 , 
 n57489 , n57490 , n57491 , n57492 , n57493 , n57494 , n57495 , n57496 , n57497 , n57498 , 
 n57499 , n57500 , n57501 , n57502 , n57503 , n57504 , n57505 , n57506 , n57507 , n57508 , 
 n57509 , n57510 , n57511 , n57512 , n57513 , n57514 , n57515 , n57516 , n57517 , n57518 , 
 n57519 , n57520 , n57521 , n57522 , n57523 , n57524 , n57525 , n57526 , n57527 , n57528 , 
 n57529 , n57530 , n57531 , n57532 , n57533 , n57534 , n57535 , n57536 , n57537 , n57538 , 
 n57539 , n57540 , n57541 , n57542 , n57543 , n57544 , n57545 , n57546 , n57547 , n57548 , 
 n57549 , n57550 , n57551 , n57552 , n57553 , n57554 , n57555 , n57556 , n57557 , n57558 , 
 n57559 , n57560 , n57561 , n57562 , n57563 , n57564 , n57565 , n57566 , n57567 , n57568 , 
 n57569 , n57570 , n57571 , n57572 , n57573 , n57574 , n57575 , n57576 , n57577 , n57578 , 
 n57579 , n57580 , n57581 , n57582 , n57583 , n57584 , n57585 , n57586 , n57587 , n57588 , 
 n57589 , n57590 , n57591 , n57592 , n57593 , n57594 , n57595 , n57596 , n57597 , n57598 , 
 n57599 , n57600 , n57601 , n57602 , n57603 , n57604 , n57605 , n57606 , n57607 , n57608 , 
 n57609 , n57610 , n57611 , n57612 , n57613 , n57614 , n57615 , n57616 , n57617 , n57618 , 
 n57619 , n57620 , n57621 , n57622 , n57623 , n57624 , n57625 , n57626 , n57627 , n57628 , 
 n57629 , n57630 , n57631 , n57632 , n57633 , n57634 , n57635 , n57636 , n57637 , n57638 , 
 n57639 , n57640 , n57641 , n57642 , n57643 , n57644 , n57645 , n57646 , n57647 , n57648 , 
 n57649 , n57650 , n57651 , n57652 , n57653 , n57654 , n57655 , n57656 , n57657 , n57658 , 
 n57659 , n57660 , n57661 , n57662 , n57663 , n57664 , n57665 , n57666 , n57667 , n57668 , 
 n57669 , n57670 , n57671 , n57672 , n57673 , n57674 , n57675 , n57676 , n57677 , n57678 , 
 n57679 , n57680 , n57681 , n57682 , n57683 , n57684 , n57685 , n57686 , n57687 , n57688 , 
 n57689 , n57690 , n57691 , n57692 , n57693 , n57694 , n57695 , n57696 , n57697 , n57698 , 
 n57699 , n57700 , n57701 , n57702 , n57703 , n57704 , n57705 , n57706 , n57707 , n57708 , 
 n57709 , n57710 , n57711 , n57712 , n57713 , n57714 , n57715 , n57716 , n57717 , n57718 , 
 n57719 , n57720 , n57721 , n57722 , n57723 , n57724 , n57725 , n57726 , n57727 , n57728 , 
 n57729 , n57730 , n57731 , n57732 , n57733 , n57734 , n57735 , n57736 , n57737 , n57738 , 
 n57739 , n57740 , n57741 , n57742 , n57743 , n57744 , n57745 , n57746 , n57747 , n57748 , 
 n57749 , n57750 , n57751 , n57752 , n57753 , n57754 , n57755 , n57756 , n57757 , n57758 , 
 n57759 , n57760 , n57761 , n57762 , n57763 , n57764 , n57765 , n57766 , n57767 , n57768 , 
 n57769 , n57770 , n57771 , n57772 , n57773 , n57774 , n57775 , n57776 , n57777 , n57778 , 
 n57779 , n57780 , n57781 , n57782 , n57783 , n57784 , n57785 , n57786 , n57787 , n57788 , 
 n57789 , n57790 , n57791 , n57792 , n57793 , n57794 , n57795 , n57796 , n57797 , n57798 , 
 n57799 , n57800 , n57801 , n57802 , n57803 , n57804 , n57805 , n57806 , n57807 , n57808 , 
 n57809 , n57810 , n57811 , n57812 , n57813 , n57814 , n57815 , n57816 , n57817 , n57818 , 
 n57819 , n57820 , n57821 , n57822 , n57823 , n57824 , n57825 , n57826 , n57827 , n57828 , 
 n57829 , n57830 , n57831 , n57832 , n57833 , n57834 , n57835 , n57836 , n57837 , n57838 , 
 n57839 , n57840 , n57841 , n57842 , n57843 , n57844 , n57845 , n57846 , n57847 , n57848 , 
 n57849 , n57850 , n57851 , n57852 , n57853 , n57854 , n57855 , n57856 , n57857 , n57858 , 
 n57859 , n57860 , n57861 , n57862 , n57863 , n57864 , n57865 , n57866 , n57867 , n57868 , 
 n57869 , n57870 , n57871 , n57872 , n57873 , n57874 , n57875 , n57876 , n57877 , n57878 , 
 n57879 , n57880 , n57881 , n57882 , n57883 , n57884 , n57885 , n57886 , n57887 , n57888 , 
 n57889 , n57890 , n57891 , n57892 , n57893 , n57894 , n57895 , n57896 , n57897 , n57898 , 
 n57899 , n57900 , n57901 , n57902 , n57903 , n57904 , n57905 , n57906 , n57907 , n57908 , 
 n57909 , n57910 , n57911 , n57912 , n57913 , n57914 , n57915 , n57916 , n57917 , n57918 , 
 n57919 , n57920 , n57921 , n57922 , n57923 , n57924 , n57925 , n57926 , n57927 , n57928 , 
 n57929 , n57930 , n57931 , n57932 , n57933 , n57934 , n57935 , n57936 , n57937 , n57938 , 
 n57939 , n57940 , n57941 , n57942 , n57943 , n57944 , n57945 , n57946 , n57947 , n57948 , 
 n57949 , n57950 , n57951 , n57952 , n57953 , n57954 , n57955 , n57956 , n57957 , n57958 , 
 n57959 , n57960 , n57961 , n57962 , n57963 , n57964 , n57965 , n57966 , n57967 , n57968 , 
 n57969 , n57970 , n57971 , n57972 , n57973 , n57974 , n57975 , n57976 , n57977 , n57978 , 
 n57979 , n57980 , n57981 , n57982 , n57983 , n57984 , n57985 , n57986 , n57987 , n57988 , 
 n57989 , n57990 , n57991 , n57992 , n57993 , n57994 , n57995 , n57996 , n57997 , n57998 , 
 n57999 , n58000 , n58001 , n58002 , n58003 , n58004 , n58005 , n58006 , n58007 , n58008 , 
 n58009 , n58010 , n58011 , n58012 , n58013 , n58014 , n58015 , n58016 , n58017 , n58018 , 
 n58019 , n58020 , n58021 , n58022 , n58023 , n58024 , n58025 , n58026 , n58027 , n58028 , 
 n58029 , n58030 , n58031 , n58032 , n58033 , n58034 , n58035 , n58036 , n58037 , n58038 , 
 n58039 , n58040 , n58041 , n58042 , n58043 , n58044 , n58045 , n58046 , n58047 , n58048 , 
 n58049 , n58050 , n58051 , n58052 , n58053 , n58054 , n58055 , n58056 , n58057 , n58058 , 
 n58059 , n58060 , n58061 , n58062 , n58063 , n58064 , n58065 , n58066 , n58067 , n58068 , 
 n58069 , n58070 , n58071 , n58072 , n58073 , n58074 , n58075 , n58076 , n58077 , n58078 , 
 n58079 , n58080 , n58081 , n58082 , n58083 , n58084 , n58085 , n58086 , n58087 , n58088 , 
 n58089 , n58090 , n58091 , n58092 , n58093 , n58094 , n58095 , n58096 , n58097 , n58098 , 
 n58099 , n58100 , n58101 , n58102 , n58103 , n58104 , n58105 , n58106 , n58107 , n58108 , 
 n58109 , n58110 , n58111 , n58112 , n58113 , n58114 , n58115 , n58116 , n58117 , n58118 , 
 n58119 , n58120 , n58121 , n58122 , n58123 , n58124 , n58125 , n58126 , n58127 , n58128 , 
 n58129 , n58130 , n58131 , n58132 , n58133 , n58134 , n58135 , n58136 , n58137 , n58138 , 
 n58139 , n58140 , n58141 , n58142 , n58143 , n58144 , n58145 , n58146 , n58147 , n58148 , 
 n58149 , n58150 , n58151 , n58152 , n58153 , n58154 , n58155 , n58156 , n58157 , n58158 , 
 n58159 , n58160 , n58161 , n58162 , n58163 , n58164 , n58165 , n58166 , n58167 , n58168 , 
 n58169 , n58170 , n58171 , n58172 , n58173 , n58174 , n58175 , n58176 , n58177 , n58178 , 
 n58179 , n58180 , n58181 , n58182 , n58183 , n58184 , n58185 , n58186 , n58187 , n58188 , 
 n58189 , n58190 , n58191 , n58192 , n58193 , n58194 , n58195 , n58196 , n58197 , n58198 , 
 n58199 , n58200 , n58201 , n58202 , n58203 , n58204 , n58205 , n58206 , n58207 , n58208 , 
 n58209 , n58210 , n58211 , n58212 , n58213 , n58214 , n58215 , n58216 , n58217 , n58218 , 
 n58219 , n58220 , n58221 , n58222 , n58223 , n58224 , n58225 , n58226 , n58227 , n58228 , 
 n58229 , n58230 , n58231 , n58232 , n58233 , n58234 , n58235 , n58236 , n58237 , n58238 , 
 n58239 , n58240 , n58241 , n58242 , n58243 , n58244 , n58245 , n58246 , n58247 , n58248 , 
 n58249 , n58250 , n58251 , n58252 , n58253 , n58254 , n58255 , n58256 , n58257 , n58258 , 
 n58259 , n58260 , n58261 , n58262 , n58263 , n58264 , n58265 , n58266 , n58267 , n58268 , 
 n58269 , n58270 , n58271 , n58272 , n58273 , n58274 , n58275 , n58276 , n58277 , n58278 , 
 n58279 , n58280 , n58281 , n58282 , n58283 , n58284 , n58285 , n58286 , n58287 , n58288 , 
 n58289 , n58290 , n58291 , n58292 , n58293 , n58294 , n58295 , n58296 , n58297 , n58298 , 
 n58299 , n58300 , n58301 , n58302 , n58303 , n58304 , n58305 , n58306 , n58307 , n58308 , 
 n58309 , n58310 , n58311 , n58312 , n58313 , n58314 , n58315 , n58316 , n58317 , n58318 , 
 n58319 , n58320 , n58321 , n58322 , n58323 , n58324 , n58325 , n58326 , n58327 , n58328 , 
 n58329 , n58330 , n58331 , n58332 , n58333 , n58334 , n58335 , n58336 , n58337 , n58338 , 
 n58339 , n58340 , n58341 , n58342 , n58343 , n58344 , n58345 , n58346 , n58347 , n58348 , 
 n58349 , n58350 , n58351 , n58352 , n58353 , n58354 , n58355 , n58356 , n58357 , n58358 , 
 n58359 , n58360 , n58361 , n58362 , n58363 , n58364 , n58365 , n58366 , n58367 , n58368 , 
 n58369 , n58370 , n58371 , n58372 , n58373 , n58374 , n58375 , n58376 , n58377 , n58378 , 
 n58379 , n58380 , n58381 , n58382 , n58383 , n58384 , n58385 , n58386 , n58387 , n58388 , 
 n58389 , n58390 , n58391 , n58392 , n58393 , n58394 , n58395 , n58396 , n58397 , n58398 , 
 n58399 , n58400 , n58401 , n58402 , n58403 , n58404 , n58405 , n58406 , n58407 , n58408 , 
 n58409 , n58410 , n58411 , n58412 , n58413 , n58414 , n58415 , n58416 , n58417 , n58418 , 
 n58419 , n58420 , n58421 , n58422 , n58423 , n58424 , n58425 , n58426 , n58427 , n58428 , 
 n58429 , n58430 , n58431 , n58432 , n58433 , n58434 , n58435 , n58436 , n58437 , n58438 , 
 n58439 , n58440 , n58441 , n58442 , n58443 , n58444 , n58445 , n58446 , n58447 , n58448 , 
 n58449 , n58450 , n58451 , n58452 , n58453 , n58454 , n58455 , n58456 , n58457 , n58458 , 
 n58459 , n58460 , n58461 , n58462 , n58463 , n58464 , n58465 , n58466 , n58467 , n58468 , 
 n58469 , n58470 , n58471 , n58472 , n58473 , n58474 , n58475 , n58476 , n58477 , n58478 , 
 n58479 , n58480 , n58481 , n58482 , n58483 , n58484 , n58485 , n58486 , n58487 , n58488 , 
 n58489 , n58490 , n58491 , n58492 , n58493 , n58494 , n58495 , n58496 , n58497 , n58498 , 
 n58499 , n58500 , n58501 , n58502 , n58503 , n58504 , n58505 , n58506 , n58507 , n58508 , 
 n58509 , n58510 , n58511 , n58512 , n58513 , n58514 , n58515 , n58516 , n58517 , n58518 , 
 n58519 , n58520 , n58521 , n58522 , n58523 , n58524 , n58525 , n58526 , n58527 , n58528 , 
 n58529 , n58530 , n58531 , n58532 , n58533 , n58534 , n58535 , n58536 , n58537 , n58538 , 
 n58539 , n58540 , n58541 , n58542 , n58543 , n58544 , n58545 , n58546 , n58547 , n58548 , 
 n58549 , n58550 , n58551 , n58552 , n58553 , n58554 , n58555 , n58556 , n58557 , n58558 , 
 n58559 , n58560 , n58561 , n58562 , n58563 , n58564 , n58565 , n58566 , n58567 , n58568 , 
 n58569 , n58570 , n58571 , n58572 , n58573 , n58574 , n58575 , n58576 , n58577 , n58578 , 
 n58579 , n58580 , n58581 , n58582 , n58583 , n58584 , n58585 , n58586 , n58587 , n58588 , 
 n58589 , n58590 , n58591 , n58592 , n58593 , n58594 , n58595 , n58596 , n58597 , n58598 , 
 n58599 , n58600 , n58601 , n58602 , n58603 , n58604 , n58605 , n58606 , n58607 , n58608 , 
 n58609 , n58610 , n58611 , n58612 , n58613 , n58614 , n58615 , n58616 , n58617 , n58618 , 
 n58619 , n58620 , n58621 , n58622 , n58623 , n58624 , n58625 , n58626 , n58627 , n58628 , 
 n58629 , n58630 , n58631 , n58632 , n58633 , n58634 , n58635 , n58636 , n58637 , n58638 , 
 n58639 , n58640 , n58641 , n58642 , n58643 , n58644 , n58645 , n58646 , n58647 , n58648 , 
 n58649 , n58650 , n58651 , n58652 , n58653 , n58654 , n58655 , n58656 , n58657 , n58658 , 
 n58659 , n58660 , n58661 , n58662 , n58663 , n58664 , n58665 , n58666 , n58667 , n58668 , 
 n58669 , n58670 , n58671 , n58672 , n58673 , n58674 , n58675 , n58676 , n58677 , n58678 , 
 n58679 , n58680 , n58681 , n58682 , n58683 , n58684 , n58685 , n58686 , n58687 , n58688 , 
 n58689 , n58690 , n58691 , n58692 , n58693 , n58694 , n58695 , n58696 , n58697 , n58698 , 
 n58699 , n58700 , n58701 , n58702 , n58703 , n58704 , n58705 , n58706 , n58707 , n58708 , 
 n58709 , n58710 , n58711 , n58712 , n58713 , n58714 , n58715 , n58716 , n58717 , n58718 , 
 n58719 , n58720 , n58721 , n58722 , n58723 , n58724 , n58725 , n58726 , n58727 , n58728 , 
 n58729 , n58730 , n58731 , n58732 , n58733 , n58734 , n58735 , n58736 , n58737 , n58738 , 
 n58739 , n58740 , n58741 , n58742 , n58743 , n58744 , n58745 , n58746 , n58747 , n58748 , 
 n58749 , n58750 , n58751 , n58752 , n58753 , n58754 , n58755 , n58756 , n58757 , n58758 , 
 n58759 , n58760 , n58761 , n58762 , n58763 , n58764 , n58765 , n58766 , n58767 , n58768 , 
 n58769 , n58770 , n58771 , n58772 , n58773 , n58774 , n58775 , n58776 , n58777 , n58778 , 
 n58779 , n58780 , n58781 , n58782 , n58783 , n58784 , n58785 , n58786 , n58787 , n58788 , 
 n58789 , n58790 , n58791 , n58792 , n58793 , n58794 , n58795 , n58796 , n58797 , n58798 , 
 n58799 , n58800 , n58801 , n58802 , n58803 , n58804 , n58805 , n58806 , n58807 , n58808 , 
 n58809 , n58810 , n58811 , n58812 , n58813 , n58814 , n58815 , n58816 , n58817 , n58818 , 
 n58819 , n58820 , n58821 , n58822 , n58823 , n58824 , n58825 , n58826 , n58827 , n58828 , 
 n58829 , n58830 , n58831 , n58832 , n58833 , n58834 , n58835 , n58836 , n58837 , n58838 , 
 n58839 , n58840 , n58841 , n58842 , n58843 , n58844 , n58845 , n58846 , n58847 , n58848 , 
 n58849 , n58850 , n58851 , n58852 , n58853 , n58854 , n58855 , n58856 , n58857 , n58858 , 
 n58859 , n58860 , n58861 , n58862 , n58863 , n58864 , n58865 , n58866 , n58867 , n58868 , 
 n58869 , n58870 , n58871 , n58872 , n58873 , n58874 , n58875 , n58876 , n58877 , n58878 , 
 n58879 , n58880 , n58881 , n58882 , n58883 , n58884 , n58885 , n58886 , n58887 , n58888 , 
 n58889 , n58890 , n58891 , n58892 , n58893 , n58894 , n58895 , n58896 , n58897 , n58898 , 
 n58899 , n58900 , n58901 , n58902 , n58903 , n58904 , n58905 , n58906 , n58907 , n58908 , 
 n58909 , n58910 , n58911 , n58912 , n58913 , n58914 , n58915 , n58916 , n58917 , n58918 , 
 n58919 , n58920 , n58921 , n58922 , n58923 , n58924 , n58925 , n58926 , n58927 , n58928 , 
 n58929 , n58930 , n58931 , n58932 , n58933 , n58934 , n58935 , n58936 , n58937 , n58938 , 
 n58939 , n58940 , n58941 , n58942 , n58943 , n58944 , n58945 , n58946 , n58947 , n58948 , 
 n58949 , n58950 , n58951 , n58952 , n58953 , n58954 , n58955 , n58956 , n58957 , n58958 , 
 n58959 , n58960 , n58961 , n58962 , n58963 , n58964 , n58965 , n58966 , n58967 , n58968 , 
 n58969 , n58970 , n58971 , n58972 , n58973 , n58974 , n58975 , n58976 , n58977 , n58978 , 
 n58979 , n58980 , n58981 , n58982 , n58983 , n58984 , n58985 , n58986 , n58987 , n58988 , 
 n58989 , n58990 , n58991 , n58992 , n58993 , n58994 , n58995 , n58996 , n58997 , n58998 , 
 n58999 , n59000 , n59001 , n59002 , n59003 , n59004 , n59005 , n59006 , n59007 , n59008 , 
 n59009 , n59010 , n59011 , n59012 , n59013 , n59014 , n59015 , n59016 , n59017 , n59018 , 
 n59019 , n59020 , n59021 , n59022 , n59023 , n59024 , n59025 , n59026 , n59027 , n59028 , 
 n59029 , n59030 , n59031 , n59032 , n59033 , n59034 , n59035 , n59036 , n59037 , n59038 , 
 n59039 , n59040 , n59041 , n59042 , n59043 , n59044 , n59045 , n59046 , n59047 , n59048 , 
 n59049 , n59050 , n59051 , n59052 , n59053 , n59054 , n59055 , n59056 , n59057 , n59058 , 
 n59059 , n59060 , n59061 , n59062 , n59063 , n59064 , n59065 , n59066 , n59067 , n59068 , 
 n59069 , n59070 , n59071 , n59072 , n59073 , n59074 , n59075 , n59076 , n59077 , n59078 , 
 n59079 , n59080 , n59081 , n59082 , n59083 , n59084 , n59085 , n59086 , n59087 , n59088 , 
 n59089 , n59090 , n59091 , n59092 , n59093 , n59094 , n59095 , n59096 , n59097 , n59098 , 
 n59099 , n59100 , n59101 , n59102 , n59103 , n59104 , n59105 , n59106 , n59107 , n59108 , 
 n59109 , n59110 , n59111 , n59112 , n59113 , n59114 , n59115 , n59116 , n59117 , n59118 , 
 n59119 , n59120 , n59121 , n59122 , n59123 , n59124 , n59125 , n59126 , n59127 , n59128 , 
 n59129 , n59130 , n59131 , n59132 , n59133 , n59134 , n59135 , n59136 , n59137 , n59138 , 
 n59139 , n59140 , n59141 , n59142 , n59143 , n59144 , n59145 , n59146 , n59147 , n59148 , 
 n59149 , n59150 , n59151 , n59152 , n59153 , n59154 , n59155 , n59156 , n59157 , n59158 , 
 n59159 , n59160 , n59161 , n59162 , n59163 , n59164 , n59165 , n59166 , n59167 , n59168 , 
 n59169 , n59170 , n59171 , n59172 , n59173 , n59174 , n59175 , n59176 , n59177 , n59178 , 
 n59179 , n59180 , n59181 , n59182 , n59183 , n59184 , n59185 , n59186 , n59187 , n59188 , 
 n59189 , n59190 , n59191 , n59192 , n59193 , n59194 , n59195 , n59196 , n59197 , n59198 , 
 n59199 , n59200 , n59201 , n59202 , n59203 , n59204 , n59205 , n59206 , n59207 , n59208 , 
 n59209 , n59210 , n59211 , n59212 , n59213 , n59214 , n59215 , n59216 , n59217 , n59218 , 
 n59219 , n59220 , n59221 , n59222 , n59223 , n59224 , n59225 , n59226 , n59227 , n59228 , 
 n59229 , n59230 , n59231 , n59232 , n59233 , n59234 , n59235 , n59236 , n59237 , n59238 , 
 n59239 , n59240 , n59241 , n59242 , n59243 , n59244 , n59245 , n59246 , n59247 , n59248 , 
 n59249 , n59250 , n59251 , n59252 , n59253 , n59254 , n59255 , n59256 , n59257 , n59258 , 
 n59259 , n59260 , n59261 , n59262 , n59263 , n59264 , n59265 , n59266 , n59267 , n59268 , 
 n59269 , n59270 , n59271 , n59272 , n59273 , n59274 , n59275 , n59276 , n59277 , n59278 , 
 n59279 , n59280 , n59281 , n59282 , n59283 , n59284 , n59285 , n59286 , n59287 , n59288 , 
 n59289 , n59290 , n59291 , n59292 , n59293 , n59294 , n59295 , n59296 , n59297 , n59298 , 
 n59299 , n59300 , n59301 , n59302 , n59303 , n59304 , n59305 , n59306 , n59307 , n59308 , 
 n59309 , n59310 , n59311 , n59312 , n59313 , n59314 , n59315 , n59316 , n59317 , n59318 , 
 n59319 , n59320 , n59321 , n59322 , n59323 , n59324 , n59325 , n59326 , n59327 , n59328 , 
 n59329 , n59330 , n59331 , n59332 , n59333 , n59334 , n59335 , n59336 , n59337 , n59338 , 
 n59339 , n59340 , n59341 , n59342 , n59343 , n59344 , n59345 , n59346 , n59347 , n59348 , 
 n59349 , n59350 , n59351 , n59352 , n59353 , n59354 , n59355 , n59356 , n59357 , n59358 , 
 n59359 , n59360 , n59361 , n59362 , n59363 , n59364 , n59365 , n59366 , n59367 , n59368 , 
 n59369 , n59370 , n59371 , n59372 , n59373 , n59374 , n59375 , n59376 , n59377 , n59378 , 
 n59379 , n59380 , n59381 , n59382 , n59383 , n59384 , n59385 , n59386 , n59387 , n59388 , 
 n59389 , n59390 , n59391 , n59392 , n59393 , n59394 , n59395 , n59396 , n59397 , n59398 , 
 n59399 , n59400 , n59401 , n59402 , n59403 , n59404 , n59405 , n59406 , n59407 , n59408 , 
 n59409 , n59410 , n59411 , n59412 , n59413 , n59414 , n59415 , n59416 , n59417 , n59418 , 
 n59419 , n59420 , n59421 , n59422 , n59423 , n59424 , n59425 , n59426 , n59427 , n59428 , 
 n59429 , n59430 , n59431 , n59432 , n59433 , n59434 , n59435 , n59436 , n59437 , n59438 , 
 n59439 , n59440 , n59441 , n59442 , n59443 , n59444 , n59445 , n59446 , n59447 , n59448 , 
 n59449 , n59450 , n59451 , n59452 , n59453 , n59454 , n59455 , n59456 , n59457 , n59458 , 
 n59459 , n59460 , n59461 , n59462 , n59463 , n59464 , n59465 , n59466 , n59467 , n59468 , 
 n59469 , n59470 , n59471 , n59472 , n59473 , n59474 , n59475 , n59476 , n59477 , n59478 , 
 n59479 , n59480 , n59481 , n59482 , n59483 , n59484 , n59485 , n59486 , n59487 , n59488 , 
 n59489 , n59490 , n59491 , n59492 , n59493 , n59494 , n59495 , n59496 , n59497 , n59498 , 
 n59499 , n59500 , n59501 , n59502 , n59503 , n59504 , n59505 , n59506 , n59507 , n59508 , 
 n59509 , n59510 , n59511 , n59512 , n59513 , n59514 , n59515 , n59516 , n59517 , n59518 , 
 n59519 , n59520 , n59521 , n59522 , n59523 , n59524 , n59525 , n59526 , n59527 , n59528 , 
 n59529 , n59530 , n59531 , n59532 , n59533 , n59534 , n59535 , n59536 , n59537 , n59538 , 
 n59539 , n59540 , n59541 , n59542 , n59543 , n59544 , n59545 , n59546 , n59547 , n59548 , 
 n59549 , n59550 , n59551 , n59552 , n59553 , n59554 , n59555 , n59556 , n59557 , n59558 , 
 n59559 , n59560 , n59561 , n59562 , n59563 , n59564 , n59565 , n59566 , n59567 , n59568 , 
 n59569 , n59570 , n59571 , n59572 , n59573 , n59574 , n59575 , n59576 , n59577 , n59578 , 
 n59579 , n59580 , n59581 , n59582 , n59583 , n59584 , n59585 , n59586 , n59587 , n59588 , 
 n59589 , n59590 , n59591 , n59592 , n59593 , n59594 , n59595 , n59596 , n59597 , n59598 , 
 n59599 , n59600 , n59601 , n59602 , n59603 , n59604 , n59605 , n59606 , n59607 , n59608 , 
 n59609 , n59610 , n59611 , n59612 , n59613 , n59614 , n59615 , n59616 , n59617 , n59618 , 
 n59619 , n59620 , n59621 , n59622 , n59623 , n59624 , n59625 , n59626 , n59627 , n59628 , 
 n59629 , n59630 , n59631 , n59632 , n59633 , n59634 , n59635 , n59636 , n59637 , n59638 , 
 n59639 , n59640 , n59641 , n59642 , n59643 , n59644 , n59645 , n59646 , n59647 , n59648 , 
 n59649 , n59650 , n59651 , n59652 , n59653 , n59654 , n59655 , n59656 , n59657 , n59658 , 
 n59659 , n59660 , n59661 , n59662 , n59663 , n59664 , n59665 , n59666 , n59667 , n59668 , 
 n59669 , n59670 , n59671 , n59672 , n59673 , n59674 , n59675 , n59676 , n59677 , n59678 , 
 n59679 , n59680 , n59681 , n59682 , n59683 , n59684 , n59685 , n59686 , n59687 , n59688 , 
 n59689 , n59690 , n59691 , n59692 , n59693 , n59694 , n59695 , n59696 , n59697 , n59698 , 
 n59699 , n59700 , n59701 , n59702 , n59703 , n59704 , n59705 , n59706 , n59707 , n59708 , 
 n59709 , n59710 , n59711 , n59712 , n59713 , n59714 , n59715 , n59716 , n59717 , n59718 , 
 n59719 , n59720 , n59721 , n59722 , n59723 , n59724 , n59725 , n59726 , n59727 , n59728 , 
 n59729 , n59730 , n59731 , n59732 , n59733 , n59734 , n59735 , n59736 , n59737 , n59738 , 
 n59739 , n59740 , n59741 , n59742 , n59743 , n59744 , n59745 , n59746 , n59747 , n59748 , 
 n59749 , n59750 , n59751 , n59752 , n59753 , n59754 , n59755 , n59756 , n59757 , n59758 , 
 n59759 , n59760 , n59761 , n59762 , n59763 , n59764 , n59765 , n59766 , n59767 , n59768 , 
 n59769 , n59770 , n59771 , n59772 , n59773 , n59774 , n59775 , n59776 , n59777 , n59778 , 
 n59779 , n59780 , n59781 , n59782 , n59783 , n59784 , n59785 , n59786 , n59787 , n59788 , 
 n59789 , n59790 , n59791 , n59792 , n59793 , n59794 , n59795 , n59796 , n59797 , n59798 , 
 n59799 , n59800 , n59801 , n59802 , n59803 , n59804 , n59805 , n59806 , n59807 , n59808 , 
 n59809 , n59810 , n59811 , n59812 , n59813 , n59814 , n59815 , n59816 , n59817 , n59818 , 
 n59819 , n59820 , n59821 , n59822 , n59823 , n59824 , n59825 , n59826 , n59827 , n59828 , 
 n59829 , n59830 , n59831 , n59832 , n59833 , n59834 , n59835 , n59836 , n59837 , n59838 , 
 n59839 , n59840 , n59841 , n59842 , n59843 , n59844 , n59845 , n59846 , n59847 , n59848 , 
 n59849 , n59850 , n59851 , n59852 , n59853 , n59854 , n59855 , n59856 , n59857 , n59858 , 
 n59859 , n59860 , n59861 , n59862 , n59863 , n59864 , n59865 , n59866 , n59867 , n59868 , 
 n59869 , n59870 , n59871 , n59872 , n59873 , n59874 , n59875 , n59876 , n59877 , n59878 , 
 n59879 , n59880 , n59881 , n59882 , n59883 , n59884 , n59885 , n59886 , n59887 , n59888 , 
 n59889 , n59890 , n59891 , n59892 , n59893 , n59894 , n59895 , n59896 , n59897 , n59898 , 
 n59899 , n59900 , n59901 , n59902 , n59903 , n59904 , n59905 , n59906 , n59907 , n59908 , 
 n59909 , n59910 , n59911 , n59912 , n59913 , n59914 , n59915 , n59916 , n59917 , n59918 , 
 n59919 , n59920 , n59921 , n59922 , n59923 , n59924 , n59925 , n59926 , n59927 , n59928 , 
 n59929 , n59930 , n59931 , n59932 , n59933 , n59934 , n59935 , n59936 , n59937 , n59938 , 
 n59939 , n59940 , n59941 , n59942 , n59943 , n59944 , n59945 , n59946 , n59947 , n59948 , 
 n59949 , n59950 , n59951 , n59952 , n59953 , n59954 , n59955 , n59956 , n59957 , n59958 , 
 n59959 , n59960 , n59961 , n59962 , n59963 , n59964 , n59965 , n59966 , n59967 , n59968 , 
 n59969 , n59970 , n59971 , n59972 , n59973 , n59974 , n59975 , n59976 , n59977 , n59978 , 
 n59979 , n59980 , n59981 , n59982 , n59983 , n59984 , n59985 , n59986 , n59987 , n59988 , 
 n59989 , n59990 , n59991 , n59992 , n59993 , n59994 , n59995 , n59996 , n59997 , n59998 , 
 n59999 , n60000 , n60001 , n60002 , n60003 , n60004 , n60005 , n60006 , n60007 , n60008 , 
 n60009 , n60010 , n60011 , n60012 , n60013 , n60014 , n60015 , n60016 , n60017 , n60018 , 
 n60019 , n60020 , n60021 , n60022 , n60023 , n60024 , n60025 , n60026 , n60027 , n60028 , 
 n60029 , n60030 , n60031 , n60032 , n60033 , n60034 , n60035 , n60036 , n60037 , n60038 , 
 n60039 , n60040 , n60041 , n60042 , n60043 , n60044 , n60045 , n60046 , n60047 , n60048 , 
 n60049 , n60050 , n60051 , n60052 , n60053 , n60054 , n60055 , n60056 , n60057 , n60058 , 
 n60059 , n60060 , n60061 , n60062 , n60063 , n60064 , n60065 , n60066 , n60067 , n60068 , 
 n60069 , n60070 , n60071 , n60072 , n60073 , n60074 , n60075 , n60076 , n60077 , n60078 , 
 n60079 , n60080 , n60081 , n60082 , n60083 , n60084 , n60085 , n60086 , n60087 , n60088 , 
 n60089 , n60090 , n60091 , n60092 , n60093 , n60094 , n60095 , n60096 , n60097 , n60098 , 
 n60099 , n60100 , n60101 , n60102 , n60103 , n60104 , n60105 , n60106 , n60107 , n60108 , 
 n60109 , n60110 , n60111 , n60112 , n60113 , n60114 , n60115 , n60116 , n60117 , n60118 , 
 n60119 , n60120 , n60121 , n60122 , n60123 , n60124 , n60125 , n60126 , n60127 , n60128 , 
 n60129 , n60130 , n60131 , n60132 , n60133 , n60134 , n60135 , n60136 , n60137 , n60138 , 
 n60139 , n60140 , n60141 , n60142 , n60143 , n60144 , n60145 , n60146 , n60147 , n60148 , 
 n60149 , n60150 , n60151 , n60152 , n60153 , n60154 , n60155 , n60156 , n60157 , n60158 , 
 n60159 , n60160 , n60161 , n60162 , n60163 , n60164 , n60165 , n60166 , n60167 , n60168 , 
 n60169 , n60170 , n60171 , n60172 , n60173 , n60174 , n60175 , n60176 , n60177 , n60178 , 
 n60179 , n60180 , n60181 , n60182 , n60183 , n60184 , n60185 , n60186 , n60187 , n60188 , 
 n60189 , n60190 , n60191 , n60192 , n60193 , n60194 , n60195 , n60196 , n60197 , n60198 , 
 n60199 , n60200 , n60201 , n60202 , n60203 , n60204 , n60205 , n60206 , n60207 , n60208 , 
 n60209 , n60210 , n60211 , n60212 , n60213 , n60214 , n60215 , n60216 , n60217 , n60218 , 
 n60219 , n60220 , n60221 , n60222 , n60223 , n60224 , n60225 , n60226 , n60227 , n60228 , 
 n60229 , n60230 , n60231 , n60232 , n60233 , n60234 , n60235 , n60236 , n60237 , n60238 , 
 n60239 , n60240 , n60241 , n60242 , n60243 , n60244 , n60245 , n60246 , n60247 , n60248 , 
 n60249 , n60250 , n60251 , n60252 , n60253 , n60254 , n60255 , n60256 , n60257 , n60258 , 
 n60259 , n60260 , n60261 , n60262 , n60263 , n60264 , n60265 , n60266 , n60267 , n60268 , 
 n60269 , n60270 , n60271 , n60272 , n60273 , n60274 , n60275 , n60276 , n60277 , n60278 , 
 n60279 , n60280 , n60281 , n60282 , n60283 , n60284 , n60285 , n60286 , n60287 , n60288 , 
 n60289 , n60290 , n60291 , n60292 , n60293 , n60294 , n60295 , n60296 , n60297 , n60298 , 
 n60299 , n60300 , n60301 , n60302 , n60303 , n60304 , n60305 , n60306 , n60307 , n60308 , 
 n60309 , n60310 , n60311 , n60312 , n60313 , n60314 , n60315 , n60316 , n60317 , n60318 , 
 n60319 , n60320 , n60321 , n60322 , n60323 , n60324 , n60325 , n60326 , n60327 , n60328 , 
 n60329 , n60330 , n60331 , n60332 , n60333 , n60334 , n60335 , n60336 , n60337 , n60338 , 
 n60339 , n60340 , n60341 , n60342 , n60343 , n60344 , n60345 , n60346 , n60347 , n60348 , 
 n60349 , n60350 , n60351 , n60352 , n60353 , n60354 , n60355 , n60356 , n60357 , n60358 , 
 n60359 , n60360 , n60361 , n60362 , n60363 , n60364 , n60365 , n60366 , n60367 , n60368 , 
 n60369 , n60370 , n60371 , n60372 , n60373 , n60374 , n60375 , n60376 , n60377 , n60378 , 
 n60379 , n60380 , n60381 , n60382 , n60383 , n60384 , n60385 , n60386 , n60387 , n60388 , 
 n60389 , n60390 , n60391 , n60392 , n60393 , n60394 , n60395 , n60396 , n60397 , n60398 , 
 n60399 , n60400 , n60401 , n60402 , n60403 , n60404 , n60405 , n60406 , n60407 , n60408 , 
 n60409 , n60410 , n60411 , n60412 , n60413 , n60414 , n60415 , n60416 , n60417 , n60418 , 
 n60419 , n60420 , n60421 , n60422 , n60423 , n60424 , n60425 , n60426 , n60427 , n60428 , 
 n60429 , n60430 , n60431 , n60432 , n60433 , n60434 , n60435 , n60436 , n60437 , n60438 , 
 n60439 , n60440 , n60441 , n60442 , n60443 , n60444 , n60445 , n60446 , n60447 , n60448 , 
 n60449 , n60450 , n60451 , n60452 , n60453 , n60454 , n60455 , n60456 , n60457 , n60458 , 
 n60459 , n60460 , n60461 , n60462 , n60463 , n60464 , n60465 , n60466 , n60467 , n60468 , 
 n60469 , n60470 , n60471 , n60472 , n60473 , n60474 , n60475 , n60476 , n60477 , n60478 , 
 n60479 , n60480 , n60481 , n60482 , n60483 , n60484 , n60485 , n60486 , n60487 , n60488 , 
 n60489 , n60490 , n60491 , n60492 , n60493 , n60494 , n60495 , n60496 , n60497 , n60498 , 
 n60499 , n60500 , n60501 , n60502 , n60503 , n60504 , n60505 , n60506 , n60507 , n60508 , 
 n60509 , n60510 , n60511 , n60512 , n60513 , n60514 , n60515 , n60516 , n60517 , n60518 , 
 n60519 , n60520 , n60521 , n60522 , n60523 , n60524 , n60525 , n60526 , n60527 , n60528 , 
 n60529 , n60530 , n60531 , n60532 , n60533 , n60534 , n60535 , n60536 , n60537 , n60538 , 
 n60539 , n60540 , n60541 , n60542 , n60543 , n60544 , n60545 , n60546 , n60547 , n60548 , 
 n60549 , n60550 , n60551 , n60552 , n60553 , n60554 , n60555 , n60556 , n60557 , n60558 , 
 n60559 , n60560 , n60561 , n60562 , n60563 , n60564 , n60565 , n60566 , n60567 , n60568 , 
 n60569 , n60570 , n60571 , n60572 , n60573 , n60574 , n60575 , n60576 , n60577 , n60578 , 
 n60579 , n60580 , n60581 , n60582 , n60583 , n60584 , n60585 , n60586 , n60587 , n60588 , 
 n60589 , n60590 , n60591 , n60592 , n60593 , n60594 , n60595 , n60596 , n60597 , n60598 , 
 n60599 , n60600 , n60601 , n60602 , n60603 , n60604 , n60605 , n60606 , n60607 , n60608 , 
 n60609 , n60610 , n60611 , n60612 , n60613 , n60614 , n60615 , n60616 , n60617 , n60618 , 
 n60619 , n60620 , n60621 , n60622 , n60623 , n60624 , n60625 , n60626 , n60627 , n60628 , 
 n60629 , n60630 , n60631 , n60632 , n60633 , n60634 , n60635 , n60636 , n60637 , n60638 , 
 n60639 , n60640 , n60641 , n60642 , n60643 , n60644 , n60645 , n60646 , n60647 , n60648 , 
 n60649 , n60650 , n60651 , n60652 , n60653 , n60654 , n60655 , n60656 , n60657 , n60658 , 
 n60659 , n60660 , n60661 , n60662 , n60663 , n60664 , n60665 , n60666 , n60667 , n60668 , 
 n60669 , n60670 , n60671 , n60672 , n60673 , n60674 , n60675 , n60676 , n60677 , n60678 , 
 n60679 , n60680 , n60681 , n60682 , n60683 , n60684 , n60685 , n60686 , n60687 , n60688 , 
 n60689 , n60690 , n60691 , n60692 , n60693 , n60694 , n60695 , n60696 , n60697 , n60698 , 
 n60699 , n60700 , n60701 , n60702 , n60703 , n60704 , n60705 , n60706 , n60707 , n60708 , 
 n60709 , n60710 , n60711 , n60712 , n60713 , n60714 , n60715 , n60716 , n60717 , n60718 , 
 n60719 , n60720 , n60721 , n60722 , n60723 , n60724 , n60725 , n60726 , n60727 , n60728 , 
 n60729 , n60730 , n60731 , n60732 , n60733 , n60734 , n60735 , n60736 , n60737 , n60738 , 
 n60739 , n60740 , n60741 , n60742 , n60743 , n60744 , n60745 , n60746 , n60747 , n60748 , 
 n60749 , n60750 , n60751 , n60752 , n60753 , n60754 , n60755 , n60756 , n60757 , n60758 , 
 n60759 , n60760 , n60761 , n60762 , n60763 , n60764 , n60765 , n60766 , n60767 , n60768 , 
 n60769 , n60770 , n60771 , n60772 , n60773 , n60774 , n60775 , n60776 , n60777 , n60778 , 
 n60779 , n60780 , n60781 , n60782 , n60783 , n60784 , n60785 , n60786 , n60787 , n60788 , 
 n60789 , n60790 , n60791 , n60792 , n60793 , n60794 , n60795 , n60796 , n60797 , n60798 , 
 n60799 , n60800 , n60801 , n60802 , n60803 , n60804 , n60805 , n60806 , n60807 , n60808 , 
 n60809 , n60810 , n60811 , n60812 , n60813 , n60814 , n60815 , n60816 , n60817 , n60818 , 
 n60819 , n60820 , n60821 , n60822 , n60823 , n60824 , n60825 , n60826 , n60827 , n60828 , 
 n60829 , n60830 , n60831 , n60832 , n60833 , n60834 , n60835 , n60836 , n60837 , n60838 , 
 n60839 , n60840 , n60841 , n60842 , n60843 , n60844 , n60845 , n60846 , n60847 , n60848 , 
 n60849 , n60850 , n60851 , n60852 , n60853 , n60854 , n60855 , n60856 , n60857 , n60858 , 
 n60859 , n60860 , n60861 , n60862 , n60863 , n60864 , n60865 , n60866 , n60867 , n60868 , 
 n60869 , n60870 , n60871 , n60872 , n60873 , n60874 , n60875 , n60876 , n60877 , n60878 , 
 n60879 , n60880 , n60881 , n60882 , n60883 , n60884 , n60885 , n60886 , n60887 , n60888 , 
 n60889 , n60890 , n60891 , n60892 , n60893 , n60894 , n60895 , n60896 , n60897 , n60898 , 
 n60899 , n60900 , n60901 , n60902 , n60903 , n60904 , n60905 , n60906 , n60907 , n60908 , 
 n60909 , n60910 , n60911 , n60912 , n60913 , n60914 , n60915 , n60916 , n60917 , n60918 , 
 n60919 , n60920 , n60921 , n60922 , n60923 , n60924 , n60925 , n60926 , n60927 , n60928 , 
 n60929 , n60930 , n60931 , n60932 , n60933 , n60934 , n60935 , n60936 , n60937 , n60938 , 
 n60939 , n60940 , n60941 , n60942 , n60943 , n60944 , n60945 , n60946 , n60947 , n60948 , 
 n60949 , n60950 , n60951 , n60952 , n60953 , n60954 , n60955 , n60956 , n60957 , n60958 , 
 n60959 , n60960 , n60961 , n60962 , n60963 , n60964 , n60965 , n60966 , n60967 , n60968 , 
 n60969 , n60970 , n60971 , n60972 , n60973 , n60974 , n60975 , n60976 , n60977 , n60978 , 
 n60979 , n60980 , n60981 , n60982 , n60983 , n60984 , n60985 , n60986 , n60987 , n60988 , 
 n60989 , n60990 , n60991 , n60992 , n60993 , n60994 , n60995 , n60996 , n60997 , n60998 , 
 n60999 , n61000 , n61001 , n61002 , n61003 , n61004 , n61005 , n61006 , n61007 , n61008 , 
 n61009 , n61010 , n61011 , n61012 , n61013 , n61014 , n61015 , n61016 , n61017 , n61018 , 
 n61019 , n61020 , n61021 , n61022 , n61023 , n61024 , n61025 , n61026 , n61027 , n61028 , 
 n61029 , n61030 , n61031 , n61032 , n61033 , n61034 , n61035 , n61036 , n61037 , n61038 , 
 n61039 , n61040 , n61041 , n61042 , n61043 , n61044 , n61045 , n61046 , n61047 , n61048 , 
 n61049 , n61050 , n61051 , n61052 , n61053 , n61054 , n61055 , n61056 , n61057 , n61058 , 
 n61059 , n61060 , n61061 , n61062 , n61063 , n61064 , n61065 , n61066 , n61067 , n61068 , 
 n61069 , n61070 , n61071 , n61072 , n61073 , n61074 , n61075 , n61076 , n61077 , n61078 , 
 n61079 , n61080 , n61081 , n61082 , n61083 , n61084 , n61085 , n61086 , n61087 , n61088 , 
 n61089 , n61090 , n61091 , n61092 , n61093 , n61094 , n61095 , n61096 , n61097 , n61098 , 
 n61099 , n61100 , n61101 , n61102 , n61103 , n61104 , n61105 , n61106 , n61107 , n61108 , 
 n61109 , n61110 , n61111 , n61112 , n61113 , n61114 , n61115 , n61116 , n61117 , n61118 , 
 n61119 , n61120 , n61121 , n61122 , n61123 , n61124 , n61125 , n61126 , n61127 , n61128 , 
 n61129 , n61130 , n61131 , n61132 , n61133 , n61134 , n61135 , n61136 , n61137 , n61138 , 
 n61139 , n61140 , n61141 , n61142 , n61143 , n61144 , n61145 , n61146 , n61147 , n61148 , 
 n61149 , n61150 , n61151 , n61152 , n61153 , n61154 , n61155 , n61156 , n61157 , n61158 , 
 n61159 , n61160 , n61161 , n61162 , n61163 , n61164 , n61165 , n61166 , n61167 , n61168 , 
 n61169 , n61170 , n61171 , n61172 , n61173 , n61174 , n61175 , n61176 , n61177 , n61178 , 
 n61179 , n61180 , n61181 , n61182 , n61183 , n61184 , n61185 , n61186 , n61187 , n61188 , 
 n61189 , n61190 , n61191 , n61192 , n61193 , n61194 , n61195 , n61196 , n61197 , n61198 , 
 n61199 , n61200 , n61201 , n61202 , n61203 , n61204 , n61205 , n61206 , n61207 , n61208 , 
 n61209 , n61210 , n61211 , n61212 , n61213 , n61214 , n61215 , n61216 , n61217 , n61218 , 
 n61219 , n61220 , n61221 , n61222 , n61223 , n61224 , n61225 , n61226 , n61227 , n61228 , 
 n61229 , n61230 , n61231 , n61232 , n61233 , n61234 , n61235 , n61236 , n61237 , n61238 , 
 n61239 , n61240 , n61241 , n61242 , n61243 , n61244 , n61245 , n61246 , n61247 , n61248 , 
 n61249 , n61250 , n61251 , n61252 , n61253 , n61254 , n61255 , n61256 , n61257 , n61258 , 
 n61259 , n61260 , n61261 , n61262 , n61263 , n61264 , n61265 , n61266 , n61267 , n61268 , 
 n61269 , n61270 , n61271 , n61272 , n61273 , n61274 , n61275 , n61276 , n61277 , n61278 , 
 n61279 , n61280 , n61281 , n61282 , n61283 , n61284 , n61285 , n61286 , n61287 , n61288 , 
 n61289 , n61290 , n61291 , n61292 , n61293 , n61294 , n61295 , n61296 , n61297 , n61298 , 
 n61299 , n61300 , n61301 , n61302 , n61303 , n61304 , n61305 , n61306 , n61307 , n61308 , 
 n61309 , n61310 , n61311 , n61312 , n61313 , n61314 , n61315 , n61316 , n61317 , n61318 , 
 n61319 , n61320 , n61321 , n61322 , n61323 , n61324 , n61325 , n61326 , n61327 , n61328 , 
 n61329 , n61330 , n61331 , n61332 , n61333 , n61334 , n61335 , n61336 , n61337 , n61338 , 
 n61339 , n61340 , n61341 , n61342 , n61343 , n61344 , n61345 , n61346 , n61347 , n61348 , 
 n61349 , n61350 , n61351 , n61352 , n61353 , n61354 , n61355 , n61356 , n61357 , n61358 , 
 n61359 , n61360 , n61361 , n61362 , n61363 , n61364 , n61365 , n61366 , n61367 , n61368 , 
 n61369 , n61370 , n61371 , n61372 , n61373 , n61374 , n61375 , n61376 , n61377 , n61378 , 
 n61379 , n61380 , n61381 , n61382 , n61383 , n61384 , n61385 , n61386 , n61387 , n61388 , 
 n61389 , n61390 , n61391 , n61392 , n61393 , n61394 , n61395 , n61396 , n61397 , n61398 , 
 n61399 , n61400 , n61401 , n61402 , n61403 , n61404 , n61405 , n61406 , n61407 , n61408 , 
 n61409 , n61410 , n61411 , n61412 , n61413 , n61414 , n61415 , n61416 , n61417 , n61418 , 
 n61419 , n61420 , n61421 , n61422 , n61423 , n61424 , n61425 , n61426 , n61427 , n61428 , 
 n61429 , n61430 , n61431 , n61432 , n61433 , n61434 , n61435 , n61436 , n61437 , n61438 , 
 n61439 , n61440 , n61441 , n61442 , n61443 , n61444 , n61445 , n61446 , n61447 , n61448 , 
 n61449 , n61450 , n61451 , n61452 , n61453 , n61454 , n61455 , n61456 , n61457 , n61458 , 
 n61459 , n61460 , n61461 , n61462 , n61463 , n61464 , n61465 , n61466 , n61467 , n61468 , 
 n61469 , n61470 , n61471 , n61472 , n61473 , n61474 , n61475 , n61476 , n61477 , n61478 , 
 n61479 , n61480 , n61481 , n61482 , n61483 , n61484 , n61485 , n61486 , n61487 , n61488 , 
 n61489 , n61490 , n61491 , n61492 , n61493 , n61494 , n61495 , n61496 , n61497 , n61498 , 
 n61499 , n61500 , n61501 , n61502 , n61503 , n61504 , n61505 , n61506 , n61507 , n61508 , 
 n61509 , n61510 , n61511 , n61512 , n61513 , n61514 , n61515 , n61516 , n61517 , n61518 , 
 n61519 , n61520 , n61521 , n61522 , n61523 , n61524 , n61525 , n61526 , n61527 , n61528 , 
 n61529 , n61530 , n61531 , n61532 , n61533 , n61534 , n61535 , n61536 , n61537 , n61538 , 
 n61539 , n61540 , n61541 , n61542 , n61543 , n61544 , n61545 , n61546 , n61547 , n61548 , 
 n61549 , n61550 , n61551 , n61552 , n61553 , n61554 , n61555 , n61556 , n61557 , n61558 , 
 n61559 , n61560 , n61561 , n61562 , n61563 , n61564 , n61565 , n61566 , n61567 , n61568 , 
 n61569 , n61570 , n61571 , n61572 , n61573 , n61574 , n61575 , n61576 , n61577 , n61578 , 
 n61579 , n61580 , n61581 , n61582 , n61583 , n61584 , n61585 , n61586 , n61587 , n61588 , 
 n61589 , n61590 , n61591 , n61592 , n61593 , n61594 , n61595 , n61596 , n61597 , n61598 , 
 n61599 , n61600 , n61601 , n61602 , n61603 , n61604 , n61605 , n61606 , n61607 , n61608 , 
 n61609 , n61610 , n61611 , n61612 , n61613 , n61614 , n61615 , n61616 , n61617 , n61618 , 
 n61619 , n61620 , n61621 , n61622 , n61623 , n61624 , n61625 , n61626 , n61627 , n61628 , 
 n61629 , n61630 , n61631 , n61632 , n61633 , n61634 , n61635 , n61636 , n61637 , n61638 , 
 n61639 , n61640 , n61641 , n61642 , n61643 , n61644 , n61645 , n61646 , n61647 , n61648 , 
 n61649 , n61650 , n61651 , n61652 , n61653 , n61654 , n61655 , n61656 , n61657 , n61658 , 
 n61659 , n61660 , n61661 , n61662 , n61663 , n61664 , n61665 , n61666 , n61667 , n61668 , 
 n61669 , n61670 , n61671 , n61672 , n61673 , n61674 , n61675 , n61676 , n61677 , n61678 , 
 n61679 , n61680 , n61681 , n61682 , n61683 , n61684 , n61685 , n61686 , n61687 , n61688 , 
 n61689 , n61690 , n61691 , n61692 , n61693 , n61694 , n61695 , n61696 , n61697 , n61698 , 
 n61699 , n61700 , n61701 , n61702 , n61703 , n61704 , n61705 , n61706 , n61707 , n61708 , 
 n61709 , n61710 , n61711 , n61712 , n61713 , n61714 , n61715 , n61716 , n61717 , n61718 , 
 n61719 , n61720 , n61721 , n61722 , n61723 , n61724 , n61725 , n61726 , n61727 , n61728 , 
 n61729 , n61730 , n61731 , n61732 , n61733 , n61734 , n61735 , n61736 , n61737 , n61738 , 
 n61739 , n61740 , n61741 , n61742 , n61743 , n61744 , n61745 , n61746 , n61747 , n61748 , 
 n61749 , n61750 , n61751 , n61752 , n61753 , n61754 , n61755 , n61756 , n61757 , n61758 , 
 n61759 , n61760 , n61761 , n61762 , n61763 , n61764 , n61765 , n61766 , n61767 , n61768 , 
 n61769 , n61770 , n61771 , n61772 , n61773 , n61774 , n61775 , n61776 , n61777 , n61778 , 
 n61779 , n61780 , n61781 , n61782 , n61783 , n61784 , n61785 , n61786 , n61787 , n61788 , 
 n61789 , n61790 , n61791 , n61792 , n61793 , n61794 , n61795 , n61796 , n61797 , n61798 , 
 n61799 , n61800 , n61801 , n61802 , n61803 , n61804 , n61805 , n61806 , n61807 , n61808 , 
 n61809 , n61810 , n61811 , n61812 , n61813 , n61814 , n61815 , n61816 , n61817 , n61818 , 
 n61819 , n61820 , n61821 , n61822 , n61823 , n61824 , n61825 , n61826 , n61827 , n61828 , 
 n61829 , n61830 , n61831 , n61832 , n61833 , n61834 , n61835 , n61836 , n61837 , n61838 , 
 n61839 , n61840 , n61841 , n61842 , n61843 , n61844 , n61845 , n61846 , n61847 , n61848 , 
 n61849 , n61850 , n61851 , n61852 , n61853 , n61854 , n61855 , n61856 , n61857 , n61858 , 
 n61859 , n61860 , n61861 , n61862 , n61863 , n61864 , n61865 , n61866 , n61867 , n61868 , 
 n61869 , n61870 , n61871 , n61872 , n61873 , n61874 , n61875 , n61876 , n61877 , n61878 , 
 n61879 , n61880 , n61881 , n61882 , n61883 , n61884 , n61885 , n61886 , n61887 , n61888 , 
 n61889 , n61890 , n61891 , n61892 , n61893 , n61894 , n61895 , n61896 , n61897 , n61898 , 
 n61899 , n61900 , n61901 , n61902 , n61903 , n61904 , n61905 , n61906 , n61907 , n61908 , 
 n61909 , n61910 , n61911 , n61912 , n61913 , n61914 , n61915 , n61916 , n61917 , n61918 , 
 n61919 , n61920 , n61921 , n61922 , n61923 , n61924 , n61925 , n61926 , n61927 , n61928 , 
 n61929 , n61930 , n61931 , n61932 , n61933 , n61934 , n61935 , n61936 , n61937 , n61938 , 
 n61939 , n61940 , n61941 , n61942 , n61943 , n61944 , n61945 , n61946 , n61947 , n61948 , 
 n61949 , n61950 , n61951 , n61952 , n61953 , n61954 , n61955 , n61956 , n61957 , n61958 , 
 n61959 , n61960 , n61961 , n61962 , n61963 , n61964 , n61965 , n61966 , n61967 , n61968 , 
 n61969 , n61970 , n61971 , n61972 , n61973 , n61974 , n61975 , n61976 , n61977 , n61978 , 
 n61979 , n61980 , n61981 , n61982 , n61983 , n61984 , n61985 , n61986 , n61987 , n61988 , 
 n61989 , n61990 , n61991 , n61992 , n61993 , n61994 , n61995 , n61996 , n61997 , n61998 , 
 n61999 , n62000 , n62001 , n62002 , n62003 , n62004 , n62005 , n62006 , n62007 , n62008 , 
 n62009 , n62010 , n62011 , n62012 , n62013 , n62014 , n62015 , n62016 , n62017 , n62018 , 
 n62019 , n62020 , n62021 , n62022 , n62023 , n62024 , n62025 , n62026 , n62027 , n62028 , 
 n62029 , n62030 , n62031 , n62032 , n62033 , n62034 , n62035 , n62036 , n62037 , n62038 , 
 n62039 , n62040 , n62041 , n62042 , n62043 , n62044 , n62045 , n62046 , n62047 , n62048 , 
 n62049 , n62050 , n62051 , n62052 , n62053 , n62054 , n62055 , n62056 , n62057 , n62058 , 
 n62059 , n62060 , n62061 , n62062 , n62063 , n62064 , n62065 , n62066 , n62067 , n62068 , 
 n62069 , n62070 , n62071 , n62072 , n62073 , n62074 , n62075 , n62076 , n62077 , n62078 , 
 n62079 , n62080 , n62081 , n62082 , n62083 , n62084 , n62085 , n62086 , n62087 , n62088 , 
 n62089 , n62090 , n62091 , n62092 , n62093 , n62094 , n62095 , n62096 , n62097 , n62098 , 
 n62099 , n62100 , n62101 , n62102 , n62103 , n62104 , n62105 , n62106 , n62107 , n62108 , 
 n62109 , n62110 , n62111 , n62112 , n62113 , n62114 , n62115 , n62116 , n62117 , n62118 , 
 n62119 , n62120 , n62121 , n62122 , n62123 , n62124 , n62125 , n62126 , n62127 , n62128 , 
 n62129 , n62130 , n62131 , n62132 , n62133 , n62134 , n62135 , n62136 , n62137 , n62138 , 
 n62139 , n62140 , n62141 , n62142 , n62143 , n62144 , n62145 , n62146 , n62147 , n62148 , 
 n62149 , n62150 , n62151 , n62152 , n62153 , n62154 , n62155 , n62156 , n62157 , n62158 , 
 n62159 , n62160 , n62161 , n62162 , n62163 , n62164 , n62165 , n62166 , n62167 , n62168 , 
 n62169 , n62170 , n62171 , n62172 , n62173 , n62174 , n62175 , n62176 , n62177 , n62178 , 
 n62179 , n62180 , n62181 , n62182 , n62183 , n62184 , n62185 , n62186 , n62187 , n62188 , 
 n62189 , n62190 , n62191 , n62192 , n62193 , n62194 , n62195 , n62196 , n62197 , n62198 , 
 n62199 , n62200 , n62201 , n62202 , n62203 , n62204 , n62205 , n62206 , n62207 , n62208 , 
 n62209 , n62210 , n62211 , n62212 , n62213 , n62214 , n62215 , n62216 , n62217 , n62218 , 
 n62219 , n62220 , n62221 , n62222 , n62223 , n62224 , n62225 , n62226 , n62227 , n62228 , 
 n62229 , n62230 , n62231 , n62232 , n62233 , n62234 , n62235 , n62236 , n62237 , n62238 , 
 n62239 , n62240 , n62241 , n62242 , n62243 , n62244 , n62245 , n62246 , n62247 , n62248 , 
 n62249 , n62250 , n62251 , n62252 , n62253 , n62254 , n62255 , n62256 , n62257 , n62258 , 
 n62259 , n62260 , n62261 , n62262 , n62263 , n62264 , n62265 , n62266 , n62267 , n62268 , 
 n62269 , n62270 , n62271 , n62272 , n62273 , n62274 , n62275 , n62276 , n62277 , n62278 , 
 n62279 , n62280 , n62281 , n62282 , n62283 , n62284 , n62285 , n62286 , n62287 , n62288 , 
 n62289 , n62290 , n62291 , n62292 , n62293 , n62294 , n62295 , n62296 , n62297 , n62298 , 
 n62299 , n62300 , n62301 , n62302 , n62303 , n62304 , n62305 , n62306 , n62307 , n62308 , 
 n62309 , n62310 , n62311 , n62312 , n62313 , n62314 , n62315 , n62316 , n62317 , n62318 , 
 n62319 , n62320 , n62321 , n62322 , n62323 , n62324 , n62325 , n62326 , n62327 , n62328 , 
 n62329 , n62330 , n62331 , n62332 , n62333 , n62334 , n62335 , n62336 , n62337 , n62338 , 
 n62339 , n62340 , n62341 , n62342 , n62343 , n62344 , n62345 , n62346 , n62347 , n62348 , 
 n62349 , n62350 , n62351 , n62352 , n62353 , n62354 , n62355 , n62356 , n62357 , n62358 , 
 n62359 , n62360 , n62361 , n62362 , n62363 , n62364 , n62365 , n62366 , n62367 , n62368 , 
 n62369 , n62370 , n62371 , n62372 , n62373 , n62374 , n62375 , n62376 , n62377 , n62378 , 
 n62379 , n62380 , n62381 , n62382 , n62383 , n62384 , n62385 , n62386 , n62387 , n62388 , 
 n62389 , n62390 , n62391 , n62392 , n62393 , n62394 , n62395 , n62396 , n62397 , n62398 , 
 n62399 , n62400 , n62401 , n62402 , n62403 , n62404 , n62405 , n62406 , n62407 , n62408 , 
 n62409 , n62410 , n62411 , n62412 , n62413 , n62414 , n62415 , n62416 , n62417 , n62418 , 
 n62419 , n62420 , n62421 , n62422 , n62423 , n62424 , n62425 , n62426 , n62427 , n62428 , 
 n62429 , n62430 , n62431 , n62432 , n62433 , n62434 , n62435 , n62436 , n62437 , n62438 , 
 n62439 , n62440 , n62441 , n62442 , n62443 , n62444 , n62445 , n62446 , n62447 , n62448 , 
 n62449 , n62450 , n62451 , n62452 , n62453 , n62454 , n62455 , n62456 , n62457 , n62458 , 
 n62459 , n62460 , n62461 , n62462 , n62463 , n62464 , n62465 , n62466 , n62467 , n62468 , 
 n62469 , n62470 , n62471 , n62472 , n62473 , n62474 , n62475 , n62476 , n62477 , n62478 , 
 n62479 , n62480 , n62481 , n62482 , n62483 , n62484 , n62485 , n62486 , n62487 , n62488 , 
 n62489 , n62490 , n62491 , n62492 , n62493 , n62494 , n62495 , n62496 , n62497 , n62498 , 
 n62499 , n62500 , n62501 , n62502 , n62503 , n62504 , n62505 , n62506 , n62507 , n62508 , 
 n62509 , n62510 , n62511 , n62512 , n62513 , n62514 , n62515 , n62516 , n62517 , n62518 , 
 n62519 , n62520 , n62521 , n62522 , n62523 , n62524 , n62525 , n62526 , n62527 , n62528 , 
 n62529 , n62530 , n62531 , n62532 , n62533 , n62534 , n62535 , n62536 , n62537 , n62538 , 
 n62539 , n62540 , n62541 , n62542 , n62543 , n62544 , n62545 , n62546 , n62547 , n62548 , 
 n62549 , n62550 , n62551 , n62552 , n62553 , n62554 , n62555 , n62556 , n62557 , n62558 , 
 n62559 , n62560 , n62561 , n62562 , n62563 , n62564 , n62565 , n62566 , n62567 , n62568 , 
 n62569 , n62570 , n62571 , n62572 , n62573 , n62574 , n62575 , n62576 , n62577 , n62578 , 
 n62579 , n62580 , n62581 , n62582 , n62583 , n62584 , n62585 , n62586 , n62587 , n62588 , 
 n62589 , n62590 , n62591 , n62592 , n62593 , n62594 , n62595 , n62596 , n62597 , n62598 , 
 n62599 , n62600 , n62601 , n62602 , n62603 , n62604 , n62605 , n62606 , n62607 , n62608 , 
 n62609 , n62610 , n62611 , n62612 , n62613 , n62614 , n62615 , n62616 , n62617 , n62618 , 
 n62619 , n62620 , n62621 , n62622 , n62623 , n62624 , n62625 , n62626 , n62627 , n62628 , 
 n62629 , n62630 , n62631 , n62632 , n62633 , n62634 , n62635 , n62636 , n62637 , n62638 , 
 n62639 , n62640 , n62641 , n62642 , n62643 , n62644 , n62645 , n62646 , n62647 , n62648 , 
 n62649 , n62650 , n62651 , n62652 , n62653 , n62654 , n62655 , n62656 , n62657 , n62658 , 
 n62659 , n62660 , n62661 , n62662 , n62663 , n62664 , n62665 , n62666 , n62667 , n62668 , 
 n62669 , n62670 , n62671 , n62672 , n62673 , n62674 , n62675 , n62676 , n62677 , n62678 , 
 n62679 , n62680 , n62681 , n62682 , n62683 , n62684 , n62685 , n62686 , n62687 , n62688 , 
 n62689 , n62690 , n62691 , n62692 , n62693 , n62694 , n62695 , n62696 , n62697 , n62698 , 
 n62699 , n62700 , n62701 , n62702 , n62703 , n62704 , n62705 , n62706 , n62707 , n62708 , 
 n62709 , n62710 , n62711 , n62712 , n62713 , n62714 , n62715 , n62716 , n62717 , n62718 , 
 n62719 , n62720 , n62721 , n62722 , n62723 , n62724 , n62725 , n62726 , n62727 , n62728 , 
 n62729 , n62730 , n62731 , n62732 , n62733 , n62734 , n62735 , n62736 , n62737 , n62738 , 
 n62739 , n62740 , n62741 , n62742 , n62743 , n62744 , n62745 , n62746 , n62747 , n62748 , 
 n62749 , n62750 , n62751 , n62752 , n62753 , n62754 , n62755 , n62756 , n62757 , n62758 , 
 n62759 , n62760 , n62761 , n62762 , n62763 , n62764 , n62765 , n62766 , n62767 , n62768 , 
 n62769 , n62770 , n62771 , n62772 , n62773 , n62774 , n62775 , n62776 , n62777 , n62778 , 
 n62779 , n62780 , n62781 , n62782 , n62783 , n62784 , n62785 , n62786 , n62787 , n62788 , 
 n62789 , n62790 , n62791 , n62792 , n62793 , n62794 , n62795 , n62796 , n62797 , n62798 , 
 n62799 , n62800 , n62801 , n62802 , n62803 , n62804 , n62805 , n62806 , n62807 , n62808 , 
 n62809 , n62810 , n62811 , n62812 , n62813 , n62814 , n62815 , n62816 , n62817 , n62818 , 
 n62819 , n62820 , n62821 , n62822 , n62823 , n62824 , n62825 , n62826 , n62827 , n62828 , 
 n62829 , n62830 , n62831 , n62832 , n62833 , n62834 , n62835 , n62836 , n62837 , n62838 , 
 n62839 , n62840 , n62841 , n62842 , n62843 , n62844 , n62845 , n62846 , n62847 , n62848 , 
 n62849 , n62850 , n62851 , n62852 , n62853 , n62854 , n62855 , n62856 , n62857 , n62858 , 
 n62859 , n62860 , n62861 , n62862 , n62863 , n62864 , n62865 , n62866 , n62867 , n62868 , 
 n62869 , n62870 , n62871 , n62872 , n62873 , n62874 , n62875 , n62876 , n62877 , n62878 , 
 n62879 , n62880 , n62881 , n62882 , n62883 , n62884 , n62885 , n62886 , n62887 , n62888 , 
 n62889 , n62890 , n62891 , n62892 , n62893 , n62894 , n62895 , n62896 , n62897 , n62898 , 
 n62899 , n62900 , n62901 , n62902 , n62903 , n62904 , n62905 , n62906 , n62907 , n62908 , 
 n62909 , n62910 , n62911 , n62912 , n62913 , n62914 , n62915 , n62916 , n62917 , n62918 , 
 n62919 , n62920 , n62921 , n62922 , n62923 , n62924 , n62925 , n62926 , n62927 , n62928 , 
 n62929 , n62930 , n62931 , n62932 , n62933 , n62934 , n62935 , n62936 , n62937 , n62938 , 
 n62939 , n62940 , n62941 , n62942 , n62943 , n62944 , n62945 , n62946 , n62947 , n62948 , 
 n62949 , n62950 , n62951 , n62952 , n62953 , n62954 , n62955 , n62956 , n62957 , n62958 , 
 n62959 , n62960 , n62961 , n62962 , n62963 , n62964 , n62965 , n62966 , n62967 , n62968 , 
 n62969 , n62970 , n62971 , n62972 , n62973 , n62974 , n62975 , n62976 , n62977 , n62978 , 
 n62979 , n62980 , n62981 , n62982 , n62983 , n62984 , n62985 , n62986 , n62987 , n62988 , 
 n62989 , n62990 , n62991 , n62992 , n62993 , n62994 , n62995 , n62996 , n62997 , n62998 , 
 n62999 , n63000 , n63001 , n63002 , n63003 , n63004 , n63005 , n63006 , n63007 , n63008 , 
 n63009 , n63010 , n63011 , n63012 , n63013 , n63014 , n63015 , n63016 , n63017 , n63018 , 
 n63019 , n63020 , n63021 , n63022 , n63023 , n63024 , n63025 , n63026 , n63027 , n63028 , 
 n63029 , n63030 , n63031 , n63032 , n63033 , n63034 , n63035 , n63036 , n63037 , n63038 , 
 n63039 , n63040 , n63041 , n63042 , n63043 , n63044 , n63045 , n63046 , n63047 , n63048 , 
 n63049 , n63050 , n63051 , n63052 , n63053 , n63054 , n63055 , n63056 , n63057 , n63058 , 
 n63059 , n63060 , n63061 , n63062 , n63063 , n63064 , n63065 , n63066 , n63067 , n63068 , 
 n63069 , n63070 , n63071 , n63072 , n63073 , n63074 , n63075 , n63076 , n63077 , n63078 , 
 n63079 , n63080 , n63081 , n63082 , n63083 , n63084 , n63085 , n63086 , n63087 , n63088 , 
 n63089 , n63090 , n63091 , n63092 , n63093 , n63094 , n63095 , n63096 , n63097 , n63098 , 
 n63099 , n63100 , n63101 , n63102 , n63103 , n63104 , n63105 , n63106 , n63107 , n63108 , 
 n63109 , n63110 , n63111 , n63112 , n63113 , n63114 , n63115 , n63116 , n63117 , n63118 , 
 n63119 , n63120 , n63121 , n63122 , n63123 , n63124 , n63125 , n63126 , n63127 , n63128 , 
 n63129 , n63130 , n63131 , n63132 , n63133 , n63134 , n63135 , n63136 , n63137 , n63138 , 
 n63139 , n63140 , n63141 , n63142 , n63143 , n63144 , n63145 , n63146 , n63147 , n63148 , 
 n63149 , n63150 , n63151 , n63152 , n63153 , n63154 , n63155 , n63156 , n63157 , n63158 , 
 n63159 , n63160 , n63161 , n63162 , n63163 , n63164 , n63165 , n63166 , n63167 , n63168 , 
 n63169 , n63170 , n63171 , n63172 , n63173 , n63174 , n63175 , n63176 , n63177 , n63178 , 
 n63179 , n63180 , n63181 , n63182 , n63183 , n63184 , n63185 , n63186 , n63187 , n63188 , 
 n63189 , n63190 , n63191 , n63192 , n63193 , n63194 , n63195 , n63196 , n63197 , n63198 , 
 n63199 , n63200 , n63201 , n63202 , n63203 , n63204 , n63205 , n63206 , n63207 , n63208 , 
 n63209 , n63210 , n63211 , n63212 , n63213 , n63214 , n63215 , n63216 , n63217 , n63218 , 
 n63219 , n63220 , n63221 , n63222 , n63223 , n63224 , n63225 , n63226 , n63227 , n63228 , 
 n63229 , n63230 , n63231 , n63232 , n63233 , n63234 , n63235 , n63236 , n63237 , n63238 , 
 n63239 , n63240 , n63241 , n63242 , n63243 , n63244 , n63245 , n63246 , n63247 , n63248 , 
 n63249 , n63250 , n63251 , n63252 , n63253 , n63254 , n63255 , n63256 , n63257 , n63258 , 
 n63259 , n63260 , n63261 , n63262 , n63263 , n63264 , n63265 , n63266 , n63267 , n63268 , 
 n63269 , n63270 , n63271 , n63272 , n63273 , n63274 , n63275 , n63276 , n63277 , n63278 , 
 n63279 , n63280 , n63281 , n63282 , n63283 , n63284 , n63285 , n63286 , n63287 , n63288 , 
 n63289 , n63290 , n63291 , n63292 , n63293 , n63294 , n63295 , n63296 , n63297 , n63298 , 
 n63299 , n63300 , n63301 , n63302 , n63303 , n63304 , n63305 , n63306 , n63307 , n63308 , 
 n63309 , n63310 , n63311 , n63312 , n63313 , n63314 , n63315 , n63316 , n63317 , n63318 , 
 n63319 , n63320 , n63321 , n63322 , n63323 , n63324 , n63325 , n63326 , n63327 , n63328 , 
 n63329 , n63330 , n63331 , n63332 , n63333 , n63334 , n63335 , n63336 , n63337 , n63338 , 
 n63339 , n63340 , n63341 , n63342 , n63343 , n63344 , n63345 , n63346 , n63347 , n63348 , 
 n63349 , n63350 , n63351 , n63352 , n63353 , n63354 , n63355 , n63356 , n63357 , n63358 , 
 n63359 , n63360 , n63361 , n63362 , n63363 , n63364 , n63365 , n63366 , n63367 , n63368 , 
 n63369 , n63370 , n63371 , n63372 , n63373 , n63374 , n63375 , n63376 , n63377 , n63378 , 
 n63379 , n63380 , n63381 , n63382 , n63383 , n63384 , n63385 , n63386 , n63387 , n63388 , 
 n63389 , n63390 , n63391 , n63392 , n63393 , n63394 , n63395 , n63396 , n63397 , n63398 , 
 n63399 , n63400 , n63401 , n63402 , n63403 , n63404 , n63405 , n63406 , n63407 , n63408 , 
 n63409 , n63410 , n63411 , n63412 , n63413 , n63414 , n63415 , n63416 , n63417 , n63418 , 
 n63419 , n63420 , n63421 , n63422 , n63423 , n63424 , n63425 , n63426 , n63427 , n63428 , 
 n63429 , n63430 , n63431 , n63432 , n63433 , n63434 , n63435 , n63436 , n63437 , n63438 , 
 n63439 , n63440 , n63441 , n63442 , n63443 , n63444 , n63445 , n63446 , n63447 , n63448 , 
 n63449 , n63450 , n63451 , n63452 , n63453 , n63454 , n63455 , n63456 , n63457 , n63458 , 
 n63459 , n63460 , n63461 , n63462 , n63463 , n63464 , n63465 , n63466 , n63467 , n63468 , 
 n63469 , n63470 , n63471 , n63472 , n63473 , n63474 , n63475 , n63476 , n63477 , n63478 , 
 n63479 , n63480 , n63481 , n63482 , n63483 , n63484 , n63485 , n63486 , n63487 , n63488 , 
 n63489 , n63490 , n63491 , n63492 , n63493 , n63494 , n63495 , n63496 , n63497 , n63498 , 
 n63499 , n63500 , n63501 , n63502 , n63503 , n63504 , n63505 , n63506 , n63507 , n63508 , 
 n63509 , n63510 , n63511 , n63512 , n63513 , n63514 , n63515 , n63516 , n63517 , n63518 , 
 n63519 , n63520 , n63521 , n63522 , n63523 , n63524 , n63525 , n63526 , n63527 , n63528 , 
 n63529 , n63530 , n63531 , n63532 , n63533 , n63534 , n63535 , n63536 , n63537 , n63538 , 
 n63539 , n63540 , n63541 , n63542 , n63543 , n63544 , n63545 , n63546 , n63547 , n63548 , 
 n63549 , n63550 , n63551 , n63552 , n63553 , n63554 , n63555 , n63556 , n63557 , n63558 , 
 n63559 , n63560 , n63561 , n63562 , n63563 , n63564 , n63565 , n63566 , n63567 , n63568 , 
 n63569 , n63570 , n63571 , n63572 , n63573 , n63574 , n63575 , n63576 , n63577 , n63578 , 
 n63579 , n63580 , n63581 , n63582 , n63583 , n63584 , n63585 , n63586 , n63587 , n63588 , 
 n63589 , n63590 , n63591 , n63592 , n63593 , n63594 , n63595 , n63596 , n63597 , n63598 , 
 n63599 , n63600 , n63601 , n63602 , n63603 , n63604 , n63605 , n63606 , n63607 , n63608 , 
 n63609 , n63610 , n63611 , n63612 , n63613 , n63614 , n63615 , n63616 , n63617 , n63618 , 
 n63619 , n63620 , n63621 , n63622 , n63623 , n63624 , n63625 , n63626 , n63627 , n63628 , 
 n63629 , n63630 , n63631 , n63632 , n63633 , n63634 , n63635 , n63636 , n63637 , n63638 , 
 n63639 , n63640 , n63641 , n63642 , n63643 , n63644 , n63645 , n63646 , n63647 , n63648 , 
 n63649 , n63650 , n63651 , n63652 , n63653 , n63654 , n63655 , n63656 , n63657 , n63658 , 
 n63659 , n63660 , n63661 , n63662 , n63663 , n63664 , n63665 , n63666 , n63667 , n63668 , 
 n63669 , n63670 , n63671 , n63672 , n63673 , n63674 , n63675 , n63676 , n63677 , n63678 , 
 n63679 , n63680 , n63681 , n63682 , n63683 , n63684 , n63685 , n63686 , n63687 , n63688 , 
 n63689 , n63690 , n63691 , n63692 , n63693 , n63694 , n63695 , n63696 , n63697 , n63698 , 
 n63699 , n63700 , n63701 , n63702 , n63703 , n63704 , n63705 , n63706 , n63707 , n63708 , 
 n63709 , n63710 , n63711 , n63712 , n63713 , n63714 , n63715 , n63716 , n63717 , n63718 , 
 n63719 , n63720 , n63721 , n63722 , n63723 , n63724 , n63725 , n63726 , n63727 , n63728 , 
 n63729 , n63730 , n63731 , n63732 , n63733 , n63734 , n63735 , n63736 , n63737 , n63738 , 
 n63739 , n63740 , n63741 , n63742 , n63743 , n63744 , n63745 , n63746 , n63747 , n63748 , 
 n63749 , n63750 , n63751 , n63752 , n63753 , n63754 , n63755 , n63756 , n63757 , n63758 , 
 n63759 , n63760 , n63761 , n63762 , n63763 , n63764 , n63765 , n63766 , n63767 , n63768 , 
 n63769 , n63770 , n63771 , n63772 , n63773 , n63774 , n63775 , n63776 , n63777 , n63778 , 
 n63779 , n63780 , n63781 , n63782 , n63783 , n63784 , n63785 , n63786 , n63787 , n63788 , 
 n63789 , n63790 , n63791 , n63792 , n63793 , n63794 , n63795 , n63796 , n63797 , n63798 , 
 n63799 , n63800 , n63801 , n63802 , n63803 , n63804 , n63805 , n63806 , n63807 , n63808 , 
 n63809 , n63810 , n63811 , n63812 , n63813 , n63814 , n63815 , n63816 , n63817 , n63818 , 
 n63819 , n63820 , n63821 , n63822 , n63823 , n63824 , n63825 , n63826 , n63827 , n63828 , 
 n63829 , n63830 , n63831 , n63832 , n63833 , n63834 , n63835 , n63836 , n63837 , n63838 , 
 n63839 , n63840 , n63841 , n63842 , n63843 , n63844 , n63845 , n63846 , n63847 , n63848 , 
 n63849 , n63850 , n63851 , n63852 , n63853 , n63854 , n63855 , n63856 , n63857 , n63858 , 
 n63859 , n63860 , n63861 , n63862 , n63863 , n63864 , n63865 , n63866 , n63867 , n63868 , 
 n63869 , n63870 , n63871 , n63872 , n63873 , n63874 , n63875 , n63876 , n63877 , n63878 , 
 n63879 , n63880 , n63881 , n63882 , n63883 , n63884 , n63885 , n63886 , n63887 , n63888 , 
 n63889 , n63890 , n63891 , n63892 , n63893 , n63894 , n63895 , n63896 , n63897 , n63898 , 
 n63899 , n63900 , n63901 , n63902 , n63903 , n63904 , n63905 , n63906 , n63907 , n63908 , 
 n63909 , n63910 , n63911 , n63912 , n63913 , n63914 , n63915 , n63916 , n63917 , n63918 , 
 n63919 , n63920 , n63921 , n63922 , n63923 , n63924 , n63925 , n63926 , n63927 , n63928 , 
 n63929 , n63930 , n63931 , n63932 , n63933 , n63934 , n63935 , n63936 , n63937 , n63938 , 
 n63939 , n63940 , n63941 , n63942 , n63943 , n63944 , n63945 , n63946 , n63947 , n63948 , 
 n63949 , n63950 , n63951 , n63952 , n63953 , n63954 , n63955 , n63956 , n63957 , n63958 , 
 n63959 , n63960 , n63961 , n63962 , n63963 , n63964 , n63965 , n63966 , n63967 , n63968 , 
 n63969 , n63970 , n63971 , n63972 , n63973 , n63974 , n63975 , n63976 , n63977 , n63978 , 
 n63979 , n63980 , n63981 , n63982 , n63983 , n63984 , n63985 , n63986 , n63987 , n63988 , 
 n63989 , n63990 , n63991 , n63992 , n63993 , n63994 , n63995 , n63996 , n63997 , n63998 , 
 n63999 , n64000 , n64001 , n64002 , n64003 , n64004 , n64005 , n64006 , n64007 , n64008 , 
 n64009 , n64010 , n64011 , n64012 , n64013 , n64014 , n64015 , n64016 , n64017 , n64018 , 
 n64019 , n64020 , n64021 , n64022 , n64023 , n64024 , n64025 , n64026 , n64027 , n64028 , 
 n64029 , n64030 , n64031 , n64032 , n64033 , n64034 , n64035 , n64036 , n64037 , n64038 , 
 n64039 , n64040 , n64041 , n64042 , n64043 , n64044 , n64045 , n64046 , n64047 , n64048 , 
 n64049 , n64050 , n64051 , n64052 , n64053 , n64054 , n64055 , n64056 , n64057 , n64058 , 
 n64059 , n64060 , n64061 , n64062 , n64063 , n64064 , n64065 , n64066 , n64067 , n64068 , 
 n64069 , n64070 , n64071 , n64072 , n64073 , n64074 , n64075 , n64076 , n64077 , n64078 , 
 n64079 , n64080 , n64081 , n64082 , n64083 , n64084 , n64085 , n64086 , n64087 , n64088 , 
 n64089 , n64090 , n64091 , n64092 , n64093 , n64094 , n64095 , n64096 , n64097 , n64098 , 
 n64099 , n64100 , n64101 , n64102 , n64103 , n64104 , n64105 , n64106 , n64107 , n64108 , 
 n64109 , n64110 , n64111 , n64112 , n64113 , n64114 , n64115 , n64116 , n64117 , n64118 , 
 n64119 , n64120 , n64121 , n64122 , n64123 , n64124 , n64125 , n64126 , n64127 , n64128 , 
 n64129 , n64130 , n64131 , n64132 , n64133 , n64134 , n64135 , n64136 , n64137 , n64138 , 
 n64139 , n64140 , n64141 , n64142 , n64143 , n64144 , n64145 , n64146 , n64147 , n64148 , 
 n64149 , n64150 , n64151 , n64152 , n64153 , n64154 , n64155 , n64156 , n64157 , n64158 , 
 n64159 , n64160 , n64161 , n64162 , n64163 , n64164 , n64165 , n64166 , n64167 , n64168 , 
 n64169 , n64170 , n64171 , n64172 , n64173 , n64174 , n64175 , n64176 , n64177 , n64178 , 
 n64179 , n64180 , n64181 , n64182 , n64183 , n64184 , n64185 , n64186 , n64187 , n64188 , 
 n64189 , n64190 , n64191 , n64192 , n64193 , n64194 , n64195 , n64196 , n64197 , n64198 , 
 n64199 , n64200 , n64201 , n64202 , n64203 , n64204 , n64205 , n64206 , n64207 , n64208 , 
 n64209 , n64210 , n64211 , n64212 , n64213 , n64214 , n64215 , n64216 , n64217 , n64218 , 
 n64219 , n64220 , n64221 , n64222 , n64223 , n64224 , n64225 , n64226 , n64227 , n64228 , 
 n64229 , n64230 , n64231 , n64232 , n64233 , n64234 , n64235 , n64236 , n64237 , n64238 , 
 n64239 , n64240 , n64241 , n64242 , n64243 , n64244 , n64245 , n64246 , n64247 , n64248 , 
 n64249 , n64250 , n64251 , n64252 , n64253 , n64254 , n64255 , n64256 , n64257 , n64258 , 
 n64259 , n64260 , n64261 , n64262 , n64263 , n64264 , n64265 , n64266 , n64267 , n64268 , 
 n64269 , n64270 , n64271 , n64272 , n64273 , n64274 , n64275 , n64276 , n64277 , n64278 , 
 n64279 , n64280 , n64281 , n64282 , n64283 , n64284 , n64285 , n64286 , n64287 , n64288 , 
 n64289 , n64290 , n64291 , n64292 , n64293 , n64294 , n64295 , n64296 , n64297 , n64298 , 
 n64299 , n64300 , n64301 , n64302 , n64303 , n64304 , n64305 , n64306 , n64307 , n64308 , 
 n64309 , n64310 , n64311 , n64312 , n64313 , n64314 , n64315 , n64316 , n64317 , n64318 , 
 n64319 , n64320 , n64321 , n64322 , n64323 , n64324 , n64325 , n64326 , n64327 , n64328 , 
 n64329 , n64330 , n64331 , n64332 , n64333 , n64334 , n64335 , n64336 , n64337 , n64338 , 
 n64339 , n64340 , n64341 , n64342 , n64343 , n64344 , n64345 , n64346 , n64347 , n64348 , 
 n64349 , n64350 , n64351 , n64352 , n64353 , n64354 , n64355 , n64356 , n64357 , n64358 , 
 n64359 , n64360 , n64361 , n64362 , n64363 , n64364 , n64365 , n64366 , n64367 , n64368 , 
 n64369 , n64370 , n64371 , n64372 , n64373 , n64374 , n64375 , n64376 , n64377 , n64378 , 
 n64379 , n64380 , n64381 , n64382 , n64383 , n64384 , n64385 , n64386 , n64387 , n64388 , 
 n64389 , n64390 , n64391 , n64392 , n64393 , n64394 , n64395 , n64396 , n64397 , n64398 , 
 n64399 , n64400 , n64401 , n64402 , n64403 , n64404 , n64405 , n64406 , n64407 , n64408 , 
 n64409 , n64410 , n64411 , n64412 , n64413 , n64414 , n64415 , n64416 , n64417 , n64418 , 
 n64419 , n64420 , n64421 , n64422 , n64423 , n64424 , n64425 , n64426 , n64427 , n64428 , 
 n64429 , n64430 , n64431 , n64432 , n64433 , n64434 , n64435 , n64436 , n64437 , n64438 , 
 n64439 , n64440 , n64441 , n64442 , n64443 , n64444 , n64445 , n64446 , n64447 , n64448 , 
 n64449 , n64450 , n64451 , n64452 , n64453 , n64454 , n64455 , n64456 , n64457 , n64458 , 
 n64459 , n64460 , n64461 , n64462 , n64463 , n64464 , n64465 , n64466 , n64467 , n64468 , 
 n64469 , n64470 , n64471 , n64472 , n64473 , n64474 , n64475 , n64476 , n64477 , n64478 , 
 n64479 , n64480 , n64481 , n64482 , n64483 , n64484 , n64485 , n64486 , n64487 , n64488 , 
 n64489 , n64490 , n64491 , n64492 , n64493 , n64494 , n64495 , n64496 , n64497 , n64498 , 
 n64499 , n64500 , n64501 , n64502 , n64503 , n64504 , n64505 , n64506 , n64507 , n64508 , 
 n64509 , n64510 , n64511 , n64512 , n64513 , n64514 , n64515 , n64516 , n64517 , n64518 , 
 n64519 , n64520 , n64521 , n64522 , n64523 , n64524 , n64525 , n64526 , n64527 , n64528 , 
 n64529 , n64530 , n64531 , n64532 , n64533 , n64534 , n64535 , n64536 , n64537 , n64538 , 
 n64539 , n64540 , n64541 , n64542 , n64543 , n64544 , n64545 , n64546 , n64547 , n64548 , 
 n64549 , n64550 , n64551 , n64552 , n64553 , n64554 , n64555 , n64556 , n64557 , n64558 , 
 n64559 , n64560 , n64561 , n64562 , n64563 , n64564 , n64565 , n64566 , n64567 , n64568 , 
 n64569 , n64570 , n64571 , n64572 , n64573 , n64574 , n64575 , n64576 , n64577 , n64578 , 
 n64579 , n64580 , n64581 , n64582 , n64583 , n64584 , n64585 , n64586 , n64587 , n64588 , 
 n64589 , n64590 , n64591 , n64592 , n64593 , n64594 , n64595 , n64596 , n64597 , n64598 , 
 n64599 , n64600 , n64601 , n64602 , n64603 , n64604 , n64605 , n64606 , n64607 , n64608 , 
 n64609 , n64610 , n64611 , n64612 , n64613 , n64614 , n64615 , n64616 , n64617 , n64618 , 
 n64619 , n64620 , n64621 , n64622 , n64623 , n64624 , n64625 , n64626 , n64627 , n64628 , 
 n64629 , n64630 , n64631 , n64632 , n64633 , n64634 , n64635 , n64636 , n64637 , n64638 , 
 n64639 , n64640 , n64641 , n64642 , n64643 , n64644 , n64645 , n64646 , n64647 , n64648 , 
 n64649 , n64650 , n64651 , n64652 , n64653 , n64654 , n64655 , n64656 , n64657 , n64658 , 
 n64659 , n64660 , n64661 , n64662 , n64663 , n64664 , n64665 , n64666 , n64667 , n64668 , 
 n64669 , n64670 , n64671 , n64672 , n64673 , n64674 , n64675 , n64676 , n64677 , n64678 , 
 n64679 , n64680 , n64681 , n64682 , n64683 , n64684 , n64685 , n64686 , n64687 , n64688 , 
 n64689 , n64690 , n64691 , n64692 , n64693 , n64694 , n64695 , n64696 , n64697 , n64698 , 
 n64699 , n64700 , n64701 , n64702 , n64703 , n64704 , n64705 , n64706 , n64707 , n64708 , 
 n64709 , n64710 , n64711 , n64712 , n64713 , n64714 , n64715 , n64716 , n64717 , n64718 , 
 n64719 , n64720 , n64721 , n64722 , n64723 , n64724 , n64725 , n64726 , n64727 , n64728 , 
 n64729 , n64730 , n64731 , n64732 , n64733 , n64734 , n64735 , n64736 , n64737 , n64738 , 
 n64739 , n64740 , n64741 , n64742 , n64743 , n64744 , n64745 , n64746 , n64747 , n64748 , 
 n64749 , n64750 , n64751 , n64752 , n64753 , n64754 , n64755 , n64756 , n64757 , n64758 , 
 n64759 , n64760 , n64761 , n64762 , n64763 , n64764 , n64765 , n64766 , n64767 , n64768 , 
 n64769 , n64770 , n64771 , n64772 , n64773 , n64774 , n64775 , n64776 , n64777 , n64778 , 
 n64779 , n64780 , n64781 , n64782 , n64783 , n64784 , n64785 , n64786 , n64787 , n64788 , 
 n64789 , n64790 , n64791 , n64792 , n64793 , n64794 , n64795 , n64796 , n64797 , n64798 , 
 n64799 , n64800 , n64801 , n64802 , n64803 , n64804 , n64805 , n64806 , n64807 , n64808 , 
 n64809 , n64810 , n64811 , n64812 , n64813 , n64814 , n64815 , n64816 , n64817 , n64818 , 
 n64819 , n64820 , n64821 , n64822 , n64823 , n64824 , n64825 , n64826 , n64827 , n64828 , 
 n64829 , n64830 , n64831 , n64832 , n64833 , n64834 , n64835 , n64836 , n64837 , n64838 , 
 n64839 , n64840 , n64841 , n64842 , n64843 , n64844 , n64845 , n64846 , n64847 , n64848 , 
 n64849 , n64850 , n64851 , n64852 , n64853 , n64854 , n64855 , n64856 , n64857 , n64858 , 
 n64859 , n64860 , n64861 , n64862 , n64863 , n64864 , n64865 , n64866 , n64867 , n64868 , 
 n64869 , n64870 , n64871 , n64872 , n64873 , n64874 , n64875 , n64876 , n64877 , n64878 , 
 n64879 , n64880 , n64881 , n64882 , n64883 , n64884 , n64885 , n64886 , n64887 , n64888 , 
 n64889 , n64890 , n64891 , n64892 , n64893 , n64894 , n64895 , n64896 , n64897 , n64898 , 
 n64899 , n64900 , n64901 , n64902 , n64903 , n64904 , n64905 , n64906 , n64907 , n64908 , 
 n64909 , n64910 , n64911 , n64912 , n64913 , n64914 , n64915 , n64916 , n64917 , n64918 , 
 n64919 , n64920 , n64921 , n64922 , n64923 , n64924 , n64925 , n64926 , n64927 , n64928 , 
 n64929 , n64930 , n64931 , n64932 , n64933 , n64934 , n64935 , n64936 , n64937 , n64938 , 
 n64939 , n64940 , n64941 , n64942 , n64943 , n64944 , n64945 , n64946 , n64947 , n64948 , 
 n64949 , n64950 , n64951 , n64952 , n64953 , n64954 , n64955 , n64956 , n64957 , n64958 , 
 n64959 , n64960 , n64961 , n64962 , n64963 , n64964 , n64965 , n64966 , n64967 , n64968 , 
 n64969 , n64970 , n64971 , n64972 , n64973 , n64974 , n64975 , n64976 , n64977 , n64978 , 
 n64979 , n64980 , n64981 , n64982 , n64983 , n64984 , n64985 , n64986 , n64987 , n64988 , 
 n64989 , n64990 , n64991 , n64992 , n64993 , n64994 , n64995 , n64996 , n64997 , n64998 , 
 n64999 , n65000 , n65001 , n65002 , n65003 , n65004 , n65005 , n65006 , n65007 , n65008 , 
 n65009 , n65010 , n65011 , n65012 , n65013 , n65014 , n65015 , n65016 , n65017 , n65018 , 
 n65019 , n65020 , n65021 , n65022 , n65023 , n65024 , n65025 , n65026 , n65027 , n65028 , 
 n65029 , n65030 , n65031 , n65032 , n65033 , n65034 , n65035 , n65036 , n65037 , n65038 , 
 n65039 , n65040 , n65041 , n65042 , n65043 , n65044 , n65045 , n65046 , n65047 , n65048 , 
 n65049 , n65050 , n65051 , n65052 , n65053 , n65054 , n65055 , n65056 , n65057 , n65058 , 
 n65059 , n65060 , n65061 , n65062 , n65063 , n65064 , n65065 , n65066 , n65067 , n65068 , 
 n65069 , n65070 , n65071 , n65072 , n65073 , n65074 , n65075 , n65076 , n65077 , n65078 , 
 n65079 , n65080 , n65081 , n65082 , n65083 , n65084 , n65085 , n65086 , n65087 , n65088 , 
 n65089 , n65090 , n65091 , n65092 , n65093 , n65094 , n65095 , n65096 , n65097 , n65098 , 
 n65099 , n65100 , n65101 , n65102 , n65103 , n65104 , n65105 , n65106 , n65107 , n65108 , 
 n65109 , n65110 , n65111 , n65112 , n65113 , n65114 , n65115 , n65116 , n65117 , n65118 , 
 n65119 , n65120 , n65121 , n65122 , n65123 , n65124 , n65125 , n65126 , n65127 , n65128 , 
 n65129 , n65130 , n65131 , n65132 , n65133 , n65134 , n65135 , n65136 , n65137 , n65138 , 
 n65139 , n65140 , n65141 , n65142 , n65143 , n65144 , n65145 , n65146 , n65147 , n65148 , 
 n65149 , n65150 , n65151 , n65152 , n65153 , n65154 , n65155 , n65156 , n65157 , n65158 , 
 n65159 , n65160 , n65161 , n65162 , n65163 , n65164 , n65165 , n65166 , n65167 , n65168 , 
 n65169 , n65170 , n65171 , n65172 , n65173 , n65174 , n65175 , n65176 , n65177 , n65178 , 
 n65179 , n65180 , n65181 , n65182 , n65183 , n65184 , n65185 , n65186 , n65187 , n65188 , 
 n65189 , n65190 , n65191 , n65192 , n65193 , n65194 , n65195 , n65196 , n65197 , n65198 , 
 n65199 , n65200 , n65201 , n65202 , n65203 , n65204 , n65205 , n65206 , n65207 , n65208 , 
 n65209 , n65210 , n65211 , n65212 , n65213 , n65214 , n65215 , n65216 , n65217 , n65218 , 
 n65219 , n65220 , n65221 , n65222 , n65223 , n65224 , n65225 , n65226 , n65227 , n65228 , 
 n65229 , n65230 , n65231 , n65232 , n65233 , n65234 , n65235 , n65236 , n65237 , n65238 , 
 n65239 , n65240 , n65241 , n65242 , n65243 , n65244 , n65245 , n65246 , n65247 , n65248 , 
 n65249 , n65250 , n65251 , n65252 , n65253 , n65254 , n65255 , n65256 , n65257 , n65258 , 
 n65259 , n65260 , n65261 , n65262 , n65263 , n65264 , n65265 , n65266 , n65267 , n65268 , 
 n65269 , n65270 , n65271 , n65272 , n65273 , n65274 , n65275 , n65276 , n65277 , n65278 , 
 n65279 , n65280 , n65281 , n65282 , n65283 , n65284 , n65285 , n65286 , n65287 , n65288 , 
 n65289 , n65290 , n65291 , n65292 , n65293 , n65294 , n65295 , n65296 , n65297 , n65298 , 
 n65299 , n65300 , n65301 , n65302 , n65303 , n65304 , n65305 , n65306 , n65307 , n65308 , 
 n65309 , n65310 , n65311 , n65312 , n65313 , n65314 , n65315 , n65316 , n65317 , n65318 , 
 n65319 , n65320 , n65321 , n65322 , n65323 , n65324 , n65325 , n65326 , n65327 , n65328 , 
 n65329 , n65330 , n65331 , n65332 , n65333 , n65334 , n65335 , n65336 , n65337 , n65338 , 
 n65339 , n65340 , n65341 , n65342 , n65343 , n65344 , n65345 , n65346 , n65347 , n65348 , 
 n65349 , n65350 , n65351 , n65352 , n65353 , n65354 , n65355 , n65356 , n65357 , n65358 , 
 n65359 , n65360 , n65361 , n65362 , n65363 , n65364 , n65365 , n65366 , n65367 , n65368 , 
 n65369 , n65370 , n65371 , n65372 , n65373 , n65374 , n65375 , n65376 , n65377 , n65378 , 
 n65379 , n65380 , n65381 , n65382 , n65383 , n65384 , n65385 , n65386 , n65387 , n65388 , 
 n65389 , n65390 , n65391 , n65392 , n65393 , n65394 , n65395 , n65396 , n65397 , n65398 , 
 n65399 , n65400 , n65401 , n65402 , n65403 , n65404 , n65405 , n65406 , n65407 , n65408 , 
 n65409 , n65410 , n65411 , n65412 , n65413 , n65414 , n65415 , n65416 , n65417 , n65418 , 
 n65419 , n65420 , n65421 , n65422 , n65423 , n65424 , n65425 , n65426 , n65427 , n65428 , 
 n65429 , n65430 , n65431 , n65432 , n65433 , n65434 , n65435 , n65436 , n65437 , n65438 , 
 n65439 , n65440 , n65441 , n65442 , n65443 , n65444 , n65445 , n65446 , n65447 , n65448 , 
 n65449 , n65450 , n65451 , n65452 , n65453 , n65454 , n65455 , n65456 , n65457 , n65458 , 
 n65459 , n65460 , n65461 , n65462 , n65463 , n65464 , n65465 , n65466 , n65467 , n65468 , 
 n65469 , n65470 , n65471 , n65472 , n65473 , n65474 , n65475 , n65476 , n65477 , n65478 , 
 n65479 , n65480 , n65481 , n65482 , n65483 , n65484 , n65485 , n65486 , n65487 , n65488 , 
 n65489 , n65490 , n65491 , n65492 , n65493 , n65494 , n65495 , n65496 , n65497 , n65498 , 
 n65499 , n65500 , n65501 , n65502 , n65503 , n65504 , n65505 , n65506 , n65507 , n65508 , 
 n65509 , n65510 , n65511 , n65512 , n65513 , n65514 , n65515 , n65516 , n65517 , n65518 , 
 n65519 , n65520 , n65521 , n65522 , n65523 , n65524 , n65525 , n65526 , n65527 , n65528 , 
 n65529 , n65530 , n65531 , n65532 , n65533 , n65534 , n65535 , n65536 , n65537 , n65538 , 
 n65539 , n65540 , n65541 , n65542 , n65543 , n65544 , n65545 , n65546 , n65547 , n65548 , 
 n65549 , n65550 , n65551 , n65552 , n65553 , n65554 , n65555 , n65556 , n65557 , n65558 , 
 n65559 , n65560 , n65561 , n65562 , n65563 , n65564 , n65565 , n65566 , n65567 , n65568 , 
 n65569 , n65570 , n65571 , n65572 , n65573 , n65574 , n65575 , n65576 , n65577 , n65578 , 
 n65579 , n65580 , n65581 , n65582 , n65583 , n65584 , n65585 , n65586 , n65587 , n65588 , 
 n65589 , n65590 , n65591 , n65592 , n65593 , n65594 , n65595 , n65596 , n65597 , n65598 , 
 n65599 , n65600 , n65601 , n65602 , n65603 , n65604 , n65605 , n65606 , n65607 , n65608 , 
 n65609 , n65610 , n65611 , n65612 , n65613 , n65614 , n65615 , n65616 , n65617 , n65618 , 
 n65619 , n65620 , n65621 , n65622 , n65623 , n65624 , n65625 , n65626 , n65627 , n65628 , 
 n65629 , n65630 , n65631 , n65632 , n65633 , n65634 , n65635 , n65636 , n65637 , n65638 , 
 n65639 , n65640 , n65641 , n65642 , n65643 , n65644 , n65645 , n65646 , n65647 , n65648 , 
 n65649 , n65650 , n65651 , n65652 , n65653 , n65654 , n65655 , n65656 , n65657 , n65658 , 
 n65659 , n65660 , n65661 , n65662 , n65663 , n65664 , n65665 , n65666 , n65667 , n65668 , 
 n65669 , n65670 , n65671 , n65672 , n65673 , n65674 , n65675 , n65676 , n65677 , n65678 , 
 n65679 , n65680 , n65681 , n65682 , n65683 , n65684 , n65685 , n65686 , n65687 , n65688 , 
 n65689 , n65690 , n65691 , n65692 , n65693 , n65694 , n65695 , n65696 , n65697 , n65698 , 
 n65699 , n65700 , n65701 , n65702 , n65703 , n65704 , n65705 , n65706 , n65707 , n65708 , 
 n65709 , n65710 , n65711 , n65712 , n65713 , n65714 , n65715 , n65716 , n65717 , n65718 , 
 n65719 , n65720 , n65721 , n65722 , n65723 , n65724 , n65725 , n65726 , n65727 , n65728 , 
 n65729 , n65730 , n65731 , n65732 , n65733 , n65734 , n65735 , n65736 , n65737 , n65738 , 
 n65739 , n65740 , n65741 , n65742 , n65743 , n65744 , n65745 , n65746 , n65747 , n65748 , 
 n65749 , n65750 , n65751 , n65752 , n65753 , n65754 , n65755 , n65756 , n65757 , n65758 , 
 n65759 , n65760 , n65761 , n65762 , n65763 , n65764 , n65765 , n65766 , n65767 , n65768 , 
 n65769 , n65770 , n65771 , n65772 , n65773 , n65774 , n65775 , n65776 , n65777 , n65778 , 
 n65779 , n65780 , n65781 , n65782 , n65783 , n65784 , n65785 , n65786 , n65787 , n65788 , 
 n65789 , n65790 , n65791 , n65792 , n65793 , n65794 , n65795 , n65796 , n65797 , n65798 , 
 n65799 , n65800 , n65801 , n65802 , n65803 , n65804 , n65805 , n65806 , n65807 , n65808 , 
 n65809 , n65810 , n65811 , n65812 , n65813 , n65814 , n65815 , n65816 , n65817 , n65818 , 
 n65819 , n65820 , n65821 , n65822 , n65823 , n65824 , n65825 , n65826 , n65827 , n65828 , 
 n65829 , n65830 , n65831 , n65832 , n65833 , n65834 , n65835 , n65836 , n65837 , n65838 , 
 n65839 , n65840 , n65841 , n65842 , n65843 , n65844 , n65845 , n65846 , n65847 , n65848 , 
 n65849 , n65850 , n65851 , n65852 , n65853 , n65854 , n65855 , n65856 , n65857 , n65858 , 
 n65859 , n65860 , n65861 , n65862 , n65863 , n65864 , n65865 , n65866 , n65867 , n65868 , 
 n65869 , n65870 , n65871 , n65872 , n65873 , n65874 , n65875 , n65876 , n65877 , n65878 , 
 n65879 , n65880 , n65881 , n65882 , n65883 , n65884 , n65885 , n65886 , n65887 , n65888 , 
 n65889 , n65890 , n65891 , n65892 , n65893 , n65894 , n65895 , n65896 , n65897 , n65898 , 
 n65899 , n65900 , n65901 , n65902 , n65903 , n65904 , n65905 , n65906 , n65907 , n65908 , 
 n65909 , n65910 , n65911 , n65912 , n65913 , n65914 , n65915 , n65916 , n65917 , n65918 , 
 n65919 , n65920 , n65921 , n65922 , n65923 , n65924 , n65925 , n65926 , n65927 , n65928 , 
 n65929 , n65930 , n65931 , n65932 , n65933 , n65934 , n65935 , n65936 , n65937 , n65938 , 
 n65939 , n65940 , n65941 , n65942 , n65943 , n65944 , n65945 , n65946 , n65947 , n65948 , 
 n65949 , n65950 , n65951 , n65952 , n65953 , n65954 , n65955 , n65956 , n65957 , n65958 , 
 n65959 , n65960 , n65961 , n65962 , n65963 , n65964 , n65965 , n65966 , n65967 , n65968 , 
 n65969 , n65970 , n65971 , n65972 , n65973 , n65974 , n65975 , n65976 , n65977 , n65978 , 
 n65979 , n65980 , n65981 , n65982 , n65983 , n65984 , n65985 , n65986 , n65987 , n65988 , 
 n65989 , n65990 , n65991 , n65992 , n65993 , n65994 , n65995 , n65996 , n65997 , n65998 , 
 n65999 , n66000 , n66001 , n66002 , n66003 , n66004 , n66005 , n66006 , n66007 , n66008 , 
 n66009 , n66010 , n66011 , n66012 , n66013 , n66014 , n66015 , n66016 , n66017 , n66018 , 
 n66019 , n66020 , n66021 , n66022 , n66023 , n66024 , n66025 , n66026 , n66027 , n66028 , 
 n66029 , n66030 , n66031 , n66032 , n66033 , n66034 , n66035 , n66036 , n66037 , n66038 , 
 n66039 , n66040 , n66041 , n66042 , n66043 , n66044 , n66045 , n66046 , n66047 , n66048 , 
 n66049 , n66050 , n66051 , n66052 , n66053 , n66054 , n66055 , n66056 , n66057 , n66058 , 
 n66059 , n66060 , n66061 , n66062 , n66063 , n66064 , n66065 , n66066 , n66067 , n66068 , 
 n66069 , n66070 , n66071 , n66072 , n66073 , n66074 , n66075 , n66076 , n66077 , n66078 , 
 n66079 , n66080 , n66081 , n66082 , n66083 , n66084 , n66085 , n66086 , n66087 , n66088 , 
 n66089 , n66090 , n66091 , n66092 , n66093 , n66094 , n66095 , n66096 , n66097 , n66098 , 
 n66099 , n66100 , n66101 , n66102 , n66103 , n66104 , n66105 , n66106 , n66107 , n66108 , 
 n66109 , n66110 , n66111 , n66112 , n66113 , n66114 , n66115 , n66116 , n66117 , n66118 , 
 n66119 , n66120 , n66121 , n66122 , n66123 , n66124 , n66125 , n66126 , n66127 , n66128 , 
 n66129 , n66130 , n66131 , n66132 , n66133 , n66134 , n66135 , n66136 , n66137 , n66138 , 
 n66139 , n66140 , n66141 , n66142 , n66143 , n66144 , n66145 , n66146 , n66147 , n66148 , 
 n66149 , n66150 , n66151 , n66152 , n66153 , n66154 , n66155 , n66156 , n66157 , n66158 , 
 n66159 , n66160 , n66161 , n66162 , n66163 , n66164 , n66165 , n66166 , n66167 , n66168 , 
 n66169 , n66170 , n66171 , n66172 , n66173 , n66174 , n66175 , n66176 , n66177 , n66178 , 
 n66179 , n66180 , n66181 , n66182 , n66183 , n66184 , n66185 , n66186 , n66187 , n66188 , 
 n66189 , n66190 , n66191 , n66192 , n66193 , n66194 , n66195 , n66196 , n66197 , n66198 , 
 n66199 , n66200 , n66201 , n66202 , n66203 , n66204 , n66205 , n66206 , n66207 , n66208 , 
 n66209 , n66210 , n66211 , n66212 , n66213 , n66214 , n66215 , n66216 , n66217 , n66218 , 
 n66219 , n66220 , n66221 , n66222 , n66223 , n66224 , n66225 , n66226 , n66227 , n66228 , 
 n66229 , n66230 , n66231 , n66232 , n66233 , n66234 , n66235 , n66236 , n66237 , n66238 , 
 n66239 , n66240 , n66241 , n66242 , n66243 , n66244 , n66245 , n66246 , n66247 , n66248 , 
 n66249 , n66250 , n66251 , n66252 , n66253 , n66254 , n66255 , n66256 , n66257 , n66258 , 
 n66259 , n66260 , n66261 , n66262 , n66263 , n66264 , n66265 , n66266 , n66267 , n66268 , 
 n66269 , n66270 , n66271 , n66272 , n66273 , n66274 , n66275 , n66276 , n66277 , n66278 , 
 n66279 , n66280 , n66281 , n66282 , n66283 , n66284 , n66285 , n66286 , n66287 , n66288 , 
 n66289 , n66290 , n66291 , n66292 , n66293 , n66294 , n66295 , n66296 , n66297 , n66298 , 
 n66299 , n66300 , n66301 , n66302 , n66303 , n66304 , n66305 , n66306 , n66307 , n66308 , 
 n66309 , n66310 , n66311 , n66312 , n66313 , n66314 , n66315 , n66316 , n66317 , n66318 , 
 n66319 , n66320 , n66321 , n66322 , n66323 , n66324 , n66325 , n66326 , n66327 , n66328 , 
 n66329 , n66330 , n66331 , n66332 , n66333 , n66334 , n66335 , n66336 , n66337 , n66338 , 
 n66339 , n66340 , n66341 , n66342 , n66343 , n66344 , n66345 , n66346 , n66347 , n66348 , 
 n66349 , n66350 , n66351 , n66352 , n66353 , n66354 , n66355 , n66356 , n66357 , n66358 , 
 n66359 , n66360 , n66361 , n66362 , n66363 , n66364 , n66365 , n66366 , n66367 , n66368 , 
 n66369 , n66370 , n66371 , n66372 , n66373 , n66374 , n66375 , n66376 , n66377 , n66378 , 
 n66379 , n66380 , n66381 , n66382 , n66383 , n66384 , n66385 , n66386 , n66387 , n66388 , 
 n66389 , n66390 , n66391 , n66392 , n66393 , n66394 , n66395 , n66396 , n66397 , n66398 , 
 n66399 , n66400 , n66401 , n66402 , n66403 , n66404 , n66405 , n66406 , n66407 , n66408 , 
 n66409 , n66410 , n66411 , n66412 , n66413 , n66414 , n66415 , n66416 , n66417 , n66418 , 
 n66419 , n66420 , n66421 , n66422 , n66423 , n66424 , n66425 , n66426 , n66427 , n66428 , 
 n66429 , n66430 , n66431 , n66432 , n66433 , n66434 , n66435 , n66436 , n66437 , n66438 , 
 n66439 , n66440 , n66441 , n66442 , n66443 , n66444 , n66445 , n66446 , n66447 , n66448 , 
 n66449 , n66450 , n66451 , n66452 , n66453 , n66454 , n66455 , n66456 , n66457 , n66458 , 
 n66459 , n66460 , n66461 , n66462 , n66463 , n66464 , n66465 , n66466 , n66467 , n66468 , 
 n66469 , n66470 , n66471 , n66472 , n66473 , n66474 , n66475 , n66476 , n66477 , n66478 , 
 n66479 , n66480 , n66481 , n66482 , n66483 , n66484 , n66485 , n66486 , n66487 , n66488 , 
 n66489 , n66490 , n66491 , n66492 , n66493 , n66494 , n66495 , n66496 , n66497 , n66498 , 
 n66499 , n66500 , n66501 , n66502 , n66503 , n66504 , n66505 , n66506 , n66507 , n66508 , 
 n66509 , n66510 , n66511 , n66512 , n66513 , n66514 , n66515 , n66516 , n66517 , n66518 , 
 n66519 , n66520 , n66521 , n66522 , n66523 , n66524 , n66525 , n66526 , n66527 , n66528 , 
 n66529 , n66530 , n66531 , n66532 , n66533 , n66534 , n66535 , n66536 , n66537 , n66538 , 
 n66539 , n66540 , n66541 , n66542 , n66543 , n66544 , n66545 , n66546 , n66547 , n66548 , 
 n66549 , n66550 , n66551 , n66552 , n66553 , n66554 , n66555 , n66556 , n66557 , n66558 , 
 n66559 , n66560 , n66561 , n66562 , n66563 , n66564 , n66565 , n66566 , n66567 , n66568 , 
 n66569 , n66570 , n66571 , n66572 , n66573 , n66574 , n66575 , n66576 , n66577 , n66578 , 
 n66579 , n66580 , n66581 , n66582 , n66583 , n66584 , n66585 , n66586 , n66587 , n66588 , 
 n66589 , n66590 , n66591 , n66592 , n66593 , n66594 , n66595 , n66596 , n66597 , n66598 , 
 n66599 , n66600 , n66601 , n66602 , n66603 , n66604 , n66605 , n66606 , n66607 , n66608 , 
 n66609 , n66610 , n66611 , n66612 , n66613 , n66614 , n66615 , n66616 , n66617 , n66618 , 
 n66619 , n66620 , n66621 , n66622 , n66623 , n66624 , n66625 , n66626 , n66627 , n66628 , 
 n66629 , n66630 , n66631 , n66632 , n66633 , n66634 , n66635 , n66636 , n66637 , n66638 , 
 n66639 , n66640 , n66641 , n66642 , n66643 , n66644 , n66645 , n66646 , n66647 , n66648 , 
 n66649 , n66650 , n66651 , n66652 , n66653 , n66654 , n66655 , n66656 , n66657 , n66658 , 
 n66659 , n66660 , n66661 , n66662 , n66663 , n66664 , n66665 , n66666 , n66667 , n66668 , 
 n66669 , n66670 , n66671 , n66672 , n66673 , n66674 , n66675 , n66676 , n66677 , n66678 , 
 n66679 , n66680 , n66681 , n66682 , n66683 , n66684 , n66685 , n66686 , n66687 , n66688 , 
 n66689 , n66690 , n66691 , n66692 , n66693 , n66694 , n66695 , n66696 , n66697 , n66698 , 
 n66699 , n66700 , n66701 , n66702 , n66703 , n66704 , n66705 , n66706 , n66707 , n66708 , 
 n66709 , n66710 , n66711 , n66712 , n66713 , n66714 , n66715 , n66716 , n66717 , n66718 , 
 n66719 , n66720 , n66721 , n66722 , n66723 , n66724 , n66725 , n66726 , n66727 , n66728 , 
 n66729 , n66730 , n66731 , n66732 , n66733 , n66734 , n66735 , n66736 , n66737 , n66738 , 
 n66739 , n66740 , n66741 , n66742 , n66743 , n66744 , n66745 , n66746 , n66747 , n66748 , 
 n66749 , n66750 , n66751 , n66752 , n66753 , n66754 , n66755 , n66756 , n66757 , n66758 , 
 n66759 , n66760 , n66761 , n66762 , n66763 , n66764 , n66765 , n66766 , n66767 , n66768 , 
 n66769 , n66770 , n66771 , n66772 , n66773 , n66774 , n66775 , n66776 , n66777 , n66778 , 
 n66779 , n66780 , n66781 , n66782 , n66783 , n66784 , n66785 , n66786 , n66787 , n66788 , 
 n66789 , n66790 , n66791 , n66792 , n66793 , n66794 , n66795 , n66796 , n66797 , n66798 , 
 n66799 , n66800 , n66801 , n66802 , n66803 , n66804 , n66805 , n66806 , n66807 , n66808 , 
 n66809 , n66810 , n66811 , n66812 , n66813 , n66814 , n66815 , n66816 , n66817 , n66818 , 
 n66819 , n66820 , n66821 , n66822 , n66823 , n66824 , n66825 , n66826 , n66827 , n66828 , 
 n66829 , n66830 , n66831 , n66832 , n66833 , n66834 , n66835 , n66836 , n66837 , n66838 , 
 n66839 , n66840 , n66841 , n66842 , n66843 , n66844 , n66845 , n66846 , n66847 , n66848 , 
 n66849 , n66850 , n66851 , n66852 , n66853 , n66854 , n66855 , n66856 , n66857 , n66858 , 
 n66859 , n66860 , n66861 , n66862 , n66863 , n66864 , n66865 , n66866 , n66867 , n66868 , 
 n66869 , n66870 , n66871 , n66872 , n66873 , n66874 , n66875 , n66876 , n66877 , n66878 , 
 n66879 , n66880 , n66881 , n66882 , n66883 , n66884 , n66885 , n66886 , n66887 , n66888 , 
 n66889 , n66890 , n66891 , n66892 , n66893 , n66894 , n66895 , n66896 , n66897 , n66898 , 
 n66899 , n66900 , n66901 , n66902 , n66903 , n66904 , n66905 , n66906 , n66907 , n66908 , 
 n66909 , n66910 , n66911 , n66912 , n66913 , n66914 , n66915 , n66916 , n66917 , n66918 , 
 n66919 , n66920 , n66921 , n66922 , n66923 , n66924 , n66925 , n66926 , n66927 , n66928 , 
 n66929 , n66930 , n66931 , n66932 , n66933 , n66934 , n66935 , n66936 , n66937 , n66938 , 
 n66939 , n66940 , n66941 , n66942 , n66943 , n66944 , n66945 , n66946 , n66947 , n66948 , 
 n66949 , n66950 , n66951 , n66952 , n66953 , n66954 , n66955 , n66956 , n66957 , n66958 , 
 n66959 , n66960 , n66961 , n66962 , n66963 , n66964 , n66965 , n66966 , n66967 , n66968 , 
 n66969 , n66970 , n66971 , n66972 , n66973 , n66974 , n66975 , n66976 , n66977 , n66978 , 
 n66979 , n66980 , n66981 , n66982 , n66983 , n66984 , n66985 , n66986 , n66987 , n66988 , 
 n66989 , n66990 , n66991 , n66992 , n66993 , n66994 , n66995 , n66996 , n66997 , n66998 , 
 n66999 , n67000 , n67001 , n67002 , n67003 , n67004 , n67005 , n67006 , n67007 , n67008 , 
 n67009 , n67010 , n67011 , n67012 , n67013 , n67014 , n67015 , n67016 , n67017 , n67018 , 
 n67019 , n67020 , n67021 , n67022 , n67023 , n67024 , n67025 , n67026 , n67027 , n67028 , 
 n67029 , n67030 , n67031 , n67032 , n67033 , n67034 , n67035 , n67036 , n67037 , n67038 , 
 n67039 , n67040 , n67041 , n67042 , n67043 , n67044 , n67045 , n67046 , n67047 , n67048 , 
 n67049 , n67050 , n67051 , n67052 , n67053 , n67054 , n67055 , n67056 , n67057 , n67058 , 
 n67059 , n67060 , n67061 , n67062 , n67063 , n67064 , n67065 , n67066 , n67067 , n67068 , 
 n67069 , n67070 , n67071 , n67072 , n67073 , n67074 , n67075 , n67076 , n67077 , n67078 , 
 n67079 , n67080 , n67081 , n67082 , n67083 , n67084 , n67085 , n67086 , n67087 , n67088 , 
 n67089 , n67090 , n67091 , n67092 , n67093 , n67094 , n67095 , n67096 , n67097 , n67098 , 
 n67099 , n67100 , n67101 , n67102 , n67103 , n67104 , n67105 , n67106 , n67107 , n67108 , 
 n67109 , n67110 , n67111 , n67112 , n67113 , n67114 , n67115 , n67116 , n67117 , n67118 , 
 n67119 , n67120 , n67121 , n67122 , n67123 , n67124 , n67125 , n67126 , n67127 , n67128 , 
 n67129 , n67130 , n67131 , n67132 , n67133 , n67134 , n67135 , n67136 , n67137 , n67138 , 
 n67139 , n67140 , n67141 , n67142 , n67143 , n67144 , n67145 , n67146 , n67147 , n67148 , 
 n67149 , n67150 , n67151 , n67152 , n67153 , n67154 , n67155 , n67156 , n67157 , n67158 , 
 n67159 , n67160 , n67161 , n67162 , n67163 , n67164 , n67165 , n67166 , n67167 , n67168 , 
 n67169 , n67170 , n67171 , n67172 , n67173 , n67174 , n67175 , n67176 , n67177 , n67178 , 
 n67179 , n67180 , n67181 , n67182 , n67183 , n67184 , n67185 , n67186 , n67187 , n67188 , 
 n67189 , n67190 , n67191 , n67192 , n67193 , n67194 , n67195 , n67196 , n67197 , n67198 , 
 n67199 , n67200 , n67201 , n67202 , n67203 , n67204 , n67205 , n67206 , n67207 , n67208 , 
 n67209 , n67210 , n67211 , n67212 , n67213 , n67214 , n67215 , n67216 , n67217 , n67218 , 
 n67219 , n67220 , n67221 , n67222 , n67223 , n67224 , n67225 , n67226 , n67227 , n67228 , 
 n67229 , n67230 , n67231 , n67232 , n67233 , n67234 , n67235 , n67236 , n67237 , n67238 , 
 n67239 , n67240 , n67241 , n67242 , n67243 , n67244 , n67245 , n67246 , n67247 , n67248 , 
 n67249 , n67250 , n67251 , n67252 , n67253 , n67254 , n67255 , n67256 , n67257 , n67258 , 
 n67259 , n67260 , n67261 , n67262 , n67263 , n67264 , n67265 , n67266 , n67267 , n67268 , 
 n67269 , n67270 , n67271 , n67272 , n67273 , n67274 , n67275 , n67276 , n67277 , n67278 , 
 n67279 , n67280 , n67281 , n67282 , n67283 , n67284 , n67285 , n67286 , n67287 , n67288 , 
 n67289 , n67290 , n67291 , n67292 , n67293 , n67294 , n67295 , n67296 , n67297 , n67298 , 
 n67299 , n67300 , n67301 , n67302 , n67303 , n67304 , n67305 , n67306 , n67307 , n67308 , 
 n67309 , n67310 , n67311 , n67312 , n67313 , n67314 , n67315 , n67316 , n67317 , n67318 , 
 n67319 , n67320 , n67321 , n67322 , n67323 , n67324 , n67325 , n67326 , n67327 , n67328 , 
 n67329 , n67330 , n67331 , n67332 , n67333 , n67334 , n67335 , n67336 , n67337 , n67338 , 
 n67339 , n67340 , n67341 , n67342 , n67343 , n67344 , n67345 , n67346 , n67347 , n67348 , 
 n67349 , n67350 , n67351 , n67352 , n67353 , n67354 , n67355 , n67356 , n67357 , n67358 , 
 n67359 , n67360 , n67361 , n67362 , n67363 , n67364 , n67365 , n67366 , n67367 , n67368 , 
 n67369 , n67370 , n67371 , n67372 , n67373 , n67374 , n67375 , n67376 , n67377 , n67378 , 
 n67379 , n67380 , n67381 , n67382 , n67383 , n67384 , n67385 , n67386 , n67387 , n67388 , 
 n67389 , n67390 , n67391 , n67392 , n67393 , n67394 , n67395 , n67396 , n67397 , n67398 , 
 n67399 , n67400 , n67401 , n67402 , n67403 , n67404 , n67405 , n67406 , n67407 , n67408 , 
 n67409 , n67410 , n67411 , n67412 , n67413 , n67414 , n67415 , n67416 , n67417 , n67418 , 
 n67419 , n67420 , n67421 , n67422 , n67423 , n67424 , n67425 , n67426 , n67427 , n67428 , 
 n67429 , n67430 , n67431 , n67432 , n67433 , n67434 , n67435 , n67436 , n67437 , n67438 , 
 n67439 , n67440 , n67441 , n67442 , n67443 , n67444 , n67445 , n67446 , n67447 , n67448 , 
 n67449 , n67450 , n67451 , n67452 , n67453 , n67454 , n67455 , n67456 , n67457 , n67458 , 
 n67459 , n67460 , n67461 , n67462 , n67463 , n67464 , n67465 , n67466 , n67467 , n67468 , 
 n67469 , n67470 , n67471 , n67472 , n67473 , n67474 , n67475 , n67476 , n67477 , n67478 , 
 n67479 , n67480 , n67481 , n67482 , n67483 , n67484 , n67485 , n67486 , n67487 , n67488 , 
 n67489 , n67490 , n67491 , n67492 , n67493 , n67494 , n67495 , n67496 , n67497 , n67498 , 
 n67499 , n67500 , n67501 , n67502 , n67503 , n67504 , n67505 , n67506 , n67507 , n67508 , 
 n67509 , n67510 , n67511 , n67512 , n67513 , n67514 , n67515 , n67516 , n67517 , n67518 , 
 n67519 , n67520 , n67521 , n67522 , n67523 , n67524 , n67525 , n67526 , n67527 , n67528 , 
 n67529 , n67530 , n67531 , n67532 , n67533 , n67534 , n67535 , n67536 , n67537 , n67538 , 
 n67539 , n67540 , n67541 , n67542 , n67543 , n67544 , n67545 , n67546 , n67547 , n67548 , 
 n67549 , n67550 , n67551 , n67552 , n67553 , n67554 , n67555 , n67556 , n67557 , n67558 , 
 n67559 , n67560 , n67561 , n67562 , n67563 , n67564 , n67565 , n67566 , n67567 , n67568 , 
 n67569 , n67570 , n67571 , n67572 , n67573 , n67574 , n67575 , n67576 , n67577 , n67578 , 
 n67579 , n67580 , n67581 , n67582 , n67583 , n67584 , n67585 , n67586 , n67587 , n67588 , 
 n67589 , n67590 , n67591 , n67592 , n67593 , n67594 , n67595 , n67596 , n67597 , n67598 , 
 n67599 , n67600 , n67601 , n67602 , n67603 , n67604 , n67605 , n67606 , n67607 , n67608 , 
 n67609 , n67610 , n67611 , n67612 , n67613 , n67614 , n67615 , n67616 , n67617 , n67618 , 
 n67619 , n67620 , n67621 , n67622 , n67623 , n67624 , n67625 , n67626 , n67627 , n67628 , 
 n67629 , n67630 , n67631 , n67632 , n67633 , n67634 , n67635 , n67636 , n67637 , n67638 , 
 n67639 , n67640 , n67641 , n67642 , n67643 , n67644 , n67645 , n67646 , n67647 , n67648 , 
 n67649 , n67650 , n67651 , n67652 , n67653 , n67654 , n67655 , n67656 , n67657 , n67658 , 
 n67659 , n67660 , n67661 , n67662 , n67663 , n67664 , n67665 , n67666 , n67667 , n67668 , 
 n67669 , n67670 , n67671 , n67672 , n67673 , n67674 , n67675 , n67676 , n67677 , n67678 , 
 n67679 , n67680 , n67681 , n67682 , n67683 , n67684 , n67685 , n67686 , n67687 , n67688 , 
 n67689 , n67690 , n67691 , n67692 , n67693 , n67694 , n67695 , n67696 , n67697 , n67698 , 
 n67699 , n67700 , n67701 , n67702 , n67703 , n67704 , n67705 , n67706 , n67707 , n67708 , 
 n67709 , n67710 , n67711 , n67712 , n67713 , n67714 , n67715 , n67716 , n67717 , n67718 , 
 n67719 , n67720 , n67721 , n67722 , n67723 , n67724 , n67725 , n67726 , n67727 , n67728 , 
 n67729 , n67730 , n67731 , n67732 , n67733 , n67734 , n67735 , n67736 , n67737 , n67738 , 
 n67739 , n67740 , n67741 , n67742 , n67743 , n67744 , n67745 , n67746 , n67747 , n67748 , 
 n67749 , n67750 , n67751 , n67752 , n67753 , n67754 , n67755 , n67756 , n67757 , n67758 , 
 n67759 , n67760 , n67761 , n67762 , n67763 , n67764 , n67765 , n67766 , n67767 , n67768 , 
 n67769 , n67770 , n67771 , n67772 , n67773 , n67774 , n67775 , n67776 , n67777 , n67778 , 
 n67779 , n67780 , n67781 , n67782 , n67783 , n67784 , n67785 , n67786 , n67787 , n67788 , 
 n67789 , n67790 , n67791 , n67792 , n67793 , n67794 , n67795 , n67796 , n67797 , n67798 , 
 n67799 , n67800 , n67801 , n67802 , n67803 , n67804 , n67805 , n67806 , n67807 , n67808 , 
 n67809 , n67810 , n67811 , n67812 , n67813 , n67814 , n67815 , n67816 , n67817 , n67818 , 
 n67819 , n67820 , n67821 , n67822 , n67823 , n67824 , n67825 , n67826 , n67827 , n67828 , 
 n67829 , n67830 , n67831 , n67832 , n67833 , n67834 , n67835 , n67836 , n67837 , n67838 , 
 n67839 , n67840 , n67841 , n67842 , n67843 , n67844 , n67845 , n67846 , n67847 , n67848 , 
 n67849 , n67850 , n67851 , n67852 , n67853 , n67854 , n67855 , n67856 , n67857 , n67858 , 
 n67859 , n67860 , n67861 , n67862 , n67863 , n67864 , n67865 , n67866 , n67867 , n67868 , 
 n67869 , n67870 , n67871 , n67872 , n67873 , n67874 , n67875 , n67876 , n67877 , n67878 , 
 n67879 , n67880 , n67881 , n67882 , n67883 , n67884 , n67885 , n67886 , n67887 , n67888 , 
 n67889 , n67890 , n67891 , n67892 , n67893 , n67894 , n67895 , n67896 , n67897 , n67898 , 
 n67899 , n67900 , n67901 , n67902 , n67903 , n67904 , n67905 , n67906 , n67907 , n67908 , 
 n67909 , n67910 , n67911 , n67912 , n67913 , n67914 , n67915 , n67916 , n67917 , n67918 , 
 n67919 , n67920 , n67921 , n67922 , n67923 , n67924 , n67925 , n67926 , n67927 , n67928 , 
 n67929 , n67930 , n67931 , n67932 , n67933 , n67934 , n67935 , n67936 , n67937 , n67938 , 
 n67939 , n67940 , n67941 , n67942 , n67943 , n67944 , n67945 , n67946 , n67947 , n67948 , 
 n67949 , n67950 , n67951 , n67952 , n67953 , n67954 , n67955 , n67956 , n67957 , n67958 , 
 n67959 , n67960 , n67961 , n67962 , n67963 , n67964 , n67965 , n67966 , n67967 , n67968 , 
 n67969 , n67970 , n67971 , n67972 , n67973 , n67974 , n67975 , n67976 , n67977 , n67978 , 
 n67979 , n67980 , n67981 , n67982 , n67983 , n67984 , n67985 , n67986 , n67987 , n67988 , 
 n67989 , n67990 , n67991 , n67992 , n67993 , n67994 , n67995 , n67996 , n67997 , n67998 , 
 n67999 , n68000 , n68001 , n68002 , n68003 , n68004 , n68005 , n68006 , n68007 , n68008 , 
 n68009 , n68010 , n68011 , n68012 , n68013 , n68014 , n68015 , n68016 , n68017 , n68018 , 
 n68019 , n68020 , n68021 , n68022 , n68023 , n68024 , n68025 , n68026 , n68027 , n68028 , 
 n68029 , n68030 , n68031 , n68032 , n68033 , n68034 , n68035 , n68036 , n68037 , n68038 , 
 n68039 , n68040 , n68041 , n68042 , n68043 , n68044 , n68045 , n68046 , n68047 , n68048 , 
 n68049 , n68050 , n68051 , n68052 , n68053 , n68054 , n68055 , n68056 , n68057 , n68058 , 
 n68059 , n68060 , n68061 , n68062 , n68063 , n68064 , n68065 , n68066 , n68067 , n68068 , 
 n68069 , n68070 , n68071 , n68072 , n68073 , n68074 , n68075 , n68076 , n68077 , n68078 , 
 n68079 , n68080 , n68081 , n68082 , n68083 , n68084 , n68085 , n68086 , n68087 , n68088 , 
 n68089 , n68090 , n68091 , n68092 , n68093 , n68094 , n68095 , n68096 , n68097 , n68098 , 
 n68099 , n68100 , n68101 , n68102 , n68103 , n68104 , n68105 , n68106 , n68107 , n68108 , 
 n68109 , n68110 , n68111 , n68112 , n68113 , n68114 , n68115 , n68116 , n68117 , n68118 , 
 n68119 , n68120 , n68121 , n68122 , n68123 , n68124 , n68125 , n68126 , n68127 , n68128 , 
 n68129 , n68130 , n68131 , n68132 , n68133 , n68134 , n68135 , n68136 , n68137 , n68138 , 
 n68139 , n68140 , n68141 , n68142 , n68143 , n68144 , n68145 , n68146 , n68147 , n68148 , 
 n68149 , n68150 , n68151 , n68152 , n68153 , n68154 , n68155 , n68156 , n68157 , n68158 , 
 n68159 , n68160 , n68161 , n68162 , n68163 , n68164 , n68165 , n68166 , n68167 , n68168 , 
 n68169 , n68170 , n68171 , n68172 , n68173 , n68174 , n68175 , n68176 , n68177 , n68178 , 
 n68179 , n68180 , n68181 , n68182 , n68183 , n68184 , n68185 , n68186 , n68187 , n68188 , 
 n68189 , n68190 , n68191 , n68192 , n68193 , n68194 , n68195 , n68196 , n68197 , n68198 , 
 n68199 , n68200 , n68201 , n68202 , n68203 , n68204 , n68205 , n68206 , n68207 , n68208 , 
 n68209 , n68210 , n68211 , n68212 , n68213 , n68214 , n68215 , n68216 , n68217 , n68218 , 
 n68219 , n68220 , n68221 , n68222 , n68223 , n68224 , n68225 , n68226 , n68227 , n68228 , 
 n68229 , n68230 , n68231 , n68232 , n68233 , n68234 , n68235 , n68236 , n68237 , n68238 , 
 n68239 , n68240 , n68241 , n68242 , n68243 , n68244 , n68245 , n68246 , n68247 , n68248 , 
 n68249 , n68250 , n68251 , n68252 , n68253 , n68254 , n68255 , n68256 , n68257 , n68258 , 
 n68259 , n68260 , n68261 , n68262 , n68263 , n68264 , n68265 , n68266 , n68267 , n68268 , 
 n68269 , n68270 , n68271 , n68272 , n68273 , n68274 , n68275 , n68276 , n68277 , n68278 , 
 n68279 , n68280 , n68281 , n68282 , n68283 , n68284 , n68285 , n68286 , n68287 , n68288 , 
 n68289 , n68290 , n68291 , n68292 , n68293 , n68294 , n68295 , n68296 , n68297 , n68298 , 
 n68299 , n68300 , n68301 , n68302 , n68303 , n68304 , n68305 , n68306 , n68307 , n68308 , 
 n68309 , n68310 , n68311 , n68312 , n68313 , n68314 , n68315 , n68316 , n68317 , n68318 , 
 n68319 , n68320 , n68321 , n68322 , n68323 , n68324 , n68325 , n68326 , n68327 , n68328 , 
 n68329 , n68330 , n68331 , n68332 , n68333 , n68334 , n68335 , n68336 , n68337 , n68338 , 
 n68339 , n68340 , n68341 , n68342 , n68343 , n68344 , n68345 , n68346 , n68347 , n68348 , 
 n68349 , n68350 , n68351 , n68352 , n68353 , n68354 , n68355 , n68356 , n68357 , n68358 , 
 n68359 , n68360 , n68361 , n68362 , n68363 , n68364 , n68365 , n68366 , n68367 , n68368 , 
 n68369 , n68370 , n68371 , n68372 , n68373 , n68374 , n68375 , n68376 , n68377 , n68378 , 
 n68379 , n68380 , n68381 , n68382 , n68383 , n68384 , n68385 , n68386 , n68387 , n68388 , 
 n68389 , n68390 , n68391 , n68392 , n68393 , n68394 , n68395 , n68396 , n68397 , n68398 , 
 n68399 , n68400 , n68401 , n68402 , n68403 , n68404 , n68405 , n68406 , n68407 , n68408 , 
 n68409 , n68410 , n68411 , n68412 , n68413 , n68414 , n68415 , n68416 , n68417 , n68418 , 
 n68419 , n68420 , n68421 , n68422 , n68423 , n68424 , n68425 , n68426 , n68427 , n68428 , 
 n68429 , n68430 , n68431 , n68432 , n68433 , n68434 , n68435 , n68436 , n68437 , n68438 , 
 n68439 , n68440 , n68441 , n68442 , n68443 , n68444 , n68445 , n68446 , n68447 , n68448 , 
 n68449 , n68450 , n68451 , n68452 , n68453 , n68454 , n68455 , n68456 , n68457 , n68458 , 
 n68459 , n68460 , n68461 , n68462 , n68463 , n68464 , n68465 , n68466 , n68467 , n68468 , 
 n68469 , n68470 , n68471 , n68472 , n68473 , n68474 , n68475 , n68476 , n68477 , n68478 , 
 n68479 , n68480 , n68481 , n68482 , n68483 , n68484 , n68485 , n68486 , n68487 , n68488 , 
 n68489 , n68490 , n68491 , n68492 , n68493 , n68494 , n68495 , n68496 , n68497 , n68498 , 
 n68499 , n68500 , n68501 , n68502 , n68503 , n68504 , n68505 , n68506 , n68507 , n68508 , 
 n68509 , n68510 , n68511 , n68512 , n68513 , n68514 , n68515 , n68516 , n68517 , n68518 , 
 n68519 , n68520 , n68521 , n68522 , n68523 , n68524 , n68525 , n68526 , n68527 , n68528 , 
 n68529 , n68530 , n68531 , n68532 , n68533 , n68534 , n68535 , n68536 , n68537 , n68538 , 
 n68539 , n68540 , n68541 , n68542 , n68543 , n68544 , n68545 , n68546 , n68547 , n68548 , 
 n68549 , n68550 , n68551 , n68552 , n68553 , n68554 , n68555 , n68556 , n68557 , n68558 , 
 n68559 , n68560 , n68561 , n68562 , n68563 , n68564 , n68565 , n68566 , n68567 , n68568 , 
 n68569 , n68570 , n68571 , n68572 , n68573 , n68574 , n68575 , n68576 , n68577 , n68578 , 
 n68579 , n68580 , n68581 , n68582 , n68583 , n68584 , n68585 , n68586 , n68587 , n68588 , 
 n68589 , n68590 , n68591 , n68592 , n68593 , n68594 , n68595 , n68596 , n68597 , n68598 , 
 n68599 , n68600 , n68601 , n68602 , n68603 , n68604 , n68605 , n68606 , n68607 , n68608 , 
 n68609 , n68610 , n68611 , n68612 , n68613 , n68614 , n68615 , n68616 , n68617 , n68618 , 
 n68619 , n68620 , n68621 , n68622 , n68623 , n68624 , n68625 , n68626 , n68627 , n68628 , 
 n68629 , n68630 , n68631 , n68632 , n68633 , n68634 , n68635 , n68636 , n68637 , n68638 , 
 n68639 , n68640 , n68641 , n68642 , n68643 , n68644 , n68645 , n68646 , n68647 , n68648 , 
 n68649 , n68650 , n68651 , n68652 , n68653 , n68654 , n68655 , n68656 , n68657 , n68658 , 
 n68659 , n68660 , n68661 , n68662 , n68663 , n68664 , n68665 , n68666 , n68667 , n68668 , 
 n68669 , n68670 , n68671 , n68672 , n68673 , n68674 , n68675 , n68676 , n68677 , n68678 , 
 n68679 , n68680 , n68681 , n68682 , n68683 , n68684 , n68685 , n68686 , n68687 , n68688 , 
 n68689 , n68690 , n68691 , n68692 , n68693 , n68694 , n68695 , n68696 , n68697 , n68698 , 
 n68699 , n68700 , n68701 , n68702 , n68703 , n68704 , n68705 , n68706 , n68707 , n68708 , 
 n68709 , n68710 , n68711 , n68712 , n68713 , n68714 , n68715 , n68716 , n68717 , n68718 , 
 n68719 , n68720 , n68721 , n68722 , n68723 , n68724 , n68725 , n68726 , n68727 , n68728 , 
 n68729 , n68730 , n68731 , n68732 , n68733 , n68734 , n68735 , n68736 , n68737 , n68738 , 
 n68739 , n68740 , n68741 , n68742 , n68743 , n68744 , n68745 , n68746 , n68747 , n68748 , 
 n68749 , n68750 , n68751 , n68752 , n68753 , n68754 , n68755 , n68756 , n68757 , n68758 , 
 n68759 , n68760 , n68761 , n68762 , n68763 , n68764 , n68765 , n68766 , n68767 , n68768 , 
 n68769 , n68770 , n68771 , n68772 , n68773 , n68774 , n68775 , n68776 , n68777 , n68778 , 
 n68779 , n68780 , n68781 , n68782 , n68783 , n68784 , n68785 , n68786 , n68787 , n68788 , 
 n68789 , n68790 , n68791 , n68792 , n68793 , n68794 , n68795 , n68796 , n68797 , n68798 , 
 n68799 , n68800 , n68801 , n68802 , n68803 , n68804 , n68805 , n68806 , n68807 , n68808 , 
 n68809 , n68810 , n68811 , n68812 , n68813 , n68814 , n68815 , n68816 , n68817 , n68818 , 
 n68819 , n68820 , n68821 , n68822 , n68823 , n68824 , n68825 , n68826 , n68827 , n68828 , 
 n68829 , n68830 , n68831 , n68832 , n68833 , n68834 , n68835 , n68836 , n68837 , n68838 , 
 n68839 , n68840 , n68841 , n68842 , n68843 , n68844 , n68845 , n68846 , n68847 , n68848 , 
 n68849 , n68850 , n68851 , n68852 , n68853 , n68854 , n68855 , n68856 , n68857 , n68858 , 
 n68859 , n68860 , n68861 , n68862 , n68863 , n68864 , n68865 , n68866 , n68867 , n68868 , 
 n68869 , n68870 , n68871 , n68872 , n68873 , n68874 , n68875 , n68876 , n68877 , n68878 , 
 n68879 , n68880 , n68881 , n68882 , n68883 , n68884 , n68885 , n68886 , n68887 , n68888 , 
 n68889 , n68890 , n68891 , n68892 , n68893 , n68894 , n68895 , n68896 , n68897 , n68898 , 
 n68899 , n68900 , n68901 , n68902 , n68903 , n68904 , n68905 , n68906 , n68907 , n68908 , 
 n68909 , n68910 , n68911 , n68912 , n68913 , n68914 , n68915 , n68916 , n68917 , n68918 , 
 n68919 , n68920 , n68921 , n68922 , n68923 , n68924 , n68925 , n68926 , n68927 , n68928 , 
 n68929 , n68930 , n68931 , n68932 , n68933 , n68934 , n68935 , n68936 , n68937 , n68938 , 
 n68939 , n68940 , n68941 , n68942 , n68943 , n68944 , n68945 , n68946 , n68947 , n68948 , 
 n68949 , n68950 , n68951 , n68952 , n68953 , n68954 , n68955 , n68956 , n68957 , n68958 , 
 n68959 , n68960 , n68961 , n68962 , n68963 , n68964 , n68965 , n68966 , n68967 , n68968 , 
 n68969 , n68970 , n68971 , n68972 , n68973 , n68974 , n68975 , n68976 , n68977 , n68978 , 
 n68979 , n68980 , n68981 , n68982 , n68983 , n68984 , n68985 , n68986 , n68987 , n68988 , 
 n68989 , n68990 , n68991 , n68992 , n68993 , n68994 , n68995 , n68996 , n68997 , n68998 , 
 n68999 , n69000 , n69001 , n69002 , n69003 , n69004 , n69005 , n69006 , n69007 , n69008 , 
 n69009 , n69010 , n69011 , n69012 , n69013 , n69014 , n69015 , n69016 , n69017 , n69018 , 
 n69019 , n69020 , n69021 , n69022 , n69023 , n69024 , n69025 , n69026 , n69027 , n69028 , 
 n69029 , n69030 , n69031 , n69032 , n69033 , n69034 , n69035 , n69036 , n69037 , n69038 , 
 n69039 , n69040 , n69041 , n69042 , n69043 , n69044 , n69045 , n69046 , n69047 , n69048 , 
 n69049 , n69050 , n69051 , n69052 , n69053 , n69054 , n69055 , n69056 , n69057 , n69058 , 
 n69059 , n69060 , n69061 , n69062 , n69063 , n69064 , n69065 , n69066 , n69067 , n69068 , 
 n69069 , n69070 , n69071 , n69072 , n69073 , n69074 , n69075 , n69076 , n69077 , n69078 , 
 n69079 , n69080 , n69081 , n69082 , n69083 , n69084 , n69085 , n69086 , n69087 , n69088 , 
 n69089 , n69090 , n69091 , n69092 , n69093 , n69094 , n69095 , n69096 , n69097 , n69098 , 
 n69099 , n69100 , n69101 , n69102 , n69103 , n69104 , n69105 , n69106 , n69107 , n69108 , 
 n69109 , n69110 , n69111 , n69112 , n69113 , n69114 , n69115 , n69116 , n69117 , n69118 , 
 n69119 , n69120 , n69121 , n69122 , n69123 , n69124 , n69125 , n69126 , n69127 , n69128 , 
 n69129 , n69130 , n69131 , n69132 , n69133 , n69134 , n69135 , n69136 , n69137 , n69138 , 
 n69139 , n69140 , n69141 , n69142 , n69143 , n69144 , n69145 , n69146 , n69147 , n69148 , 
 n69149 , n69150 , n69151 , n69152 , n69153 , n69154 , n69155 , n69156 , n69157 , n69158 , 
 n69159 , n69160 , n69161 , n69162 , n69163 , n69164 , n69165 , n69166 , n69167 , n69168 , 
 n69169 , n69170 , n69171 , n69172 , n69173 , n69174 , n69175 , n69176 , n69177 , n69178 , 
 n69179 , n69180 , n69181 , n69182 , n69183 , n69184 , n69185 , n69186 , n69187 , n69188 , 
 n69189 , n69190 , n69191 , n69192 , n69193 , n69194 , n69195 , n69196 , n69197 , n69198 , 
 n69199 , n69200 , n69201 , n69202 , n69203 , n69204 , n69205 , n69206 , n69207 , n69208 , 
 n69209 , n69210 , n69211 , n69212 , n69213 , n69214 , n69215 , n69216 , n69217 , n69218 , 
 n69219 , n69220 , n69221 , n69222 , n69223 , n69224 , n69225 , n69226 , n69227 , n69228 , 
 n69229 , n69230 , n69231 , n69232 , n69233 , n69234 , n69235 , n69236 , n69237 , n69238 , 
 n69239 , n69240 , n69241 , n69242 , n69243 , n69244 , n69245 , n69246 , n69247 , n69248 , 
 n69249 , n69250 , n69251 , n69252 , n69253 , n69254 , n69255 , n69256 , n69257 , n69258 , 
 n69259 , n69260 , n69261 , n69262 , n69263 , n69264 , n69265 , n69266 , n69267 , n69268 , 
 n69269 , n69270 , n69271 , n69272 , n69273 , n69274 , n69275 , n69276 , n69277 , n69278 , 
 n69279 , n69280 , n69281 , n69282 , n69283 , n69284 , n69285 , n69286 , n69287 , n69288 , 
 n69289 , n69290 , n69291 , n69292 , n69293 , n69294 , n69295 , n69296 , n69297 , n69298 , 
 n69299 , n69300 , n69301 , n69302 , n69303 , n69304 , n69305 , n69306 , n69307 , n69308 , 
 n69309 , n69310 , n69311 , n69312 , n69313 , n69314 , n69315 , n69316 , n69317 , n69318 , 
 n69319 , n69320 , n69321 , n69322 , n69323 , n69324 , n69325 , n69326 , n69327 , n69328 , 
 n69329 , n69330 , n69331 , n69332 , n69333 , n69334 , n69335 , n69336 , n69337 , n69338 , 
 n69339 , n69340 , n69341 , n69342 , n69343 , n69344 , n69345 , n69346 , n69347 , n69348 , 
 n69349 , n69350 , n69351 , n69352 , n69353 , n69354 , n69355 , n69356 , n69357 , n69358 , 
 n69359 , n69360 , n69361 , n69362 , n69363 , n69364 , n69365 , n69366 , n69367 , n69368 , 
 n69369 , n69370 , n69371 , n69372 , n69373 , n69374 , n69375 , n69376 , n69377 , n69378 , 
 n69379 , n69380 , n69381 , n69382 , n69383 , n69384 , n69385 , n69386 , n69387 , n69388 , 
 n69389 , n69390 , n69391 , n69392 , n69393 , n69394 , n69395 , n69396 , n69397 , n69398 , 
 n69399 , n69400 , n69401 , n69402 , n69403 , n69404 , n69405 , n69406 , n69407 , n69408 , 
 n69409 , n69410 , n69411 , n69412 , n69413 , n69414 , n69415 , n69416 , n69417 , n69418 , 
 n69419 , n69420 , n69421 , n69422 , n69423 , n69424 , n69425 , n69426 , n69427 , n69428 , 
 n69429 , n69430 , n69431 , n69432 , n69433 , n69434 , n69435 , n69436 , n69437 , n69438 , 
 n69439 , n69440 , n69441 , n69442 , n69443 , n69444 , n69445 , n69446 , n69447 , n69448 , 
 n69449 , n69450 , n69451 , n69452 , n69453 , n69454 , n69455 , n69456 , n69457 , n69458 , 
 n69459 , n69460 , n69461 , n69462 , n69463 , n69464 , n69465 , n69466 , n69467 , n69468 , 
 n69469 , n69470 , n69471 , n69472 , n69473 , n69474 , n69475 , n69476 , n69477 , n69478 , 
 n69479 , n69480 , n69481 , n69482 , n69483 , n69484 , n69485 , n69486 , n69487 , n69488 , 
 n69489 , n69490 , n69491 , n69492 , n69493 , n69494 , n69495 , n69496 , n69497 , n69498 , 
 n69499 , n69500 , n69501 , n69502 , n69503 , n69504 , n69505 , n69506 , n69507 , n69508 , 
 n69509 , n69510 , n69511 , n69512 , n69513 , n69514 , n69515 , n69516 , n69517 , n69518 , 
 n69519 , n69520 , n69521 , n69522 , n69523 , n69524 , n69525 , n69526 , n69527 , n69528 , 
 n69529 , n69530 , n69531 , n69532 , n69533 , n69534 , n69535 , n69536 , n69537 , n69538 , 
 n69539 , n69540 , n69541 , n69542 , n69543 , n69544 , n69545 , n69546 , n69547 , n69548 , 
 n69549 , n69550 , n69551 , n69552 , n69553 , n69554 , n69555 , n69556 , n69557 , n69558 , 
 n69559 , n69560 , n69561 , n69562 , n69563 , n69564 , n69565 , n69566 , n69567 , n69568 , 
 n69569 , n69570 , n69571 , n69572 , n69573 , n69574 , n69575 , n69576 , n69577 , n69578 , 
 n69579 , n69580 , n69581 , n69582 , n69583 , n69584 , n69585 , n69586 , n69587 , n69588 , 
 n69589 , n69590 , n69591 , n69592 , n69593 , n69594 , n69595 , n69596 , n69597 , n69598 , 
 n69599 , n69600 , n69601 , n69602 , n69603 , n69604 , n69605 , n69606 , n69607 , n69608 , 
 n69609 , n69610 , n69611 , n69612 , n69613 , n69614 , n69615 , n69616 , n69617 , n69618 , 
 n69619 , n69620 , n69621 , n69622 , n69623 , n69624 , n69625 , n69626 , n69627 , n69628 , 
 n69629 , n69630 , n69631 , n69632 , n69633 , n69634 , n69635 , n69636 , n69637 , n69638 , 
 n69639 , n69640 , n69641 , n69642 , n69643 , n69644 , n69645 , n69646 , n69647 , n69648 , 
 n69649 , n69650 , n69651 , n69652 , n69653 , n69654 , n69655 , n69656 , n69657 , n69658 , 
 n69659 , n69660 , n69661 , n69662 , n69663 , n69664 , n69665 , n69666 , n69667 , n69668 , 
 n69669 , n69670 , n69671 , n69672 , n69673 , n69674 , n69675 , n69676 , n69677 , n69678 , 
 n69679 , n69680 , n69681 , n69682 , n69683 , n69684 , n69685 , n69686 , n69687 , n69688 , 
 n69689 , n69690 , n69691 , n69692 , n69693 , n69694 , n69695 , n69696 , n69697 , n69698 , 
 n69699 , n69700 , n69701 , n69702 , n69703 , n69704 , n69705 , n69706 , n69707 , n69708 , 
 n69709 , n69710 , n69711 , n69712 , n69713 , n69714 , n69715 , n69716 , n69717 , n69718 , 
 n69719 , n69720 , n69721 , n69722 , n69723 , n69724 , n69725 , n69726 , n69727 , n69728 , 
 n69729 , n69730 , n69731 , n69732 , n69733 , n69734 , n69735 , n69736 , n69737 , n69738 , 
 n69739 , n69740 , n69741 , n69742 , n69743 , n69744 , n69745 , n69746 , n69747 , n69748 , 
 n69749 , n69750 , n69751 , n69752 , n69753 , n69754 , n69755 , n69756 , n69757 , n69758 , 
 n69759 , n69760 , n69761 , n69762 , n69763 , n69764 , n69765 , n69766 , n69767 , n69768 , 
 n69769 , n69770 , n69771 , n69772 , n69773 , n69774 , n69775 , n69776 , n69777 , n69778 , 
 n69779 , n69780 , n69781 , n69782 , n69783 , n69784 , n69785 , n69786 , n69787 , n69788 , 
 n69789 , n69790 , n69791 , n69792 , n69793 , n69794 , n69795 , n69796 , n69797 , n69798 , 
 n69799 , n69800 , n69801 , n69802 , n69803 , n69804 , n69805 , n69806 , n69807 , n69808 , 
 n69809 , n69810 , n69811 , n69812 , n69813 , n69814 , n69815 , n69816 , n69817 , n69818 , 
 n69819 , n69820 , n69821 , n69822 , n69823 , n69824 , n69825 , n69826 , n69827 , n69828 , 
 n69829 , n69830 , n69831 , n69832 , n69833 , n69834 , n69835 , n69836 , n69837 , n69838 , 
 n69839 , n69840 , n69841 , n69842 , n69843 , n69844 , n69845 , n69846 , n69847 , n69848 , 
 n69849 , n69850 , n69851 , n69852 , n69853 , n69854 , n69855 , n69856 , n69857 , n69858 , 
 n69859 , n69860 , n69861 , n69862 , n69863 , n69864 , n69865 , n69866 , n69867 , n69868 , 
 n69869 , n69870 , n69871 , n69872 , n69873 , n69874 , n69875 , n69876 , n69877 , n69878 , 
 n69879 , n69880 , n69881 , n69882 , n69883 , n69884 , n69885 , n69886 , n69887 , n69888 , 
 n69889 , n69890 , n69891 , n69892 , n69893 , n69894 , n69895 , n69896 , n69897 , n69898 , 
 n69899 , n69900 , n69901 , n69902 , n69903 , n69904 , n69905 , n69906 , n69907 , n69908 , 
 n69909 , n69910 , n69911 , n69912 , n69913 , n69914 , n69915 , n69916 , n69917 , n69918 , 
 n69919 , n69920 , n69921 , n69922 , n69923 , n69924 , n69925 , n69926 , n69927 , n69928 , 
 n69929 , n69930 , n69931 , n69932 , n69933 , n69934 , n69935 , n69936 , n69937 , n69938 , 
 n69939 , n69940 , n69941 , n69942 , n69943 , n69944 , n69945 , n69946 , n69947 , n69948 , 
 n69949 , n69950 , n69951 , n69952 , n69953 , n69954 , n69955 , n69956 , n69957 , n69958 , 
 n69959 , n69960 , n69961 , n69962 , n69963 , n69964 , n69965 , n69966 , n69967 , n69968 , 
 n69969 , n69970 , n69971 , n69972 , n69973 , n69974 , n69975 , n69976 , n69977 , n69978 , 
 n69979 , n69980 , n69981 , n69982 , n69983 , n69984 , n69985 , n69986 , n69987 , n69988 , 
 n69989 , n69990 , n69991 , n69992 , n69993 , n69994 , n69995 , n69996 , n69997 , n69998 , 
 n69999 , n70000 , n70001 , n70002 , n70003 , n70004 , n70005 , n70006 , n70007 , n70008 , 
 n70009 , n70010 , n70011 , n70012 , n70013 , n70014 , n70015 , n70016 , n70017 , n70018 , 
 n70019 , n70020 , n70021 , n70022 , n70023 , n70024 , n70025 , n70026 , n70027 , n70028 , 
 n70029 , n70030 , n70031 , n70032 , n70033 , n70034 , n70035 , n70036 , n70037 , n70038 , 
 n70039 , n70040 , n70041 , n70042 , n70043 , n70044 , n70045 , n70046 , n70047 , n70048 , 
 n70049 , n70050 , n70051 , n70052 , n70053 , n70054 , n70055 , n70056 , n70057 , n70058 , 
 n70059 , n70060 , n70061 , n70062 , n70063 , n70064 , n70065 , n70066 , n70067 , n70068 , 
 n70069 , n70070 , n70071 , n70072 , n70073 , n70074 , n70075 , n70076 , n70077 , n70078 , 
 n70079 , n70080 , n70081 , n70082 , n70083 , n70084 , n70085 , n70086 , n70087 , n70088 , 
 n70089 , n70090 , n70091 , n70092 , n70093 , n70094 , n70095 , n70096 , n70097 , n70098 , 
 n70099 , n70100 , n70101 , n70102 , n70103 , n70104 , n70105 , n70106 , n70107 , n70108 , 
 n70109 , n70110 , n70111 , n70112 , n70113 , n70114 , n70115 , n70116 , n70117 , n70118 , 
 n70119 , n70120 , n70121 , n70122 , n70123 , n70124 , n70125 , n70126 , n70127 , n70128 , 
 n70129 , n70130 , n70131 , n70132 , n70133 , n70134 , n70135 , n70136 , n70137 , n70138 , 
 n70139 , n70140 , n70141 , n70142 , n70143 , n70144 , n70145 , n70146 , n70147 , n70148 , 
 n70149 , n70150 , n70151 , n70152 , n70153 , n70154 , n70155 , n70156 , n70157 , n70158 , 
 n70159 , n70160 , n70161 , n70162 , n70163 , n70164 , n70165 , n70166 , n70167 , n70168 , 
 n70169 , n70170 , n70171 , n70172 , n70173 , n70174 , n70175 , n70176 , n70177 , n70178 , 
 n70179 , n70180 , n70181 , n70182 , n70183 , n70184 , n70185 , n70186 , n70187 , n70188 , 
 n70189 , n70190 , n70191 , n70192 , n70193 , n70194 , n70195 , n70196 , n70197 , n70198 , 
 n70199 , n70200 , n70201 , n70202 , n70203 , n70204 , n70205 , n70206 , n70207 , n70208 , 
 n70209 , n70210 , n70211 , n70212 , n70213 , n70214 , n70215 , n70216 , n70217 , n70218 , 
 n70219 , n70220 , n70221 , n70222 , n70223 , n70224 , n70225 , n70226 , n70227 , n70228 , 
 n70229 , n70230 , n70231 , n70232 , n70233 , n70234 , n70235 , n70236 , n70237 , n70238 , 
 n70239 , n70240 , n70241 , n70242 , n70243 , n70244 , n70245 , n70246 , n70247 , n70248 , 
 n70249 , n70250 , n70251 , n70252 , n70253 , n70254 , n70255 , n70256 , n70257 , n70258 , 
 n70259 , n70260 , n70261 , n70262 , n70263 , n70264 , n70265 , n70266 , n70267 , n70268 , 
 n70269 , n70270 , n70271 , n70272 , n70273 , n70274 , n70275 , n70276 , n70277 , n70278 , 
 n70279 , n70280 , n70281 , n70282 , n70283 , n70284 , n70285 , n70286 , n70287 , n70288 , 
 n70289 , n70290 , n70291 , n70292 , n70293 , n70294 , n70295 , n70296 , n70297 , n70298 , 
 n70299 , n70300 , n70301 , n70302 , n70303 , n70304 , n70305 , n70306 , n70307 , n70308 , 
 n70309 , n70310 , n70311 , n70312 , n70313 , n70314 , n70315 , n70316 , n70317 , n70318 , 
 n70319 , n70320 , n70321 , n70322 , n70323 , n70324 , n70325 , n70326 , n70327 , n70328 , 
 n70329 , n70330 , n70331 , n70332 , n70333 , n70334 , n70335 , n70336 , n70337 , n70338 , 
 n70339 , n70340 , n70341 , n70342 , n70343 , n70344 , n70345 , n70346 , n70347 , n70348 , 
 n70349 , n70350 , n70351 , n70352 , n70353 , n70354 , n70355 , n70356 , n70357 , n70358 , 
 n70359 , n70360 , n70361 , n70362 , n70363 , n70364 , n70365 , n70366 , n70367 , n70368 , 
 n70369 , n70370 , n70371 , n70372 , n70373 , n70374 , n70375 , n70376 , n70377 , n70378 , 
 n70379 , n70380 , n70381 , n70382 , n70383 , n70384 , n70385 , n70386 , n70387 , n70388 , 
 n70389 , n70390 , n70391 , n70392 , n70393 , n70394 , n70395 , n70396 , n70397 , n70398 , 
 n70399 , n70400 , n70401 , n70402 , n70403 , n70404 , n70405 , n70406 , n70407 , n70408 , 
 n70409 , n70410 , n70411 , n70412 , n70413 , n70414 , n70415 , n70416 , n70417 , n70418 , 
 n70419 , n70420 , n70421 , n70422 , n70423 , n70424 , n70425 , n70426 , n70427 , n70428 , 
 n70429 , n70430 , n70431 , n70432 , n70433 , n70434 , n70435 , n70436 , n70437 , n70438 , 
 n70439 , n70440 , n70441 , n70442 , n70443 , n70444 , n70445 , n70446 , n70447 , n70448 , 
 n70449 , n70450 , n70451 , n70452 , n70453 , n70454 , n70455 , n70456 , n70457 , n70458 , 
 n70459 , n70460 , n70461 , n70462 , n70463 , n70464 , n70465 , n70466 , n70467 , n70468 , 
 n70469 , n70470 , n70471 , n70472 , n70473 , n70474 , n70475 , n70476 , n70477 , n70478 , 
 n70479 , n70480 , n70481 , n70482 , n70483 , n70484 , n70485 , n70486 , n70487 , n70488 , 
 n70489 , n70490 , n70491 , n70492 , n70493 , n70494 , n70495 , n70496 , n70497 , n70498 , 
 n70499 , n70500 , n70501 , n70502 , n70503 , n70504 , n70505 , n70506 , n70507 , n70508 , 
 n70509 , n70510 , n70511 , n70512 , n70513 , n70514 , n70515 , n70516 , n70517 , n70518 , 
 n70519 , n70520 , n70521 , n70522 , n70523 , n70524 , n70525 , n70526 , n70527 , n70528 , 
 n70529 , n70530 , n70531 , n70532 , n70533 , n70534 , n70535 , n70536 , n70537 , n70538 , 
 n70539 , n70540 , n70541 , n70542 , n70543 , n70544 , n70545 , n70546 , n70547 , n70548 , 
 n70549 , n70550 , n70551 , n70552 , n70553 , n70554 , n70555 , n70556 , n70557 , n70558 , 
 n70559 , n70560 , n70561 , n70562 , n70563 , n70564 , n70565 , n70566 , n70567 , n70568 , 
 n70569 , n70570 , n70571 , n70572 , n70573 , n70574 , n70575 , n70576 , n70577 , n70578 , 
 n70579 , n70580 , n70581 , n70582 , n70583 , n70584 , n70585 , n70586 , n70587 , n70588 , 
 n70589 , n70590 , n70591 , n70592 , n70593 , n70594 , n70595 , n70596 , n70597 , n70598 , 
 n70599 , n70600 , n70601 , n70602 , n70603 , n70604 , n70605 , n70606 , n70607 , n70608 , 
 n70609 , n70610 , n70611 , n70612 , n70613 , n70614 , n70615 , n70616 , n70617 , n70618 , 
 n70619 , n70620 , n70621 , n70622 , n70623 , n70624 , n70625 , n70626 , n70627 , n70628 , 
 n70629 , n70630 , n70631 , n70632 , n70633 , n70634 , n70635 , n70636 , n70637 , n70638 , 
 n70639 , n70640 , n70641 , n70642 , n70643 , n70644 , n70645 , n70646 , n70647 , n70648 , 
 n70649 , n70650 , n70651 , n70652 , n70653 , n70654 , n70655 , n70656 , n70657 , n70658 , 
 n70659 , n70660 , n70661 , n70662 , n70663 , n70664 , n70665 , n70666 , n70667 , n70668 , 
 n70669 , n70670 , n70671 , n70672 , n70673 , n70674 , n70675 , n70676 , n70677 , n70678 , 
 n70679 , n70680 , n70681 , n70682 , n70683 , n70684 , n70685 , n70686 , n70687 , n70688 , 
 n70689 , n70690 , n70691 , n70692 , n70693 , n70694 , n70695 , n70696 , n70697 , n70698 , 
 n70699 , n70700 , n70701 , n70702 , n70703 , n70704 , n70705 , n70706 , n70707 , n70708 , 
 n70709 , n70710 , n70711 , n70712 , n70713 , n70714 , n70715 , n70716 , n70717 , n70718 , 
 n70719 , n70720 , n70721 , n70722 , n70723 , n70724 , n70725 , n70726 , n70727 , n70728 , 
 n70729 , n70730 , n70731 , n70732 , n70733 , n70734 , n70735 , n70736 , n70737 , n70738 , 
 n70739 , n70740 , n70741 , n70742 , n70743 , n70744 , n70745 , n70746 , n70747 , n70748 , 
 n70749 , n70750 , n70751 , n70752 , n70753 , n70754 , n70755 , n70756 , n70757 , n70758 , 
 n70759 , n70760 , n70761 , n70762 , n70763 , n70764 , n70765 , n70766 , n70767 , n70768 , 
 n70769 , n70770 , n70771 , n70772 , n70773 , n70774 , n70775 , n70776 , n70777 , n70778 , 
 n70779 , n70780 , n70781 , n70782 , n70783 , n70784 , n70785 , n70786 , n70787 , n70788 , 
 n70789 , n70790 , n70791 , n70792 , n70793 , n70794 , n70795 , n70796 , n70797 , n70798 , 
 n70799 , n70800 , n70801 , n70802 , n70803 , n70804 , n70805 , n70806 , n70807 , n70808 , 
 n70809 , n70810 , n70811 , n70812 , n70813 , n70814 , n70815 , n70816 , n70817 , n70818 , 
 n70819 , n70820 , n70821 , n70822 , n70823 , n70824 , n70825 , n70826 , n70827 , n70828 , 
 n70829 , n70830 , n70831 , n70832 , n70833 , n70834 , n70835 , n70836 , n70837 , n70838 , 
 n70839 , n70840 , n70841 , n70842 , n70843 , n70844 , n70845 , n70846 , n70847 , n70848 , 
 n70849 , n70850 , n70851 , n70852 , n70853 , n70854 , n70855 , n70856 , n70857 , n70858 , 
 n70859 , n70860 , n70861 , n70862 , n70863 , n70864 , n70865 , n70866 , n70867 , n70868 , 
 n70869 , n70870 , n70871 , n70872 , n70873 , n70874 , n70875 , n70876 , n70877 , n70878 , 
 n70879 , n70880 , n70881 , n70882 , n70883 , n70884 , n70885 , n70886 , n70887 , n70888 , 
 n70889 , n70890 , n70891 , n70892 , n70893 , n70894 , n70895 , n70896 , n70897 , n70898 , 
 n70899 , n70900 , n70901 , n70902 , n70903 , n70904 , n70905 , n70906 , n70907 , n70908 , 
 n70909 , n70910 , n70911 , n70912 , n70913 , n70914 , n70915 , n70916 , n70917 , n70918 , 
 n70919 , n70920 , n70921 , n70922 , n70923 , n70924 , n70925 , n70926 , n70927 , n70928 , 
 n70929 , n70930 , n70931 , n70932 , n70933 , n70934 , n70935 , n70936 , n70937 , n70938 , 
 n70939 , n70940 , n70941 , n70942 , n70943 , n70944 , n70945 , n70946 , n70947 , n70948 , 
 n70949 , n70950 , n70951 , n70952 , n70953 , n70954 , n70955 , n70956 , n70957 , n70958 , 
 n70959 , n70960 , n70961 , n70962 , n70963 , n70964 , n70965 , n70966 , n70967 , n70968 , 
 n70969 , n70970 , n70971 , n70972 , n70973 , n70974 , n70975 , n70976 , n70977 , n70978 , 
 n70979 , n70980 , n70981 , n70982 , n70983 , n70984 , n70985 , n70986 , n70987 , n70988 , 
 n70989 , n70990 , n70991 , n70992 , n70993 , n70994 , n70995 , n70996 , n70997 , n70998 , 
 n70999 , n71000 , n71001 , n71002 , n71003 , n71004 , n71005 , n71006 , n71007 , n71008 , 
 n71009 , n71010 , n71011 , n71012 , n71013 , n71014 , n71015 , n71016 , n71017 , n71018 , 
 n71019 , n71020 , n71021 , n71022 , n71023 , n71024 , n71025 , n71026 , n71027 , n71028 , 
 n71029 , n71030 , n71031 , n71032 , n71033 , n71034 , n71035 , n71036 , n71037 , n71038 , 
 n71039 , n71040 , n71041 , n71042 , n71043 , n71044 , n71045 , n71046 , n71047 , n71048 , 
 n71049 , n71050 , n71051 , n71052 , n71053 , n71054 , n71055 , n71056 , n71057 , n71058 , 
 n71059 , n71060 , n71061 , n71062 , n71063 , n71064 , n71065 , n71066 , n71067 , n71068 , 
 n71069 , n71070 , n71071 , n71072 , n71073 , n71074 , n71075 , n71076 , n71077 , n71078 , 
 n71079 , n71080 , n71081 , n71082 , n71083 , n71084 , n71085 , n71086 , n71087 , n71088 , 
 n71089 , n71090 , n71091 , n71092 , n71093 , n71094 , n71095 , n71096 , n71097 , n71098 , 
 n71099 , n71100 , n71101 , n71102 , n71103 , n71104 , n71105 , n71106 , n71107 , n71108 , 
 n71109 , n71110 , n71111 , n71112 , n71113 , n71114 , n71115 , n71116 , n71117 , n71118 , 
 n71119 , n71120 , n71121 , n71122 , n71123 , n71124 , n71125 , n71126 , n71127 , n71128 , 
 n71129 , n71130 , n71131 , n71132 , n71133 , n71134 , n71135 , n71136 , n71137 , n71138 , 
 n71139 , n71140 , n71141 , n71142 , n71143 , n71144 , n71145 , n71146 , n71147 , n71148 , 
 n71149 , n71150 , n71151 , n71152 , n71153 , n71154 , n71155 , n71156 , n71157 , n71158 , 
 n71159 , n71160 , n71161 , n71162 , n71163 , n71164 , n71165 , n71166 , n71167 , n71168 , 
 n71169 , n71170 , n71171 , n71172 , n71173 , n71174 , n71175 , n71176 , n71177 , n71178 , 
 n71179 , n71180 , n71181 , n71182 , n71183 , n71184 , n71185 , n71186 , n71187 , n71188 , 
 n71189 , n71190 , n71191 , n71192 , n71193 , n71194 , n71195 , n71196 , n71197 , n71198 , 
 n71199 , n71200 , n71201 , n71202 , n71203 , n71204 , n71205 , n71206 , n71207 , n71208 , 
 n71209 , n71210 , n71211 , n71212 , n71213 , n71214 , n71215 , n71216 , n71217 , n71218 , 
 n71219 , n71220 , n71221 , n71222 , n71223 , n71224 , n71225 , n71226 , n71227 , n71228 , 
 n71229 , n71230 , n71231 , n71232 , n71233 , n71234 , n71235 , n71236 , n71237 , n71238 , 
 n71239 , n71240 , n71241 , n71242 , n71243 , n71244 , n71245 , n71246 , n71247 , n71248 , 
 n71249 , n71250 , n71251 , n71252 , n71253 , n71254 , n71255 , n71256 , n71257 , n71258 , 
 n71259 , n71260 , n71261 , n71262 , n71263 , n71264 , n71265 , n71266 , n71267 , n71268 , 
 n71269 , n71270 , n71271 , n71272 , n71273 , n71274 , n71275 , n71276 , n71277 , n71278 , 
 n71279 , n71280 , n71281 , n71282 , n71283 , n71284 , n71285 , n71286 , n71287 , n71288 , 
 n71289 , n71290 , n71291 , n71292 , n71293 , n71294 , n71295 , n71296 , n71297 , n71298 , 
 n71299 , n71300 , n71301 , n71302 , n71303 , n71304 , n71305 , n71306 , n71307 , n71308 , 
 n71309 , n71310 , n71311 , n71312 , n71313 , n71314 , n71315 , n71316 , n71317 , n71318 , 
 n71319 , n71320 , n71321 , n71322 , n71323 , n71324 , n71325 , n71326 , n71327 , n71328 , 
 n71329 , n71330 , n71331 , n71332 , n71333 , n71334 , n71335 , n71336 , n71337 , n71338 , 
 n71339 , n71340 , n71341 , n71342 , n71343 , n71344 , n71345 , n71346 , n71347 , n71348 , 
 n71349 , n71350 , n71351 , n71352 , n71353 , n71354 , n71355 , n71356 , n71357 , n71358 , 
 n71359 , n71360 , n71361 , n71362 , n71363 , n71364 , n71365 , n71366 , n71367 , n71368 , 
 n71369 , n71370 , n71371 , n71372 , n71373 , n71374 , n71375 , n71376 , n71377 , n71378 , 
 n71379 , n71380 , n71381 , n71382 , n71383 , n71384 , n71385 , n71386 , n71387 , n71388 , 
 n71389 , n71390 , n71391 , n71392 , n71393 , n71394 , n71395 , n71396 , n71397 , n71398 , 
 n71399 , n71400 , n71401 , n71402 , n71403 , n71404 , n71405 , n71406 , n71407 , n71408 , 
 n71409 , n71410 , n71411 , n71412 , n71413 , n71414 , n71415 , n71416 , n71417 , n71418 , 
 n71419 , n71420 , n71421 , n71422 , n71423 , n71424 , n71425 , n71426 , n71427 , n71428 , 
 n71429 , n71430 , n71431 , n71432 , n71433 , n71434 , n71435 , n71436 , n71437 , n71438 , 
 n71439 , n71440 , n71441 , n71442 , n71443 , n71444 , n71445 , n71446 , n71447 , n71448 , 
 n71449 , n71450 , n71451 , n71452 , n71453 , n71454 , n71455 , n71456 , n71457 , n71458 , 
 n71459 , n71460 , n71461 , n71462 , n71463 , n71464 , n71465 , n71466 , n71467 , n71468 , 
 n71469 , n71470 , n71471 , n71472 , n71473 , n71474 , n71475 , n71476 , n71477 , n71478 , 
 n71479 , n71480 , n71481 , n71482 , n71483 , n71484 , n71485 , n71486 , n71487 , n71488 , 
 n71489 , n71490 , n71491 , n71492 , n71493 , n71494 , n71495 , n71496 , n71497 , n71498 , 
 n71499 , n71500 , n71501 , n71502 , n71503 , n71504 , n71505 , n71506 , n71507 , n71508 , 
 n71509 , n71510 , n71511 , n71512 , n71513 , n71514 , n71515 , n71516 , n71517 , n71518 , 
 n71519 , n71520 , n71521 , n71522 , n71523 , n71524 , n71525 , n71526 , n71527 , n71528 , 
 n71529 , n71530 , n71531 , n71532 , n71533 , n71534 , n71535 , n71536 , n71537 , n71538 , 
 n71539 , n71540 , n71541 , n71542 , n71543 , n71544 , n71545 , n71546 , n71547 , n71548 , 
 n71549 , n71550 , n71551 , n71552 , n71553 , n71554 , n71555 , n71556 , n71557 , n71558 , 
 n71559 , n71560 , n71561 , n71562 , n71563 , n71564 , n71565 , n71566 , n71567 , n71568 , 
 n71569 , n71570 , n71571 , n71572 , n71573 , n71574 , n71575 , n71576 , n71577 , n71578 , 
 n71579 , n71580 , n71581 , n71582 , n71583 , n71584 , n71585 , n71586 , n71587 , n71588 , 
 n71589 , n71590 , n71591 , n71592 , n71593 , n71594 , n71595 , n71596 , n71597 , n71598 , 
 n71599 , n71600 , n71601 , n71602 , n71603 , n71604 , n71605 , n71606 , n71607 , n71608 , 
 n71609 , n71610 , n71611 , n71612 , n71613 , n71614 , n71615 , n71616 , n71617 , n71618 , 
 n71619 , n71620 , n71621 , n71622 , n71623 , n71624 , n71625 , n71626 , n71627 , n71628 , 
 n71629 , n71630 , n71631 , n71632 , n71633 , n71634 , n71635 , n71636 , n71637 , n71638 , 
 n71639 , n71640 , n71641 , n71642 , n71643 , n71644 , n71645 , n71646 , n71647 , n71648 , 
 n71649 , n71650 , n71651 , n71652 , n71653 , n71654 , n71655 , n71656 , n71657 , n71658 , 
 n71659 , n71660 , n71661 , n71662 , n71663 , n71664 , n71665 , n71666 , n71667 , n71668 , 
 n71669 , n71670 , n71671 , n71672 , n71673 , n71674 , n71675 , n71676 , n71677 , n71678 , 
 n71679 , n71680 , n71681 , n71682 , n71683 , n71684 , n71685 , n71686 , n71687 , n71688 , 
 n71689 , n71690 , n71691 , n71692 , n71693 , n71694 , n71695 , n71696 , n71697 , n71698 , 
 n71699 , n71700 , n71701 , n71702 , n71703 , n71704 , n71705 , n71706 , n71707 , n71708 , 
 n71709 , n71710 , n71711 , n71712 , n71713 , n71714 , n71715 , n71716 , n71717 , n71718 , 
 n71719 , n71720 , n71721 , n71722 , n71723 , n71724 , n71725 , n71726 , n71727 , n71728 , 
 n71729 , n71730 , n71731 , n71732 , n71733 , n71734 , n71735 , n71736 , n71737 , n71738 , 
 n71739 , n71740 , n71741 , n71742 , n71743 , n71744 , n71745 , n71746 , n71747 , n71748 , 
 n71749 , n71750 , n71751 , n71752 , n71753 , n71754 , n71755 , n71756 , n71757 , n71758 , 
 n71759 , n71760 , n71761 , n71762 , n71763 , n71764 , n71765 , n71766 , n71767 , n71768 , 
 n71769 , n71770 , n71771 , n71772 , n71773 , n71774 , n71775 , n71776 , n71777 , n71778 , 
 n71779 , n71780 , n71781 , n71782 , n71783 , n71784 , n71785 , n71786 , n71787 , n71788 , 
 n71789 , n71790 , n71791 , n71792 , n71793 , n71794 , n71795 , n71796 , n71797 , n71798 , 
 n71799 , n71800 , n71801 , n71802 , n71803 , n71804 , n71805 , n71806 , n71807 , n71808 , 
 n71809 , n71810 , n71811 , n71812 , n71813 , n71814 , n71815 , n71816 , n71817 , n71818 , 
 n71819 , n71820 , n71821 , n71822 , n71823 , n71824 , n71825 , n71826 , n71827 , n71828 , 
 n71829 , n71830 , n71831 , n71832 , n71833 , n71834 , n71835 , n71836 , n71837 , n71838 , 
 n71839 , n71840 , n71841 , n71842 , n71843 , n71844 , n71845 , n71846 , n71847 , n71848 , 
 n71849 , n71850 , n71851 , n71852 , n71853 , n71854 , n71855 , n71856 , n71857 , n71858 , 
 n71859 , n71860 , n71861 , n71862 , n71863 , n71864 , n71865 , n71866 , n71867 , n71868 , 
 n71869 , n71870 , n71871 , n71872 , n71873 , n71874 , n71875 , n71876 , n71877 , n71878 , 
 n71879 , n71880 , n71881 , n71882 , n71883 , n71884 , n71885 , n71886 , n71887 , n71888 , 
 n71889 , n71890 , n71891 , n71892 , n71893 , n71894 , n71895 , n71896 , n71897 , n71898 , 
 n71899 , n71900 , n71901 , n71902 , n71903 , n71904 , n71905 , n71906 , n71907 , n71908 , 
 n71909 , n71910 , n71911 , n71912 , n71913 , n71914 , n71915 , n71916 , n71917 , n71918 , 
 n71919 , n71920 , n71921 , n71922 , n71923 , n71924 , n71925 , n71926 , n71927 , n71928 , 
 n71929 , n71930 , n71931 , n71932 , n71933 , n71934 , n71935 , n71936 , n71937 , n71938 , 
 n71939 , n71940 , n71941 , n71942 , n71943 , n71944 , n71945 , n71946 , n71947 , n71948 , 
 n71949 , n71950 , n71951 , n71952 , n71953 , n71954 , n71955 , n71956 , n71957 , n71958 , 
 n71959 , n71960 , n71961 , n71962 , n71963 , n71964 , n71965 , n71966 , n71967 , n71968 , 
 n71969 , n71970 , n71971 , n71972 , n71973 , n71974 , n71975 , n71976 , n71977 , n71978 , 
 n71979 , n71980 , n71981 , n71982 , n71983 , n71984 , n71985 , n71986 , n71987 , n71988 , 
 n71989 , n71990 , n71991 , n71992 , n71993 , n71994 , n71995 , n71996 , n71997 , n71998 , 
 n71999 , n72000 , n72001 , n72002 , n72003 , n72004 , n72005 , n72006 , n72007 , n72008 , 
 n72009 , n72010 , n72011 , n72012 , n72013 , n72014 , n72015 , n72016 , n72017 , n72018 , 
 n72019 , n72020 , n72021 , n72022 , n72023 , n72024 , n72025 , n72026 , n72027 , n72028 , 
 n72029 , n72030 , n72031 , n72032 , n72033 , n72034 , n72035 , n72036 , n72037 , n72038 , 
 n72039 , n72040 , n72041 , n72042 , n72043 , n72044 , n72045 , n72046 , n72047 , n72048 , 
 n72049 , n72050 , n72051 , n72052 , n72053 , n72054 , n72055 , n72056 , n72057 , n72058 , 
 n72059 , n72060 , n72061 , n72062 , n72063 , n72064 , n72065 , n72066 , n72067 , n72068 , 
 n72069 , n72070 , n72071 , n72072 , n72073 , n72074 , n72075 , n72076 , n72077 , n72078 , 
 n72079 , n72080 , n72081 , n72082 , n72083 , n72084 , n72085 , n72086 , n72087 , n72088 , 
 n72089 , n72090 , n72091 , n72092 , n72093 , n72094 , n72095 , n72096 , n72097 , n72098 , 
 n72099 , n72100 , n72101 , n72102 , n72103 , n72104 , n72105 , n72106 , n72107 , n72108 , 
 n72109 , n72110 , n72111 , n72112 , n72113 , n72114 , n72115 , n72116 , n72117 , n72118 , 
 n72119 , n72120 , n72121 , n72122 , n72123 , n72124 , n72125 , n72126 , n72127 , n72128 , 
 n72129 , n72130 , n72131 , n72132 , n72133 , n72134 , n72135 , n72136 , n72137 , n72138 , 
 n72139 , n72140 , n72141 , n72142 , n72143 , n72144 , n72145 , n72146 , n72147 , n72148 , 
 n72149 , n72150 , n72151 , n72152 , n72153 , n72154 , n72155 , n72156 , n72157 , n72158 , 
 n72159 , n72160 , n72161 , n72162 , n72163 , n72164 , n72165 , n72166 , n72167 , n72168 , 
 n72169 , n72170 , n72171 , n72172 , n72173 , n72174 , n72175 , n72176 , n72177 , n72178 , 
 n72179 , n72180 , n72181 , n72182 , n72183 , n72184 , n72185 , n72186 , n72187 , n72188 , 
 n72189 , n72190 , n72191 , n72192 , n72193 , n72194 , n72195 , n72196 , n72197 , n72198 , 
 n72199 , n72200 , n72201 , n72202 , n72203 , n72204 , n72205 , n72206 , n72207 , n72208 , 
 n72209 , n72210 , n72211 , n72212 , n72213 , n72214 , n72215 , n72216 , n72217 , n72218 , 
 n72219 , n72220 , n72221 , n72222 , n72223 , n72224 , n72225 , n72226 , n72227 , n72228 , 
 n72229 , n72230 , n72231 , n72232 , n72233 , n72234 , n72235 , n72236 , n72237 , n72238 , 
 n72239 , n72240 , n72241 , n72242 , n72243 , n72244 , n72245 , n72246 , n72247 , n72248 , 
 n72249 , n72250 , n72251 , n72252 , n72253 , n72254 , n72255 , n72256 , n72257 , n72258 , 
 n72259 , n72260 , n72261 , n72262 , n72263 , n72264 , n72265 , n72266 , n72267 , n72268 , 
 n72269 , n72270 , n72271 , n72272 , n72273 , n72274 , n72275 , n72276 , n72277 , n72278 , 
 n72279 , n72280 , n72281 , n72282 , n72283 , n72284 , n72285 , n72286 , n72287 , n72288 , 
 n72289 , n72290 , n72291 , n72292 , n72293 , n72294 , n72295 , n72296 , n72297 , n72298 , 
 n72299 , n72300 , n72301 , n72302 , n72303 , n72304 , n72305 , n72306 , n72307 , n72308 , 
 n72309 , n72310 , n72311 , n72312 , n72313 , n72314 , n72315 , n72316 , n72317 , n72318 , 
 n72319 , n72320 , n72321 , n72322 , n72323 , n72324 , n72325 , n72326 , n72327 , n72328 , 
 n72329 , n72330 , n72331 , n72332 , n72333 , n72334 , n72335 , n72336 , n72337 , n72338 , 
 n72339 , n72340 , n72341 , n72342 , n72343 , n72344 , n72345 , n72346 , n72347 , n72348 , 
 n72349 , n72350 , n72351 , n72352 , n72353 , n72354 , n72355 , n72356 , n72357 , n72358 , 
 n72359 , n72360 , n72361 , n72362 , n72363 , n72364 , n72365 , n72366 , n72367 , n72368 , 
 n72369 , n72370 , n72371 , n72372 , n72373 , n72374 , n72375 , n72376 , n72377 , n72378 , 
 n72379 , n72380 , n72381 , n72382 , n72383 , n72384 , n72385 , n72386 , n72387 , n72388 , 
 n72389 , n72390 , n72391 , n72392 , n72393 , n72394 , n72395 , n72396 , n72397 , n72398 , 
 n72399 , n72400 , n72401 , n72402 , n72403 , n72404 , n72405 , n72406 , n72407 , n72408 , 
 n72409 , n72410 , n72411 , n72412 , n72413 , n72414 , n72415 , n72416 , n72417 , n72418 , 
 n72419 , n72420 , n72421 , n72422 , n72423 , n72424 , n72425 , n72426 , n72427 , n72428 , 
 n72429 , n72430 , n72431 , n72432 , n72433 , n72434 , n72435 , n72436 , n72437 , n72438 , 
 n72439 , n72440 , n72441 , n72442 , n72443 , n72444 , n72445 , n72446 , n72447 , n72448 , 
 n72449 , n72450 , n72451 , n72452 , n72453 , n72454 , n72455 , n72456 , n72457 , n72458 , 
 n72459 , n72460 , n72461 , n72462 , n72463 , n72464 , n72465 , n72466 , n72467 , n72468 , 
 n72469 , n72470 , n72471 , n72472 , n72473 , n72474 , n72475 , n72476 , n72477 , n72478 , 
 n72479 , n72480 , n72481 , n72482 , n72483 , n72484 , n72485 , n72486 , n72487 , n72488 , 
 n72489 , n72490 , n72491 , n72492 , n72493 , n72494 , n72495 , n72496 , n72497 , n72498 , 
 n72499 , n72500 , n72501 , n72502 , n72503 , n72504 , n72505 , n72506 , n72507 , n72508 , 
 n72509 , n72510 , n72511 , n72512 , n72513 , n72514 , n72515 , n72516 , n72517 , n72518 , 
 n72519 , n72520 , n72521 , n72522 , n72523 , n72524 , n72525 , n72526 , n72527 , n72528 , 
 n72529 , n72530 , n72531 , n72532 , n72533 , n72534 , n72535 , n72536 , n72537 , n72538 , 
 n72539 , n72540 , n72541 , n72542 , n72543 , n72544 , n72545 , n72546 , n72547 , n72548 , 
 n72549 , n72550 , n72551 , n72552 , n72553 , n72554 , n72555 , n72556 , n72557 , n72558 , 
 n72559 , n72560 , n72561 , n72562 , n72563 , n72564 , n72565 , n72566 , n72567 , n72568 , 
 n72569 , n72570 , n72571 , n72572 , n72573 , n72574 , n72575 , n72576 , n72577 , n72578 , 
 n72579 , n72580 , n72581 , n72582 , n72583 , n72584 , n72585 , n72586 , n72587 , n72588 , 
 n72589 , n72590 , n72591 , n72592 , n72593 , n72594 , n72595 , n72596 , n72597 , n72598 , 
 n72599 , n72600 , n72601 , n72602 , n72603 , n72604 , n72605 , n72606 , n72607 , n72608 , 
 n72609 , n72610 , n72611 , n72612 , n72613 , n72614 , n72615 , n72616 , n72617 , n72618 , 
 n72619 , n72620 , n72621 , n72622 , n72623 , n72624 , n72625 , n72626 , n72627 , n72628 , 
 n72629 , n72630 , n72631 , n72632 , n72633 , n72634 , n72635 , n72636 , n72637 , n72638 , 
 n72639 , n72640 , n72641 , n72642 , n72643 , n72644 , n72645 , n72646 , n72647 , n72648 , 
 n72649 , n72650 , n72651 , n72652 , n72653 , n72654 , n72655 , n72656 , n72657 , n72658 , 
 n72659 , n72660 , n72661 , n72662 , n72663 , n72664 , n72665 , n72666 , n72667 , n72668 , 
 n72669 , n72670 , n72671 , n72672 , n72673 , n72674 , n72675 , n72676 , n72677 , n72678 , 
 n72679 , n72680 , n72681 , n72682 , n72683 , n72684 , n72685 , n72686 , n72687 , n72688 , 
 n72689 , n72690 , n72691 , n72692 , n72693 , n72694 , n72695 , n72696 , n72697 , n72698 , 
 n72699 , n72700 , n72701 , n72702 , n72703 , n72704 , n72705 , n72706 , n72707 , n72708 , 
 n72709 , n72710 , n72711 , n72712 , n72713 , n72714 , n72715 , n72716 , n72717 , n72718 , 
 n72719 , n72720 , n72721 , n72722 , n72723 , n72724 , n72725 , n72726 , n72727 , n72728 , 
 n72729 , n72730 , n72731 , n72732 , n72733 , n72734 , n72735 , n72736 , n72737 , n72738 , 
 n72739 , n72740 , n72741 , n72742 , n72743 , n72744 , n72745 , n72746 , n72747 , n72748 , 
 n72749 , n72750 , n72751 , n72752 , n72753 , n72754 , n72755 , n72756 , n72757 , n72758 , 
 n72759 , n72760 , n72761 , n72762 , n72763 , n72764 , n72765 , n72766 , n72767 , n72768 , 
 n72769 , n72770 , n72771 , n72772 , n72773 , n72774 , n72775 , n72776 , n72777 , n72778 , 
 n72779 , n72780 , n72781 , n72782 , n72783 , n72784 , n72785 , n72786 , n72787 , n72788 , 
 n72789 , n72790 , n72791 , n72792 , n72793 , n72794 , n72795 , n72796 , n72797 , n72798 , 
 n72799 , n72800 , n72801 , n72802 , n72803 , n72804 , n72805 , n72806 , n72807 , n72808 , 
 n72809 , n72810 , n72811 , n72812 , n72813 , n72814 , n72815 , n72816 , n72817 , n72818 , 
 n72819 , n72820 , n72821 , n72822 , n72823 , n72824 , n72825 , n72826 , n72827 , n72828 , 
 n72829 , n72830 , n72831 , n72832 , n72833 , n72834 , n72835 , n72836 , n72837 , n72838 , 
 n72839 , n72840 , n72841 , n72842 , n72843 , n72844 , n72845 , n72846 , n72847 , n72848 , 
 n72849 , n72850 , n72851 , n72852 , n72853 , n72854 , n72855 , n72856 , n72857 , n72858 , 
 n72859 , n72860 , n72861 , n72862 , n72863 , n72864 , n72865 , n72866 , n72867 , n72868 , 
 n72869 , n72870 , n72871 , n72872 , n72873 , n72874 , n72875 , n72876 , n72877 , n72878 , 
 n72879 , n72880 , n72881 , n72882 , n72883 , n72884 , n72885 , n72886 , n72887 , n72888 , 
 n72889 , n72890 , n72891 , n72892 , n72893 , n72894 , n72895 , n72896 , n72897 , n72898 , 
 n72899 , n72900 , n72901 , n72902 , n72903 , n72904 , n72905 , n72906 , n72907 , n72908 , 
 n72909 , n72910 , n72911 , n72912 , n72913 , n72914 , n72915 , n72916 , n72917 , n72918 , 
 n72919 , n72920 , n72921 , n72922 , n72923 , n72924 , n72925 , n72926 , n72927 , n72928 , 
 n72929 , n72930 , n72931 , n72932 , n72933 , n72934 , n72935 , n72936 , n72937 , n72938 , 
 n72939 , n72940 , n72941 , n72942 , n72943 , n72944 , n72945 , n72946 , n72947 , n72948 , 
 n72949 , n72950 , n72951 , n72952 , n72953 , n72954 , n72955 , n72956 , n72957 , n72958 , 
 n72959 , n72960 , n72961 , n72962 , n72963 , n72964 , n72965 , n72966 , n72967 , n72968 , 
 n72969 , n72970 , n72971 , n72972 , n72973 , n72974 , n72975 , n72976 , n72977 , n72978 , 
 n72979 , n72980 , n72981 , n72982 , n72983 , n72984 , n72985 , n72986 , n72987 , n72988 , 
 n72989 , n72990 , n72991 , n72992 , n72993 , n72994 , n72995 , n72996 , n72997 , n72998 , 
 n72999 , n73000 , n73001 , n73002 , n73003 , n73004 , n73005 , n73006 , n73007 , n73008 , 
 n73009 , n73010 , n73011 , n73012 , n73013 , n73014 , n73015 , n73016 , n73017 , n73018 , 
 n73019 , n73020 , n73021 , n73022 , n73023 , n73024 , n73025 , n73026 , n73027 , n73028 , 
 n73029 , n73030 , n73031 , n73032 , n73033 , n73034 , n73035 , n73036 , n73037 , n73038 , 
 n73039 , n73040 , n73041 , n73042 , n73043 , n73044 , n73045 , n73046 , n73047 , n73048 , 
 n73049 , n73050 , n73051 , n73052 , n73053 , n73054 , n73055 , n73056 , n73057 , n73058 , 
 n73059 , n73060 , n73061 , n73062 , n73063 , n73064 , n73065 , n73066 , n73067 , n73068 , 
 n73069 , n73070 , n73071 , n73072 , n73073 , n73074 , n73075 , n73076 , n73077 , n73078 , 
 n73079 , n73080 , n73081 , n73082 , n73083 , n73084 , n73085 , n73086 , n73087 , n73088 , 
 n73089 , n73090 , n73091 , n73092 , n73093 , n73094 , n73095 , n73096 , n73097 , n73098 , 
 n73099 , n73100 , n73101 , n73102 , n73103 , n73104 , n73105 , n73106 , n73107 , n73108 , 
 n73109 , n73110 , n73111 , n73112 , n73113 , n73114 , n73115 , n73116 , n73117 , n73118 , 
 n73119 , n73120 , n73121 , n73122 , n73123 , n73124 , n73125 , n73126 , n73127 , n73128 , 
 n73129 , n73130 , n73131 , n73132 , n73133 , n73134 , n73135 , n73136 , n73137 , n73138 , 
 n73139 , n73140 , n73141 , n73142 , n73143 , n73144 , n73145 , n73146 , n73147 , n73148 , 
 n73149 , n73150 , n73151 , n73152 , n73153 , n73154 , n73155 , n73156 , n73157 , n73158 , 
 n73159 , n73160 , n73161 , n73162 , n73163 , n73164 , n73165 , n73166 , n73167 , n73168 , 
 n73169 , n73170 , n73171 , n73172 , n73173 , n73174 , n73175 , n73176 , n73177 , n73178 , 
 n73179 , n73180 , n73181 , n73182 , n73183 , n73184 , n73185 , n73186 , n73187 , n73188 , 
 n73189 , n73190 , n73191 , n73192 , n73193 , n73194 , n73195 , n73196 , n73197 , n73198 , 
 n73199 , n73200 , n73201 , n73202 , n73203 , n73204 , n73205 , n73206 , n73207 , n73208 , 
 n73209 , n73210 , n73211 , n73212 , n73213 , n73214 , n73215 , n73216 , n73217 , n73218 , 
 n73219 , n73220 , n73221 , n73222 , n73223 , n73224 , n73225 , n73226 , n73227 , n73228 , 
 n73229 , n73230 , n73231 , n73232 , n73233 , n73234 , n73235 , n73236 , n73237 , n73238 , 
 n73239 , n73240 , n73241 , n73242 , n73243 , n73244 , n73245 , n73246 , n73247 , n73248 , 
 n73249 , n73250 , n73251 , n73252 , n73253 , n73254 , n73255 , n73256 , n73257 , n73258 , 
 n73259 , n73260 , n73261 , n73262 , n73263 , n73264 , n73265 , n73266 , n73267 , n73268 , 
 n73269 , n73270 , n73271 , n73272 , n73273 , n73274 , n73275 , n73276 , n73277 , n73278 , 
 n73279 , n73280 , n73281 , n73282 , n73283 , n73284 , n73285 , n73286 , n73287 , n73288 , 
 n73289 , n73290 , n73291 , n73292 , n73293 , n73294 , n73295 , n73296 , n73297 , n73298 , 
 n73299 , n73300 , n73301 , n73302 , n73303 , n73304 , n73305 , n73306 , n73307 , n73308 , 
 n73309 , n73310 , n73311 , n73312 , n73313 , n73314 , n73315 , n73316 , n73317 , n73318 , 
 n73319 , n73320 , n73321 , n73322 , n73323 , n73324 , n73325 , n73326 , n73327 , n73328 , 
 n73329 , n73330 , n73331 , n73332 , n73333 , n73334 , n73335 , n73336 , n73337 , n73338 , 
 n73339 , n73340 , n73341 , n73342 , n73343 , n73344 , n73345 , n73346 , n73347 , n73348 , 
 n73349 , n73350 , n73351 , n73352 , n73353 , n73354 , n73355 , n73356 , n73357 , n73358 , 
 n73359 , n73360 , n73361 , n73362 , n73363 , n73364 , n73365 , n73366 , n73367 , n73368 , 
 n73369 , n73370 , n73371 , n73372 , n73373 , n73374 , n73375 , n73376 , n73377 , n73378 , 
 n73379 , n73380 , n73381 , n73382 , n73383 , n73384 , n73385 , n73386 , n73387 , n73388 , 
 n73389 , n73390 , n73391 , n73392 , n73393 , n73394 , n73395 , n73396 , n73397 , n73398 , 
 n73399 , n73400 , n73401 , n73402 , n73403 , n73404 , n73405 , n73406 , n73407 , n73408 , 
 n73409 , n73410 , n73411 , n73412 , n73413 , n73414 , n73415 , n73416 , n73417 , n73418 , 
 n73419 , n73420 , n73421 , n73422 , n73423 , n73424 , n73425 , n73426 , n73427 , n73428 , 
 n73429 , n73430 , n73431 , n73432 , n73433 , n73434 , n73435 , n73436 , n73437 , n73438 , 
 n73439 , n73440 , n73441 , n73442 , n73443 , n73444 , n73445 , n73446 , n73447 , n73448 , 
 n73449 , n73450 , n73451 , n73452 , n73453 , n73454 , n73455 , n73456 , n73457 , n73458 , 
 n73459 , n73460 , n73461 , n73462 , n73463 , n73464 , n73465 , n73466 , n73467 , n73468 , 
 n73469 , n73470 , n73471 , n73472 , n73473 , n73474 , n73475 , n73476 , n73477 , n73478 , 
 n73479 , n73480 , n73481 , n73482 , n73483 , n73484 , n73485 , n73486 , n73487 , n73488 , 
 n73489 , n73490 , n73491 , n73492 , n73493 , n73494 , n73495 , n73496 , n73497 , n73498 , 
 n73499 , n73500 , n73501 , n73502 , n73503 , n73504 , n73505 , n73506 , n73507 , n73508 , 
 n73509 , n73510 , n73511 , n73512 , n73513 , n73514 , n73515 , n73516 , n73517 , n73518 , 
 n73519 , n73520 , n73521 , n73522 , n73523 , n73524 , n73525 , n73526 , n73527 , n73528 , 
 n73529 , n73530 , n73531 , n73532 , n73533 , n73534 , n73535 , n73536 , n73537 , n73538 , 
 n73539 , n73540 , n73541 , n73542 , n73543 , n73544 , n73545 , n73546 , n73547 , n73548 , 
 n73549 , n73550 , n73551 , n73552 , n73553 , n73554 , n73555 , n73556 , n73557 , n73558 , 
 n73559 , n73560 , n73561 , n73562 , n73563 , n73564 , n73565 , n73566 , n73567 , n73568 , 
 n73569 , n73570 , n73571 , n73572 , n73573 , n73574 , n73575 , n73576 , n73577 , n73578 , 
 n73579 , n73580 , n73581 , n73582 , n73583 , n73584 , n73585 , n73586 , n73587 , n73588 , 
 n73589 , n73590 , n73591 , n73592 , n73593 , n73594 , n73595 , n73596 , n73597 , n73598 , 
 n73599 , n73600 , n73601 , n73602 , n73603 , n73604 , n73605 , n73606 , n73607 , n73608 , 
 n73609 , n73610 , n73611 , n73612 , n73613 , n73614 , n73615 , n73616 , n73617 , n73618 , 
 n73619 , n73620 , n73621 , n73622 , n73623 , n73624 , n73625 , n73626 , n73627 , n73628 , 
 n73629 , n73630 , n73631 , n73632 , n73633 , n73634 , n73635 , n73636 , n73637 , n73638 , 
 n73639 , n73640 , n73641 , n73642 , n73643 , n73644 , n73645 , n73646 , n73647 , n73648 , 
 n73649 , n73650 , n73651 , n73652 , n73653 , n73654 , n73655 , n73656 , n73657 , n73658 , 
 n73659 , n73660 , n73661 , n73662 , n73663 , n73664 , n73665 , n73666 , n73667 , n73668 , 
 n73669 , n73670 , n73671 , n73672 , n73673 , n73674 , n73675 , n73676 , n73677 , n73678 , 
 n73679 , n73680 , n73681 , n73682 , n73683 , n73684 , n73685 , n73686 , n73687 , n73688 , 
 n73689 , n73690 , n73691 , n73692 , n73693 , n73694 , n73695 , n73696 , n73697 , n73698 , 
 n73699 , n73700 , n73701 , n73702 , n73703 , n73704 , n73705 , n73706 , n73707 , n73708 , 
 n73709 , n73710 , n73711 , n73712 , n73713 , n73714 , n73715 , n73716 , n73717 , n73718 , 
 n73719 , n73720 , n73721 , n73722 , n73723 , n73724 , n73725 , n73726 , n73727 , n73728 , 
 n73729 , n73730 , n73731 , n73732 , n73733 , n73734 , n73735 , n73736 , n73737 , n73738 , 
 n73739 , n73740 , n73741 , n73742 , n73743 , n73744 , n73745 , n73746 , n73747 , n73748 , 
 n73749 , n73750 , n73751 , n73752 , n73753 , n73754 , n73755 , n73756 , n73757 , n73758 , 
 n73759 , n73760 , n73761 , n73762 , n73763 , n73764 , n73765 , n73766 , n73767 , n73768 , 
 n73769 , n73770 , n73771 , n73772 , n73773 , n73774 , n73775 , n73776 , n73777 , n73778 , 
 n73779 , n73780 , n73781 , n73782 , n73783 , n73784 , n73785 , n73786 , n73787 , n73788 , 
 n73789 , n73790 , n73791 , n73792 , n73793 , n73794 , n73795 , n73796 , n73797 , n73798 , 
 n73799 , n73800 , n73801 , n73802 , n73803 , n73804 , n73805 , n73806 , n73807 , n73808 , 
 n73809 , n73810 , n73811 , n73812 , n73813 , n73814 , n73815 , n73816 , n73817 , n73818 , 
 n73819 , n73820 , n73821 , n73822 , n73823 , n73824 , n73825 , n73826 , n73827 , n73828 , 
 n73829 , n73830 , n73831 , n73832 , n73833 , n73834 , n73835 , n73836 , n73837 , n73838 , 
 n73839 , n73840 , n73841 , n73842 , n73843 , n73844 , n73845 , n73846 , n73847 , n73848 , 
 n73849 , n73850 , n73851 , n73852 , n73853 , n73854 , n73855 , n73856 , n73857 , n73858 , 
 n73859 , n73860 , n73861 , n73862 , n73863 , n73864 , n73865 , n73866 , n73867 , n73868 , 
 n73869 , n73870 , n73871 , n73872 , n73873 , n73874 , n73875 , n73876 , n73877 , n73878 , 
 n73879 , n73880 , n73881 , n73882 , n73883 , n73884 , n73885 , n73886 , n73887 , n73888 , 
 n73889 , n73890 , n73891 , n73892 , n73893 , n73894 , n73895 , n73896 , n73897 , n73898 , 
 n73899 , n73900 , n73901 , n73902 , n73903 , n73904 , n73905 , n73906 , n73907 , n73908 , 
 n73909 , n73910 , n73911 , n73912 , n73913 , n73914 , n73915 , n73916 , n73917 , n73918 , 
 n73919 , n73920 , n73921 , n73922 , n73923 , n73924 , n73925 , n73926 , n73927 , n73928 , 
 n73929 , n73930 , n73931 , n73932 , n73933 , n73934 , n73935 , n73936 , n73937 , n73938 , 
 n73939 , n73940 , n73941 , n73942 , n73943 , n73944 , n73945 , n73946 , n73947 , n73948 , 
 n73949 , n73950 , n73951 , n73952 , n73953 , n73954 , n73955 , n73956 , n73957 , n73958 , 
 n73959 , n73960 , n73961 , n73962 , n73963 , n73964 , n73965 , n73966 , n73967 , n73968 , 
 n73969 , n73970 , n73971 , n73972 , n73973 , n73974 , n73975 , n73976 , n73977 , n73978 , 
 n73979 , n73980 , n73981 , n73982 , n73983 , n73984 , n73985 , n73986 , n73987 , n73988 , 
 n73989 , n73990 , n73991 , n73992 , n73993 , n73994 , n73995 , n73996 , n73997 , n73998 , 
 n73999 , n74000 , n74001 , n74002 , n74003 , n74004 , n74005 , n74006 , n74007 , n74008 , 
 n74009 , n74010 , n74011 , n74012 , n74013 , n74014 , n74015 , n74016 , n74017 , n74018 , 
 n74019 , n74020 , n74021 , n74022 , n74023 , n74024 , n74025 , n74026 , n74027 , n74028 , 
 n74029 , n74030 , n74031 , n74032 , n74033 , n74034 , n74035 , n74036 , n74037 , n74038 , 
 n74039 , n74040 , n74041 , n74042 , n74043 , n74044 , n74045 , n74046 , n74047 , n74048 , 
 n74049 , n74050 , n74051 , n74052 , n74053 , n74054 , n74055 , n74056 , n74057 , n74058 , 
 n74059 , n74060 , n74061 , n74062 , n74063 , n74064 , n74065 , n74066 , n74067 , n74068 , 
 n74069 , n74070 , n74071 , n74072 , n74073 , n74074 , n74075 , n74076 , n74077 , n74078 , 
 n74079 , n74080 , n74081 , n74082 , n74083 , n74084 , n74085 , n74086 , n74087 , n74088 , 
 n74089 , n74090 , n74091 , n74092 , n74093 , n74094 , n74095 , n74096 , n74097 , n74098 , 
 n74099 , n74100 , n74101 , n74102 , n74103 , n74104 , n74105 , n74106 , n74107 , n74108 , 
 n74109 , n74110 , n74111 , n74112 , n74113 , n74114 , n74115 , n74116 , n74117 , n74118 , 
 n74119 , n74120 , n74121 , n74122 , n74123 , n74124 , n74125 , n74126 , n74127 , n74128 , 
 n74129 , n74130 , n74131 , n74132 , n74133 , n74134 , n74135 , n74136 , n74137 , n74138 , 
 n74139 , n74140 , n74141 , n74142 , n74143 , n74144 , n74145 , n74146 , n74147 , n74148 , 
 n74149 , n74150 , n74151 , n74152 , n74153 , n74154 , n74155 , n74156 , n74157 , n74158 , 
 n74159 , n74160 , n74161 , n74162 , n74163 , n74164 , n74165 , n74166 , n74167 , n74168 , 
 n74169 , n74170 , n74171 , n74172 , n74173 , n74174 , n74175 , n74176 , n74177 , n74178 , 
 n74179 , n74180 , n74181 , n74182 , n74183 , n74184 , n74185 , n74186 , n74187 , n74188 , 
 n74189 , n74190 , n74191 , n74192 , n74193 , n74194 , n74195 , n74196 , n74197 , n74198 , 
 n74199 , n74200 , n74201 , n74202 , n74203 , n74204 , n74205 , n74206 , n74207 , n74208 , 
 n74209 , n74210 , n74211 , n74212 , n74213 , n74214 , n74215 , n74216 , n74217 , n74218 , 
 n74219 , n74220 , n74221 , n74222 , n74223 , n74224 , n74225 , n74226 , n74227 , n74228 , 
 n74229 , n74230 , n74231 , n74232 , n74233 , n74234 , n74235 , n74236 , n74237 , n74238 , 
 n74239 , n74240 , n74241 , n74242 , n74243 , n74244 , n74245 , n74246 , n74247 , n74248 , 
 n74249 , n74250 , n74251 , n74252 , n74253 , n74254 , n74255 , n74256 , n74257 , n74258 , 
 n74259 , n74260 , n74261 , n74262 , n74263 , n74264 , n74265 , n74266 , n74267 , n74268 , 
 n74269 , n74270 , n74271 , n74272 , n74273 , n74274 , n74275 , n74276 , n74277 , n74278 , 
 n74279 , n74280 , n74281 , n74282 , n74283 , n74284 , n74285 , n74286 , n74287 , n74288 , 
 n74289 , n74290 , n74291 , n74292 , n74293 , n74294 , n74295 , n74296 , n74297 , n74298 , 
 n74299 , n74300 , n74301 , n74302 , n74303 , n74304 , n74305 , n74306 , n74307 , n74308 , 
 n74309 , n74310 , n74311 , n74312 , n74313 , n74314 , n74315 , n74316 , n74317 , n74318 , 
 n74319 , n74320 , n74321 , n74322 , n74323 , n74324 , n74325 , n74326 , n74327 , n74328 , 
 n74329 , n74330 , n74331 , n74332 , n74333 , n74334 , n74335 , n74336 , n74337 , n74338 , 
 n74339 , n74340 , n74341 , n74342 , n74343 , n74344 , n74345 , n74346 , n74347 , n74348 , 
 n74349 , n74350 , n74351 , n74352 , n74353 , n74354 , n74355 , n74356 , n74357 , n74358 , 
 n74359 , n74360 , n74361 , n74362 , n74363 , n74364 , n74365 , n74366 , n74367 , n74368 , 
 n74369 , n74370 , n74371 , n74372 , n74373 , n74374 , n74375 , n74376 , n74377 , n74378 , 
 n74379 , n74380 , n74381 , n74382 , n74383 , n74384 , n74385 , n74386 , n74387 , n74388 , 
 n74389 , n74390 , n74391 , n74392 , n74393 , n74394 , n74395 , n74396 , n74397 , n74398 , 
 n74399 , n74400 , n74401 , n74402 , n74403 , n74404 , n74405 , n74406 , n74407 , n74408 , 
 n74409 , n74410 , n74411 , n74412 , n74413 , n74414 , n74415 , n74416 , n74417 , n74418 , 
 n74419 , n74420 , n74421 , n74422 , n74423 , n74424 , n74425 , n74426 , n74427 , n74428 , 
 n74429 , n74430 , n74431 , n74432 , n74433 , n74434 , n74435 , n74436 , n74437 , n74438 , 
 n74439 , n74440 , n74441 , n74442 , n74443 , n74444 , n74445 , n74446 , n74447 , n74448 , 
 n74449 , n74450 , n74451 , n74452 , n74453 , n74454 , n74455 , n74456 , n74457 , n74458 , 
 n74459 , n74460 , n74461 , n74462 , n74463 , n74464 , n74465 , n74466 , n74467 , n74468 , 
 n74469 , n74470 , n74471 , n74472 , n74473 , n74474 , n74475 , n74476 , n74477 , n74478 , 
 n74479 , n74480 , n74481 , n74482 , n74483 , n74484 , n74485 , n74486 , n74487 , n74488 , 
 n74489 , n74490 , n74491 , n74492 , n74493 , n74494 , n74495 , n74496 , n74497 , n74498 , 
 n74499 , n74500 , n74501 , n74502 , n74503 , n74504 , n74505 , n74506 , n74507 , n74508 , 
 n74509 , n74510 , n74511 , n74512 , n74513 , n74514 , n74515 , n74516 , n74517 , n74518 , 
 n74519 , n74520 , n74521 , n74522 , n74523 , n74524 , n74525 , n74526 , n74527 , n74528 , 
 n74529 , n74530 , n74531 , n74532 , n74533 , n74534 , n74535 , n74536 , n74537 , n74538 , 
 n74539 , n74540 , n74541 , n74542 , n74543 , n74544 , n74545 , n74546 , n74547 , n74548 , 
 n74549 , n74550 , n74551 , n74552 , n74553 , n74554 , n74555 , n74556 , n74557 , n74558 , 
 n74559 , n74560 , n74561 , n74562 , n74563 , n74564 , n74565 , n74566 , n74567 , n74568 , 
 n74569 , n74570 , n74571 , n74572 , n74573 , n74574 , n74575 , n74576 , n74577 , n74578 , 
 n74579 , n74580 , n74581 , n74582 , n74583 , n74584 , n74585 , n74586 , n74587 , n74588 , 
 n74589 , n74590 , n74591 , n74592 , n74593 , n74594 , n74595 , n74596 , n74597 , n74598 , 
 n74599 , n74600 , n74601 , n74602 , n74603 , n74604 , n74605 , n74606 , n74607 , n74608 , 
 n74609 , n74610 , n74611 , n74612 , n74613 , n74614 , n74615 , n74616 , n74617 , n74618 , 
 n74619 , n74620 , n74621 , n74622 , n74623 , n74624 , n74625 , n74626 , n74627 , n74628 , 
 n74629 , n74630 , n74631 , n74632 , n74633 , n74634 , n74635 , n74636 , n74637 , n74638 , 
 n74639 , n74640 , n74641 , n74642 , n74643 , n74644 , n74645 , n74646 , n74647 , n74648 , 
 n74649 , n74650 , n74651 , n74652 , n74653 , n74654 , n74655 , n74656 , n74657 , n74658 , 
 n74659 , n74660 , n74661 , n74662 , n74663 , n74664 , n74665 , n74666 , n74667 , n74668 , 
 n74669 , n74670 , n74671 , n74672 , n74673 , n74674 , n74675 , n74676 , n74677 , n74678 , 
 n74679 , n74680 , n74681 , n74682 , n74683 , n74684 , n74685 , n74686 , n74687 , n74688 , 
 n74689 , n74690 , n74691 , n74692 , n74693 , n74694 , n74695 , n74696 , n74697 , n74698 , 
 n74699 , n74700 , n74701 , n74702 , n74703 , n74704 , n74705 , n74706 , n74707 , n74708 , 
 n74709 , n74710 , n74711 , n74712 , n74713 , n74714 , n74715 , n74716 , n74717 , n74718 , 
 n74719 , n74720 , n74721 , n74722 , n74723 , n74724 , n74725 , n74726 , n74727 , n74728 , 
 n74729 , n74730 , n74731 , n74732 , n74733 , n74734 , n74735 , n74736 , n74737 , n74738 , 
 n74739 , n74740 , n74741 , n74742 , n74743 , n74744 , n74745 , n74746 , n74747 , n74748 , 
 n74749 , n74750 , n74751 , n74752 , n74753 , n74754 , n74755 , n74756 , n74757 , n74758 , 
 n74759 , n74760 , n74761 , n74762 , n74763 , n74764 , n74765 , n74766 , n74767 , n74768 , 
 n74769 , n74770 , n74771 , n74772 , n74773 , n74774 , n74775 , n74776 , n74777 , n74778 , 
 n74779 , n74780 , n74781 , n74782 , n74783 , n74784 , n74785 , n74786 , n74787 , n74788 , 
 n74789 , n74790 , n74791 , n74792 , n74793 , n74794 , n74795 , n74796 , n74797 , n74798 , 
 n74799 , n74800 , n74801 , n74802 , n74803 , n74804 , n74805 , n74806 , n74807 , n74808 , 
 n74809 , n74810 , n74811 , n74812 , n74813 , n74814 , n74815 , n74816 , n74817 , n74818 , 
 n74819 , n74820 , n74821 , n74822 , n74823 , n74824 , n74825 , n74826 , n74827 , n74828 , 
 n74829 , n74830 , n74831 , n74832 , n74833 , n74834 , n74835 , n74836 , n74837 , n74838 , 
 n74839 , n74840 , n74841 , n74842 , n74843 , n74844 , n74845 , n74846 , n74847 , n74848 , 
 n74849 , n74850 , n74851 , n74852 , n74853 , n74854 , n74855 , n74856 , n74857 , n74858 , 
 n74859 , n74860 , n74861 , n74862 , n74863 , n74864 , n74865 , n74866 , n74867 , n74868 , 
 n74869 , n74870 , n74871 , n74872 , n74873 , n74874 , n74875 , n74876 , n74877 , n74878 , 
 n74879 , n74880 , n74881 , n74882 , n74883 , n74884 , n74885 , n74886 , n74887 , n74888 , 
 n74889 , n74890 , n74891 , n74892 , n74893 , n74894 , n74895 , n74896 , n74897 , n74898 , 
 n74899 , n74900 , n74901 , n74902 , n74903 , n74904 , n74905 , n74906 , n74907 , n74908 , 
 n74909 , n74910 , n74911 , n74912 , n74913 , n74914 , n74915 , n74916 , n74917 , n74918 , 
 n74919 , n74920 , n74921 , n74922 , n74923 , n74924 , n74925 , n74926 , n74927 , n74928 , 
 n74929 , n74930 , n74931 , n74932 , n74933 , n74934 , n74935 , n74936 , n74937 , n74938 , 
 n74939 , n74940 , n74941 , n74942 , n74943 , n74944 , n74945 , n74946 , n74947 , n74948 , 
 n74949 , n74950 , n74951 , n74952 , n74953 , n74954 , n74955 , n74956 , n74957 , n74958 , 
 n74959 , n74960 , n74961 , n74962 , n74963 , n74964 , n74965 , n74966 , n74967 , n74968 , 
 n74969 , n74970 , n74971 , n74972 , n74973 , n74974 , n74975 , n74976 , n74977 , n74978 , 
 n74979 , n74980 , n74981 , n74982 , n74983 , n74984 , n74985 , n74986 , n74987 , n74988 , 
 n74989 , n74990 , n74991 , n74992 , n74993 , n74994 , n74995 , n74996 , n74997 , n74998 , 
 n74999 , n75000 , n75001 , n75002 , n75003 , n75004 , n75005 , n75006 , n75007 , n75008 , 
 n75009 , n75010 , n75011 , n75012 , n75013 , n75014 , n75015 , n75016 , n75017 , n75018 , 
 n75019 , n75020 , n75021 , n75022 , n75023 , n75024 , n75025 , n75026 , n75027 , n75028 , 
 n75029 , n75030 , n75031 , n75032 , n75033 , n75034 , n75035 , n75036 , n75037 , n75038 , 
 n75039 , n75040 , n75041 , n75042 , n75043 , n75044 , n75045 , n75046 , n75047 , n75048 , 
 n75049 , n75050 , n75051 , n75052 , n75053 , n75054 , n75055 , n75056 , n75057 , n75058 , 
 n75059 , n75060 , n75061 , n75062 , n75063 , n75064 , n75065 , n75066 , n75067 , n75068 , 
 n75069 , n75070 , n75071 , n75072 , n75073 , n75074 , n75075 , n75076 , n75077 , n75078 , 
 n75079 , n75080 , n75081 , n75082 , n75083 , n75084 , n75085 , n75086 , n75087 , n75088 , 
 n75089 , n75090 , n75091 , n75092 , n75093 , n75094 , n75095 , n75096 , n75097 , n75098 , 
 n75099 , n75100 , n75101 , n75102 , n75103 , n75104 , n75105 , n75106 , n75107 , n75108 , 
 n75109 , n75110 , n75111 , n75112 , n75113 , n75114 , n75115 , n75116 , n75117 , n75118 , 
 n75119 , n75120 , n75121 , n75122 , n75123 , n75124 , n75125 , n75126 , n75127 , n75128 , 
 n75129 , n75130 , n75131 , n75132 , n75133 , n75134 , n75135 , n75136 , n75137 , n75138 , 
 n75139 , n75140 , n75141 , n75142 , n75143 , n75144 , n75145 , n75146 , n75147 , n75148 , 
 n75149 , n75150 , n75151 , n75152 , n75153 , n75154 , n75155 , n75156 , n75157 , n75158 , 
 n75159 , n75160 , n75161 , n75162 , n75163 , n75164 , n75165 , n75166 , n75167 , n75168 , 
 n75169 , n75170 , n75171 , n75172 , n75173 , n75174 , n75175 , n75176 , n75177 , n75178 , 
 n75179 , n75180 , n75181 , n75182 , n75183 , n75184 , n75185 , n75186 , n75187 , n75188 , 
 n75189 , n75190 , n75191 , n75192 , n75193 , n75194 , n75195 , n75196 , n75197 , n75198 , 
 n75199 , n75200 , n75201 , n75202 , n75203 , n75204 , n75205 , n75206 , n75207 , n75208 , 
 n75209 , n75210 , n75211 , n75212 , n75213 , n75214 , n75215 , n75216 , n75217 , n75218 , 
 n75219 , n75220 , n75221 , n75222 , n75223 , n75224 , n75225 , n75226 , n75227 , n75228 , 
 n75229 , n75230 , n75231 , n75232 , n75233 , n75234 , n75235 , n75236 , n75237 , n75238 , 
 n75239 , n75240 , n75241 , n75242 , n75243 , n75244 , n75245 , n75246 , n75247 , n75248 , 
 n75249 , n75250 , n75251 , n75252 , n75253 , n75254 , n75255 , n75256 , n75257 , n75258 , 
 n75259 , n75260 , n75261 , n75262 , n75263 , n75264 , n75265 , n75266 , n75267 , n75268 , 
 n75269 , n75270 , n75271 , n75272 , n75273 , n75274 , n75275 , n75276 , n75277 , n75278 , 
 n75279 , n75280 , n75281 , n75282 , n75283 , n75284 , n75285 , n75286 , n75287 , n75288 , 
 n75289 , n75290 , n75291 , n75292 , n75293 , n75294 , n75295 , n75296 , n75297 , n75298 , 
 n75299 , n75300 , n75301 , n75302 , n75303 , n75304 , n75305 , n75306 , n75307 , n75308 , 
 n75309 , n75310 , n75311 , n75312 , n75313 , n75314 , n75315 , n75316 , n75317 , n75318 , 
 n75319 , n75320 , n75321 , n75322 , n75323 , n75324 , n75325 , n75326 , n75327 , n75328 , 
 n75329 , n75330 , n75331 , n75332 , n75333 , n75334 , n75335 , n75336 , n75337 , n75338 , 
 n75339 , n75340 , n75341 , n75342 , n75343 , n75344 , n75345 , n75346 , n75347 , n75348 , 
 n75349 , n75350 , n75351 , n75352 , n75353 , n75354 , n75355 , n75356 , n75357 , n75358 , 
 n75359 , n75360 , n75361 , n75362 , n75363 , n75364 , n75365 , n75366 , n75367 , n75368 , 
 n75369 , n75370 , n75371 , n75372 , n75373 , n75374 , n75375 , n75376 , n75377 , n75378 , 
 n75379 , n75380 , n75381 , n75382 , n75383 , n75384 , n75385 , n75386 , n75387 , n75388 , 
 n75389 , n75390 , n75391 , n75392 , n75393 , n75394 , n75395 , n75396 , n75397 , n75398 , 
 n75399 , n75400 , n75401 , n75402 , n75403 , n75404 , n75405 , n75406 , n75407 , n75408 , 
 n75409 , n75410 , n75411 , n75412 , n75413 , n75414 , n75415 , n75416 , n75417 , n75418 , 
 n75419 , n75420 , n75421 , n75422 , n75423 , n75424 , n75425 , n75426 , n75427 , n75428 , 
 n75429 , n75430 , n75431 , n75432 , n75433 , n75434 , n75435 , n75436 , n75437 , n75438 , 
 n75439 , n75440 , n75441 , n75442 , n75443 , n75444 , n75445 , n75446 , n75447 , n75448 , 
 n75449 , n75450 , n75451 , n75452 , n75453 , n75454 , n75455 , n75456 , n75457 , n75458 , 
 n75459 , n75460 , n75461 , n75462 , n75463 , n75464 , n75465 , n75466 , n75467 , n75468 , 
 n75469 , n75470 , n75471 , n75472 , n75473 , n75474 , n75475 , n75476 , n75477 , n75478 , 
 n75479 , n75480 , n75481 , n75482 , n75483 , n75484 , n75485 , n75486 , n75487 , n75488 , 
 n75489 , n75490 , n75491 , n75492 , n75493 , n75494 , n75495 , n75496 , n75497 , n75498 , 
 n75499 , n75500 , n75501 , n75502 , n75503 , n75504 , n75505 , n75506 , n75507 , n75508 , 
 n75509 , n75510 , n75511 , n75512 , n75513 , n75514 , n75515 , n75516 , n75517 , n75518 , 
 n75519 , n75520 , n75521 , n75522 , n75523 , n75524 , n75525 , n75526 , n75527 , n75528 , 
 n75529 , n75530 , n75531 , n75532 , n75533 , n75534 , n75535 , n75536 , n75537 , n75538 , 
 n75539 , n75540 , n75541 , n75542 , n75543 , n75544 , n75545 , n75546 , n75547 , n75548 , 
 n75549 , n75550 , n75551 , n75552 , n75553 , n75554 , n75555 , n75556 , n75557 , n75558 , 
 n75559 , n75560 , n75561 , n75562 , n75563 , n75564 , n75565 , n75566 , n75567 , n75568 , 
 n75569 , n75570 , n75571 , n75572 , n75573 , n75574 , n75575 , n75576 , n75577 , n75578 , 
 n75579 , n75580 , n75581 , n75582 , n75583 , n75584 , n75585 , n75586 , n75587 , n75588 , 
 n75589 , n75590 , n75591 , n75592 , n75593 , n75594 , n75595 , n75596 , n75597 , n75598 , 
 n75599 , n75600 , n75601 , n75602 , n75603 , n75604 , n75605 , n75606 , n75607 , n75608 , 
 n75609 , n75610 , n75611 , n75612 , n75613 , n75614 , n75615 , n75616 , n75617 , n75618 , 
 n75619 , n75620 , n75621 , n75622 , n75623 , n75624 , n75625 , n75626 , n75627 , n75628 , 
 n75629 , n75630 , n75631 , n75632 , n75633 , n75634 , n75635 , n75636 , n75637 , n75638 , 
 n75639 , n75640 , n75641 , n75642 , n75643 , n75644 , n75645 , n75646 , n75647 , n75648 , 
 n75649 , n75650 , n75651 , n75652 , n75653 , n75654 , n75655 , n75656 , n75657 , n75658 , 
 n75659 , n75660 , n75661 , n75662 , n75663 , n75664 , n75665 , n75666 , n75667 , n75668 , 
 n75669 , n75670 , n75671 , n75672 , n75673 , n75674 , n75675 , n75676 , n75677 , n75678 , 
 n75679 , n75680 , n75681 , n75682 , n75683 , n75684 , n75685 , n75686 , n75687 , n75688 , 
 n75689 , n75690 , n75691 , n75692 , n75693 , n75694 , n75695 , n75696 , n75697 , n75698 , 
 n75699 , n75700 , n75701 , n75702 , n75703 , n75704 , n75705 , n75706 , n75707 , n75708 , 
 n75709 , n75710 , n75711 , n75712 , n75713 , n75714 , n75715 , n75716 , n75717 , n75718 , 
 n75719 , n75720 , n75721 , n75722 , n75723 , n75724 , n75725 , n75726 , n75727 , n75728 , 
 n75729 , n75730 , n75731 , n75732 , n75733 , n75734 , n75735 , n75736 , n75737 , n75738 , 
 n75739 , n75740 , n75741 , n75742 , n75743 , n75744 , n75745 , n75746 , n75747 , n75748 , 
 n75749 , n75750 , n75751 , n75752 , n75753 , n75754 , n75755 , n75756 , n75757 , n75758 , 
 n75759 , n75760 , n75761 , n75762 , n75763 , n75764 , n75765 , n75766 , n75767 , n75768 , 
 n75769 , n75770 , n75771 , n75772 , n75773 , n75774 , n75775 , n75776 , n75777 , n75778 , 
 n75779 , n75780 , n75781 , n75782 , n75783 , n75784 , n75785 , n75786 , n75787 , n75788 , 
 n75789 , n75790 , n75791 , n75792 , n75793 , n75794 , n75795 , n75796 , n75797 , n75798 , 
 n75799 , n75800 , n75801 , n75802 , n75803 , n75804 , n75805 , n75806 , n75807 , n75808 , 
 n75809 , n75810 , n75811 , n75812 , n75813 , n75814 , n75815 , n75816 , n75817 , n75818 , 
 n75819 , n75820 , n75821 , n75822 , n75823 , n75824 , n75825 , n75826 , n75827 , n75828 , 
 n75829 , n75830 , n75831 , n75832 , n75833 , n75834 , n75835 , n75836 , n75837 , n75838 , 
 n75839 , n75840 , n75841 , n75842 , n75843 , n75844 , n75845 , n75846 , n75847 , n75848 , 
 n75849 , n75850 , n75851 , n75852 , n75853 , n75854 , n75855 , n75856 , n75857 , n75858 , 
 n75859 , n75860 , n75861 , n75862 , n75863 , n75864 , n75865 , n75866 , n75867 , n75868 , 
 n75869 , n75870 , n75871 , n75872 , n75873 , n75874 , n75875 , n75876 , n75877 , n75878 , 
 n75879 , n75880 , n75881 , n75882 , n75883 , n75884 , n75885 , n75886 , n75887 , n75888 , 
 n75889 , n75890 , n75891 , n75892 , n75893 , n75894 , n75895 , n75896 , n75897 , n75898 , 
 n75899 , n75900 , n75901 , n75902 , n75903 , n75904 , n75905 , n75906 , n75907 , n75908 , 
 n75909 , n75910 , n75911 , n75912 , n75913 , n75914 , n75915 , n75916 , n75917 , n75918 , 
 n75919 , n75920 , n75921 , n75922 , n75923 , n75924 , n75925 , n75926 , n75927 , n75928 , 
 n75929 , n75930 , n75931 , n75932 , n75933 , n75934 , n75935 , n75936 , n75937 , n75938 , 
 n75939 , n75940 , n75941 , n75942 , n75943 , n75944 , n75945 , n75946 , n75947 , n75948 , 
 n75949 , n75950 , n75951 , n75952 , n75953 , n75954 , n75955 , n75956 , n75957 , n75958 , 
 n75959 , n75960 , n75961 , n75962 , n75963 , n75964 , n75965 , n75966 , n75967 , n75968 , 
 n75969 , n75970 , n75971 , n75972 , n75973 , n75974 , n75975 , n75976 , n75977 , n75978 , 
 n75979 , n75980 , n75981 , n75982 , n75983 , n75984 , n75985 , n75986 , n75987 , n75988 , 
 n75989 , n75990 , n75991 , n75992 , n75993 , n75994 , n75995 , n75996 , n75997 , n75998 , 
 n75999 , n76000 , n76001 , n76002 , n76003 , n76004 , n76005 , n76006 , n76007 , n76008 , 
 n76009 , n76010 , n76011 , n76012 , n76013 , n76014 , n76015 , n76016 , n76017 , n76018 , 
 n76019 , n76020 , n76021 , n76022 , n76023 , n76024 , n76025 , n76026 , n76027 , n76028 , 
 n76029 , n76030 , n76031 , n76032 , n76033 , n76034 , n76035 , n76036 , n76037 , n76038 , 
 n76039 , n76040 , n76041 , n76042 , n76043 , n76044 , n76045 , n76046 , n76047 , n76048 , 
 n76049 , n76050 , n76051 , n76052 , n76053 , n76054 , n76055 , n76056 , n76057 , n76058 , 
 n76059 , n76060 , n76061 , n76062 , n76063 , n76064 , n76065 , n76066 , n76067 , n76068 , 
 n76069 , n76070 , n76071 , n76072 , n76073 , n76074 , n76075 , n76076 , n76077 , n76078 , 
 n76079 , n76080 , n76081 , n76082 , n76083 , n76084 , n76085 , n76086 , n76087 , n76088 , 
 n76089 , n76090 , n76091 , n76092 , n76093 , n76094 , n76095 , n76096 , n76097 , n76098 , 
 n76099 , n76100 , n76101 , n76102 , n76103 , n76104 , n76105 , n76106 , n76107 , n76108 , 
 n76109 , n76110 , n76111 , n76112 , n76113 , n76114 , n76115 , n76116 , n76117 , n76118 , 
 n76119 , n76120 , n76121 , n76122 , n76123 , n76124 , n76125 , n76126 , n76127 , n76128 , 
 n76129 , n76130 , n76131 , n76132 , n76133 , n76134 , n76135 , n76136 , n76137 , n76138 , 
 n76139 , n76140 , n76141 , n76142 , n76143 , n76144 , n76145 , n76146 , n76147 , n76148 , 
 n76149 , n76150 , n76151 , n76152 , n76153 , n76154 , n76155 , n76156 , n76157 , n76158 , 
 n76159 , n76160 , n76161 , n76162 , n76163 , n76164 , n76165 , n76166 , n76167 , n76168 , 
 n76169 , n76170 , n76171 , n76172 , n76173 , n76174 , n76175 , n76176 , n76177 , n76178 , 
 n76179 , n76180 , n76181 , n76182 , n76183 , n76184 , n76185 , n76186 , n76187 , n76188 , 
 n76189 , n76190 , n76191 , n76192 , n76193 , n76194 , n76195 , n76196 , n76197 , n76198 , 
 n76199 , n76200 , n76201 , n76202 , n76203 , n76204 , n76205 , n76206 , n76207 , n76208 , 
 n76209 , n76210 , n76211 , n76212 , n76213 , n76214 , n76215 , n76216 , n76217 , n76218 , 
 n76219 , n76220 , n76221 , n76222 , n76223 , n76224 , n76225 , n76226 , n76227 , n76228 , 
 n76229 , n76230 , n76231 , n76232 , n76233 , n76234 , n76235 , n76236 , n76237 , n76238 , 
 n76239 , n76240 , n76241 , n76242 , n76243 , n76244 , n76245 , n76246 , n76247 , n76248 , 
 n76249 , n76250 , n76251 , n76252 , n76253 , n76254 , n76255 , n76256 , n76257 , n76258 , 
 n76259 , n76260 , n76261 , n76262 , n76263 , n76264 , n76265 , n76266 , n76267 , n76268 , 
 n76269 , n76270 , n76271 , n76272 , n76273 , n76274 , n76275 , n76276 , n76277 , n76278 , 
 n76279 , n76280 , n76281 , n76282 , n76283 , n76284 , n76285 , n76286 , n76287 , n76288 , 
 n76289 , n76290 , n76291 , n76292 , n76293 , n76294 , n76295 , n76296 , n76297 , n76298 , 
 n76299 , n76300 , n76301 , n76302 , n76303 , n76304 , n76305 , n76306 , n76307 , n76308 , 
 n76309 , n76310 , n76311 , n76312 , n76313 , n76314 , n76315 , n76316 , n76317 , n76318 , 
 n76319 , n76320 , n76321 , n76322 , n76323 , n76324 , n76325 , n76326 , n76327 , n76328 , 
 n76329 , n76330 , n76331 , n76332 , n76333 , n76334 , n76335 , n76336 , n76337 , n76338 , 
 n76339 , n76340 , n76341 , n76342 , n76343 , n76344 , n76345 , n76346 , n76347 , n76348 , 
 n76349 , n76350 , n76351 , n76352 , n76353 , n76354 , n76355 , n76356 , n76357 , n76358 , 
 n76359 , n76360 , n76361 , n76362 , n76363 , n76364 , n76365 , n76366 , n76367 , n76368 , 
 n76369 , n76370 , n76371 , n76372 , n76373 , n76374 , n76375 , n76376 , n76377 , n76378 , 
 n76379 , n76380 , n76381 , n76382 , n76383 , n76384 , n76385 , n76386 , n76387 , n76388 , 
 n76389 , n76390 , n76391 , n76392 , n76393 , n76394 , n76395 , n76396 , n76397 , n76398 , 
 n76399 , n76400 , n76401 , n76402 , n76403 , n76404 , n76405 , n76406 , n76407 , n76408 , 
 n76409 , n76410 , n76411 , n76412 , n76413 , n76414 , n76415 , n76416 , n76417 , n76418 , 
 n76419 , n76420 , n76421 , n76422 , n76423 , n76424 , n76425 , n76426 , n76427 , n76428 , 
 n76429 , n76430 , n76431 , n76432 , n76433 , n76434 , n76435 , n76436 , n76437 , n76438 , 
 n76439 , n76440 , n76441 , n76442 , n76443 , n76444 , n76445 , n76446 , n76447 , n76448 , 
 n76449 , n76450 , n76451 , n76452 , n76453 , n76454 , n76455 , n76456 , n76457 , n76458 , 
 n76459 , n76460 , n76461 , n76462 , n76463 , n76464 , n76465 , n76466 , n76467 , n76468 , 
 n76469 , n76470 , n76471 , n76472 , n76473 , n76474 , n76475 , n76476 , n76477 , n76478 , 
 n76479 , n76480 , n76481 , n76482 , n76483 , n76484 , n76485 , n76486 , n76487 , n76488 , 
 n76489 , n76490 , n76491 , n76492 , n76493 , n76494 , n76495 , n76496 , n76497 , n76498 , 
 n76499 , n76500 , n76501 , n76502 , n76503 , n76504 , n76505 , n76506 , n76507 , n76508 , 
 n76509 , n76510 , n76511 , n76512 , n76513 , n76514 , n76515 , n76516 , n76517 , n76518 , 
 n76519 , n76520 , n76521 , n76522 , n76523 , n76524 , n76525 , n76526 , n76527 , n76528 , 
 n76529 , n76530 , n76531 , n76532 , n76533 , n76534 , n76535 , n76536 , n76537 , n76538 , 
 n76539 , n76540 , n76541 , n76542 , n76543 , n76544 , n76545 , n76546 , n76547 , n76548 , 
 n76549 , n76550 , n76551 , n76552 , n76553 , n76554 , n76555 , n76556 , n76557 , n76558 , 
 n76559 , n76560 , n76561 , n76562 , n76563 , n76564 , n76565 , n76566 , n76567 , n76568 , 
 n76569 , n76570 , n76571 , n76572 , n76573 , n76574 , n76575 , n76576 , n76577 , n76578 , 
 n76579 , n76580 , n76581 , n76582 , n76583 , n76584 , n76585 , n76586 , n76587 , n76588 , 
 n76589 , n76590 , n76591 , n76592 , n76593 , n76594 , n76595 , n76596 , n76597 , n76598 , 
 n76599 , n76600 , n76601 , n76602 , n76603 , n76604 , n76605 , n76606 , n76607 , n76608 , 
 n76609 , n76610 , n76611 , n76612 , n76613 , n76614 , n76615 , n76616 , n76617 , n76618 , 
 n76619 , n76620 , n76621 , n76622 , n76623 , n76624 , n76625 , n76626 , n76627 , n76628 , 
 n76629 , n76630 , n76631 , n76632 , n76633 , n76634 , n76635 , n76636 , n76637 , n76638 , 
 n76639 , n76640 , n76641 , n76642 , n76643 , n76644 , n76645 , n76646 , n76647 , n76648 , 
 n76649 , n76650 , n76651 , n76652 , n76653 , n76654 , n76655 , n76656 , n76657 , n76658 , 
 n76659 , n76660 , n76661 , n76662 , n76663 , n76664 , n76665 , n76666 , n76667 , n76668 , 
 n76669 , n76670 , n76671 , n76672 , n76673 , n76674 , n76675 , n76676 , n76677 , n76678 , 
 n76679 , n76680 , n76681 , n76682 , n76683 , n76684 , n76685 , n76686 , n76687 , n76688 , 
 n76689 , n76690 , n76691 , n76692 , n76693 , n76694 , n76695 , n76696 , n76697 , n76698 , 
 n76699 , n76700 , n76701 , n76702 , n76703 , n76704 , n76705 , n76706 , n76707 , n76708 , 
 n76709 , n76710 , n76711 , n76712 , n76713 , n76714 , n76715 , n76716 , n76717 , n76718 , 
 n76719 , n76720 , n76721 , n76722 , n76723 , n76724 , n76725 , n76726 , n76727 , n76728 , 
 n76729 , n76730 , n76731 , n76732 , n76733 , n76734 , n76735 , n76736 , n76737 , n76738 , 
 n76739 , n76740 , n76741 , n76742 , n76743 , n76744 , n76745 , n76746 , n76747 , n76748 , 
 n76749 , n76750 , n76751 , n76752 , n76753 , n76754 , n76755 , n76756 , n76757 , n76758 , 
 n76759 , n76760 , n76761 , n76762 , n76763 , n76764 , n76765 , n76766 , n76767 , n76768 , 
 n76769 , n76770 , n76771 , n76772 , n76773 , n76774 , n76775 , n76776 , n76777 , n76778 , 
 n76779 , n76780 , n76781 , n76782 , n76783 , n76784 , n76785 , n76786 , n76787 , n76788 , 
 n76789 , n76790 , n76791 , n76792 , n76793 , n76794 , n76795 , n76796 , n76797 , n76798 , 
 n76799 , n76800 , n76801 , n76802 , n76803 , n76804 , n76805 , n76806 , n76807 , n76808 , 
 n76809 , n76810 , n76811 , n76812 , n76813 , n76814 , n76815 , n76816 , n76817 , n76818 , 
 n76819 , n76820 , n76821 , n76822 , n76823 , n76824 , n76825 , n76826 , n76827 , n76828 , 
 n76829 , n76830 , n76831 , n76832 , n76833 , n76834 , n76835 , n76836 , n76837 , n76838 , 
 n76839 , n76840 , n76841 , n76842 , n76843 , n76844 , n76845 , n76846 , n76847 , n76848 , 
 n76849 , n76850 , n76851 , n76852 , n76853 , n76854 , n76855 , n76856 , n76857 , n76858 , 
 n76859 , n76860 , n76861 , n76862 , n76863 , n76864 , n76865 , n76866 , n76867 , n76868 , 
 n76869 , n76870 , n76871 , n76872 , n76873 , n76874 , n76875 , n76876 , n76877 , n76878 , 
 n76879 , n76880 , n76881 , n76882 , n76883 , n76884 , n76885 , n76886 , n76887 , n76888 , 
 n76889 , n76890 , n76891 , n76892 , n76893 , n76894 , n76895 , n76896 , n76897 , n76898 , 
 n76899 , n76900 , n76901 , n76902 , n76903 , n76904 , n76905 , n76906 , n76907 , n76908 , 
 n76909 , n76910 , n76911 , n76912 , n76913 , n76914 , n76915 , n76916 , n76917 , n76918 , 
 n76919 , n76920 , n76921 , n76922 , n76923 , n76924 , n76925 , n76926 , n76927 , n76928 , 
 n76929 , n76930 , n76931 , n76932 , n76933 , n76934 , n76935 , n76936 , n76937 , n76938 , 
 n76939 , n76940 , n76941 , n76942 , n76943 , n76944 , n76945 , n76946 , n76947 , n76948 , 
 n76949 , n76950 , n76951 , n76952 , n76953 , n76954 , n76955 , n76956 , n76957 , n76958 , 
 n76959 , n76960 , n76961 , n76962 , n76963 , n76964 , n76965 , n76966 , n76967 , n76968 , 
 n76969 , n76970 , n76971 , n76972 , n76973 , n76974 , n76975 , n76976 , n76977 , n76978 , 
 n76979 , n76980 , n76981 , n76982 , n76983 , n76984 , n76985 , n76986 , n76987 , n76988 , 
 n76989 , n76990 , n76991 , n76992 , n76993 , n76994 , n76995 , n76996 , n76997 , n76998 , 
 n76999 , n77000 , n77001 , n77002 , n77003 , n77004 , n77005 , n77006 , n77007 , n77008 , 
 n77009 , n77010 , n77011 , n77012 , n77013 , n77014 , n77015 , n77016 , n77017 , n77018 , 
 n77019 , n77020 , n77021 , n77022 , n77023 , n77024 , n77025 , n77026 , n77027 , n77028 , 
 n77029 , n77030 , n77031 , n77032 , n77033 , n77034 , n77035 , n77036 , n77037 , n77038 , 
 n77039 , n77040 , n77041 , n77042 , n77043 , n77044 , n77045 , n77046 , n77047 , n77048 , 
 n77049 , n77050 , n77051 , n77052 , n77053 , n77054 , n77055 , n77056 , n77057 , n77058 , 
 n77059 , n77060 , n77061 , n77062 , n77063 , n77064 , n77065 , n77066 , n77067 , n77068 , 
 n77069 , n77070 , n77071 , n77072 , n77073 , n77074 , n77075 , n77076 , n77077 , n77078 , 
 n77079 , n77080 , n77081 , n77082 , n77083 , n77084 , n77085 , n77086 , n77087 , n77088 , 
 n77089 , n77090 , n77091 , n77092 , n77093 , n77094 , n77095 , n77096 , n77097 , n77098 , 
 n77099 , n77100 , n77101 , n77102 , n77103 , n77104 , n77105 , n77106 , n77107 , n77108 , 
 n77109 , n77110 , n77111 , n77112 , n77113 , n77114 , n77115 , n77116 , n77117 , n77118 , 
 n77119 , n77120 , n77121 , n77122 , n77123 , n77124 , n77125 , n77126 , n77127 , n77128 , 
 n77129 , n77130 , n77131 , n77132 , n77133 , n77134 , n77135 , n77136 , n77137 , n77138 , 
 n77139 , n77140 , n77141 , n77142 , n77143 , n77144 , n77145 , n77146 , n77147 , n77148 , 
 n77149 , n77150 , n77151 , n77152 , n77153 , n77154 , n77155 , n77156 , n77157 , n77158 , 
 n77159 , n77160 , n77161 , n77162 , n77163 , n77164 , n77165 , n77166 , n77167 , n77168 , 
 n77169 , n77170 , n77171 , n77172 , n77173 , n77174 , n77175 , n77176 , n77177 , n77178 , 
 n77179 , n77180 , n77181 , n77182 , n77183 , n77184 , n77185 , n77186 , n77187 , n77188 , 
 n77189 , n77190 , n77191 , n77192 , n77193 , n77194 , n77195 , n77196 , n77197 , n77198 , 
 n77199 , n77200 , n77201 , n77202 , n77203 , n77204 , n77205 , n77206 , n77207 , n77208 , 
 n77209 , n77210 , n77211 , n77212 , n77213 , n77214 , n77215 , n77216 , n77217 , n77218 , 
 n77219 , n77220 , n77221 , n77222 , n77223 , n77224 , n77225 , n77226 , n77227 , n77228 , 
 n77229 , n77230 , n77231 , n77232 , n77233 , n77234 , n77235 , n77236 , n77237 , n77238 , 
 n77239 , n77240 , n77241 , n77242 , n77243 , n77244 , n77245 , n77246 , n77247 , n77248 , 
 n77249 , n77250 , n77251 , n77252 , n77253 , n77254 , n77255 , n77256 , n77257 , n77258 , 
 n77259 , n77260 , n77261 , n77262 , n77263 , n77264 , n77265 , n77266 , n77267 , n77268 , 
 n77269 , n77270 , n77271 , n77272 , n77273 , n77274 , n77275 , n77276 , n77277 , n77278 , 
 n77279 , n77280 , n77281 , n77282 , n77283 , n77284 , n77285 , n77286 , n77287 , n77288 , 
 n77289 , n77290 , n77291 , n77292 , n77293 , n77294 , n77295 , n77296 , n77297 , n77298 , 
 n77299 , n77300 , n77301 , n77302 , n77303 , n77304 , n77305 , n77306 , n77307 , n77308 , 
 n77309 , n77310 , n77311 , n77312 , n77313 , n77314 , n77315 , n77316 , n77317 , n77318 , 
 n77319 , n77320 , n77321 , n77322 , n77323 , n77324 , n77325 , n77326 , n77327 , n77328 , 
 n77329 , n77330 , n77331 , n77332 , n77333 , n77334 , n77335 , n77336 , n77337 , n77338 , 
 n77339 , n77340 , n77341 , n77342 , n77343 , n77344 , n77345 , n77346 , n77347 , n77348 , 
 n77349 , n77350 , n77351 , n77352 , n77353 , n77354 , n77355 , n77356 , n77357 , n77358 , 
 n77359 , n77360 , n77361 , n77362 , n77363 , n77364 , n77365 , n77366 , n77367 , n77368 , 
 n77369 , n77370 , n77371 , n77372 , n77373 , n77374 , n77375 , n77376 , n77377 , n77378 , 
 n77379 , n77380 , n77381 , n77382 , n77383 , n77384 , n77385 , n77386 , n77387 , n77388 , 
 n77389 , n77390 , n77391 , n77392 , n77393 , n77394 , n77395 , n77396 , n77397 , n77398 , 
 n77399 , n77400 , n77401 , n77402 , n77403 , n77404 , n77405 , n77406 , n77407 , n77408 , 
 n77409 , n77410 , n77411 , n77412 , n77413 , n77414 , n77415 , n77416 , n77417 , n77418 , 
 n77419 , n77420 , n77421 , n77422 , n77423 , n77424 , n77425 , n77426 , n77427 , n77428 , 
 n77429 , n77430 , n77431 , n77432 , n77433 , n77434 , n77435 , n77436 , n77437 , n77438 , 
 n77439 , n77440 , n77441 , n77442 , n77443 , n77444 , n77445 , n77446 , n77447 , n77448 , 
 n77449 , n77450 , n77451 , n77452 , n77453 , n77454 , n77455 , n77456 , n77457 , n77458 , 
 n77459 , n77460 , n77461 , n77462 , n77463 , n77464 , n77465 , n77466 , n77467 , n77468 , 
 n77469 , n77470 , n77471 , n77472 , n77473 , n77474 , n77475 , n77476 , n77477 , n77478 , 
 n77479 , n77480 , n77481 , n77482 , n77483 , n77484 , n77485 , n77486 , n77487 , n77488 , 
 n77489 , n77490 , n77491 , n77492 , n77493 , n77494 , n77495 , n77496 , n77497 , n77498 , 
 n77499 , n77500 , n77501 , n77502 , n77503 , n77504 , n77505 , n77506 , n77507 , n77508 , 
 n77509 , n77510 , n77511 , n77512 , n77513 , n77514 , n77515 , n77516 , n77517 , n77518 , 
 n77519 , n77520 , n77521 , n77522 , n77523 , n77524 , n77525 , n77526 , n77527 , n77528 , 
 n77529 , n77530 , n77531 , n77532 , n77533 , n77534 , n77535 , n77536 , n77537 , n77538 , 
 n77539 , n77540 , n77541 , n77542 , n77543 , n77544 , n77545 , n77546 , n77547 , n77548 , 
 n77549 , n77550 , n77551 , n77552 , n77553 , n77554 , n77555 , n77556 , n77557 , n77558 , 
 n77559 , n77560 , n77561 , n77562 , n77563 , n77564 , n77565 , n77566 , n77567 , n77568 , 
 n77569 , n77570 , n77571 , n77572 , n77573 , n77574 , n77575 , n77576 , n77577 , n77578 , 
 n77579 , n77580 , n77581 , n77582 , n77583 , n77584 , n77585 , n77586 , n77587 , n77588 , 
 n77589 , n77590 , n77591 , n77592 , n77593 , n77594 , n77595 , n77596 , n77597 , n77598 , 
 n77599 , n77600 , n77601 , n77602 , n77603 , n77604 , n77605 , n77606 , n77607 , n77608 , 
 n77609 , n77610 , n77611 , n77612 , n77613 , n77614 , n77615 , n77616 , n77617 , n77618 , 
 n77619 , n77620 , n77621 , n77622 , n77623 , n77624 , n77625 , n77626 , n77627 , n77628 , 
 n77629 , n77630 , n77631 , n77632 , n77633 , n77634 , n77635 , n77636 , n77637 , n77638 , 
 n77639 , n77640 , n77641 , n77642 , n77643 , n77644 , n77645 , n77646 , n77647 , n77648 , 
 n77649 , n77650 , n77651 , n77652 , n77653 , n77654 , n77655 , n77656 , n77657 , n77658 , 
 n77659 , n77660 , n77661 , n77662 , n77663 , n77664 , n77665 , n77666 , n77667 , n77668 , 
 n77669 , n77670 , n77671 , n77672 , n77673 , n77674 , n77675 , n77676 , n77677 , n77678 , 
 n77679 , n77680 , n77681 , n77682 , n77683 , n77684 , n77685 , n77686 , n77687 , n77688 , 
 n77689 , n77690 , n77691 , n77692 , n77693 , n77694 , n77695 , n77696 , n77697 , n77698 , 
 n77699 , n77700 , n77701 , n77702 , n77703 , n77704 , n77705 , n77706 , n77707 , n77708 , 
 n77709 , n77710 , n77711 , n77712 , n77713 , n77714 , n77715 , n77716 , n77717 , n77718 , 
 n77719 , n77720 , n77721 , n77722 , n77723 , n77724 , n77725 , n77726 , n77727 , n77728 , 
 n77729 , n77730 , n77731 , n77732 , n77733 , n77734 , n77735 , n77736 , n77737 , n77738 , 
 n77739 , n77740 , n77741 , n77742 , n77743 , n77744 , n77745 , n77746 , n77747 , n77748 , 
 n77749 , n77750 , n77751 , n77752 , n77753 , n77754 , n77755 , n77756 , n77757 , n77758 , 
 n77759 , n77760 , n77761 , n77762 , n77763 , n77764 , n77765 , n77766 , n77767 , n77768 , 
 n77769 , n77770 , n77771 , n77772 , n77773 , n77774 , n77775 , n77776 , n77777 , n77778 , 
 n77779 , n77780 , n77781 , n77782 , n77783 , n77784 , n77785 , n77786 , n77787 , n77788 , 
 n77789 , n77790 , n77791 , n77792 , n77793 , n77794 , n77795 , n77796 , n77797 , n77798 , 
 n77799 , n77800 , n77801 , n77802 , n77803 , n77804 , n77805 , n77806 , n77807 , n77808 , 
 n77809 , n77810 , n77811 , n77812 , n77813 , n77814 , n77815 , n77816 , n77817 , n77818 , 
 n77819 , n77820 , n77821 , n77822 , n77823 , n77824 , n77825 , n77826 , n77827 , n77828 , 
 n77829 , n77830 , n77831 , n77832 , n77833 , n77834 , n77835 , n77836 , n77837 , n77838 , 
 n77839 , n77840 , n77841 , n77842 , n77843 , n77844 , n77845 , n77846 , n77847 , n77848 , 
 n77849 , n77850 , n77851 , n77852 , n77853 , n77854 , n77855 , n77856 , n77857 , n77858 , 
 n77859 , n77860 , n77861 , n77862 , n77863 , n77864 , n77865 , n77866 , n77867 , n77868 , 
 n77869 , n77870 , n77871 , n77872 , n77873 , n77874 , n77875 , n77876 , n77877 , n77878 , 
 n77879 , n77880 , n77881 , n77882 , n77883 , n77884 , n77885 , n77886 , n77887 , n77888 , 
 n77889 , n77890 , n77891 , n77892 , n77893 , n77894 , n77895 , n77896 , n77897 , n77898 , 
 n77899 , n77900 , n77901 , n77902 , n77903 , n77904 , n77905 , n77906 , n77907 , n77908 , 
 n77909 , n77910 , n77911 , n77912 , n77913 , n77914 , n77915 , n77916 , n77917 , n77918 , 
 n77919 , n77920 , n77921 , n77922 , n77923 , n77924 , n77925 , n77926 , n77927 , n77928 , 
 n77929 , n77930 , n77931 , n77932 , n77933 , n77934 , n77935 , n77936 , n77937 , n77938 , 
 n77939 , n77940 , n77941 , n77942 , n77943 , n77944 , n77945 , n77946 , n77947 , n77948 , 
 n77949 , n77950 , n77951 , n77952 , n77953 , n77954 , n77955 , n77956 , n77957 , n77958 , 
 n77959 , n77960 , n77961 , n77962 , n77963 , n77964 , n77965 , n77966 , n77967 , n77968 , 
 n77969 , n77970 , n77971 , n77972 , n77973 , n77974 , n77975 , n77976 , n77977 , n77978 , 
 n77979 , n77980 , n77981 , n77982 , n77983 , n77984 , n77985 , n77986 , n77987 , n77988 , 
 n77989 , n77990 , n77991 , n77992 , n77993 , n77994 , n77995 , n77996 , n77997 , n77998 , 
 n77999 , n78000 , n78001 , n78002 , n78003 , n78004 , n78005 , n78006 , n78007 , n78008 , 
 n78009 , n78010 , n78011 , n78012 , n78013 , n78014 , n78015 , n78016 , n78017 , n78018 , 
 n78019 , n78020 , n78021 , n78022 , n78023 , n78024 , n78025 , n78026 , n78027 , n78028 , 
 n78029 , n78030 , n78031 , n78032 , n78033 , n78034 , n78035 , n78036 , n78037 , n78038 , 
 n78039 , n78040 , n78041 , n78042 , n78043 , n78044 , n78045 , n78046 , n78047 , n78048 , 
 n78049 , n78050 , n78051 , n78052 , n78053 , n78054 , n78055 , n78056 , n78057 , n78058 , 
 n78059 , n78060 , n78061 , n78062 , n78063 , n78064 , n78065 , n78066 , n78067 , n78068 , 
 n78069 , n78070 , n78071 , n78072 , n78073 , n78074 , n78075 , n78076 , n78077 , n78078 , 
 n78079 , n78080 , n78081 , n78082 , n78083 , n78084 , n78085 , n78086 , n78087 , n78088 , 
 n78089 , n78090 , n78091 , n78092 , n78093 , n78094 , n78095 , n78096 , n78097 , n78098 , 
 n78099 , n78100 , n78101 , n78102 , n78103 , n78104 , n78105 , n78106 , n78107 , n78108 , 
 n78109 , n78110 , n78111 , n78112 , n78113 , n78114 , n78115 , n78116 , n78117 , n78118 , 
 n78119 , n78120 , n78121 , n78122 , n78123 , n78124 , n78125 , n78126 , n78127 , n78128 , 
 n78129 , n78130 , n78131 , n78132 , n78133 , n78134 , n78135 , n78136 , n78137 , n78138 , 
 n78139 , n78140 , n78141 , n78142 , n78143 , n78144 , n78145 , n78146 , n78147 , n78148 , 
 n78149 , n78150 , n78151 , n78152 , n78153 , n78154 , n78155 , n78156 , n78157 , n78158 , 
 n78159 , n78160 , n78161 , n78162 , n78163 , n78164 , n78165 , n78166 , n78167 , n78168 , 
 n78169 , n78170 , n78171 , n78172 , n78173 , n78174 , n78175 , n78176 , n78177 , n78178 , 
 n78179 , n78180 , n78181 , n78182 , n78183 , n78184 , n78185 , n78186 , n78187 , n78188 , 
 n78189 , n78190 , n78191 , n78192 , n78193 , n78194 , n78195 , n78196 , n78197 , n78198 , 
 n78199 , n78200 , n78201 , n78202 , n78203 , n78204 , n78205 , n78206 , n78207 , n78208 , 
 n78209 , n78210 , n78211 , n78212 , n78213 , n78214 , n78215 , n78216 , n78217 , n78218 , 
 n78219 , n78220 , n78221 , n78222 , n78223 , n78224 , n78225 , n78226 , n78227 , n78228 , 
 n78229 , n78230 , n78231 , n78232 , n78233 , n78234 , n78235 , n78236 , n78237 , n78238 , 
 n78239 , n78240 , n78241 , n78242 , n78243 , n78244 , n78245 , n78246 , n78247 , n78248 , 
 n78249 , n78250 , n78251 , n78252 , n78253 , n78254 , n78255 , n78256 , n78257 , n78258 , 
 n78259 , n78260 , n78261 , n78262 , n78263 , n78264 , n78265 , n78266 , n78267 , n78268 , 
 n78269 , n78270 , n78271 , n78272 , n78273 , n78274 , n78275 , n78276 , n78277 , n78278 , 
 n78279 , n78280 , n78281 , n78282 , n78283 , n78284 , n78285 , n78286 , n78287 , n78288 , 
 n78289 , n78290 , n78291 , n78292 , n78293 , n78294 , n78295 , n78296 , n78297 , n78298 , 
 n78299 , n78300 , n78301 , n78302 , n78303 , n78304 , n78305 , n78306 , n78307 , n78308 , 
 n78309 , n78310 , n78311 , n78312 , n78313 , n78314 , n78315 , n78316 , n78317 , n78318 , 
 n78319 , n78320 , n78321 , n78322 , n78323 , n78324 , n78325 , n78326 , n78327 , n78328 , 
 n78329 , n78330 , n78331 , n78332 , n78333 , n78334 , n78335 , n78336 , n78337 , n78338 , 
 n78339 , n78340 , n78341 , n78342 , n78343 , n78344 , n78345 , n78346 , n78347 , n78348 , 
 n78349 , n78350 , n78351 , n78352 , n78353 , n78354 , n78355 , n78356 , n78357 , n78358 , 
 n78359 , n78360 , n78361 , n78362 , n78363 , n78364 , n78365 , n78366 , n78367 , n78368 , 
 n78369 , n78370 , n78371 , n78372 , n78373 , n78374 , n78375 , n78376 , n78377 , n78378 , 
 n78379 , n78380 , n78381 , n78382 , n78383 , n78384 , n78385 , n78386 , n78387 , n78388 , 
 n78389 , n78390 , n78391 , n78392 , n78393 , n78394 , n78395 , n78396 , n78397 , n78398 , 
 n78399 , n78400 , n78401 , n78402 , n78403 , n78404 , n78405 , n78406 , n78407 , n78408 , 
 n78409 , n78410 , n78411 , n78412 , n78413 , n78414 , n78415 , n78416 , n78417 , n78418 , 
 n78419 , n78420 , n78421 , n78422 , n78423 , n78424 , n78425 , n78426 , n78427 , n78428 , 
 n78429 , n78430 , n78431 , n78432 , n78433 , n78434 , n78435 , n78436 , n78437 , n78438 , 
 n78439 , n78440 , n78441 , n78442 , n78443 , n78444 , n78445 , n78446 , n78447 , n78448 , 
 n78449 , n78450 , n78451 , n78452 , n78453 , n78454 , n78455 , n78456 , n78457 , n78458 , 
 n78459 , n78460 , n78461 , n78462 , n78463 , n78464 , n78465 , n78466 , n78467 , n78468 , 
 n78469 , n78470 , n78471 , n78472 , n78473 , n78474 , n78475 , n78476 , n78477 , n78478 , 
 n78479 , n78480 , n78481 , n78482 , n78483 , n78484 , n78485 , n78486 , n78487 , n78488 , 
 n78489 , n78490 , n78491 , n78492 , n78493 , n78494 , n78495 , n78496 , n78497 , n78498 , 
 n78499 , n78500 , n78501 , n78502 , n78503 , n78504 , n78505 , n78506 , n78507 , n78508 , 
 n78509 , n78510 , n78511 , n78512 , n78513 , n78514 , n78515 , n78516 , n78517 , n78518 , 
 n78519 , n78520 , n78521 , n78522 , n78523 , n78524 , n78525 , n78526 , n78527 , n78528 , 
 n78529 , n78530 , n78531 , n78532 , n78533 , n78534 , n78535 , n78536 , n78537 , n78538 , 
 n78539 , n78540 , n78541 , n78542 , n78543 , n78544 , n78545 , n78546 , n78547 , n78548 , 
 n78549 , n78550 , n78551 , n78552 , n78553 , n78554 , n78555 , n78556 , n78557 , n78558 , 
 n78559 , n78560 , n78561 , n78562 , n78563 , n78564 , n78565 , n78566 , n78567 , n78568 , 
 n78569 , n78570 , n78571 , n78572 , n78573 , n78574 , n78575 , n78576 , n78577 , n78578 , 
 n78579 , n78580 , n78581 , n78582 , n78583 , n78584 , n78585 , n78586 , n78587 , n78588 , 
 n78589 , n78590 , n78591 , n78592 , n78593 , n78594 , n78595 , n78596 , n78597 , n78598 , 
 n78599 , n78600 , n78601 , n78602 , n78603 , n78604 , n78605 , n78606 , n78607 , n78608 , 
 n78609 , n78610 , n78611 , n78612 , n78613 , n78614 , n78615 , n78616 , n78617 , n78618 , 
 n78619 , n78620 , n78621 , n78622 , n78623 , n78624 , n78625 , n78626 , n78627 , n78628 , 
 n78629 , n78630 , n78631 , n78632 , n78633 , n78634 , n78635 , n78636 , n78637 , n78638 , 
 n78639 , n78640 , n78641 , n78642 , n78643 , n78644 , n78645 , n78646 , n78647 , n78648 , 
 n78649 , n78650 , n78651 , n78652 , n78653 , n78654 , n78655 , n78656 , n78657 , n78658 , 
 n78659 , n78660 , n78661 , n78662 , n78663 , n78664 , n78665 , n78666 , n78667 , n78668 , 
 n78669 , n78670 , n78671 , n78672 , n78673 , n78674 , n78675 , n78676 , n78677 , n78678 , 
 n78679 , n78680 , n78681 , n78682 , n78683 , n78684 , n78685 , n78686 , n78687 , n78688 , 
 n78689 , n78690 , n78691 , n78692 , n78693 , n78694 , n78695 , n78696 , n78697 , n78698 , 
 n78699 , n78700 , n78701 , n78702 , n78703 , n78704 , n78705 , n78706 , n78707 , n78708 , 
 n78709 , n78710 , n78711 , n78712 , n78713 , n78714 , n78715 , n78716 , n78717 , n78718 , 
 n78719 , n78720 , n78721 , n78722 , n78723 , n78724 , n78725 , n78726 , n78727 , n78728 , 
 n78729 , n78730 , n78731 , n78732 , n78733 , n78734 , n78735 , n78736 , n78737 , n78738 , 
 n78739 , n78740 , n78741 , n78742 , n78743 , n78744 , n78745 , n78746 , n78747 , n78748 , 
 n78749 , n78750 , n78751 , n78752 , n78753 , n78754 , n78755 , n78756 , n78757 , n78758 , 
 n78759 , n78760 , n78761 , n78762 , n78763 , n78764 , n78765 , n78766 , n78767 , n78768 , 
 n78769 , n78770 , n78771 , n78772 , n78773 , n78774 , n78775 , n78776 , n78777 , n78778 , 
 n78779 , n78780 , n78781 , n78782 , n78783 , n78784 , n78785 , n78786 , n78787 , n78788 , 
 n78789 , n78790 , n78791 , n78792 , n78793 , n78794 , n78795 , n78796 , n78797 , n78798 , 
 n78799 , n78800 , n78801 , n78802 , n78803 , n78804 , n78805 , n78806 , n78807 , n78808 , 
 n78809 , n78810 , n78811 , n78812 , n78813 , n78814 , n78815 , n78816 , n78817 , n78818 , 
 n78819 , n78820 , n78821 , n78822 , n78823 , n78824 , n78825 , n78826 , n78827 , n78828 , 
 n78829 , n78830 , n78831 , n78832 , n78833 , n78834 , n78835 , n78836 , n78837 , n78838 , 
 n78839 , n78840 , n78841 , n78842 , n78843 , n78844 , n78845 , n78846 , n78847 , n78848 , 
 n78849 , n78850 , n78851 , n78852 , n78853 , n78854 , n78855 , n78856 , n78857 , n78858 , 
 n78859 , n78860 , n78861 , n78862 , n78863 , n78864 , n78865 , n78866 , n78867 , n78868 , 
 n78869 , n78870 , n78871 , n78872 , n78873 , n78874 , n78875 , n78876 , n78877 , n78878 , 
 n78879 , n78880 , n78881 , n78882 , n78883 , n78884 , n78885 , n78886 , n78887 , n78888 , 
 n78889 , n78890 , n78891 , n78892 , n78893 , n78894 , n78895 , n78896 , n78897 , n78898 , 
 n78899 , n78900 , n78901 , n78902 , n78903 , n78904 , n78905 , n78906 , n78907 , n78908 , 
 n78909 , n78910 , n78911 , n78912 , n78913 , n78914 , n78915 , n78916 , n78917 , n78918 , 
 n78919 , n78920 , n78921 , n78922 , n78923 , n78924 , n78925 , n78926 , n78927 , n78928 , 
 n78929 , n78930 , n78931 , n78932 , n78933 , n78934 , n78935 , n78936 , n78937 , n78938 , 
 n78939 , n78940 , n78941 , n78942 , n78943 , n78944 , n78945 , n78946 , n78947 , n78948 , 
 n78949 , n78950 , n78951 , n78952 , n78953 , n78954 , n78955 , n78956 , n78957 , n78958 , 
 n78959 , n78960 , n78961 , n78962 , n78963 , n78964 , n78965 , n78966 , n78967 , n78968 , 
 n78969 , n78970 , n78971 , n78972 , n78973 , n78974 , n78975 , n78976 , n78977 , n78978 , 
 n78979 , n78980 , n78981 , n78982 , n78983 , n78984 , n78985 , n78986 , n78987 , n78988 , 
 n78989 , n78990 , n78991 , n78992 , n78993 , n78994 , n78995 , n78996 , n78997 , n78998 , 
 n78999 , n79000 , n79001 , n79002 , n79003 , n79004 , n79005 , n79006 , n79007 , n79008 , 
 n79009 , n79010 , n79011 , n79012 , n79013 , n79014 , n79015 , n79016 , n79017 , n79018 , 
 n79019 , n79020 , n79021 , n79022 , n79023 , n79024 , n79025 , n79026 , n79027 , n79028 , 
 n79029 , n79030 , n79031 , n79032 , n79033 , n79034 , n79035 , n79036 , n79037 , n79038 , 
 n79039 , n79040 , n79041 , n79042 , n79043 , n79044 , n79045 , n79046 , n79047 , n79048 , 
 n79049 , n79050 , n79051 , n79052 , n79053 , n79054 , n79055 , n79056 , n79057 , n79058 , 
 n79059 , n79060 , n79061 , n79062 , n79063 , n79064 , n79065 , n79066 , n79067 , n79068 , 
 n79069 , n79070 , n79071 , n79072 , n79073 , n79074 , n79075 , n79076 , n79077 , n79078 , 
 n79079 , n79080 , n79081 , n79082 , n79083 , n79084 , n79085 , n79086 , n79087 , n79088 , 
 n79089 , n79090 , n79091 , n79092 , n79093 , n79094 , n79095 , n79096 , n79097 , n79098 , 
 n79099 , n79100 , n79101 , n79102 , n79103 , n79104 , n79105 , n79106 , n79107 , n79108 , 
 n79109 , n79110 , n79111 , n79112 , n79113 , n79114 , n79115 , n79116 , n79117 , n79118 , 
 n79119 , n79120 , n79121 , n79122 , n79123 , n79124 , n79125 , n79126 , n79127 , n79128 , 
 n79129 , n79130 , n79131 , n79132 , n79133 , n79134 , n79135 , n79136 , n79137 , n79138 , 
 n79139 , n79140 , n79141 , n79142 , n79143 , n79144 , n79145 , n79146 , n79147 , n79148 , 
 n79149 , n79150 , n79151 , n79152 , n79153 , n79154 , n79155 , n79156 , n79157 , n79158 , 
 n79159 , n79160 , n79161 , n79162 , n79163 , n79164 , n79165 , n79166 , n79167 , n79168 , 
 n79169 , n79170 , n79171 , n79172 , n79173 , n79174 , n79175 , n79176 , n79177 , n79178 , 
 n79179 , n79180 , n79181 , n79182 , n79183 , n79184 , n79185 , n79186 , n79187 , n79188 , 
 n79189 , n79190 , n79191 , n79192 , n79193 , n79194 , n79195 , n79196 , n79197 , n79198 , 
 n79199 , n79200 , n79201 , n79202 , n79203 , n79204 , n79205 , n79206 , n79207 , n79208 , 
 n79209 , n79210 , n79211 , n79212 , n79213 , n79214 , n79215 , n79216 , n79217 , n79218 , 
 n79219 , n79220 , n79221 , n79222 , n79223 , n79224 , n79225 , n79226 , n79227 , n79228 , 
 n79229 , n79230 , n79231 , n79232 , n79233 , n79234 , n79235 , n79236 , n79237 , n79238 , 
 n79239 , n79240 , n79241 , n79242 , n79243 , n79244 , n79245 , n79246 , n79247 , n79248 , 
 n79249 , n79250 , n79251 , n79252 , n79253 , n79254 , n79255 , n79256 , n79257 , n79258 , 
 n79259 , n79260 , n79261 , n79262 , n79263 , n79264 , n79265 , n79266 , n79267 , n79268 , 
 n79269 , n79270 , n79271 , n79272 , n79273 , n79274 , n79275 , n79276 , n79277 , n79278 , 
 n79279 , n79280 , n79281 , n79282 , n79283 , n79284 , n79285 , n79286 , n79287 , n79288 , 
 n79289 , n79290 , n79291 , n79292 , n79293 , n79294 , n79295 , n79296 , n79297 , n79298 , 
 n79299 , n79300 , n79301 , n79302 , n79303 , n79304 , n79305 , n79306 , n79307 , n79308 , 
 n79309 , n79310 , n79311 , n79312 , n79313 , n79314 , n79315 , n79316 , n79317 , n79318 , 
 n79319 , n79320 , n79321 , n79322 , n79323 , n79324 , n79325 , n79326 , n79327 , n79328 , 
 n79329 , n79330 , n79331 , n79332 , n79333 , n79334 , n79335 , n79336 , n79337 , n79338 , 
 n79339 , n79340 , n79341 , n79342 , n79343 , n79344 , n79345 , n79346 , n79347 , n79348 , 
 n79349 , n79350 , n79351 , n79352 , n79353 , n79354 , n79355 , n79356 , n79357 , n79358 , 
 n79359 , n79360 , n79361 , n79362 , n79363 , n79364 , n79365 , n79366 , n79367 , n79368 , 
 n79369 , n79370 , n79371 , n79372 , n79373 , n79374 , n79375 , n79376 , n79377 , n79378 , 
 n79379 , n79380 , n79381 , n79382 , n79383 , n79384 , n79385 , n79386 , n79387 , n79388 , 
 n79389 , n79390 , n79391 , n79392 , n79393 , n79394 , n79395 , n79396 , n79397 , n79398 , 
 n79399 , n79400 , n79401 , n79402 , n79403 , n79404 , n79405 , n79406 , n79407 , n79408 , 
 n79409 , n79410 , n79411 , n79412 , n79413 , n79414 , n79415 , n79416 , n79417 , n79418 , 
 n79419 , n79420 , n79421 , n79422 , n79423 , n79424 , n79425 , n79426 , n79427 , n79428 , 
 n79429 , n79430 , n79431 , n79432 , n79433 , n79434 , n79435 , n79436 , n79437 , n79438 , 
 n79439 , n79440 , n79441 , n79442 , n79443 , n79444 , n79445 , n79446 , n79447 , n79448 , 
 n79449 , n79450 , n79451 , n79452 , n79453 , n79454 , n79455 , n79456 , n79457 , n79458 , 
 n79459 , n79460 , n79461 , n79462 , n79463 , n79464 , n79465 , n79466 , n79467 , n79468 , 
 n79469 , n79470 , n79471 , n79472 , n79473 , n79474 , n79475 , n79476 , n79477 , n79478 , 
 n79479 , n79480 , n79481 , n79482 , n79483 , n79484 , n79485 , n79486 , n79487 , n79488 , 
 n79489 , n79490 , n79491 , n79492 , n79493 , n79494 , n79495 , n79496 , n79497 , n79498 , 
 n79499 , n79500 , n79501 , n79502 , n79503 , n79504 , n79505 , n79506 , n79507 , n79508 , 
 n79509 , n79510 , n79511 , n79512 , n79513 , n79514 , n79515 , n79516 , n79517 , n79518 , 
 n79519 , n79520 , n79521 , n79522 , n79523 , n79524 , n79525 , n79526 , n79527 , n79528 , 
 n79529 , n79530 , n79531 , n79532 , n79533 , n79534 , n79535 , n79536 , n79537 , n79538 , 
 n79539 , n79540 , n79541 , n79542 , n79543 , n79544 , n79545 , n79546 , n79547 , n79548 , 
 n79549 , n79550 , n79551 , n79552 , n79553 , n79554 , n79555 , n79556 , n79557 , n79558 , 
 n79559 , n79560 , n79561 , n79562 , n79563 , n79564 , n79565 , n79566 , n79567 , n79568 , 
 n79569 , n79570 , n79571 , n79572 , n79573 , n79574 , n79575 , n79576 , n79577 , n79578 , 
 n79579 , n79580 , n79581 , n79582 , n79583 , n79584 , n79585 , n79586 , n79587 , n79588 , 
 n79589 , n79590 , n79591 , n79592 , n79593 , n79594 , n79595 , n79596 , n79597 , n79598 , 
 n79599 , n79600 , n79601 , n79602 , n79603 , n79604 , n79605 , n79606 , n79607 , n79608 , 
 n79609 , n79610 , n79611 , n79612 , n79613 , n79614 , n79615 , n79616 , n79617 , n79618 , 
 n79619 , n79620 , n79621 , n79622 , n79623 , n79624 , n79625 , n79626 , n79627 , n79628 , 
 n79629 , n79630 , n79631 , n79632 , n79633 , n79634 , n79635 , n79636 , n79637 , n79638 , 
 n79639 , n79640 , n79641 , n79642 , n79643 , n79644 , n79645 , n79646 , n79647 , n79648 , 
 n79649 , n79650 , n79651 , n79652 , n79653 , n79654 , n79655 , n79656 , n79657 , n79658 , 
 n79659 , n79660 , n79661 , n79662 , n79663 , n79664 , n79665 , n79666 , n79667 , n79668 , 
 n79669 , n79670 , n79671 , n79672 , n79673 , n79674 , n79675 , n79676 , n79677 , n79678 , 
 n79679 , n79680 , n79681 , n79682 , n79683 , n79684 , n79685 , n79686 , n79687 , n79688 , 
 n79689 , n79690 , n79691 , n79692 , n79693 , n79694 , n79695 , n79696 , n79697 , n79698 , 
 n79699 , n79700 , n79701 , n79702 , n79703 , n79704 , n79705 , n79706 , n79707 , n79708 , 
 n79709 , n79710 , n79711 , n79712 , n79713 , n79714 , n79715 , n79716 , n79717 , n79718 , 
 n79719 , n79720 , n79721 , n79722 , n79723 , n79724 , n79725 , n79726 , n79727 , n79728 , 
 n79729 , n79730 , n79731 , n79732 , n79733 , n79734 , n79735 , n79736 , n79737 , n79738 , 
 n79739 , n79740 , n79741 , n79742 , n79743 , n79744 , n79745 , n79746 , n79747 , n79748 , 
 n79749 , n79750 , n79751 , n79752 , n79753 , n79754 , n79755 , n79756 , n79757 , n79758 , 
 n79759 , n79760 , n79761 , n79762 , n79763 , n79764 , n79765 , n79766 , n79767 , n79768 , 
 n79769 , n79770 , n79771 , n79772 , n79773 , n79774 , n79775 , n79776 , n79777 , n79778 , 
 n79779 , n79780 , n79781 , n79782 , n79783 , n79784 , n79785 , n79786 , n79787 , n79788 , 
 n79789 , n79790 , n79791 , n79792 , n79793 , n79794 , n79795 , n79796 , n79797 , n79798 , 
 n79799 , n79800 , n79801 , n79802 , n79803 , n79804 , n79805 , n79806 , n79807 , n79808 , 
 n79809 , n79810 , n79811 , n79812 , n79813 , n79814 , n79815 , n79816 , n79817 , n79818 , 
 n79819 , n79820 , n79821 , n79822 , n79823 , n79824 , n79825 , n79826 , n79827 , n79828 , 
 n79829 , n79830 , n79831 , n79832 , n79833 , n79834 , n79835 , n79836 , n79837 , n79838 , 
 n79839 , n79840 , n79841 , n79842 , n79843 , n79844 , n79845 , n79846 , n79847 , n79848 , 
 n79849 , n79850 , n79851 , n79852 , n79853 , n79854 , n79855 , n79856 , n79857 , n79858 , 
 n79859 , n79860 , n79861 , n79862 , n79863 , n79864 , n79865 , n79866 , n79867 , n79868 , 
 n79869 , n79870 , n79871 , n79872 , n79873 , n79874 , n79875 , n79876 , n79877 , n79878 , 
 n79879 , n79880 , n79881 , n79882 , n79883 , n79884 , n79885 , n79886 , n79887 , n79888 , 
 n79889 , n79890 , n79891 , n79892 , n79893 , n79894 , n79895 , n79896 , n79897 , n79898 , 
 n79899 , n79900 , n79901 , n79902 , n79903 , n79904 , n79905 , n79906 , n79907 , n79908 , 
 n79909 , n79910 , n79911 , n79912 , n79913 , n79914 , n79915 , n79916 , n79917 , n79918 , 
 n79919 , n79920 , n79921 , n79922 , n79923 , n79924 , n79925 , n79926 , n79927 , n79928 , 
 n79929 , n79930 , n79931 , n79932 , n79933 , n79934 , n79935 , n79936 , n79937 , n79938 , 
 n79939 , n79940 , n79941 , n79942 , n79943 , n79944 , n79945 , n79946 , n79947 , n79948 , 
 n79949 , n79950 , n79951 , n79952 , n79953 , n79954 , n79955 , n79956 , n79957 , n79958 , 
 n79959 , n79960 , n79961 , n79962 , n79963 , n79964 , n79965 , n79966 , n79967 , n79968 , 
 n79969 , n79970 , n79971 , n79972 , n79973 , n79974 , n79975 , n79976 , n79977 , n79978 , 
 n79979 , n79980 , n79981 , n79982 , n79983 , n79984 , n79985 , n79986 , n79987 , n79988 , 
 n79989 , n79990 , n79991 , n79992 , n79993 , n79994 , n79995 , n79996 , n79997 , n79998 , 
 n79999 , n80000 , n80001 , n80002 , n80003 , n80004 , n80005 , n80006 , n80007 , n80008 , 
 n80009 , n80010 , n80011 , n80012 , n80013 , n80014 , n80015 , n80016 , n80017 , n80018 , 
 n80019 , n80020 , n80021 , n80022 , n80023 , n80024 , n80025 , n80026 , n80027 , n80028 , 
 n80029 , n80030 , n80031 , n80032 , n80033 , n80034 , n80035 , n80036 , n80037 , n80038 , 
 n80039 , n80040 , n80041 , n80042 , n80043 , n80044 , n80045 , n80046 , n80047 , n80048 , 
 n80049 , n80050 , n80051 , n80052 , n80053 , n80054 , n80055 , n80056 , n80057 , n80058 , 
 n80059 , n80060 , n80061 , n80062 , n80063 , n80064 , n80065 , n80066 , n80067 , n80068 , 
 n80069 , n80070 , n80071 , n80072 , n80073 , n80074 , n80075 , n80076 , n80077 , n80078 , 
 n80079 , n80080 , n80081 , n80082 , n80083 , n80084 , n80085 , n80086 , n80087 , n80088 , 
 n80089 , n80090 , n80091 , n80092 , n80093 , n80094 , n80095 , n80096 , n80097 , n80098 , 
 n80099 , n80100 , n80101 , n80102 , n80103 , n80104 , n80105 , n80106 , n80107 , n80108 , 
 n80109 , n80110 , n80111 , n80112 , n80113 , n80114 , n80115 , n80116 , n80117 , n80118 , 
 n80119 , n80120 , n80121 , n80122 , n80123 , n80124 , n80125 , n80126 , n80127 , n80128 , 
 n80129 , n80130 , n80131 , n80132 , n80133 , n80134 , n80135 , n80136 , n80137 , n80138 , 
 n80139 , n80140 , n80141 , n80142 , n80143 , n80144 , n80145 , n80146 , n80147 , n80148 , 
 n80149 , n80150 , n80151 , n80152 , n80153 , n80154 , n80155 , n80156 , n80157 , n80158 , 
 n80159 , n80160 , n80161 , n80162 , n80163 , n80164 , n80165 , n80166 , n80167 , n80168 , 
 n80169 , n80170 , n80171 , n80172 , n80173 , n80174 , n80175 , n80176 , n80177 , n80178 , 
 n80179 , n80180 , n80181 , n80182 , n80183 , n80184 , n80185 , n80186 , n80187 , n80188 , 
 n80189 , n80190 , n80191 , n80192 , n80193 , n80194 , n80195 , n80196 , n80197 , n80198 , 
 n80199 , n80200 , n80201 , n80202 , n80203 , n80204 , n80205 , n80206 , n80207 , n80208 , 
 n80209 , n80210 , n80211 , n80212 , n80213 , n80214 , n80215 , n80216 , n80217 , n80218 , 
 n80219 , n80220 , n80221 , n80222 , n80223 , n80224 , n80225 , n80226 , n80227 , n80228 , 
 n80229 , n80230 , n80231 , n80232 , n80233 , n80234 , n80235 , n80236 , n80237 , n80238 , 
 n80239 , n80240 , n80241 , n80242 , n80243 , n80244 , n80245 , n80246 , n80247 , n80248 , 
 n80249 , n80250 , n80251 , n80252 , n80253 , n80254 , n80255 , n80256 , n80257 , n80258 , 
 n80259 , n80260 , n80261 , n80262 , n80263 , n80264 , n80265 , n80266 , n80267 , n80268 , 
 n80269 , n80270 , n80271 , n80272 , n80273 , n80274 , n80275 , n80276 , n80277 , n80278 , 
 n80279 , n80280 , n80281 , n80282 , n80283 , n80284 , n80285 , n80286 , n80287 , n80288 , 
 n80289 , n80290 , n80291 , n80292 , n80293 , n80294 , n80295 , n80296 , n80297 , n80298 , 
 n80299 , n80300 , n80301 , n80302 , n80303 , n80304 , n80305 , n80306 , n80307 , n80308 , 
 n80309 , n80310 , n80311 , n80312 , n80313 , n80314 , n80315 , n80316 , n80317 , n80318 , 
 n80319 , n80320 , n80321 , n80322 , n80323 , n80324 , n80325 , n80326 , n80327 , n80328 , 
 n80329 , n80330 , n80331 , n80332 , n80333 , n80334 , n80335 , n80336 , n80337 , n80338 , 
 n80339 , n80340 , n80341 , n80342 , n80343 , n80344 , n80345 , n80346 , n80347 , n80348 , 
 n80349 , n80350 , n80351 , n80352 , n80353 , n80354 , n80355 , n80356 , n80357 , n80358 , 
 n80359 , n80360 , n80361 , n80362 , n80363 , n80364 , n80365 , n80366 , n80367 , n80368 , 
 n80369 , n80370 , n80371 , n80372 , n80373 , n80374 , n80375 , n80376 , n80377 , n80378 , 
 n80379 , n80380 , n80381 , n80382 , n80383 , n80384 , n80385 , n80386 , n80387 , n80388 , 
 n80389 , n80390 , n80391 , n80392 , n80393 , n80394 , n80395 , n80396 , n80397 , n80398 , 
 n80399 , n80400 , n80401 , n80402 , n80403 , n80404 , n80405 , n80406 , n80407 , n80408 , 
 n80409 , n80410 , n80411 , n80412 , n80413 , n80414 , n80415 , n80416 , n80417 , n80418 , 
 n80419 , n80420 , n80421 , n80422 , n80423 , n80424 , n80425 , n80426 , n80427 , n80428 , 
 n80429 , n80430 , n80431 , n80432 , n80433 , n80434 , n80435 , n80436 , n80437 , n80438 , 
 n80439 , n80440 , n80441 , n80442 , n80443 , n80444 , n80445 , n80446 , n80447 , n80448 , 
 n80449 , n80450 , n80451 , n80452 , n80453 , n80454 , n80455 , n80456 , n80457 , n80458 , 
 n80459 , n80460 , n80461 , n80462 , n80463 , n80464 , n80465 , n80466 , n80467 , n80468 , 
 n80469 , n80470 , n80471 , n80472 , n80473 , n80474 , n80475 , n80476 , n80477 , n80478 , 
 n80479 , n80480 , n80481 , n80482 , n80483 , n80484 , n80485 , n80486 , n80487 , n80488 , 
 n80489 , n80490 , n80491 , n80492 , n80493 , n80494 , n80495 , n80496 , n80497 , n80498 , 
 n80499 , n80500 , n80501 , n80502 , n80503 , n80504 , n80505 , n80506 , n80507 , n80508 , 
 n80509 , n80510 , n80511 , n80512 , n80513 , n80514 , n80515 , n80516 , n80517 , n80518 , 
 n80519 , n80520 , n80521 , n80522 , n80523 , n80524 , n80525 , n80526 , n80527 , n80528 , 
 n80529 , n80530 , n80531 , n80532 , n80533 , n80534 , n80535 , n80536 , n80537 , n80538 , 
 n80539 , n80540 , n80541 , n80542 , n80543 , n80544 , n80545 , n80546 , n80547 , n80548 , 
 n80549 , n80550 , n80551 , n80552 , n80553 , n80554 , n80555 , n80556 , n80557 , n80558 , 
 n80559 , n80560 , n80561 , n80562 , n80563 , n80564 , n80565 , n80566 , n80567 , n80568 , 
 n80569 , n80570 , n80571 , n80572 , n80573 , n80574 , n80575 , n80576 , n80577 , n80578 , 
 n80579 , n80580 , n80581 , n80582 , n80583 , n80584 , n80585 , n80586 , n80587 , n80588 , 
 n80589 , n80590 , n80591 , n80592 , n80593 , n80594 , n80595 , n80596 , n80597 , n80598 , 
 n80599 , n80600 , n80601 , n80602 , n80603 , n80604 , n80605 , n80606 , n80607 , n80608 , 
 n80609 , n80610 , n80611 , n80612 , n80613 , n80614 , n80615 , n80616 , n80617 , n80618 , 
 n80619 , n80620 , n80621 , n80622 , n80623 , n80624 , n80625 , n80626 , n80627 , n80628 , 
 n80629 , n80630 , n80631 , n80632 , n80633 , n80634 , n80635 , n80636 , n80637 , n80638 , 
 n80639 , n80640 , n80641 , n80642 , n80643 , n80644 , n80645 , n80646 , n80647 , n80648 , 
 n80649 , n80650 , n80651 , n80652 , n80653 , n80654 , n80655 , n80656 , n80657 , n80658 , 
 n80659 , n80660 , n80661 , n80662 , n80663 , n80664 , n80665 , n80666 , n80667 , n80668 , 
 n80669 , n80670 , n80671 , n80672 , n80673 , n80674 , n80675 , n80676 , n80677 , n80678 , 
 n80679 , n80680 , n80681 , n80682 , n80683 , n80684 , n80685 , n80686 , n80687 , n80688 , 
 n80689 , n80690 , n80691 , n80692 , n80693 , n80694 , n80695 , n80696 , n80697 , n80698 , 
 n80699 , n80700 , n80701 , n80702 , n80703 , n80704 , n80705 , n80706 , n80707 , n80708 , 
 n80709 , n80710 , n80711 , n80712 , n80713 , n80714 , n80715 , n80716 , n80717 , n80718 , 
 n80719 , n80720 , n80721 , n80722 , n80723 , n80724 , n80725 , n80726 , n80727 , n80728 , 
 n80729 , n80730 , n80731 , n80732 , n80733 , n80734 , n80735 , n80736 , n80737 , n80738 , 
 n80739 , n80740 , n80741 , n80742 , n80743 , n80744 , n80745 , n80746 , n80747 , n80748 , 
 n80749 , n80750 , n80751 , n80752 , n80753 , n80754 , n80755 , n80756 , n80757 , n80758 , 
 n80759 , n80760 , n80761 , n80762 , n80763 , n80764 , n80765 , n80766 , n80767 , n80768 , 
 n80769 , n80770 , n80771 , n80772 , n80773 , n80774 , n80775 , n80776 , n80777 , n80778 , 
 n80779 , n80780 , n80781 , n80782 , n80783 , n80784 , n80785 , n80786 , n80787 , n80788 , 
 n80789 , n80790 , n80791 , n80792 , n80793 , n80794 , n80795 , n80796 , n80797 , n80798 , 
 n80799 , n80800 , n80801 , n80802 , n80803 , n80804 , n80805 , n80806 , n80807 , n80808 , 
 n80809 , n80810 , n80811 , n80812 , n80813 , n80814 , n80815 , n80816 , n80817 , n80818 , 
 n80819 , n80820 , n80821 , n80822 , n80823 , n80824 , n80825 , n80826 , n80827 , n80828 , 
 n80829 , n80830 , n80831 , n80832 , n80833 , n80834 , n80835 , n80836 , n80837 , n80838 , 
 n80839 , n80840 , n80841 , n80842 , n80843 , n80844 , n80845 , n80846 , n80847 , n80848 , 
 n80849 , n80850 , n80851 , n80852 , n80853 , n80854 , n80855 , n80856 , n80857 , n80858 , 
 n80859 , n80860 , n80861 , n80862 , n80863 , n80864 , n80865 , n80866 , n80867 , n80868 , 
 n80869 , n80870 , n80871 , n80872 , n80873 , n80874 , n80875 , n80876 , n80877 , n80878 , 
 n80879 , n80880 , n80881 , n80882 , n80883 , n80884 , n80885 , n80886 , n80887 , n80888 , 
 n80889 , n80890 , n80891 , n80892 , n80893 , n80894 , n80895 , n80896 , n80897 , n80898 , 
 n80899 , n80900 , n80901 , n80902 , n80903 , n80904 , n80905 , n80906 , n80907 , n80908 , 
 n80909 , n80910 , n80911 , n80912 , n80913 , n80914 , n80915 , n80916 , n80917 , n80918 , 
 n80919 , n80920 , n80921 , n80922 , n80923 , n80924 , n80925 , n80926 , n80927 , n80928 , 
 n80929 , n80930 , n80931 , n80932 , n80933 , n80934 , n80935 , n80936 , n80937 , n80938 , 
 n80939 , n80940 , n80941 , n80942 , n80943 , n80944 , n80945 , n80946 , n80947 , n80948 , 
 n80949 , n80950 , n80951 , n80952 , n80953 , n80954 , n80955 , n80956 , n80957 , n80958 , 
 n80959 , n80960 , n80961 , n80962 , n80963 , n80964 , n80965 , n80966 , n80967 , n80968 , 
 n80969 , n80970 , n80971 , n80972 , n80973 , n80974 , n80975 , n80976 , n80977 , n80978 , 
 n80979 , n80980 , n80981 , n80982 , n80983 , n80984 , n80985 , n80986 , n80987 , n80988 , 
 n80989 , n80990 , n80991 , n80992 , n80993 , n80994 , n80995 , n80996 , n80997 , n80998 , 
 n80999 , n81000 , n81001 , n81002 , n81003 , n81004 , n81005 , n81006 , n81007 , n81008 , 
 n81009 , n81010 , n81011 , n81012 , n81013 , n81014 , n81015 , n81016 , n81017 , n81018 , 
 n81019 , n81020 , n81021 , n81022 , n81023 , n81024 , n81025 , n81026 , n81027 , n81028 , 
 n81029 , n81030 , n81031 , n81032 , n81033 , n81034 , n81035 , n81036 , n81037 , n81038 , 
 n81039 , n81040 , n81041 , n81042 , n81043 , n81044 , n81045 , n81046 , n81047 , n81048 , 
 n81049 , n81050 , n81051 , n81052 , n81053 , n81054 , n81055 , n81056 , n81057 , n81058 , 
 n81059 , n81060 , n81061 , n81062 , n81063 , n81064 , n81065 , n81066 , n81067 , n81068 , 
 n81069 , n81070 , n81071 , n81072 , n81073 , n81074 , n81075 , n81076 , n81077 , n81078 , 
 n81079 , n81080 , n81081 , n81082 , n81083 , n81084 , n81085 , n81086 , n81087 , n81088 , 
 n81089 , n81090 , n81091 , n81092 , n81093 , n81094 , n81095 , n81096 , n81097 , n81098 , 
 n81099 , n81100 , n81101 , n81102 , n81103 , n81104 , n81105 , n81106 , n81107 , n81108 , 
 n81109 , n81110 , n81111 , n81112 , n81113 , n81114 , n81115 , n81116 , n81117 , n81118 , 
 n81119 , n81120 , n81121 , n81122 , n81123 , n81124 , n81125 , n81126 , n81127 , n81128 , 
 n81129 , n81130 , n81131 , n81132 , n81133 , n81134 , n81135 , n81136 , n81137 , n81138 , 
 n81139 , n81140 , n81141 , n81142 , n81143 , n81144 , n81145 , n81146 , n81147 , n81148 , 
 n81149 , n81150 , n81151 , n81152 , n81153 , n81154 , n81155 , n81156 , n81157 , n81158 , 
 n81159 , n81160 , n81161 , n81162 , n81163 , n81164 , n81165 , n81166 , n81167 , n81168 , 
 n81169 , n81170 , n81171 , n81172 , n81173 , n81174 , n81175 , n81176 , n81177 , n81178 , 
 n81179 , n81180 , n81181 , n81182 , n81183 , n81184 , n81185 , n81186 , n81187 , n81188 , 
 n81189 , n81190 , n81191 , n81192 , n81193 , n81194 , n81195 , n81196 , n81197 , n81198 , 
 n81199 , n81200 , n81201 , n81202 , n81203 , n81204 , n81205 , n81206 , n81207 , n81208 , 
 n81209 , n81210 , n81211 , n81212 , n81213 , n81214 , n81215 , n81216 , n81217 , n81218 , 
 n81219 , n81220 , n81221 , n81222 , n81223 , n81224 , n81225 , n81226 , n81227 , n81228 , 
 n81229 , n81230 , n81231 , n81232 , n81233 , n81234 , n81235 , n81236 , n81237 , n81238 , 
 n81239 , n81240 , n81241 , n81242 , n81243 , n81244 , n81245 , n81246 , n81247 , n81248 , 
 n81249 , n81250 , n81251 , n81252 , n81253 , n81254 , n81255 , n81256 , n81257 , n81258 , 
 n81259 , n81260 , n81261 , n81262 , n81263 , n81264 , n81265 , n81266 , n81267 , n81268 , 
 n81269 , n81270 , n81271 , n81272 , n81273 , n81274 , n81275 , n81276 , n81277 , n81278 , 
 n81279 , n81280 , n81281 , n81282 , n81283 , n81284 , n81285 , n81286 , n81287 , n81288 , 
 n81289 , n81290 , n81291 , n81292 , n81293 , n81294 , n81295 , n81296 , n81297 , n81298 , 
 n81299 , n81300 , n81301 , n81302 , n81303 , n81304 , n81305 , n81306 , n81307 , n81308 , 
 n81309 , n81310 , n81311 , n81312 , n81313 , n81314 , n81315 , n81316 , n81317 , n81318 , 
 n81319 , n81320 , n81321 , n81322 , n81323 , n81324 , n81325 , n81326 , n81327 , n81328 , 
 n81329 , n81330 , n81331 , n81332 , n81333 , n81334 , n81335 , n81336 , n81337 , n81338 , 
 n81339 , n81340 , n81341 , n81342 , n81343 , n81344 , n81345 , n81346 , n81347 , n81348 , 
 n81349 , n81350 , n81351 , n81352 , n81353 , n81354 , n81355 , n81356 , n81357 , n81358 , 
 n81359 , n81360 , n81361 , n81362 , n81363 , n81364 , n81365 , n81366 , n81367 , n81368 , 
 n81369 , n81370 , n81371 , n81372 , n81373 , n81374 , n81375 , n81376 , n81377 , n81378 , 
 n81379 , n81380 , n81381 , n81382 , n81383 , n81384 , n81385 , n81386 , n81387 , n81388 , 
 n81389 , n81390 , n81391 , n81392 , n81393 , n81394 , n81395 , n81396 , n81397 , n81398 , 
 n81399 , n81400 , n81401 , n81402 , n81403 , n81404 , n81405 , n81406 , n81407 , n81408 , 
 n81409 , n81410 , n81411 , n81412 , n81413 , n81414 , n81415 , n81416 , n81417 , n81418 , 
 n81419 , n81420 , n81421 , n81422 , n81423 , n81424 , n81425 , n81426 , n81427 , n81428 , 
 n81429 , n81430 , n81431 , n81432 , n81433 , n81434 , n81435 , n81436 , n81437 , n81438 , 
 n81439 , n81440 , n81441 , n81442 , n81443 , n81444 , n81445 , n81446 , n81447 , n81448 , 
 n81449 , n81450 , n81451 , n81452 , n81453 , n81454 , n81455 , n81456 , n81457 , n81458 , 
 n81459 , n81460 , n81461 , n81462 , n81463 , n81464 , n81465 , n81466 , n81467 , n81468 , 
 n81469 , n81470 , n81471 , n81472 , n81473 , n81474 , n81475 , n81476 , n81477 , n81478 , 
 n81479 , n81480 , n81481 , n81482 , n81483 , n81484 , n81485 , n81486 , n81487 , n81488 , 
 n81489 , n81490 , n81491 , n81492 , n81493 , n81494 , n81495 , n81496 , n81497 , n81498 , 
 n81499 , n81500 , n81501 , n81502 , n81503 , n81504 , n81505 , n81506 , n81507 , n81508 , 
 n81509 , n81510 , n81511 , n81512 , n81513 , n81514 , n81515 , n81516 , n81517 , n81518 , 
 n81519 , n81520 , n81521 , n81522 , n81523 , n81524 , n81525 , n81526 , n81527 , n81528 , 
 n81529 , n81530 , n81531 , n81532 , n81533 , n81534 , n81535 , n81536 , n81537 , n81538 , 
 n81539 , n81540 , n81541 , n81542 , n81543 , n81544 , n81545 , n81546 , n81547 , n81548 , 
 n81549 , n81550 , n81551 , n81552 , n81553 , n81554 , n81555 , n81556 , n81557 , n81558 , 
 n81559 , n81560 , n81561 , n81562 , n81563 , n81564 , n81565 , n81566 , n81567 , n81568 , 
 n81569 , n81570 , n81571 , n81572 , n81573 , n81574 , n81575 , n81576 , n81577 , n81578 , 
 n81579 , n81580 , n81581 , n81582 , n81583 , n81584 , n81585 , n81586 , n81587 , n81588 , 
 n81589 , n81590 , n81591 , n81592 , n81593 , n81594 , n81595 , n81596 , n81597 , n81598 , 
 n81599 , n81600 , n81601 , n81602 , n81603 , n81604 , n81605 , n81606 , n81607 , n81608 , 
 n81609 , n81610 , n81611 , n81612 , n81613 , n81614 , n81615 , n81616 , n81617 , n81618 , 
 n81619 , n81620 , n81621 , n81622 , n81623 , n81624 , n81625 , n81626 , n81627 , n81628 , 
 n81629 , n81630 , n81631 , n81632 , n81633 , n81634 , n81635 , n81636 , n81637 , n81638 , 
 n81639 , n81640 , n81641 , n81642 , n81643 , n81644 , n81645 , n81646 , n81647 , n81648 , 
 n81649 , n81650 , n81651 , n81652 , n81653 , n81654 , n81655 , n81656 , n81657 , n81658 , 
 n81659 , n81660 , n81661 , n81662 , n81663 , n81664 , n81665 , n81666 , n81667 , n81668 , 
 n81669 , n81670 , n81671 , n81672 , n81673 , n81674 , n81675 , n81676 , n81677 , n81678 , 
 n81679 , n81680 , n81681 , n81682 , n81683 , n81684 , n81685 , n81686 , n81687 , n81688 , 
 n81689 , n81690 , n81691 , n81692 , n81693 , n81694 , n81695 , n81696 , n81697 , n81698 , 
 n81699 , n81700 , n81701 , n81702 , n81703 , n81704 , n81705 , n81706 , n81707 , n81708 , 
 n81709 , n81710 , n81711 , n81712 , n81713 , n81714 , n81715 , n81716 , n81717 , n81718 , 
 n81719 , n81720 , n81721 , n81722 , n81723 , n81724 , n81725 , n81726 , n81727 , n81728 , 
 n81729 , n81730 , n81731 , n81732 , n81733 , n81734 , n81735 , n81736 , n81737 , n81738 , 
 n81739 , n81740 , n81741 , n81742 , n81743 , n81744 , n81745 , n81746 , n81747 , n81748 , 
 n81749 , n81750 , n81751 , n81752 , n81753 , n81754 , n81755 , n81756 , n81757 , n81758 , 
 n81759 , n81760 , n81761 , n81762 , n81763 , n81764 , n81765 , n81766 , n81767 , n81768 , 
 n81769 , n81770 , n81771 , n81772 , n81773 , n81774 , n81775 , n81776 , n81777 , n81778 , 
 n81779 , n81780 , n81781 , n81782 , n81783 , n81784 , n81785 , n81786 , n81787 , n81788 , 
 n81789 , n81790 , n81791 , n81792 , n81793 , n81794 , n81795 , n81796 , n81797 , n81798 , 
 n81799 , n81800 , n81801 , n81802 , n81803 , n81804 , n81805 , n81806 , n81807 , n81808 , 
 n81809 , n81810 , n81811 , n81812 , n81813 , n81814 , n81815 , n81816 , n81817 , n81818 , 
 n81819 , n81820 , n81821 , n81822 , n81823 , n81824 , n81825 , n81826 , n81827 , n81828 , 
 n81829 , n81830 , n81831 , n81832 , n81833 , n81834 , n81835 , n81836 , n81837 , n81838 , 
 n81839 , n81840 , n81841 , n81842 , n81843 , n81844 , n81845 , n81846 , n81847 , n81848 , 
 n81849 , n81850 , n81851 , n81852 , n81853 , n81854 , n81855 , n81856 , n81857 , n81858 , 
 n81859 , n81860 , n81861 , n81862 , n81863 , n81864 , n81865 , n81866 , n81867 , n81868 , 
 n81869 , n81870 , n81871 , n81872 , n81873 , n81874 , n81875 , n81876 , n81877 , n81878 , 
 n81879 , n81880 , n81881 , n81882 , n81883 , n81884 , n81885 , n81886 , n81887 , n81888 , 
 n81889 , n81890 , n81891 , n81892 , n81893 , n81894 , n81895 , n81896 , n81897 , n81898 , 
 n81899 , n81900 , n81901 , n81902 , n81903 , n81904 , n81905 , n81906 , n81907 , n81908 , 
 n81909 , n81910 , n81911 , n81912 , n81913 , n81914 , n81915 , n81916 , n81917 , n81918 , 
 n81919 , n81920 , n81921 , n81922 , n81923 , n81924 , n81925 , n81926 , n81927 , n81928 , 
 n81929 , n81930 , n81931 , n81932 , n81933 , n81934 , n81935 , n81936 , n81937 , n81938 , 
 n81939 , n81940 , n81941 , n81942 , n81943 , n81944 , n81945 , n81946 , n81947 , n81948 , 
 n81949 , n81950 , n81951 , n81952 , n81953 , n81954 , n81955 , n81956 , n81957 , n81958 , 
 n81959 , n81960 , n81961 , n81962 , n81963 , n81964 , n81965 , n81966 , n81967 , n81968 , 
 n81969 , n81970 , n81971 , n81972 , n81973 , n81974 , n81975 , n81976 , n81977 , n81978 , 
 n81979 , n81980 , n81981 , n81982 , n81983 , n81984 , n81985 , n81986 , n81987 , n81988 , 
 n81989 , n81990 , n81991 , n81992 , n81993 , n81994 , n81995 , n81996 , n81997 , n81998 , 
 n81999 , n82000 , n82001 , n82002 , n82003 , n82004 , n82005 , n82006 , n82007 , n82008 , 
 n82009 , n82010 , n82011 , n82012 , n82013 , n82014 , n82015 , n82016 , n82017 , n82018 , 
 n82019 , n82020 , n82021 , n82022 , n82023 , n82024 , n82025 , n82026 , n82027 , n82028 , 
 n82029 , n82030 , n82031 , n82032 , n82033 , n82034 , n82035 , n82036 , n82037 , n82038 , 
 n82039 , n82040 , n82041 , n82042 , n82043 , n82044 , n82045 , n82046 , n82047 , n82048 , 
 n82049 , n82050 , n82051 , n82052 , n82053 , n82054 , n82055 , n82056 , n82057 , n82058 , 
 n82059 , n82060 , n82061 , n82062 , n82063 , n82064 , n82065 , n82066 , n82067 , n82068 , 
 n82069 , n82070 , n82071 , n82072 , n82073 , n82074 , n82075 , n82076 , n82077 , n82078 , 
 n82079 , n82080 , n82081 , n82082 , n82083 , n82084 , n82085 , n82086 , n82087 , n82088 , 
 n82089 , n82090 , n82091 , n82092 , n82093 , n82094 , n82095 , n82096 , n82097 , n82098 , 
 n82099 , n82100 , n82101 , n82102 , n82103 , n82104 , n82105 , n82106 , n82107 , n82108 , 
 n82109 , n82110 , n82111 , n82112 , n82113 , n82114 , n82115 , n82116 , n82117 , n82118 , 
 n82119 , n82120 , n82121 , n82122 , n82123 , n82124 , n82125 , n82126 , n82127 , n82128 , 
 n82129 , n82130 , n82131 , n82132 , n82133 , n82134 , n82135 , n82136 , n82137 , n82138 , 
 n82139 , n82140 , n82141 , n82142 , n82143 , n82144 , n82145 , n82146 , n82147 , n82148 , 
 n82149 , n82150 , n82151 , n82152 , n82153 , n82154 , n82155 , n82156 , n82157 , n82158 , 
 n82159 , n82160 , n82161 , n82162 , n82163 , n82164 , n82165 , n82166 , n82167 , n82168 , 
 n82169 , n82170 , n82171 , n82172 , n82173 , n82174 , n82175 , n82176 , n82177 , n82178 , 
 n82179 , n82180 , n82181 , n82182 , n82183 , n82184 , n82185 , n82186 , n82187 , n82188 , 
 n82189 , n82190 , n82191 , n82192 , n82193 , n82194 , n82195 , n82196 , n82197 , n82198 , 
 n82199 , n82200 , n82201 , n82202 , n82203 , n82204 , n82205 , n82206 , n82207 , n82208 , 
 n82209 , n82210 , n82211 , n82212 , n82213 , n82214 , n82215 , n82216 , n82217 , n82218 , 
 n82219 , n82220 , n82221 , n82222 , n82223 , n82224 , n82225 , n82226 , n82227 , n82228 , 
 n82229 , n82230 , n82231 , n82232 , n82233 , n82234 , n82235 , n82236 , n82237 , n82238 , 
 n82239 , n82240 , n82241 , n82242 , n82243 , n82244 , n82245 , n82246 , n82247 , n82248 , 
 n82249 , n82250 , n82251 , n82252 , n82253 , n82254 , n82255 , n82256 , n82257 , n82258 , 
 n82259 , n82260 , n82261 , n82262 , n82263 , n82264 , n82265 , n82266 , n82267 , n82268 , 
 n82269 , n82270 , n82271 , n82272 , n82273 , n82274 , n82275 , n82276 , n82277 , n82278 , 
 n82279 , n82280 , n82281 , n82282 , n82283 , n82284 , n82285 , n82286 , n82287 , n82288 , 
 n82289 , n82290 , n82291 , n82292 , n82293 , n82294 , n82295 , n82296 , n82297 , n82298 , 
 n82299 , n82300 , n82301 , n82302 , n82303 , n82304 , n82305 , n82306 , n82307 , n82308 , 
 n82309 , n82310 , n82311 , n82312 , n82313 , n82314 , n82315 , n82316 , n82317 , n82318 , 
 n82319 , n82320 , n82321 , n82322 , n82323 , n82324 , n82325 , n82326 , n82327 , n82328 , 
 n82329 , n82330 , n82331 , n82332 , n82333 , n82334 , n82335 , n82336 , n82337 , n82338 , 
 n82339 , n82340 , n82341 , n82342 , n82343 , n82344 , n82345 , n82346 , n82347 , n82348 , 
 n82349 , n82350 , n82351 , n82352 , n82353 , n82354 , n82355 , n82356 , n82357 , n82358 , 
 n82359 , n82360 , n82361 , n82362 , n82363 , n82364 , n82365 , n82366 , n82367 , n82368 , 
 n82369 , n82370 , n82371 , n82372 , n82373 , n82374 , n82375 , n82376 , n82377 , n82378 , 
 n82379 , n82380 , n82381 , n82382 , n82383 , n82384 , n82385 , n82386 , n82387 , n82388 , 
 n82389 , n82390 , n82391 , n82392 , n82393 , n82394 , n82395 , n82396 , n82397 , n82398 , 
 n82399 , n82400 , n82401 , n82402 , n82403 , n82404 , n82405 , n82406 , n82407 , n82408 , 
 n82409 , n82410 , n82411 , n82412 , n82413 , n82414 , n82415 , n82416 , n82417 , n82418 , 
 n82419 , n82420 , n82421 , n82422 , n82423 , n82424 , n82425 , n82426 , n82427 , n82428 , 
 n82429 , n82430 , n82431 , n82432 , n82433 , n82434 , n82435 , n82436 , n82437 , n82438 , 
 n82439 , n82440 , n82441 , n82442 , n82443 , n82444 , n82445 , n82446 , n82447 , n82448 , 
 n82449 , n82450 , n82451 , n82452 , n82453 , n82454 , n82455 , n82456 , n82457 , n82458 , 
 n82459 , n82460 , n82461 , n82462 , n82463 , n82464 , n82465 , n82466 , n82467 , n82468 , 
 n82469 , n82470 , n82471 , n82472 , n82473 , n82474 , n82475 , n82476 , n82477 , n82478 , 
 n82479 , n82480 , n82481 , n82482 , n82483 , n82484 , n82485 , n82486 , n82487 , n82488 , 
 n82489 , n82490 , n82491 , n82492 , n82493 , n82494 , n82495 , n82496 , n82497 , n82498 , 
 n82499 , n82500 , n82501 , n82502 , n82503 , n82504 , n82505 , n82506 , n82507 , n82508 , 
 n82509 , n82510 , n82511 , n82512 , n82513 , n82514 , n82515 , n82516 , n82517 , n82518 , 
 n82519 , n82520 , n82521 , n82522 , n82523 , n82524 , n82525 , n82526 , n82527 , n82528 , 
 n82529 , n82530 , n82531 , n82532 , n82533 , n82534 , n82535 , n82536 , n82537 , n82538 , 
 n82539 , n82540 , n82541 , n82542 , n82543 , n82544 , n82545 , n82546 , n82547 , n82548 , 
 n82549 , n82550 , n82551 , n82552 , n82553 , n82554 , n82555 , n82556 , n82557 , n82558 , 
 n82559 , n82560 , n82561 , n82562 , n82563 , n82564 , n82565 , n82566 , n82567 , n82568 , 
 n82569 , n82570 , n82571 , n82572 , n82573 , n82574 , n82575 , n82576 , n82577 , n82578 , 
 n82579 , n82580 , n82581 , n82582 , n82583 , n82584 , n82585 , n82586 , n82587 , n82588 , 
 n82589 , n82590 , n82591 , n82592 , n82593 , n82594 , n82595 , n82596 , n82597 , n82598 , 
 n82599 , n82600 , n82601 , n82602 , n82603 , n82604 , n82605 , n82606 , n82607 , n82608 , 
 n82609 , n82610 , n82611 , n82612 , n82613 , n82614 , n82615 , n82616 , n82617 , n82618 , 
 n82619 , n82620 , n82621 , n82622 , n82623 , n82624 , n82625 , n82626 , n82627 , n82628 , 
 n82629 , n82630 , n82631 , n82632 , n82633 , n82634 , n82635 , n82636 , n82637 , n82638 , 
 n82639 , n82640 , n82641 , n82642 , n82643 , n82644 , n82645 , n82646 , n82647 , n82648 , 
 n82649 , n82650 , n82651 , n82652 , n82653 , n82654 , n82655 , n82656 , n82657 , n82658 , 
 n82659 , n82660 , n82661 , n82662 , n82663 , n82664 , n82665 , n82666 , n82667 , n82668 , 
 n82669 , n82670 , n82671 , n82672 , n82673 , n82674 , n82675 , n82676 , n82677 , n82678 , 
 n82679 , n82680 , n82681 , n82682 , n82683 , n82684 , n82685 , n82686 , n82687 , n82688 , 
 n82689 , n82690 , n82691 , n82692 , n82693 , n82694 , n82695 , n82696 , n82697 , n82698 , 
 n82699 , n82700 , n82701 , n82702 , n82703 , n82704 , n82705 , n82706 , n82707 , n82708 , 
 n82709 , n82710 , n82711 , n82712 , n82713 , n82714 , n82715 , n82716 , n82717 , n82718 , 
 n82719 , n82720 , n82721 , n82722 , n82723 , n82724 , n82725 , n82726 , n82727 , n82728 , 
 n82729 , n82730 , n82731 , n82732 , n82733 , n82734 , n82735 , n82736 , n82737 , n82738 , 
 n82739 , n82740 , n82741 , n82742 , n82743 , n82744 , n82745 , n82746 , n82747 , n82748 , 
 n82749 , n82750 , n82751 , n82752 , n82753 , n82754 , n82755 , n82756 , n82757 , n82758 , 
 n82759 , n82760 , n82761 , n82762 , n82763 , n82764 , n82765 , n82766 , n82767 , n82768 , 
 n82769 , n82770 , n82771 , n82772 , n82773 , n82774 , n82775 , n82776 , n82777 , n82778 , 
 n82779 , n82780 , n82781 , n82782 , n82783 , n82784 , n82785 , n82786 , n82787 , n82788 , 
 n82789 , n82790 , n82791 , n82792 , n82793 , n82794 , n82795 , n82796 , n82797 , n82798 , 
 n82799 , n82800 , n82801 , n82802 , n82803 , n82804 , n82805 , n82806 , n82807 , n82808 , 
 n82809 , n82810 , n82811 , n82812 , n82813 , n82814 , n82815 , n82816 , n82817 , n82818 , 
 n82819 , n82820 , n82821 , n82822 , n82823 , n82824 , n82825 , n82826 , n82827 , n82828 , 
 n82829 , n82830 , n82831 , n82832 , n82833 , n82834 , n82835 , n82836 , n82837 , n82838 , 
 n82839 , n82840 , n82841 , n82842 , n82843 , n82844 , n82845 , n82846 , n82847 , n82848 , 
 n82849 , n82850 , n82851 , n82852 , n82853 , n82854 , n82855 , n82856 , n82857 , n82858 , 
 n82859 , n82860 , n82861 , n82862 , n82863 , n82864 , n82865 , n82866 , n82867 , n82868 , 
 n82869 , n82870 , n82871 , n82872 , n82873 , n82874 , n82875 , n82876 , n82877 , n82878 , 
 n82879 , n82880 , n82881 , n82882 , n82883 , n82884 , n82885 , n82886 , n82887 , n82888 , 
 n82889 , n82890 , n82891 , n82892 , n82893 , n82894 , n82895 , n82896 , n82897 , n82898 , 
 n82899 , n82900 , n82901 , n82902 , n82903 , n82904 , n82905 , n82906 , n82907 , n82908 , 
 n82909 , n82910 , n82911 , n82912 , n82913 , n82914 , n82915 , n82916 , n82917 , n82918 , 
 n82919 , n82920 , n82921 , n82922 , n82923 , n82924 , n82925 , n82926 , n82927 , n82928 , 
 n82929 , n82930 , n82931 , n82932 , n82933 , n82934 , n82935 , n82936 , n82937 , n82938 , 
 n82939 , n82940 , n82941 , n82942 , n82943 , n82944 , n82945 , n82946 , n82947 , n82948 , 
 n82949 , n82950 , n82951 , n82952 , n82953 , n82954 , n82955 , n82956 , n82957 , n82958 , 
 n82959 , n82960 , n82961 , n82962 , n82963 , n82964 , n82965 , n82966 , n82967 , n82968 , 
 n82969 , n82970 , n82971 , n82972 , n82973 , n82974 , n82975 , n82976 , n82977 , n82978 , 
 n82979 , n82980 , n82981 , n82982 , n82983 , n82984 , n82985 , n82986 , n82987 , n82988 , 
 n82989 , C0n , C0 ;
buf ( n768 , n0 );
buf ( n769 , n1 );
buf ( n770 , n2 );
buf ( n771 , n3 );
buf ( n772 , n4 );
buf ( n773 , n5 );
buf ( n774 , n6 );
buf ( n775 , n7 );
buf ( n776 , n8 );
buf ( n777 , n9 );
buf ( n778 , n10 );
buf ( n779 , n11 );
buf ( n780 , n12 );
buf ( n781 , n13 );
buf ( n782 , n14 );
buf ( n783 , n15 );
buf ( n784 , n16 );
buf ( n785 , n17 );
buf ( n786 , n18 );
buf ( n787 , n19 );
buf ( n788 , n20 );
buf ( n789 , n21 );
buf ( n790 , n22 );
buf ( n791 , n23 );
buf ( n792 , n24 );
buf ( n793 , n25 );
buf ( n794 , n26 );
buf ( n795 , n27 );
buf ( n796 , n28 );
buf ( n797 , n29 );
buf ( n798 , n30 );
buf ( n799 , n31 );
buf ( n800 , n32 );
buf ( n801 , n33 );
buf ( n802 , n34 );
buf ( n803 , n35 );
buf ( n804 , n36 );
buf ( n805 , n37 );
buf ( n806 , n38 );
buf ( n807 , n39 );
buf ( n808 , n40 );
buf ( n809 , n41 );
buf ( n810 , n42 );
buf ( n811 , n43 );
buf ( n812 , n44 );
buf ( n813 , n45 );
buf ( n814 , n46 );
buf ( n815 , n47 );
buf ( n816 , n48 );
buf ( n817 , n49 );
buf ( n818 , n50 );
buf ( n819 , n51 );
buf ( n820 , n52 );
buf ( n821 , n53 );
buf ( n822 , n54 );
buf ( n823 , n55 );
buf ( n824 , n56 );
buf ( n825 , n57 );
buf ( n826 , n58 );
buf ( n827 , n59 );
buf ( n828 , n60 );
buf ( n829 , n61 );
buf ( n830 , n62 );
buf ( n831 , n63 );
buf ( n832 , n64 );
buf ( n833 , n65 );
buf ( n834 , n66 );
buf ( n835 , n67 );
buf ( n836 , n68 );
buf ( n837 , n69 );
buf ( n838 , n70 );
buf ( n839 , n71 );
buf ( n840 , n72 );
buf ( n841 , n73 );
buf ( n842 , n74 );
buf ( n843 , n75 );
buf ( n844 , n76 );
buf ( n845 , n77 );
buf ( n846 , n78 );
buf ( n847 , n79 );
buf ( n848 , n80 );
buf ( n849 , n81 );
buf ( n850 , n82 );
buf ( n851 , n83 );
buf ( n852 , n84 );
buf ( n853 , n85 );
buf ( n854 , n86 );
buf ( n855 , n87 );
buf ( n856 , n88 );
buf ( n857 , n89 );
buf ( n858 , n90 );
buf ( n859 , n91 );
buf ( n860 , n92 );
buf ( n861 , n93 );
buf ( n862 , n94 );
buf ( n863 , n95 );
buf ( n864 , n96 );
buf ( n865 , n97 );
buf ( n866 , n98 );
buf ( n867 , n99 );
buf ( n868 , n100 );
buf ( n869 , n101 );
buf ( n870 , n102 );
buf ( n871 , n103 );
buf ( n872 , n104 );
buf ( n873 , n105 );
buf ( n874 , n106 );
buf ( n875 , n107 );
buf ( n876 , n108 );
buf ( n877 , n109 );
buf ( n878 , n110 );
buf ( n879 , n111 );
buf ( n880 , n112 );
buf ( n881 , n113 );
buf ( n882 , n114 );
buf ( n883 , n115 );
buf ( n884 , n116 );
buf ( n885 , n117 );
buf ( n886 , n118 );
buf ( n887 , n119 );
buf ( n888 , n120 );
buf ( n889 , n121 );
buf ( n890 , n122 );
buf ( n891 , n123 );
buf ( n892 , n124 );
buf ( n893 , n125 );
buf ( n894 , n126 );
buf ( n895 , n127 );
buf ( n128 , n896 );
buf ( n129 , n897 );
buf ( n130 , n898 );
buf ( n131 , n899 );
buf ( n132 , n900 );
buf ( n133 , n901 );
buf ( n134 , n902 );
buf ( n135 , n903 );
buf ( n136 , n904 );
buf ( n137 , n905 );
buf ( n138 , n906 );
buf ( n139 , n907 );
buf ( n140 , n908 );
buf ( n141 , n909 );
buf ( n142 , n910 );
buf ( n143 , n911 );
buf ( n144 , n912 );
buf ( n145 , n913 );
buf ( n146 , n914 );
buf ( n147 , n915 );
buf ( n148 , n916 );
buf ( n149 , n917 );
buf ( n150 , n918 );
buf ( n151 , n919 );
buf ( n152 , n920 );
buf ( n153 , n921 );
buf ( n154 , n922 );
buf ( n155 , n923 );
buf ( n156 , n924 );
buf ( n157 , n925 );
buf ( n158 , n926 );
buf ( n159 , n927 );
buf ( n160 , n928 );
buf ( n161 , n929 );
buf ( n162 , n930 );
buf ( n163 , n931 );
buf ( n164 , n932 );
buf ( n165 , n933 );
buf ( n166 , n934 );
buf ( n167 , n935 );
buf ( n168 , n936 );
buf ( n169 , n937 );
buf ( n170 , n938 );
buf ( n171 , n939 );
buf ( n172 , n940 );
buf ( n173 , n941 );
buf ( n174 , n942 );
buf ( n175 , n943 );
buf ( n176 , n944 );
buf ( n177 , n945 );
buf ( n178 , n946 );
buf ( n179 , n947 );
buf ( n180 , n948 );
buf ( n181 , n949 );
buf ( n182 , n950 );
buf ( n183 , n951 );
buf ( n184 , n952 );
buf ( n185 , n953 );
buf ( n186 , n954 );
buf ( n187 , n955 );
buf ( n188 , n956 );
buf ( n189 , n957 );
buf ( n190 , n958 );
buf ( n191 , n959 );
buf ( n192 , n960 );
buf ( n193 , n961 );
buf ( n194 , n962 );
buf ( n195 , n963 );
buf ( n196 , n964 );
buf ( n197 , n965 );
buf ( n198 , n966 );
buf ( n199 , n967 );
buf ( n200 , n968 );
buf ( n201 , n969 );
buf ( n202 , n970 );
buf ( n203 , n971 );
buf ( n204 , n972 );
buf ( n205 , n973 );
buf ( n206 , n974 );
buf ( n207 , n975 );
buf ( n208 , n976 );
buf ( n209 , n977 );
buf ( n210 , n978 );
buf ( n211 , n979 );
buf ( n212 , n980 );
buf ( n213 , n981 );
buf ( n214 , n982 );
buf ( n215 , n983 );
buf ( n216 , n984 );
buf ( n217 , n985 );
buf ( n218 , n986 );
buf ( n219 , n987 );
buf ( n220 , n988 );
buf ( n221 , n989 );
buf ( n222 , n990 );
buf ( n223 , n991 );
buf ( n224 , n992 );
buf ( n225 , n993 );
buf ( n226 , n994 );
buf ( n227 , n995 );
buf ( n228 , n996 );
buf ( n229 , n997 );
buf ( n230 , n998 );
buf ( n231 , n999 );
buf ( n232 , n1000 );
buf ( n233 , n1001 );
buf ( n234 , n1002 );
buf ( n235 , n1003 );
buf ( n236 , n1004 );
buf ( n237 , n1005 );
buf ( n238 , n1006 );
buf ( n239 , n1007 );
buf ( n240 , n1008 );
buf ( n241 , n1009 );
buf ( n242 , n1010 );
buf ( n243 , n1011 );
buf ( n244 , n1012 );
buf ( n245 , n1013 );
buf ( n246 , n1014 );
buf ( n247 , n1015 );
buf ( n248 , n1016 );
buf ( n249 , n1017 );
buf ( n250 , n1018 );
buf ( n251 , n1019 );
buf ( n252 , n1020 );
buf ( n253 , n1021 );
buf ( n254 , n1022 );
buf ( n255 , n1023 );
buf ( n256 , n1024 );
buf ( n257 , n1025 );
buf ( n258 , n1026 );
buf ( n259 , n1027 );
buf ( n260 , n1028 );
buf ( n261 , n1029 );
buf ( n262 , n1030 );
buf ( n263 , n1031 );
buf ( n264 , n1032 );
buf ( n265 , n1033 );
buf ( n266 , n1034 );
buf ( n267 , n1035 );
buf ( n268 , n1036 );
buf ( n269 , n1037 );
buf ( n270 , n1038 );
buf ( n271 , n1039 );
buf ( n272 , n1040 );
buf ( n273 , n1041 );
buf ( n274 , n1042 );
buf ( n275 , n1043 );
buf ( n276 , n1044 );
buf ( n277 , n1045 );
buf ( n278 , n1046 );
buf ( n279 , n1047 );
buf ( n280 , n1048 );
buf ( n281 , n1049 );
buf ( n282 , n1050 );
buf ( n283 , n1051 );
buf ( n284 , n1052 );
buf ( n285 , n1053 );
buf ( n286 , n1054 );
buf ( n287 , n1055 );
buf ( n288 , n1056 );
buf ( n289 , n1057 );
buf ( n290 , n1058 );
buf ( n291 , n1059 );
buf ( n292 , n1060 );
buf ( n293 , n1061 );
buf ( n294 , n1062 );
buf ( n295 , n1063 );
buf ( n296 , n1064 );
buf ( n297 , n1065 );
buf ( n298 , n1066 );
buf ( n299 , n1067 );
buf ( n300 , n1068 );
buf ( n301 , n1069 );
buf ( n302 , n1070 );
buf ( n303 , n1071 );
buf ( n304 , n1072 );
buf ( n305 , n1073 );
buf ( n306 , n1074 );
buf ( n307 , n1075 );
buf ( n308 , n1076 );
buf ( n309 , n1077 );
buf ( n310 , n1078 );
buf ( n311 , n1079 );
buf ( n312 , n1080 );
buf ( n313 , n1081 );
buf ( n314 , n1082 );
buf ( n315 , n1083 );
buf ( n316 , n1084 );
buf ( n317 , n1085 );
buf ( n318 , n1086 );
buf ( n319 , n1087 );
buf ( n320 , n1088 );
buf ( n321 , n1089 );
buf ( n322 , n1090 );
buf ( n323 , n1091 );
buf ( n324 , n1092 );
buf ( n325 , n1093 );
buf ( n326 , n1094 );
buf ( n327 , n1095 );
buf ( n328 , n1096 );
buf ( n329 , n1097 );
buf ( n330 , n1098 );
buf ( n331 , n1099 );
buf ( n332 , n1100 );
buf ( n333 , n1101 );
buf ( n334 , n1102 );
buf ( n335 , n1103 );
buf ( n336 , n1104 );
buf ( n337 , n1105 );
buf ( n338 , n1106 );
buf ( n339 , n1107 );
buf ( n340 , n1108 );
buf ( n341 , n1109 );
buf ( n342 , n1110 );
buf ( n343 , n1111 );
buf ( n344 , n1112 );
buf ( n345 , n1113 );
buf ( n346 , n1114 );
buf ( n347 , n1115 );
buf ( n348 , n1116 );
buf ( n349 , n1117 );
buf ( n350 , n1118 );
buf ( n351 , n1119 );
buf ( n352 , n1120 );
buf ( n353 , n1121 );
buf ( n354 , n1122 );
buf ( n355 , n1123 );
buf ( n356 , n1124 );
buf ( n357 , n1125 );
buf ( n358 , n1126 );
buf ( n359 , n1127 );
buf ( n360 , n1128 );
buf ( n361 , n1129 );
buf ( n362 , n1130 );
buf ( n363 , n1131 );
buf ( n364 , n1132 );
buf ( n365 , n1133 );
buf ( n366 , n1134 );
buf ( n367 , n1135 );
buf ( n368 , n1136 );
buf ( n369 , n1137 );
buf ( n370 , n1138 );
buf ( n371 , n1139 );
buf ( n372 , n1140 );
buf ( n373 , n1141 );
buf ( n374 , n1142 );
buf ( n375 , n1143 );
buf ( n376 , n1144 );
buf ( n377 , n1145 );
buf ( n378 , n1146 );
buf ( n379 , n1147 );
buf ( n380 , n1148 );
buf ( n381 , n1149 );
buf ( n382 , n1150 );
buf ( n383 , n1151 );
buf ( n896 , n42669 );
buf ( n897 , n42673 );
buf ( n898 , n82766 );
buf ( n899 , n42677 );
buf ( n900 , n42689 );
buf ( n901 , n42695 );
buf ( n902 , n43083 );
buf ( n903 , n42722 );
buf ( n904 , n42710 );
buf ( n905 , n43069 );
buf ( n906 , n43074 );
buf ( n907 , n43075 );
buf ( n908 , n43076 );
buf ( n909 , n43072 );
buf ( n910 , n43073 );
buf ( n911 , n42806 );
buf ( n912 , n43077 );
buf ( n913 , n43078 );
buf ( n914 , n43079 );
buf ( n915 , n42812 );
buf ( n916 , n43081 );
buf ( n917 , n43082 );
buf ( n918 , n82838 );
buf ( n919 , n42831 );
buf ( n920 , n43071 );
buf ( n921 , n42800 );
buf ( n922 , n42794 );
buf ( n923 , n42837 );
buf ( n924 , n43070 );
buf ( n925 , n42825 );
buf ( n926 , n42846 );
buf ( n927 , n42863 );
buf ( n928 , n42857 );
buf ( n929 , n82969 );
buf ( n930 , n42875 );
buf ( n931 , n42891 );
buf ( n932 , n43080 );
buf ( n933 , n82622 );
buf ( n934 , n42898 );
buf ( n935 , n42929 );
buf ( n936 , n82881 );
buf ( n937 , n82626 );
buf ( n938 , n42923 );
buf ( n939 , n82895 );
buf ( n940 , n42910 );
buf ( n941 , n42935 );
buf ( n942 , n42944 );
buf ( n943 , n42950 );
buf ( n944 , n42962 );
buf ( n945 , n42968 );
buf ( n946 , n42976 );
buf ( n947 , n42994 );
buf ( n948 , n42988 );
buf ( n949 , n43000 );
buf ( n950 , n43008 );
buf ( n951 , n43014 );
buf ( n952 , n43016 );
buf ( n953 , n43022 );
buf ( n954 , n43028 );
buf ( n955 , n43034 );
buf ( n956 , n82932 );
buf ( n957 , n43040 );
buf ( n958 , n43047 );
buf ( n959 , n82963 );
buf ( n960 , n82946 );
buf ( n961 , n44804 );
buf ( n962 , n82915 );
buf ( n963 , n45680 );
buf ( n964 , n44836 );
buf ( n965 , n45591 );
buf ( n966 , n82852 );
buf ( n967 , n45684 );
buf ( n968 , n82905 );
buf ( n969 , n45688 );
buf ( n970 , n45692 );
buf ( n971 , n45704 );
buf ( n972 , n45708 );
buf ( n973 , n45712 );
buf ( n974 , n45716 );
buf ( n975 , n45720 );
buf ( n976 , n45652 );
buf ( n977 , n45676 );
buf ( n978 , n45656 );
buf ( n979 , n45604 );
buf ( n980 , n45608 );
buf ( n981 , n82810 );
buf ( n982 , n45668 );
buf ( n983 , n82975 );
buf ( n984 , n45612 );
buf ( n985 , n45648 );
buf ( n986 , n45664 );
buf ( n987 , n45624 );
buf ( n988 , n82862 );
buf ( n989 , n45628 );
buf ( n990 , n45632 );
buf ( n991 , n45096 );
buf ( n992 , n45672 );
buf ( n993 , n45600 );
buf ( n994 , n82889 );
buf ( n995 , n45636 );
buf ( n996 , n45616 );
buf ( n997 , n45660 );
buf ( n998 , n45724 );
buf ( n999 , n45140 );
buf ( n1000 , n45700 );
buf ( n1001 , n45644 );
buf ( n1002 , n45620 );
buf ( n1003 , n45195 );
buf ( n1004 , n82790 );
buf ( n1005 , n45166 );
buf ( n1006 , n45215 );
buf ( n1007 , n45256 );
buf ( n1008 , n45241 );
buf ( n1009 , n45270 );
buf ( n1010 , n45289 );
buf ( n1011 , n45332 );
buf ( n1012 , n45318 );
buf ( n1013 , n45346 );
buf ( n1014 , n45372 );
buf ( n1015 , n45386 );
buf ( n1016 , n45389 );
buf ( n1017 , n45392 );
buf ( n1018 , n45395 );
buf ( n1019 , n45398 );
buf ( n1020 , n45401 );
buf ( n1021 , n45416 );
buf ( n1022 , n45438 );
buf ( n1023 , n82974 );
buf ( n1024 , n82674 );
buf ( n1025 , n82029 );
buf ( n1026 , n82052 );
buf ( n1027 , n81717 );
buf ( n1028 , n81463 );
buf ( n1029 , n82694 );
buf ( n1030 , n82773 );
buf ( n1031 , n82074 );
buf ( n1032 , n82740 );
buf ( n1033 , n81545 );
buf ( n1034 , n81882 );
buf ( n1035 , n81740 );
buf ( n1036 , n81858 );
buf ( n1037 , n82660 );
buf ( n1038 , n81584 );
buf ( n1039 , n81872 );
buf ( n1040 , n81616 );
buf ( n1041 , n81821 );
buf ( n1042 , n81837 );
buf ( n1043 , n81627 );
buf ( n1044 , n81806 );
buf ( n1045 , n81595 );
buf ( n1046 , n82962 );
buf ( n1047 , n81478 );
buf ( n1048 , n82611 );
buf ( n1049 , n81786 );
buf ( n1050 , n82628 );
buf ( n1051 , n82989 );
buf ( n1052 , n81645 );
buf ( n1053 , n81657 );
buf ( n1054 , n82627 );
buf ( n1055 , n81773 );
buf ( n1056 , n81759 );
buf ( n1057 , n82704 );
buf ( n1058 , n81901 );
buf ( n1059 , n81913 );
buf ( n1060 , n81924 );
buf ( n1061 , n82144 );
buf ( n1062 , n81508 );
buf ( n1063 , n81930 );
buf ( n1064 , n81677 );
buf ( n1065 , n81940 );
buf ( n1066 , n81691 );
buf ( n1067 , n81950 );
buf ( n1068 , n82138 );
buf ( n1069 , n81969 );
buf ( n1070 , n82576 );
buf ( n1071 , n82132 );
buf ( n1072 , n82170 );
buf ( n1073 , n82119 );
buf ( n1074 , n82956 );
buf ( n1075 , n81996 );
buf ( n1076 , n82099 );
buf ( n1077 , n82942 );
buf ( n1078 , n82633 );
buf ( n1079 , n82177 );
buf ( n1080 , n82093 );
buf ( n1081 , n82634 );
buf ( n1082 , n82208 );
buf ( n1083 , n82214 );
buf ( n1084 , n82195 );
buf ( n1085 , n82220 );
buf ( n1086 , n82164 );
buf ( n1087 , n82226 );
buf ( n1088 , n82239 );
buf ( n1089 , n82779 );
buf ( n1090 , n82256 );
buf ( n1091 , n82279 );
buf ( n1092 , n82273 );
buf ( n1093 , n82761 );
buf ( n1094 , n82293 );
buf ( n1095 , n82719 );
buf ( n1096 , n82308 );
buf ( n1097 , n82327 );
buf ( n1098 , n82320 );
buf ( n1099 , n82335 );
buf ( n1100 , n82724 );
buf ( n1101 , n82570 );
buf ( n1102 , n82349 );
buf ( n1103 , n82363 );
buf ( n1104 , n82729 );
buf ( n1105 , n82804 );
buf ( n1106 , n82573 );
buf ( n1107 , n82574 );
buf ( n1108 , n82376 );
buf ( n1109 , n82870 );
buf ( n1110 , n82577 );
buf ( n1111 , n82751 );
buf ( n1112 , n82844 );
buf ( n1113 , n82822 );
buf ( n1114 , n82581 );
buf ( n1115 , n82582 );
buf ( n1116 , n82831 );
buf ( n1117 , n82583 );
buf ( n1118 , n82585 );
buf ( n1119 , n82586 );
buf ( n1120 , n82587 );
buf ( n1121 , n82593 );
buf ( n1122 , n82970 );
buf ( n1123 , n82599 );
buf ( n1124 , n82709 );
buf ( n1125 , n82602 );
buf ( n1126 , n82926 );
buf ( n1127 , n82603 );
buf ( n1128 , n82610 );
buf ( n1129 , n82613 );
buf ( n1130 , n82615 );
buf ( n1131 , n82614 );
buf ( n1132 , n82578 );
buf ( n1133 , n82438 );
buf ( n1134 , n82798 );
buf ( n1135 , n82457 );
buf ( n1136 , n82468 );
buf ( n1137 , n82481 );
buf ( n1138 , n82635 );
buf ( n1139 , n82502 );
buf ( n1140 , n82512 );
buf ( n1141 , n82519 );
buf ( n1142 , n82528 );
buf ( n1143 , n82537 );
buf ( n1144 , n82543 );
buf ( n1145 , n82545 );
buf ( n1146 , n82547 );
buf ( n1147 , n82554 );
buf ( n1148 , n82556 );
buf ( n1149 , n82558 );
buf ( n1150 , n82560 );
buf ( n1151 , n80883 );
not ( n1152 , n831 );
not ( n1153 , n1152 );
buf ( n1154 , n799 );
not ( n1155 , n1154 );
buf ( n1156 , n1155 );
buf ( n1157 , n1156 );
not ( n1158 , n1157 );
not ( n1159 , n831 );
nand ( n1160 , n1159 , n830 );
not ( n1161 , n1160 );
buf ( n1162 , n1161 );
not ( n1163 , n1162 );
or ( n1164 , n1158 , n1163 );
buf ( n1165 , n798 );
buf ( n1166 , n830 );
xor ( n1167 , n1165 , n1166 );
buf ( n1168 , n1167 );
buf ( n1169 , n1168 );
buf ( n1170 , n831 );
nand ( n1171 , n1169 , n1170 );
buf ( n1172 , n1171 );
buf ( n1173 , n1172 );
nand ( n1174 , n1164 , n1173 );
buf ( n1175 , n1174 );
not ( n1176 , n1175 );
buf ( n1177 , n799 );
buf ( n1178 , n831 );
nand ( n1179 , n1177 , n1178 );
buf ( n1180 , n1179 );
buf ( n1181 , n1180 );
not ( n1182 , n1181 );
buf ( n1183 , n1182 );
and ( n1184 , n1183 , n895 );
buf ( n1185 , n894 );
buf ( n1186 , n1180 );
buf ( n1187 , n830 );
and ( n1188 , n1186 , n1187 );
buf ( n1189 , n1188 );
buf ( n1190 , n1189 );
xor ( n1191 , n1185 , n1190 );
buf ( n1192 , n1191 );
not ( n1193 , n1192 );
and ( n1194 , n1184 , n1193 );
not ( n1195 , n1184 );
and ( n1196 , n1195 , n1192 );
nor ( n1197 , n1194 , n1196 );
xor ( n1198 , n1176 , n1197 );
not ( n1199 , n1198 );
or ( n1200 , n1153 , n1199 );
nand ( n1201 , n1183 , n863 );
buf ( n1202 , n862 );
buf ( n1203 , n1189 );
xor ( n1204 , n1202 , n1203 );
buf ( n1205 , n1204 );
buf ( n1206 , n1205 );
not ( n1207 , n1206 );
buf ( n1208 , n1207 );
xor ( n1209 , n1201 , n1208 );
xor ( n1210 , n1209 , n1175 );
nand ( n1211 , n1210 , n831 );
nand ( n1212 , n1200 , n1211 );
buf ( n1213 , n1212 );
buf ( n1214 , n832 );
buf ( n1215 , n801 );
buf ( n1216 , n802 );
xor ( n1217 , n1215 , n1216 );
buf ( n1218 , n1217 );
buf ( n1219 , n1218 );
buf ( n1220 , n799 );
and ( n1221 , n1219 , n1220 );
buf ( n1222 , n1221 );
buf ( n1223 , n1222 );
buf ( n1224 , n772 );
buf ( n1225 , n828 );
xor ( n1226 , n1224 , n1225 );
buf ( n1227 , n1226 );
buf ( n1228 , n1227 );
not ( n1229 , n1228 );
buf ( n1230 , n829 );
buf ( n1231 , n830 );
xnor ( n1232 , n1230 , n1231 );
buf ( n1233 , n1232 );
buf ( n1234 , n828 );
buf ( n1235 , n829 );
xor ( n1236 , n1234 , n1235 );
buf ( n1237 , n1236 );
nand ( n1238 , n1233 , n1237 );
not ( n1239 , n1238 );
buf ( n1240 , n1239 );
not ( n1241 , n1240 );
or ( n1242 , n1229 , n1241 );
buf ( n1243 , n829 );
buf ( n1244 , n830 );
xor ( n1245 , n1243 , n1244 );
buf ( n1246 , n1245 );
buf ( n1247 , n1246 );
buf ( n1248 , n1247 );
buf ( n1249 , n1248 );
buf ( n1250 , n1249 );
buf ( n1251 , n771 );
buf ( n1252 , n828 );
xor ( n1253 , n1251 , n1252 );
buf ( n1254 , n1253 );
buf ( n1255 , n1254 );
nand ( n1256 , n1250 , n1255 );
buf ( n1257 , n1256 );
buf ( n1258 , n1257 );
nand ( n1259 , n1242 , n1258 );
buf ( n1260 , n1259 );
buf ( n1261 , n1260 );
xor ( n1262 , n1223 , n1261 );
buf ( n1263 , n770 );
buf ( n1264 , n830 );
xor ( n1265 , n1263 , n1264 );
buf ( n1266 , n1265 );
buf ( n1267 , n1266 );
not ( n1268 , n1267 );
buf ( n1269 , n1161 );
not ( n1270 , n1269 );
or ( n1271 , n1268 , n1270 );
buf ( n1272 , n769 );
buf ( n1273 , n830 );
xor ( n1274 , n1272 , n1273 );
buf ( n1275 , n1274 );
buf ( n1276 , n1275 );
buf ( n1277 , n831 );
nand ( n1278 , n1276 , n1277 );
buf ( n1279 , n1278 );
buf ( n1280 , n1279 );
nand ( n1281 , n1271 , n1280 );
buf ( n1282 , n1281 );
buf ( n1283 , n1282 );
xor ( n1284 , n1262 , n1283 );
buf ( n1285 , n1284 );
buf ( n1286 , n1285 );
buf ( n1287 , n792 );
buf ( n1288 , n808 );
xor ( n1289 , n1287 , n1288 );
buf ( n1290 , n1289 );
buf ( n1291 , n1290 );
not ( n1292 , n1291 );
buf ( n1293 , n809 );
buf ( n1294 , n810 );
xor ( n1295 , n1293 , n1294 );
buf ( n1296 , n1295 );
not ( n1297 , n1296 );
buf ( n1298 , n1297 );
xor ( n1299 , n809 , n808 );
buf ( n1300 , n1299 );
nand ( n1301 , n1298 , n1300 );
buf ( n1302 , n1301 );
buf ( n1303 , n1302 );
not ( n1304 , n1303 );
buf ( n1305 , n1304 );
buf ( n1306 , n1305 );
not ( n1307 , n1306 );
or ( n1308 , n1292 , n1307 );
buf ( n1309 , n1296 );
buf ( n1310 , n1309 );
buf ( n1311 , n791 );
buf ( n1312 , n808 );
xor ( n1313 , n1311 , n1312 );
buf ( n1314 , n1313 );
buf ( n1315 , n1314 );
nand ( n1316 , n1310 , n1315 );
buf ( n1317 , n1316 );
buf ( n1318 , n1317 );
nand ( n1319 , n1308 , n1318 );
buf ( n1320 , n1319 );
not ( n1321 , n780 );
and ( n1322 , n820 , n1321 );
not ( n1323 , n820 );
and ( n1324 , n1323 , n780 );
or ( n1325 , n1322 , n1324 );
not ( n1326 , n1325 );
buf ( n1327 , n821 );
not ( n1328 , n1327 );
buf ( n1329 , n822 );
nand ( n1330 , n1328 , n1329 );
buf ( n1331 , n1330 );
xor ( n1332 , n821 , n820 );
buf ( n1333 , n822 );
not ( n1334 , n1333 );
buf ( n1335 , n821 );
nand ( n1336 , n1334 , n1335 );
buf ( n1337 , n1336 );
and ( n1338 , n1331 , n1332 , n1337 );
not ( n1339 , n1338 );
or ( n1340 , n1326 , n1339 );
buf ( n1341 , n779 );
buf ( n1342 , n820 );
xor ( n1343 , n1341 , n1342 );
buf ( n1344 , n1343 );
xor ( n1345 , n821 , n822 );
buf ( n1346 , n1345 );
nand ( n1347 , n1344 , n1346 );
nand ( n1348 , n1340 , n1347 );
xor ( n1349 , n1320 , n1348 );
not ( n1350 , n826 );
nand ( n1351 , n1350 , n827 );
not ( n1352 , n827 );
nand ( n1353 , n1352 , n826 );
nand ( n1354 , n1351 , n1353 );
xnor ( n1355 , n828 , n827 );
and ( n1356 , n1354 , n1355 );
not ( n1357 , n1356 );
buf ( n1358 , n1357 );
buf ( n1359 , n774 );
buf ( n1360 , n826 );
xor ( n1361 , n1359 , n1360 );
buf ( n1362 , n1361 );
buf ( n1363 , n1362 );
not ( n1364 , n1363 );
buf ( n1365 , n1364 );
buf ( n1366 , n1365 );
or ( n1367 , n1358 , n1366 );
buf ( n1368 , n827 );
buf ( n1369 , n828 );
xor ( n1370 , n1368 , n1369 );
buf ( n1371 , n1370 );
buf ( n1372 , n1371 );
buf ( n1373 , n1372 );
buf ( n1374 , n1373 );
buf ( n1375 , n1374 );
xor ( n1376 , n826 , n773 );
buf ( n1377 , n1376 );
nand ( n1378 , n1375 , n1377 );
buf ( n1379 , n1378 );
buf ( n1380 , n1379 );
nand ( n1381 , n1367 , n1380 );
buf ( n1382 , n1381 );
xor ( n1383 , n1349 , n1382 );
buf ( n1384 , n1383 );
xor ( n1385 , n1286 , n1384 );
buf ( n1386 , n794 );
buf ( n1387 , n806 );
xor ( n1388 , n1386 , n1387 );
buf ( n1389 , n1388 );
buf ( n1390 , n1389 );
not ( n1391 , n1390 );
xor ( n1392 , n807 , n808 );
not ( n1393 , n1392 );
buf ( n1394 , n1393 );
and ( n1395 , n806 , n807 );
nor ( n1396 , n806 , n807 );
nor ( n1397 , n1395 , n1396 );
buf ( n1398 , n1397 );
nand ( n1399 , n1394 , n1398 );
buf ( n1400 , n1399 );
buf ( n1401 , n1400 );
not ( n1402 , n1401 );
buf ( n1403 , n1402 );
buf ( n1404 , n1403 );
not ( n1405 , n1404 );
or ( n1406 , n1391 , n1405 );
buf ( n1407 , n1393 );
not ( n1408 , n1407 );
buf ( n1409 , n1408 );
buf ( n1410 , n1409 );
buf ( n1411 , n793 );
buf ( n1412 , n806 );
xor ( n1413 , n1411 , n1412 );
buf ( n1414 , n1413 );
buf ( n1415 , n1414 );
nand ( n1416 , n1410 , n1415 );
buf ( n1417 , n1416 );
buf ( n1418 , n1417 );
nand ( n1419 , n1406 , n1418 );
buf ( n1420 , n1419 );
not ( n1421 , n1420 );
not ( n1422 , n1421 );
buf ( n1423 , n796 );
buf ( n1424 , n804 );
xor ( n1425 , n1423 , n1424 );
buf ( n1426 , n1425 );
buf ( n1427 , n1426 );
not ( n1428 , n1427 );
xnor ( n1429 , n804 , n805 );
buf ( n1430 , n805 );
buf ( n1431 , n806 );
xor ( n1432 , n1430 , n1431 );
buf ( n1433 , n1432 );
nor ( n1434 , n1429 , n1433 );
buf ( n1435 , n1434 );
not ( n1436 , n1435 );
buf ( n1437 , n1436 );
buf ( n1438 , n1437 );
not ( n1439 , n1438 );
buf ( n1440 , n1439 );
buf ( n1441 , n1440 );
not ( n1442 , n1441 );
or ( n1443 , n1428 , n1442 );
buf ( n1444 , n1433 );
not ( n1445 , n1444 );
buf ( n1446 , n1445 );
buf ( n1447 , n1446 );
not ( n1448 , n1447 );
buf ( n1449 , n1448 );
buf ( n1450 , n1449 );
buf ( n1451 , n795 );
buf ( n1452 , n804 );
xor ( n1453 , n1451 , n1452 );
buf ( n1454 , n1453 );
buf ( n1455 , n1454 );
nand ( n1456 , n1450 , n1455 );
buf ( n1457 , n1456 );
buf ( n1458 , n1457 );
nand ( n1459 , n1443 , n1458 );
buf ( n1460 , n1459 );
not ( n1461 , n1460 );
or ( n1462 , n1422 , n1461 );
not ( n1463 , n1460 );
nand ( n1464 , n1463 , n1420 );
nand ( n1465 , n1462 , n1464 );
buf ( n1466 , n782 );
buf ( n1467 , n818 );
xor ( n1468 , n1466 , n1467 );
buf ( n1469 , n1468 );
buf ( n1470 , n1469 );
not ( n1471 , n1470 );
or ( n1472 , n818 , n819 );
nand ( n1473 , n818 , n819 );
nand ( n1474 , n1472 , n1473 );
buf ( n1475 , n819 );
buf ( n1476 , n820 );
xor ( n1477 , n1475 , n1476 );
buf ( n1478 , n1477 );
nor ( n1479 , n1474 , n1478 );
buf ( n1480 , n1479 );
buf ( n1481 , n1480 );
not ( n1482 , n1481 );
buf ( n1483 , n1482 );
buf ( n1484 , n1483 );
not ( n1485 , n1484 );
buf ( n1486 , n1485 );
buf ( n1487 , n1486 );
not ( n1488 , n1487 );
or ( n1489 , n1471 , n1488 );
buf ( n1490 , n819 );
buf ( n1491 , n820 );
xor ( n1492 , n1490 , n1491 );
buf ( n1493 , n1492 );
buf ( n1494 , n1493 );
buf ( n1495 , n1494 );
buf ( n1496 , n1495 );
buf ( n1497 , n1496 );
xor ( n1498 , n818 , n781 );
buf ( n1499 , n1498 );
nand ( n1500 , n1497 , n1499 );
buf ( n1501 , n1500 );
buf ( n1502 , n1501 );
nand ( n1503 , n1489 , n1502 );
buf ( n1504 , n1503 );
and ( n1505 , n1465 , n1504 );
not ( n1506 , n1465 );
not ( n1507 , n1504 );
and ( n1508 , n1506 , n1507 );
nor ( n1509 , n1505 , n1508 );
buf ( n1510 , n1509 );
xor ( n1511 , n1385 , n1510 );
buf ( n1512 , n1511 );
buf ( n1513 , n1512 );
buf ( n1514 , n797 );
buf ( n1515 , n804 );
xor ( n1516 , n1514 , n1515 );
buf ( n1517 , n1516 );
buf ( n1518 , n1517 );
not ( n1519 , n1518 );
buf ( n1520 , n1437 );
not ( n1521 , n1520 );
buf ( n1522 , n1521 );
buf ( n1523 , n1522 );
not ( n1524 , n1523 );
or ( n1525 , n1519 , n1524 );
buf ( n1526 , n1446 );
not ( n1527 , n1526 );
buf ( n1528 , n1527 );
buf ( n1529 , n1528 );
buf ( n1530 , n1426 );
nand ( n1531 , n1529 , n1530 );
buf ( n1532 , n1531 );
buf ( n1533 , n1532 );
nand ( n1534 , n1525 , n1533 );
buf ( n1535 , n1534 );
buf ( n1536 , n1535 );
buf ( n1537 , n799 );
buf ( n1538 , n802 );
xor ( n1539 , n1537 , n1538 );
buf ( n1540 , n1539 );
buf ( n1541 , n1540 );
not ( n1542 , n1541 );
xnor ( n1543 , n802 , n803 );
buf ( n1544 , n803 );
buf ( n1545 , n804 );
xor ( n1546 , n1544 , n1545 );
buf ( n1547 , n1546 );
nor ( n1548 , n1543 , n1547 );
buf ( n1549 , n1548 );
buf ( n1550 , n1549 );
buf ( n1551 , n1550 );
buf ( n1552 , n1551 );
not ( n1553 , n1552 );
or ( n1554 , n1542 , n1553 );
buf ( n1555 , n1547 );
buf ( n1556 , n1555 );
buf ( n1557 , n1556 );
buf ( n1558 , n1557 );
buf ( n1559 , n1558 );
buf ( n1560 , n1559 );
buf ( n1561 , n1560 );
buf ( n1562 , n798 );
buf ( n1563 , n802 );
xor ( n1564 , n1562 , n1563 );
buf ( n1565 , n1564 );
buf ( n1566 , n1565 );
nand ( n1567 , n1561 , n1566 );
buf ( n1568 , n1567 );
buf ( n1569 , n1568 );
nand ( n1570 , n1554 , n1569 );
buf ( n1571 , n1570 );
buf ( n1572 , n1571 );
and ( n1573 , n1536 , n1572 );
not ( n1574 , n1536 );
buf ( n1575 , n1571 );
not ( n1576 , n1575 );
buf ( n1577 , n1576 );
buf ( n1578 , n1577 );
and ( n1579 , n1574 , n1578 );
nor ( n1580 , n1573 , n1579 );
buf ( n1581 , n1580 );
buf ( n1582 , n1581 );
buf ( n1583 , n771 );
buf ( n1584 , n830 );
xor ( n1585 , n1583 , n1584 );
buf ( n1586 , n1585 );
not ( n1587 , n1586 );
not ( n1588 , n1161 );
or ( n1589 , n1587 , n1588 );
buf ( n1590 , n1266 );
buf ( n1591 , n831 );
nand ( n1592 , n1590 , n1591 );
buf ( n1593 , n1592 );
nand ( n1594 , n1589 , n1593 );
buf ( n1595 , n799 );
buf ( n1596 , n803 );
or ( n1597 , n1595 , n1596 );
buf ( n1598 , n804 );
nand ( n1599 , n1597 , n1598 );
buf ( n1600 , n1599 );
buf ( n1601 , n1600 );
buf ( n1602 , n799 );
buf ( n1603 , n803 );
nand ( n1604 , n1602 , n1603 );
buf ( n1605 , n1604 );
buf ( n1606 , n1605 );
buf ( n1607 , n802 );
nand ( n1608 , n1601 , n1606 , n1607 );
buf ( n1609 , n1608 );
buf ( n1610 , n1609 );
not ( n1611 , n1610 );
buf ( n1612 , n1611 );
and ( n1613 , n1594 , n1612 );
not ( n1614 , n1594 );
and ( n1615 , n1614 , n1609 );
nor ( n1616 , n1613 , n1615 );
buf ( n1617 , n1616 );
buf ( n1618 , n1617 );
xor ( n1619 , n1582 , n1618 );
buf ( n1620 , n1619 );
buf ( n1621 , n1620 );
not ( n1622 , n1621 );
buf ( n1623 , n772 );
buf ( n1624 , n830 );
xor ( n1625 , n1623 , n1624 );
buf ( n1626 , n1625 );
buf ( n1627 , n1626 );
not ( n1628 , n1627 );
nand ( n1629 , n1159 , n830 );
not ( n1630 , n1629 );
buf ( n1631 , n1630 );
not ( n1632 , n1631 );
or ( n1633 , n1628 , n1632 );
buf ( n1634 , n1586 );
buf ( n1635 , n831 );
nand ( n1636 , n1634 , n1635 );
buf ( n1637 , n1636 );
buf ( n1638 , n1637 );
nand ( n1639 , n1633 , n1638 );
buf ( n1640 , n1639 );
buf ( n1641 , n792 );
buf ( n1642 , n810 );
xor ( n1643 , n1641 , n1642 );
buf ( n1644 , n1643 );
buf ( n1645 , n1644 );
not ( n1646 , n1645 );
not ( n1647 , n810 );
nand ( n1648 , n1647 , n811 );
not ( n1649 , n1648 );
buf ( n1650 , n811 );
not ( n1651 , n1650 );
buf ( n1652 , n810 );
nand ( n1653 , n1651 , n1652 );
buf ( n1654 , n1653 );
not ( n1655 , n1654 );
or ( n1656 , n1649 , n1655 );
buf ( n1657 , n811 );
buf ( n1658 , n812 );
xor ( n1659 , n1657 , n1658 );
buf ( n1660 , n1659 );
buf ( n1661 , n1660 );
not ( n1662 , n1661 );
buf ( n1663 , n1662 );
nand ( n1664 , n1656 , n1663 );
buf ( n1665 , n1664 );
buf ( n1666 , n1665 );
buf ( n1667 , n1666 );
buf ( n1668 , n1667 );
not ( n1669 , n1668 );
buf ( n1670 , n1669 );
buf ( n1671 , n1670 );
not ( n1672 , n1671 );
or ( n1673 , n1646 , n1672 );
buf ( n1674 , n1663 );
buf ( n1675 , n1674 );
buf ( n1676 , n1675 );
buf ( n1677 , n1676 );
not ( n1678 , n1677 );
buf ( n1679 , n1678 );
buf ( n1680 , n1679 );
buf ( n1681 , n791 );
buf ( n1682 , n810 );
xor ( n1683 , n1681 , n1682 );
buf ( n1684 , n1683 );
buf ( n1685 , n1684 );
nand ( n1686 , n1680 , n1685 );
buf ( n1687 , n1686 );
buf ( n1688 , n1687 );
nand ( n1689 , n1673 , n1688 );
buf ( n1690 , n1689 );
xor ( n1691 , n1640 , n1690 );
xor ( n1692 , n813 , n814 );
buf ( n1693 , n1692 );
buf ( n1694 , n1693 );
not ( n1695 , n1694 );
buf ( n1696 , n789 );
buf ( n1697 , n812 );
xor ( n1698 , n1696 , n1697 );
buf ( n1699 , n1698 );
buf ( n1700 , n1699 );
not ( n1701 , n1700 );
buf ( n1702 , n1701 );
or ( n1703 , n1695 , n1702 );
not ( n1704 , n812 );
not ( n1705 , n1704 );
nand ( n1706 , n813 , n814 );
not ( n1707 , n1706 );
not ( n1708 , n1707 );
or ( n1709 , n1705 , n1708 );
nor ( n1710 , n813 , n814 );
nand ( n1711 , n1710 , n812 );
nand ( n1712 , n1709 , n1711 );
not ( n1713 , n1712 );
not ( n1714 , n1713 );
buf ( n1715 , n790 );
buf ( n1716 , n812 );
xor ( n1717 , n1715 , n1716 );
buf ( n1718 , n1717 );
nand ( n1719 , n1714 , n1718 );
nand ( n1720 , n1703 , n1719 );
xor ( n1721 , n1691 , n1720 );
buf ( n1722 , n1721 );
not ( n1723 , n1722 );
buf ( n1724 , n798 );
buf ( n1725 , n804 );
xor ( n1726 , n1724 , n1725 );
buf ( n1727 , n1726 );
buf ( n1728 , n1727 );
not ( n1729 , n1728 );
xor ( n1730 , n806 , n805 );
and ( n1731 , n804 , n805 );
not ( n1732 , n804 );
not ( n1733 , n805 );
and ( n1734 , n1732 , n1733 );
nor ( n1735 , n1731 , n1734 );
not ( n1736 , n1735 );
nor ( n1737 , n1730 , n1736 );
buf ( n1738 , n1737 );
not ( n1739 , n1738 );
or ( n1740 , n1729 , n1739 );
buf ( n1741 , n1449 );
buf ( n1742 , n1517 );
nand ( n1743 , n1741 , n1742 );
buf ( n1744 , n1743 );
buf ( n1745 , n1744 );
nand ( n1746 , n1740 , n1745 );
buf ( n1747 , n1746 );
buf ( n1748 , n784 );
buf ( n1749 , n818 );
xor ( n1750 , n1748 , n1749 );
buf ( n1751 , n1750 );
buf ( n1752 , n1751 );
not ( n1753 , n1752 );
buf ( n1754 , n1480 );
not ( n1755 , n1754 );
or ( n1756 , n1753 , n1755 );
buf ( n1757 , n1496 );
buf ( n1758 , n783 );
buf ( n1759 , n818 );
xor ( n1760 , n1758 , n1759 );
buf ( n1761 , n1760 );
buf ( n1762 , n1761 );
nand ( n1763 , n1757 , n1762 );
buf ( n1764 , n1763 );
buf ( n1765 , n1764 );
nand ( n1766 , n1756 , n1765 );
buf ( n1767 , n1766 );
xor ( n1768 , n1747 , n1767 );
buf ( n1769 , n1371 );
buf ( n1770 , n1769 );
buf ( n1771 , n1770 );
not ( n1772 , n1771 );
xor ( n1773 , n826 , n775 );
not ( n1774 , n1773 );
or ( n1775 , n1772 , n1774 );
not ( n1776 , n1353 );
not ( n1777 , n1351 );
or ( n1778 , n1776 , n1777 );
nand ( n1779 , n1778 , n1355 );
not ( n1780 , n1779 );
buf ( n1781 , n1780 );
not ( n1782 , n1781 );
buf ( n1783 , n1782 );
buf ( n1784 , n776 );
buf ( n1785 , n826 );
xnor ( n1786 , n1784 , n1785 );
buf ( n1787 , n1786 );
or ( n1788 , n1783 , n1787 );
nand ( n1789 , n1775 , n1788 );
xor ( n1790 , n1768 , n1789 );
buf ( n1791 , n1790 );
not ( n1792 , n1791 );
or ( n1793 , n1723 , n1792 );
not ( n1794 , n1790 );
not ( n1795 , n1794 );
not ( n1796 , n1721 );
not ( n1797 , n1796 );
or ( n1798 , n1795 , n1797 );
buf ( n1799 , n1557 );
buf ( n1800 , n799 );
and ( n1801 , n1799 , n1800 );
buf ( n1802 , n1801 );
buf ( n1803 , n1239 );
buf ( n1804 , n774 );
buf ( n1805 , n828 );
xor ( n1806 , n1804 , n1805 );
buf ( n1807 , n1806 );
buf ( n1808 , n1807 );
and ( n1809 , n1803 , n1808 );
buf ( n1810 , n1249 );
buf ( n1811 , n773 );
buf ( n1812 , n828 );
xor ( n1813 , n1811 , n1812 );
buf ( n1814 , n1813 );
buf ( n1815 , n1814 );
and ( n1816 , n1810 , n1815 );
nor ( n1817 , n1809 , n1816 );
buf ( n1818 , n1817 );
not ( n1819 , n1818 );
xor ( n1820 , n1802 , n1819 );
buf ( n1821 , n778 );
buf ( n1822 , n824 );
xor ( n1823 , n1821 , n1822 );
buf ( n1824 , n1823 );
buf ( n1825 , n1824 );
not ( n1826 , n1825 );
and ( n1827 , n825 , n824 );
not ( n1828 , n825 );
not ( n1829 , n824 );
and ( n1830 , n1828 , n1829 );
nor ( n1831 , n1827 , n1830 );
not ( n1832 , n826 );
and ( n1833 , n825 , n1832 );
not ( n1834 , n825 );
and ( n1835 , n1834 , n826 );
nor ( n1836 , n1833 , n1835 );
nand ( n1837 , n1831 , n1836 );
not ( n1838 , n1837 );
buf ( n1839 , n1838 );
not ( n1840 , n1839 );
buf ( n1841 , n1840 );
buf ( n1842 , n1841 );
not ( n1843 , n1842 );
buf ( n1844 , n1843 );
buf ( n1845 , n1844 );
not ( n1846 , n1845 );
or ( n1847 , n1826 , n1846 );
buf ( n1848 , n777 );
buf ( n1849 , n824 );
xor ( n1850 , n1848 , n1849 );
buf ( n1851 , n1850 );
buf ( n1852 , n1851 );
buf ( n1853 , n825 );
buf ( n1854 , n826 );
xnor ( n1855 , n1853 , n1854 );
buf ( n1856 , n1855 );
buf ( n1857 , n1856 );
not ( n1858 , n1857 );
buf ( n1859 , n1858 );
buf ( n1860 , n1859 );
nand ( n1861 , n1852 , n1860 );
buf ( n1862 , n1861 );
buf ( n1863 , n1862 );
nand ( n1864 , n1847 , n1863 );
buf ( n1865 , n1864 );
xnor ( n1866 , n1820 , n1865 );
not ( n1867 , n1866 );
nand ( n1868 , n1798 , n1867 );
buf ( n1869 , n1868 );
nand ( n1870 , n1793 , n1869 );
buf ( n1871 , n1870 );
buf ( n1872 , n1871 );
not ( n1873 , n1872 );
or ( n1874 , n1622 , n1873 );
buf ( n1875 , n1871 );
buf ( n1876 , n1620 );
or ( n1877 , n1875 , n1876 );
buf ( n1878 , n799 );
buf ( n1879 , n805 );
or ( n1880 , n1878 , n1879 );
buf ( n1881 , n806 );
nand ( n1882 , n1880 , n1881 );
buf ( n1883 , n1882 );
buf ( n1884 , n1883 );
buf ( n1885 , n799 );
buf ( n1886 , n805 );
nand ( n1887 , n1885 , n1886 );
buf ( n1888 , n1887 );
buf ( n1889 , n1888 );
buf ( n1890 , n804 );
and ( n1891 , n1884 , n1889 , n1890 );
buf ( n1892 , n1891 );
buf ( n1893 , n1892 );
buf ( n1894 , n775 );
buf ( n1895 , n828 );
xor ( n1896 , n1894 , n1895 );
buf ( n1897 , n1896 );
buf ( n1898 , n1897 );
not ( n1899 , n1898 );
nand ( n1900 , n1233 , n1237 );
not ( n1901 , n1900 );
buf ( n1902 , n1901 );
not ( n1903 , n1902 );
or ( n1904 , n1899 , n1903 );
buf ( n1905 , n1249 );
buf ( n1906 , n1807 );
nand ( n1907 , n1905 , n1906 );
buf ( n1908 , n1907 );
buf ( n1909 , n1908 );
nand ( n1910 , n1904 , n1909 );
buf ( n1911 , n1910 );
buf ( n1912 , n1911 );
nand ( n1913 , n1893 , n1912 );
buf ( n1914 , n1913 );
buf ( n1915 , n1914 );
not ( n1916 , n1915 );
buf ( n1917 , n1916 );
buf ( n1918 , n1917 );
not ( n1919 , n1918 );
buf ( n1920 , n789 );
buf ( n1921 , n814 );
xor ( n1922 , n1920 , n1921 );
buf ( n1923 , n1922 );
buf ( n1924 , n1923 );
not ( n1925 , n1924 );
xnor ( n1926 , n814 , n815 );
xor ( n1927 , n815 , n816 );
nor ( n1928 , n1926 , n1927 );
buf ( n1929 , n1928 );
buf ( n1930 , n1929 );
buf ( n1931 , n1930 );
buf ( n1932 , n1931 );
not ( n1933 , n1932 );
or ( n1934 , n1925 , n1933 );
buf ( n1935 , n1927 );
buf ( n1936 , n1935 );
buf ( n1937 , n1936 );
buf ( n1938 , n1937 );
buf ( n1939 , n1938 );
buf ( n1940 , n1939 );
buf ( n1941 , n1940 );
buf ( n1942 , n788 );
buf ( n1943 , n814 );
xor ( n1944 , n1942 , n1943 );
buf ( n1945 , n1944 );
buf ( n1946 , n1945 );
nand ( n1947 , n1941 , n1946 );
buf ( n1948 , n1947 );
buf ( n1949 , n1948 );
nand ( n1950 , n1934 , n1949 );
buf ( n1951 , n1950 );
buf ( n1952 , n1951 );
not ( n1953 , n1952 );
buf ( n1954 , n779 );
buf ( n1955 , n824 );
xor ( n1956 , n1954 , n1955 );
buf ( n1957 , n1956 );
buf ( n1958 , n1957 );
not ( n1959 , n1958 );
and ( n1960 , n825 , n1832 );
not ( n1961 , n825 );
and ( n1962 , n1961 , n826 );
nor ( n1963 , n1960 , n1962 );
nand ( n1964 , n1963 , n1831 );
not ( n1965 , n1964 );
buf ( n1966 , n1965 );
not ( n1967 , n1966 );
or ( n1968 , n1959 , n1967 );
buf ( n1969 , n1824 );
buf ( n1970 , n1859 );
nand ( n1971 , n1969 , n1970 );
buf ( n1972 , n1971 );
buf ( n1973 , n1972 );
nand ( n1974 , n1968 , n1973 );
buf ( n1975 , n1974 );
buf ( n1976 , n1975 );
not ( n1977 , n1976 );
or ( n1978 , n1953 , n1977 );
buf ( n1979 , n1951 );
not ( n1980 , n1979 );
buf ( n1981 , n1980 );
buf ( n1982 , n1981 );
not ( n1983 , n1982 );
buf ( n1984 , n1975 );
not ( n1985 , n1984 );
buf ( n1986 , n1985 );
buf ( n1987 , n1986 );
not ( n1988 , n1987 );
or ( n1989 , n1983 , n1988 );
buf ( n1990 , n787 );
buf ( n1991 , n816 );
xor ( n1992 , n1990 , n1991 );
buf ( n1993 , n1992 );
buf ( n1994 , n1993 );
not ( n1995 , n1994 );
xnor ( n1996 , n817 , n816 );
buf ( n1997 , n817 );
buf ( n1998 , n818 );
xor ( n1999 , n1997 , n1998 );
buf ( n2000 , n1999 );
nor ( n2001 , n1996 , n2000 );
buf ( n2002 , n2001 );
buf ( n2003 , n2002 );
buf ( n2004 , n2003 );
buf ( n2005 , n2004 );
not ( n2006 , n2005 );
or ( n2007 , n1995 , n2006 );
buf ( n2008 , n2000 );
buf ( n2009 , n2008 );
buf ( n2010 , n2009 );
buf ( n2011 , n2010 );
buf ( n2012 , n786 );
buf ( n2013 , n816 );
xor ( n2014 , n2012 , n2013 );
buf ( n2015 , n2014 );
buf ( n2016 , n2015 );
nand ( n2017 , n2011 , n2016 );
buf ( n2018 , n2017 );
buf ( n2019 , n2018 );
nand ( n2020 , n2007 , n2019 );
buf ( n2021 , n2020 );
buf ( n2022 , n2021 );
nand ( n2023 , n1989 , n2022 );
buf ( n2024 , n2023 );
buf ( n2025 , n2024 );
nand ( n2026 , n1978 , n2025 );
buf ( n2027 , n2026 );
buf ( n2028 , n2027 );
not ( n2029 , n2028 );
or ( n2030 , n1919 , n2029 );
buf ( n2031 , n1914 );
not ( n2032 , n2031 );
buf ( n2033 , n2027 );
not ( n2034 , n2033 );
buf ( n2035 , n2034 );
buf ( n2036 , n2035 );
not ( n2037 , n2036 );
or ( n2038 , n2032 , n2037 );
buf ( n2039 , n793 );
buf ( n2040 , n810 );
xor ( n2041 , n2039 , n2040 );
buf ( n2042 , n2041 );
buf ( n2043 , n2042 );
not ( n2044 , n2043 );
buf ( n2045 , n1670 );
not ( n2046 , n2045 );
or ( n2047 , n2044 , n2046 );
buf ( n2048 , n1679 );
buf ( n2049 , n1644 );
nand ( n2050 , n2048 , n2049 );
buf ( n2051 , n2050 );
buf ( n2052 , n2051 );
nand ( n2053 , n2047 , n2052 );
buf ( n2054 , n2053 );
buf ( n2055 , n2054 );
buf ( n2056 , n791 );
buf ( n2057 , n812 );
xor ( n2058 , n2056 , n2057 );
buf ( n2059 , n2058 );
buf ( n2060 , n2059 );
not ( n2061 , n2060 );
not ( n2062 , n1704 );
not ( n2063 , n1707 );
or ( n2064 , n2062 , n2063 );
nand ( n2065 , n2064 , n1711 );
buf ( n2066 , n2065 );
buf ( n2067 , n2066 );
not ( n2068 , n2067 );
or ( n2069 , n2061 , n2068 );
buf ( n2070 , n1694 );
buf ( n2071 , n1718 );
nand ( n2072 , n2070 , n2071 );
buf ( n2073 , n2072 );
buf ( n2074 , n2073 );
nand ( n2075 , n2069 , n2074 );
buf ( n2076 , n2075 );
buf ( n2077 , n2076 );
xor ( n2078 , n2055 , n2077 );
buf ( n2079 , n781 );
buf ( n2080 , n822 );
xor ( n2081 , n2079 , n2080 );
buf ( n2082 , n2081 );
buf ( n2083 , n2082 );
not ( n2084 , n2083 );
and ( n2085 , n823 , n822 );
not ( n2086 , n823 );
not ( n2087 , n822 );
and ( n2088 , n2086 , n2087 );
nor ( n2089 , n2085 , n2088 );
buf ( n2090 , n2089 );
not ( n2091 , n2090 );
buf ( n2092 , n2091 );
buf ( n2093 , n823 );
buf ( n2094 , n824 );
xor ( n2095 , n2093 , n2094 );
buf ( n2096 , n2095 );
nor ( n2097 , n2092 , n2096 );
buf ( n2098 , n2097 );
buf ( n2099 , n2098 );
buf ( n2100 , n2099 );
buf ( n2101 , n2100 );
buf ( n2102 , n2101 );
not ( n2103 , n2102 );
or ( n2104 , n2084 , n2103 );
buf ( n2105 , n2096 );
buf ( n2106 , n2105 );
buf ( n2107 , n2106 );
buf ( n2108 , n2107 );
not ( n2109 , n2108 );
buf ( n2110 , n2109 );
buf ( n2111 , n2110 );
not ( n2112 , n2111 );
buf ( n2113 , n2112 );
buf ( n2114 , n2113 );
buf ( n2115 , n780 );
buf ( n2116 , n822 );
xor ( n2117 , n2115 , n2116 );
buf ( n2118 , n2117 );
buf ( n2119 , n2118 );
nand ( n2120 , n2114 , n2119 );
buf ( n2121 , n2120 );
buf ( n2122 , n2121 );
nand ( n2123 , n2104 , n2122 );
buf ( n2124 , n2123 );
buf ( n2125 , n2124 );
and ( n2126 , n2078 , n2125 );
and ( n2127 , n2055 , n2077 );
or ( n2128 , n2126 , n2127 );
buf ( n2129 , n2128 );
buf ( n2130 , n2129 );
nand ( n2131 , n2038 , n2130 );
buf ( n2132 , n2131 );
buf ( n2133 , n2132 );
nand ( n2134 , n2030 , n2133 );
buf ( n2135 , n2134 );
buf ( n2136 , n2135 );
nand ( n2137 , n1877 , n2136 );
buf ( n2138 , n2137 );
buf ( n2139 , n2138 );
nand ( n2140 , n1874 , n2139 );
buf ( n2141 , n2140 );
buf ( n2142 , n2141 );
xor ( n2143 , n1513 , n2142 );
not ( n2144 , n1865 );
not ( n2145 , n1802 );
or ( n2146 , n2144 , n2145 );
buf ( n2147 , n1818 );
buf ( n2148 , n1865 );
buf ( n2149 , n1802 );
nor ( n2150 , n2148 , n2149 );
buf ( n2151 , n2150 );
or ( n2152 , n2147 , n2151 );
nand ( n2153 , n2146 , n2152 );
xor ( n2154 , n1640 , n1690 );
and ( n2155 , n2154 , n1720 );
and ( n2156 , n1640 , n1690 );
or ( n2157 , n2155 , n2156 );
xor ( n2158 , n2153 , n2157 );
not ( n2159 , n2118 );
not ( n2160 , n2101 );
or ( n2161 , n2159 , n2160 );
buf ( n2162 , n2113 );
buf ( n2163 , n779 );
buf ( n2164 , n822 );
xor ( n2165 , n2163 , n2164 );
buf ( n2166 , n2165 );
buf ( n2167 , n2166 );
nand ( n2168 , n2162 , n2167 );
buf ( n2169 , n2168 );
nand ( n2170 , n2161 , n2169 );
not ( n2171 , n1945 );
not ( n2172 , n1931 );
or ( n2173 , n2171 , n2172 );
buf ( n2174 , n1940 );
buf ( n2175 , n787 );
buf ( n2176 , n814 );
xor ( n2177 , n2175 , n2176 );
buf ( n2178 , n2177 );
buf ( n2179 , n2178 );
nand ( n2180 , n2174 , n2179 );
buf ( n2181 , n2180 );
nand ( n2182 , n2173 , n2181 );
buf ( n2183 , n2182 );
nand ( n2184 , n2170 , n2183 );
or ( n2185 , n2183 , n2170 );
buf ( n2186 , n2015 );
not ( n2187 , n2186 );
buf ( n2188 , n2004 );
not ( n2189 , n2188 );
or ( n2190 , n2187 , n2189 );
buf ( n2191 , n2010 );
buf ( n2192 , n785 );
buf ( n2193 , n816 );
xor ( n2194 , n2192 , n2193 );
buf ( n2195 , n2194 );
buf ( n2196 , n2195 );
nand ( n2197 , n2191 , n2196 );
buf ( n2198 , n2197 );
buf ( n2199 , n2198 );
nand ( n2200 , n2190 , n2199 );
buf ( n2201 , n2200 );
nand ( n2202 , n2185 , n2201 );
nand ( n2203 , n2184 , n2202 );
xor ( n2204 , n2158 , n2203 );
buf ( n2205 , n2204 );
not ( n2206 , n831 );
and ( n2207 , n2206 , n830 );
not ( n2208 , n2207 );
buf ( n2209 , n773 );
buf ( n2210 , n830 );
xor ( n2211 , n2209 , n2210 );
buf ( n2212 , n2211 );
not ( n2213 , n2212 );
or ( n2214 , n2208 , n2213 );
buf ( n2215 , n1626 );
buf ( n2216 , n831 );
nand ( n2217 , n2215 , n2216 );
buf ( n2218 , n2217 );
nand ( n2219 , n2214 , n2218 );
not ( n2220 , n2219 );
buf ( n2221 , n2220 );
not ( n2222 , n2221 );
buf ( n2223 , n795 );
buf ( n2224 , n808 );
xor ( n2225 , n2223 , n2224 );
buf ( n2226 , n2225 );
buf ( n2227 , n2226 );
not ( n2228 , n2227 );
buf ( n2229 , n1297 );
buf ( n2230 , n1299 );
nand ( n2231 , n2229 , n2230 );
buf ( n2232 , n2231 );
buf ( n2233 , n2232 );
not ( n2234 , n2233 );
buf ( n2235 , n2234 );
buf ( n2236 , n2235 );
not ( n2237 , n2236 );
or ( n2238 , n2228 , n2237 );
buf ( n2239 , n794 );
buf ( n2240 , n808 );
xor ( n2241 , n2239 , n2240 );
buf ( n2242 , n2241 );
buf ( n2243 , n2242 );
buf ( n2244 , n1309 );
nand ( n2245 , n2243 , n2244 );
buf ( n2246 , n2245 );
buf ( n2247 , n2246 );
nand ( n2248 , n2238 , n2247 );
buf ( n2249 , n2248 );
not ( n2250 , n2249 );
buf ( n2251 , n2250 );
not ( n2252 , n2251 );
or ( n2253 , n2222 , n2252 );
buf ( n2254 , n783 );
buf ( n2255 , n820 );
xor ( n2256 , n2254 , n2255 );
buf ( n2257 , n2256 );
buf ( n2258 , n2257 );
not ( n2259 , n2258 );
not ( n2260 , n820 );
nor ( n2261 , n821 , n822 );
not ( n2262 , n2261 );
or ( n2263 , n2260 , n2262 );
not ( n2264 , n820 );
nand ( n2265 , n2264 , n821 , n822 );
nand ( n2266 , n2263 , n2265 );
buf ( n2267 , n2266 );
buf ( n2268 , n2267 );
not ( n2269 , n2268 );
or ( n2270 , n2259 , n2269 );
buf ( n2271 , n1346 );
buf ( n2272 , n782 );
buf ( n2273 , n820 );
xor ( n2274 , n2272 , n2273 );
buf ( n2275 , n2274 );
buf ( n2276 , n2275 );
nand ( n2277 , n2271 , n2276 );
buf ( n2278 , n2277 );
buf ( n2279 , n2278 );
nand ( n2280 , n2270 , n2279 );
buf ( n2281 , n2280 );
buf ( n2282 , n2281 );
nand ( n2283 , n2253 , n2282 );
buf ( n2284 , n2283 );
buf ( n2285 , n2284 );
buf ( n2286 , n2220 );
not ( n2287 , n2286 );
buf ( n2288 , n2249 );
nand ( n2289 , n2287 , n2288 );
buf ( n2290 , n2289 );
buf ( n2291 , n2290 );
nand ( n2292 , n2285 , n2291 );
buf ( n2293 , n2292 );
buf ( n2294 , n2293 );
buf ( n2295 , n799 );
buf ( n2296 , n804 );
xor ( n2297 , n2295 , n2296 );
buf ( n2298 , n2297 );
buf ( n2299 , n2298 );
not ( n2300 , n2299 );
buf ( n2301 , n1522 );
not ( n2302 , n2301 );
or ( n2303 , n2300 , n2302 );
buf ( n2304 , n1528 );
buf ( n2305 , n1727 );
nand ( n2306 , n2304 , n2305 );
buf ( n2307 , n2306 );
buf ( n2308 , n2307 );
nand ( n2309 , n2303 , n2308 );
buf ( n2310 , n2309 );
buf ( n2311 , n2310 );
not ( n2312 , n2311 );
buf ( n2313 , n797 );
buf ( n2314 , n806 );
xor ( n2315 , n2313 , n2314 );
buf ( n2316 , n2315 );
buf ( n2317 , n2316 );
not ( n2318 , n2317 );
buf ( n2319 , n1393 );
buf ( n2320 , n1397 );
nand ( n2321 , n2319 , n2320 );
buf ( n2322 , n2321 );
buf ( n2323 , n2322 );
not ( n2324 , n2323 );
buf ( n2325 , n2324 );
buf ( n2326 , n2325 );
not ( n2327 , n2326 );
or ( n2328 , n2318 , n2327 );
buf ( n2329 , n1393 );
not ( n2330 , n2329 );
buf ( n2331 , n2330 );
buf ( n2332 , n2331 );
buf ( n2333 , n796 );
buf ( n2334 , n806 );
xor ( n2335 , n2333 , n2334 );
buf ( n2336 , n2335 );
buf ( n2337 , n2336 );
nand ( n2338 , n2332 , n2337 );
buf ( n2339 , n2338 );
buf ( n2340 , n2339 );
nand ( n2341 , n2328 , n2340 );
buf ( n2342 , n2341 );
buf ( n2343 , n2342 );
not ( n2344 , n2343 );
or ( n2345 , n2312 , n2344 );
buf ( n2346 , n2310 );
not ( n2347 , n2346 );
buf ( n2348 , n2347 );
buf ( n2349 , n2348 );
not ( n2350 , n2349 );
buf ( n2351 , n2342 );
not ( n2352 , n2351 );
buf ( n2353 , n2352 );
buf ( n2354 , n2353 );
not ( n2355 , n2354 );
or ( n2356 , n2350 , n2355 );
not ( n2357 , n1351 );
not ( n2358 , n1353 );
or ( n2359 , n2357 , n2358 );
xnor ( n2360 , n828 , n827 );
nand ( n2361 , n2359 , n2360 );
buf ( n2362 , n2361 );
not ( n2363 , n2362 );
buf ( n2364 , n2363 );
not ( n2365 , n2364 );
xor ( n2366 , n777 , n826 );
not ( n2367 , n2366 );
or ( n2368 , n2365 , n2367 );
buf ( n2369 , n1374 );
not ( n2370 , n2369 );
buf ( n2371 , n2370 );
or ( n2372 , n1787 , n2371 );
nand ( n2373 , n2368 , n2372 );
buf ( n2374 , n2373 );
nand ( n2375 , n2356 , n2374 );
buf ( n2376 , n2375 );
buf ( n2377 , n2376 );
nand ( n2378 , n2345 , n2377 );
buf ( n2379 , n2378 );
buf ( n2380 , n2379 );
xor ( n2381 , n2294 , n2380 );
buf ( n2382 , n2170 );
not ( n2383 , n2382 );
not ( n2384 , n2182 );
buf ( n2385 , n2384 );
not ( n2386 , n2385 );
buf ( n2387 , n2201 );
not ( n2388 , n2387 );
and ( n2389 , n2386 , n2388 );
buf ( n2390 , n2201 );
buf ( n2391 , n2384 );
and ( n2392 , n2390 , n2391 );
nor ( n2393 , n2389 , n2392 );
buf ( n2394 , n2393 );
buf ( n2395 , n2394 );
not ( n2396 , n2395 );
or ( n2397 , n2383 , n2396 );
buf ( n2398 , n2394 );
buf ( n2399 , n2170 );
or ( n2400 , n2398 , n2399 );
nand ( n2401 , n2397 , n2400 );
buf ( n2402 , n2401 );
buf ( n2403 , n2402 );
and ( n2404 , n2381 , n2403 );
and ( n2405 , n2294 , n2380 );
or ( n2406 , n2404 , n2405 );
buf ( n2407 , n2406 );
buf ( n2408 , n2407 );
xor ( n2409 , n2205 , n2408 );
buf ( n2410 , n2266 );
not ( n2411 , n2410 );
not ( n2412 , n2275 );
or ( n2413 , n2411 , n2412 );
buf ( n2414 , n1345 );
buf ( n2415 , n781 );
buf ( n2416 , n820 );
xor ( n2417 , n2415 , n2416 );
buf ( n2418 , n2417 );
buf ( n2419 , n2418 );
nand ( n2420 , n2414 , n2419 );
buf ( n2421 , n2420 );
nand ( n2422 , n2413 , n2421 );
buf ( n2423 , n2422 );
buf ( n2424 , n2242 );
not ( n2425 , n2424 );
buf ( n2426 , n2235 );
not ( n2427 , n2426 );
or ( n2428 , n2425 , n2427 );
buf ( n2429 , n1309 );
buf ( n2430 , n793 );
buf ( n2431 , n808 );
xor ( n2432 , n2430 , n2431 );
buf ( n2433 , n2432 );
buf ( n2434 , n2433 );
nand ( n2435 , n2429 , n2434 );
buf ( n2436 , n2435 );
buf ( n2437 , n2436 );
nand ( n2438 , n2428 , n2437 );
buf ( n2439 , n2438 );
buf ( n2440 , n2439 );
or ( n2441 , n2423 , n2440 );
buf ( n2442 , n2336 );
not ( n2443 , n2442 );
buf ( n2444 , n1403 );
not ( n2445 , n2444 );
or ( n2446 , n2443 , n2445 );
buf ( n2447 , n1409 );
buf ( n2448 , n2447 );
buf ( n2449 , n2448 );
buf ( n2450 , n2449 );
buf ( n2451 , n795 );
buf ( n2452 , n806 );
xor ( n2453 , n2451 , n2452 );
buf ( n2454 , n2453 );
buf ( n2455 , n2454 );
nand ( n2456 , n2450 , n2455 );
buf ( n2457 , n2456 );
buf ( n2458 , n2457 );
nand ( n2459 , n2446 , n2458 );
buf ( n2460 , n2459 );
buf ( n2461 , n2460 );
nand ( n2462 , n2441 , n2461 );
buf ( n2463 , n2462 );
buf ( n2464 , n2463 );
buf ( n2465 , n2422 );
buf ( n2466 , n2439 );
nand ( n2467 , n2465 , n2466 );
buf ( n2468 , n2467 );
buf ( n2469 , n2468 );
nand ( n2470 , n2464 , n2469 );
buf ( n2471 , n2470 );
buf ( n2472 , n2471 );
xor ( n2473 , n1747 , n1767 );
and ( n2474 , n2473 , n1789 );
and ( n2475 , n1747 , n1767 );
or ( n2476 , n2474 , n2475 );
buf ( n2477 , n2476 );
xor ( n2478 , n2472 , n2477 );
buf ( n2479 , n1851 );
not ( n2480 , n2479 );
buf ( n2481 , n1838 );
buf ( n2482 , n2481 );
buf ( n2483 , n2482 );
buf ( n2484 , n2483 );
not ( n2485 , n2484 );
or ( n2486 , n2480 , n2485 );
buf ( n2487 , n1856 );
buf ( n2488 , n2487 );
buf ( n2489 , n2488 );
buf ( n2490 , n2489 );
not ( n2491 , n2490 );
buf ( n2492 , n2491 );
buf ( n2493 , n2492 );
buf ( n2494 , n776 );
buf ( n2495 , n824 );
xor ( n2496 , n2494 , n2495 );
buf ( n2497 , n2496 );
buf ( n2498 , n2497 );
nand ( n2499 , n2493 , n2498 );
buf ( n2500 , n2499 );
buf ( n2501 , n2500 );
nand ( n2502 , n2486 , n2501 );
buf ( n2503 , n2502 );
buf ( n2504 , n2503 );
buf ( n2505 , n1814 );
not ( n2506 , n2505 );
buf ( n2507 , n1901 );
not ( n2508 , n2507 );
or ( n2509 , n2506 , n2508 );
buf ( n2510 , n1249 );
buf ( n2511 , n1227 );
nand ( n2512 , n2510 , n2511 );
buf ( n2513 , n2512 );
buf ( n2514 , n2513 );
nand ( n2515 , n2509 , n2514 );
buf ( n2516 , n2515 );
buf ( n2517 , n2516 );
xor ( n2518 , n2504 , n2517 );
buf ( n2519 , n2195 );
not ( n2520 , n2519 );
buf ( n2521 , n2001 );
buf ( n2522 , n2521 );
buf ( n2523 , n2522 );
buf ( n2524 , n2523 );
buf ( n2525 , n2524 );
buf ( n2526 , n2525 );
buf ( n2527 , n2526 );
not ( n2528 , n2527 );
or ( n2529 , n2520 , n2528 );
buf ( n2530 , n2000 );
buf ( n2531 , n2530 );
buf ( n2532 , n2531 );
buf ( n2533 , n2532 );
buf ( n2534 , n2533 );
buf ( n2535 , n2534 );
buf ( n2536 , n2535 );
buf ( n2537 , n784 );
buf ( n2538 , n816 );
xor ( n2539 , n2537 , n2538 );
buf ( n2540 , n2539 );
buf ( n2541 , n2540 );
nand ( n2542 , n2536 , n2541 );
buf ( n2543 , n2542 );
buf ( n2544 , n2543 );
nand ( n2545 , n2529 , n2544 );
buf ( n2546 , n2545 );
buf ( n2547 , n2546 );
xor ( n2548 , n2518 , n2547 );
buf ( n2549 , n2548 );
buf ( n2550 , n2549 );
xor ( n2551 , n2478 , n2550 );
buf ( n2552 , n2551 );
buf ( n2553 , n2552 );
and ( n2554 , n2409 , n2553 );
and ( n2555 , n2205 , n2408 );
or ( n2556 , n2554 , n2555 );
buf ( n2557 , n2556 );
buf ( n2558 , n2557 );
xor ( n2559 , n2143 , n2558 );
buf ( n2560 , n2559 );
buf ( n2561 , n2560 );
xor ( n2562 , n2205 , n2408 );
xor ( n2563 , n2562 , n2553 );
buf ( n2564 , n2563 );
buf ( n2565 , n2564 );
not ( n2566 , n2565 );
xor ( n2567 , n1620 , n2135 );
xnor ( n2568 , n2567 , n1871 );
buf ( n2569 , n2568 );
nand ( n2570 , n2566 , n2569 );
buf ( n2571 , n2570 );
buf ( n2572 , n2571 );
not ( n2573 , n2572 );
buf ( n2574 , n2166 );
not ( n2575 , n2574 );
xnor ( n2576 , n822 , n823 );
nor ( n2577 , n2576 , n2096 );
buf ( n2578 , n2577 );
not ( n2579 , n2578 );
or ( n2580 , n2575 , n2579 );
buf ( n2581 , n2107 );
buf ( n2582 , n778 );
buf ( n2583 , n822 );
xor ( n2584 , n2582 , n2583 );
buf ( n2585 , n2584 );
buf ( n2586 , n2585 );
nand ( n2587 , n2581 , n2586 );
buf ( n2588 , n2587 );
buf ( n2589 , n2588 );
nand ( n2590 , n2580 , n2589 );
buf ( n2591 , n2590 );
buf ( n2592 , n2591 );
buf ( n2593 , n1699 );
not ( n2594 , n2593 );
buf ( n2595 , n2066 );
not ( n2596 , n2595 );
or ( n2597 , n2594 , n2596 );
buf ( n2598 , n1693 );
xor ( n2599 , n812 , n788 );
buf ( n2600 , n2599 );
nand ( n2601 , n2598 , n2600 );
buf ( n2602 , n2601 );
buf ( n2603 , n2602 );
nand ( n2604 , n2597 , n2603 );
buf ( n2605 , n2604 );
buf ( n2606 , n2605 );
xor ( n2607 , n2592 , n2606 );
buf ( n2608 , n2178 );
not ( n2609 , n2608 );
buf ( n2610 , n1931 );
buf ( n2611 , n2610 );
buf ( n2612 , n2611 );
buf ( n2613 , n2612 );
not ( n2614 , n2613 );
or ( n2615 , n2609 , n2614 );
buf ( n2616 , n1937 );
not ( n2617 , n2616 );
buf ( n2618 , n2617 );
buf ( n2619 , n2618 );
not ( n2620 , n2619 );
buf ( n2621 , n2620 );
buf ( n2622 , n2621 );
buf ( n2623 , n786 );
buf ( n2624 , n814 );
xor ( n2625 , n2623 , n2624 );
buf ( n2626 , n2625 );
buf ( n2627 , n2626 );
nand ( n2628 , n2622 , n2627 );
buf ( n2629 , n2628 );
buf ( n2630 , n2629 );
nand ( n2631 , n2615 , n2630 );
buf ( n2632 , n2631 );
buf ( n2633 , n2632 );
xor ( n2634 , n2607 , n2633 );
buf ( n2635 , n2634 );
buf ( n2636 , n2635 );
buf ( n2637 , n1684 );
not ( n2638 , n2637 );
buf ( n2639 , n1667 );
not ( n2640 , n2639 );
buf ( n2641 , n2640 );
buf ( n2642 , n2641 );
not ( n2643 , n2642 );
or ( n2644 , n2638 , n2643 );
buf ( n2645 , n1663 );
not ( n2646 , n2645 );
buf ( n2647 , n2646 );
buf ( n2648 , n2647 );
xor ( n2649 , n810 , n790 );
buf ( n2650 , n2649 );
nand ( n2651 , n2648 , n2650 );
buf ( n2652 , n2651 );
buf ( n2653 , n2652 );
nand ( n2654 , n2644 , n2653 );
buf ( n2655 , n2654 );
buf ( n2656 , n2655 );
buf ( n2657 , n1773 );
not ( n2658 , n2657 );
buf ( n2659 , n1780 );
not ( n2660 , n2659 );
or ( n2661 , n2658 , n2660 );
buf ( n2662 , n1771 );
buf ( n2663 , n1362 );
nand ( n2664 , n2662 , n2663 );
buf ( n2665 , n2664 );
buf ( n2666 , n2665 );
nand ( n2667 , n2661 , n2666 );
buf ( n2668 , n2667 );
buf ( n2669 , n2668 );
xor ( n2670 , n2656 , n2669 );
not ( n2671 , n1345 );
not ( n2672 , n2671 );
not ( n2673 , n2672 );
not ( n2674 , n1325 );
or ( n2675 , n2673 , n2674 );
buf ( n2676 , n2267 );
not ( n2677 , n2676 );
buf ( n2678 , n2677 );
buf ( n2679 , n2678 );
buf ( n2680 , n2679 );
buf ( n2681 , n2680 );
buf ( n2682 , n2418 );
not ( n2683 , n2682 );
buf ( n2684 , n2683 );
or ( n2685 , n2681 , n2684 );
nand ( n2686 , n2675 , n2685 );
buf ( n2687 , n2686 );
xor ( n2688 , n2670 , n2687 );
buf ( n2689 , n2688 );
buf ( n2690 , n2689 );
xor ( n2691 , n2636 , n2690 );
buf ( n2692 , n2454 );
not ( n2693 , n2692 );
buf ( n2694 , n1403 );
not ( n2695 , n2694 );
or ( n2696 , n2693 , n2695 );
buf ( n2697 , n2449 );
buf ( n2698 , n1389 );
nand ( n2699 , n2697 , n2698 );
buf ( n2700 , n2699 );
buf ( n2701 , n2700 );
nand ( n2702 , n2696 , n2701 );
buf ( n2703 , n2702 );
buf ( n2704 , n2703 );
buf ( n2705 , n2433 );
not ( n2706 , n2705 );
buf ( n2707 , n2235 );
buf ( n2708 , n2707 );
buf ( n2709 , n2708 );
buf ( n2710 , n2709 );
not ( n2711 , n2710 );
or ( n2712 , n2706 , n2711 );
buf ( n2713 , n1309 );
buf ( n2714 , n2713 );
buf ( n2715 , n1290 );
nand ( n2716 , n2714 , n2715 );
buf ( n2717 , n2716 );
buf ( n2718 , n2717 );
nand ( n2719 , n2712 , n2718 );
buf ( n2720 , n2719 );
buf ( n2721 , n2720 );
xor ( n2722 , n2704 , n2721 );
buf ( n2723 , n1761 );
not ( n2724 , n2723 );
buf ( n2725 , n1480 );
buf ( n2726 , n2725 );
not ( n2727 , n2726 );
or ( n2728 , n2724 , n2727 );
buf ( n2729 , n1496 );
buf ( n2730 , n1469 );
nand ( n2731 , n2729 , n2730 );
buf ( n2732 , n2731 );
buf ( n2733 , n2732 );
nand ( n2734 , n2728 , n2733 );
buf ( n2735 , n2734 );
buf ( n2736 , n2735 );
xor ( n2737 , n2722 , n2736 );
buf ( n2738 , n2737 );
buf ( n2739 , n2738 );
xor ( n2740 , n2691 , n2739 );
buf ( n2741 , n2740 );
xor ( n2742 , n2439 , n2422 );
xor ( n2743 , n2742 , n2460 );
buf ( n2744 , n2743 );
buf ( n2745 , n785 );
buf ( n2746 , n818 );
xor ( n2747 , n2745 , n2746 );
buf ( n2748 , n2747 );
buf ( n2749 , n2748 );
not ( n2750 , n2749 );
buf ( n2751 , n1486 );
not ( n2752 , n2751 );
or ( n2753 , n2750 , n2752 );
buf ( n2754 , n1496 );
buf ( n2755 , n1751 );
nand ( n2756 , n2754 , n2755 );
buf ( n2757 , n2756 );
buf ( n2758 , n2757 );
nand ( n2759 , n2753 , n2758 );
buf ( n2760 , n2759 );
buf ( n2761 , n2760 );
xor ( n2762 , n1892 , n1911 );
buf ( n2763 , n2762 );
xor ( n2764 , n2761 , n2763 );
buf ( n2765 , n1433 );
buf ( n2766 , n799 );
and ( n2767 , n2765 , n2766 );
buf ( n2768 , n2767 );
buf ( n2769 , n2768 );
buf ( n2770 , n776 );
buf ( n2771 , n828 );
xor ( n2772 , n2770 , n2771 );
buf ( n2773 , n2772 );
buf ( n2774 , n2773 );
not ( n2775 , n2774 );
buf ( n2776 , n1901 );
not ( n2777 , n2776 );
or ( n2778 , n2775 , n2777 );
buf ( n2779 , n1249 );
buf ( n2780 , n1897 );
nand ( n2781 , n2779 , n2780 );
buf ( n2782 , n2781 );
buf ( n2783 , n2782 );
nand ( n2784 , n2778 , n2783 );
buf ( n2785 , n2784 );
buf ( n2786 , n2785 );
xor ( n2787 , n2769 , n2786 );
buf ( n2788 , n1838 );
buf ( n2789 , n2788 );
buf ( n2790 , n2789 );
buf ( n2791 , n2790 );
not ( n2792 , n2791 );
buf ( n2793 , n2792 );
buf ( n2794 , n2793 );
buf ( n2795 , n780 );
buf ( n2796 , n824 );
xor ( n2797 , n2795 , n2796 );
buf ( n2798 , n2797 );
buf ( n2799 , n2798 );
not ( n2800 , n2799 );
buf ( n2801 , n2800 );
buf ( n2802 , n2801 );
or ( n2803 , n2794 , n2802 );
buf ( n2804 , n2489 );
buf ( n2805 , n1957 );
not ( n2806 , n2805 );
buf ( n2807 , n2806 );
buf ( n2808 , n2807 );
or ( n2809 , n2804 , n2808 );
nand ( n2810 , n2803 , n2809 );
buf ( n2811 , n2810 );
buf ( n2812 , n2811 );
and ( n2813 , n2787 , n2812 );
and ( n2814 , n2769 , n2786 );
or ( n2815 , n2813 , n2814 );
buf ( n2816 , n2815 );
buf ( n2817 , n2816 );
and ( n2818 , n2764 , n2817 );
and ( n2819 , n2761 , n2763 );
or ( n2820 , n2818 , n2819 );
buf ( n2821 , n2820 );
buf ( n2822 , n2821 );
xor ( n2823 , n2744 , n2822 );
buf ( n2824 , n790 );
buf ( n2825 , n814 );
xor ( n2826 , n2824 , n2825 );
buf ( n2827 , n2826 );
buf ( n2828 , n2827 );
not ( n2829 , n2828 );
buf ( n2830 , n1931 );
not ( n2831 , n2830 );
or ( n2832 , n2829 , n2831 );
buf ( n2833 , n1937 );
buf ( n2834 , n1923 );
nand ( n2835 , n2833 , n2834 );
buf ( n2836 , n2835 );
buf ( n2837 , n2836 );
nand ( n2838 , n2832 , n2837 );
buf ( n2839 , n2838 );
buf ( n2840 , n788 );
buf ( n2841 , n816 );
xor ( n2842 , n2840 , n2841 );
buf ( n2843 , n2842 );
buf ( n2844 , n2843 );
not ( n2845 , n2844 );
buf ( n2846 , n2523 );
not ( n2847 , n2846 );
or ( n2848 , n2845 , n2847 );
buf ( n2849 , n2532 );
buf ( n2850 , n1993 );
nand ( n2851 , n2849 , n2850 );
buf ( n2852 , n2851 );
buf ( n2853 , n2852 );
nand ( n2854 , n2848 , n2853 );
buf ( n2855 , n2854 );
xor ( n2856 , n2839 , n2855 );
buf ( n2857 , n782 );
buf ( n2858 , n822 );
xor ( n2859 , n2857 , n2858 );
buf ( n2860 , n2859 );
buf ( n2861 , n2860 );
not ( n2862 , n2861 );
buf ( n2863 , n2101 );
not ( n2864 , n2863 );
or ( n2865 , n2862 , n2864 );
buf ( n2866 , n2107 );
buf ( n2867 , n2082 );
nand ( n2868 , n2866 , n2867 );
buf ( n2869 , n2868 );
buf ( n2870 , n2869 );
nand ( n2871 , n2865 , n2870 );
buf ( n2872 , n2871 );
and ( n2873 , n2856 , n2872 );
and ( n2874 , n2839 , n2855 );
or ( n2875 , n2873 , n2874 );
not ( n2876 , n2875 );
not ( n2877 , n2207 );
buf ( n2878 , n774 );
buf ( n2879 , n830 );
xor ( n2880 , n2878 , n2879 );
buf ( n2881 , n2880 );
not ( n2882 , n2881 );
or ( n2883 , n2877 , n2882 );
buf ( n2884 , n2212 );
buf ( n2885 , n831 );
nand ( n2886 , n2884 , n2885 );
buf ( n2887 , n2886 );
nand ( n2888 , n2883 , n2887 );
buf ( n2889 , n2888 );
xor ( n2890 , n810 , n794 );
buf ( n2891 , n2890 );
not ( n2892 , n2891 );
not ( n2893 , n810 );
nand ( n2894 , n2893 , n811 );
nand ( n2895 , n1654 , n2894 );
and ( n2896 , n1663 , n2895 );
buf ( n2897 , n2896 );
not ( n2898 , n2897 );
or ( n2899 , n2892 , n2898 );
buf ( n2900 , n1679 );
buf ( n2901 , n2042 );
nand ( n2902 , n2900 , n2901 );
buf ( n2903 , n2902 );
buf ( n2904 , n2903 );
nand ( n2905 , n2899 , n2904 );
buf ( n2906 , n2905 );
buf ( n2907 , n2906 );
xor ( n2908 , n2889 , n2907 );
buf ( n2909 , n792 );
buf ( n2910 , n812 );
xor ( n2911 , n2909 , n2910 );
buf ( n2912 , n2911 );
buf ( n2913 , n2912 );
not ( n2914 , n2913 );
not ( n2915 , n2065 );
not ( n2916 , n2915 );
buf ( n2917 , n2916 );
not ( n2918 , n2917 );
or ( n2919 , n2914 , n2918 );
buf ( n2920 , n1693 );
buf ( n2921 , n2059 );
nand ( n2922 , n2920 , n2921 );
buf ( n2923 , n2922 );
buf ( n2924 , n2923 );
nand ( n2925 , n2919 , n2924 );
buf ( n2926 , n2925 );
buf ( n2927 , n2926 );
and ( n2928 , n2908 , n2927 );
and ( n2929 , n2889 , n2907 );
or ( n2930 , n2928 , n2929 );
buf ( n2931 , n2930 );
not ( n2932 , n2931 );
buf ( n2933 , n796 );
buf ( n2934 , n808 );
xor ( n2935 , n2933 , n2934 );
buf ( n2936 , n2935 );
buf ( n2937 , n2936 );
not ( n2938 , n2937 );
buf ( n2939 , n2235 );
not ( n2940 , n2939 );
or ( n2941 , n2938 , n2940 );
buf ( n2942 , n1309 );
buf ( n2943 , n2226 );
nand ( n2944 , n2942 , n2943 );
buf ( n2945 , n2944 );
buf ( n2946 , n2945 );
nand ( n2947 , n2941 , n2946 );
buf ( n2948 , n2947 );
buf ( n2949 , n2948 );
not ( n2950 , n2949 );
buf ( n2951 , n784 );
buf ( n2952 , n820 );
xor ( n2953 , n2951 , n2952 );
buf ( n2954 , n2953 );
buf ( n2955 , n2954 );
not ( n2956 , n2955 );
buf ( n2957 , n2410 );
not ( n2958 , n2957 );
or ( n2959 , n2956 , n2958 );
buf ( n2960 , n2257 );
buf ( n2961 , n1346 );
nand ( n2962 , n2960 , n2961 );
buf ( n2963 , n2962 );
buf ( n2964 , n2963 );
nand ( n2965 , n2959 , n2964 );
buf ( n2966 , n2965 );
buf ( n2967 , n2966 );
not ( n2968 , n2967 );
or ( n2969 , n2950 , n2968 );
buf ( n2970 , n2966 );
buf ( n2971 , n2948 );
or ( n2972 , n2970 , n2971 );
buf ( n2973 , n798 );
buf ( n2974 , n806 );
xor ( n2975 , n2973 , n2974 );
buf ( n2976 , n2975 );
buf ( n2977 , n2976 );
not ( n2978 , n2977 );
buf ( n2979 , n1403 );
not ( n2980 , n2979 );
or ( n2981 , n2978 , n2980 );
xor ( n2982 , n807 , n808 );
buf ( n2983 , n2982 );
buf ( n2984 , n2316 );
nand ( n2985 , n2983 , n2984 );
buf ( n2986 , n2985 );
buf ( n2987 , n2986 );
nand ( n2988 , n2981 , n2987 );
buf ( n2989 , n2988 );
buf ( n2990 , n2989 );
nand ( n2991 , n2972 , n2990 );
buf ( n2992 , n2991 );
buf ( n2993 , n2992 );
nand ( n2994 , n2969 , n2993 );
buf ( n2995 , n2994 );
not ( n2996 , n2995 );
nand ( n2997 , n2932 , n2996 );
not ( n2998 , n2997 );
or ( n2999 , n2876 , n2998 );
not ( n3000 , n2996 );
nand ( n3001 , n3000 , n2931 );
nand ( n3002 , n2999 , n3001 );
buf ( n3003 , n3002 );
and ( n3004 , n2823 , n3003 );
and ( n3005 , n2744 , n2822 );
or ( n3006 , n3004 , n3005 );
buf ( n3007 , n3006 );
xor ( n3008 , n2741 , n3007 );
xor ( n3009 , n2294 , n2380 );
xor ( n3010 , n3009 , n2403 );
buf ( n3011 , n3010 );
buf ( n3012 , n3011 );
and ( n3013 , n2027 , n1914 );
not ( n3014 , n2027 );
and ( n3015 , n1911 , n1892 );
and ( n3016 , n3014 , n3015 );
nor ( n3017 , n3013 , n3016 );
xor ( n3018 , n2129 , n3017 );
buf ( n3019 , n3018 );
not ( n3020 , n3019 );
buf ( n3021 , n3020 );
buf ( n3022 , n3021 );
or ( n3023 , n3012 , n3022 );
not ( n3024 , n2281 );
xor ( n3025 , n2220 , n3024 );
xnor ( n3026 , n3025 , n2250 );
buf ( n3027 , n3026 );
not ( n3028 , n3027 );
buf ( n3029 , n2353 );
not ( n3030 , n3029 );
buf ( n3031 , n2373 );
not ( n3032 , n3031 );
or ( n3033 , n3030 , n3032 );
buf ( n3034 , n2373 );
buf ( n3035 , n2353 );
or ( n3036 , n3034 , n3035 );
nand ( n3037 , n3033 , n3036 );
buf ( n3038 , n3037 );
buf ( n3039 , n3038 );
buf ( n3040 , n2348 );
and ( n3041 , n3039 , n3040 );
not ( n3042 , n3039 );
buf ( n3043 , n2310 );
and ( n3044 , n3042 , n3043 );
nor ( n3045 , n3041 , n3044 );
buf ( n3046 , n3045 );
buf ( n3047 , n3046 );
not ( n3048 , n3047 );
buf ( n3049 , n3048 );
buf ( n3050 , n3049 );
not ( n3051 , n3050 );
or ( n3052 , n3028 , n3051 );
not ( n3053 , n3046 );
not ( n3054 , n3026 );
not ( n3055 , n3054 );
or ( n3056 , n3053 , n3055 );
buf ( n3057 , n2021 );
buf ( n3058 , n1975 );
and ( n3059 , n3057 , n3058 );
not ( n3060 , n3057 );
buf ( n3061 , n1986 );
and ( n3062 , n3060 , n3061 );
nor ( n3063 , n3059 , n3062 );
buf ( n3064 , n3063 );
buf ( n3065 , n1951 );
buf ( n3066 , n3065 );
buf ( n3067 , n3066 );
not ( n3068 , n3067 );
and ( n3069 , n3064 , n3068 );
not ( n3070 , n3064 );
and ( n3071 , n3070 , n3067 );
nor ( n3072 , n3069 , n3071 );
not ( n3073 , n3072 );
nand ( n3074 , n3056 , n3073 );
buf ( n3075 , n3074 );
nand ( n3076 , n3052 , n3075 );
buf ( n3077 , n3076 );
buf ( n3078 , n3077 );
nand ( n3079 , n3023 , n3078 );
buf ( n3080 , n3079 );
buf ( n3081 , n3080 );
buf ( n3082 , n3021 );
buf ( n3083 , n3011 );
nand ( n3084 , n3082 , n3083 );
buf ( n3085 , n3084 );
buf ( n3086 , n3085 );
nand ( n3087 , n3081 , n3086 );
buf ( n3088 , n3087 );
xor ( n3089 , n3008 , n3088 );
buf ( n3090 , n3089 );
not ( n3091 , n3090 );
or ( n3092 , n2573 , n3091 );
not ( n3093 , n2568 );
nand ( n3094 , n3093 , n2564 );
buf ( n3095 , n3094 );
nand ( n3096 , n3092 , n3095 );
buf ( n3097 , n3096 );
buf ( n3098 , n3097 );
xor ( n3099 , n2561 , n3098 );
buf ( n3100 , n1594 );
buf ( n3101 , n1612 );
and ( n3102 , n3100 , n3101 );
buf ( n3103 , n3102 );
buf ( n3104 , n3103 );
buf ( n3105 , n1565 );
not ( n3106 , n3105 );
buf ( n3107 , n1551 );
buf ( n3108 , n3107 );
buf ( n3109 , n3108 );
buf ( n3110 , n3109 );
not ( n3111 , n3110 );
or ( n3112 , n3106 , n3111 );
buf ( n3113 , n1560 );
xor ( n3114 , n802 , n797 );
buf ( n3115 , n3114 );
nand ( n3116 , n3113 , n3115 );
buf ( n3117 , n3116 );
buf ( n3118 , n3117 );
nand ( n3119 , n3112 , n3118 );
buf ( n3120 , n3119 );
buf ( n3121 , n3120 );
xor ( n3122 , n3104 , n3121 );
xor ( n3123 , n2504 , n2517 );
and ( n3124 , n3123 , n2547 );
and ( n3125 , n2504 , n2517 );
or ( n3126 , n3124 , n3125 );
buf ( n3127 , n3126 );
buf ( n3128 , n3127 );
xor ( n3129 , n3122 , n3128 );
buf ( n3130 , n3129 );
buf ( n3131 , n3130 );
xor ( n3132 , n2153 , n2157 );
and ( n3133 , n3132 , n2203 );
and ( n3134 , n2153 , n2157 );
or ( n3135 , n3133 , n3134 );
buf ( n3136 , n3135 );
xor ( n3137 , n3131 , n3136 );
xor ( n3138 , n2636 , n2690 );
and ( n3139 , n3138 , n2739 );
and ( n3140 , n2636 , n2690 );
or ( n3141 , n3139 , n3140 );
buf ( n3142 , n3141 );
buf ( n3143 , n3142 );
xor ( n3144 , n3137 , n3143 );
buf ( n3145 , n3144 );
buf ( n3146 , n3145 );
xor ( n3147 , n2472 , n2477 );
and ( n3148 , n3147 , n2550 );
and ( n3149 , n2472 , n2477 );
or ( n3150 , n3148 , n3149 );
buf ( n3151 , n3150 );
buf ( n3152 , n3151 );
xor ( n3153 , n2592 , n2606 );
and ( n3154 , n3153 , n2633 );
and ( n3155 , n2592 , n2606 );
or ( n3156 , n3154 , n3155 );
buf ( n3157 , n3156 );
buf ( n3158 , n3157 );
xor ( n3159 , n2656 , n2669 );
and ( n3160 , n3159 , n2687 );
and ( n3161 , n2656 , n2669 );
or ( n3162 , n3160 , n3161 );
buf ( n3163 , n3162 );
buf ( n3164 , n3163 );
xor ( n3165 , n3158 , n3164 );
xor ( n3166 , n2704 , n2721 );
and ( n3167 , n3166 , n2736 );
and ( n3168 , n2704 , n2721 );
or ( n3169 , n3167 , n3168 );
buf ( n3170 , n3169 );
buf ( n3171 , n3170 );
xor ( n3172 , n3165 , n3171 );
buf ( n3173 , n3172 );
buf ( n3174 , n3173 );
xor ( n3175 , n3152 , n3174 );
not ( n3176 , n1616 );
not ( n3177 , n1535 );
or ( n3178 , n3176 , n3177 );
buf ( n3179 , n1616 );
buf ( n3180 , n1535 );
nor ( n3181 , n3179 , n3180 );
buf ( n3182 , n3181 );
or ( n3183 , n3182 , n1577 );
nand ( n3184 , n3178 , n3183 );
buf ( n3185 , n3184 );
buf ( n3186 , n2585 );
not ( n3187 , n3186 );
buf ( n3188 , n2098 );
not ( n3189 , n3188 );
or ( n3190 , n3187 , n3189 );
buf ( n3191 , n2107 );
xor ( n3192 , n822 , n777 );
buf ( n3193 , n3192 );
nand ( n3194 , n3191 , n3193 );
buf ( n3195 , n3194 );
buf ( n3196 , n3195 );
nand ( n3197 , n3190 , n3196 );
buf ( n3198 , n3197 );
buf ( n3199 , n3198 );
not ( n3200 , n3199 );
buf ( n3201 , n2599 );
not ( n3202 , n3201 );
buf ( n3203 , n2066 );
not ( n3204 , n3203 );
or ( n3205 , n3202 , n3204 );
buf ( n3206 , n1693 );
xor ( n3207 , n812 , n787 );
buf ( n3208 , n3207 );
nand ( n3209 , n3206 , n3208 );
buf ( n3210 , n3209 );
buf ( n3211 , n3210 );
nand ( n3212 , n3205 , n3211 );
buf ( n3213 , n3212 );
buf ( n3214 , n3213 );
not ( n3215 , n3214 );
buf ( n3216 , n3215 );
buf ( n3217 , n3216 );
not ( n3218 , n3217 );
or ( n3219 , n3200 , n3218 );
buf ( n3220 , n3216 );
buf ( n3221 , n3198 );
or ( n3222 , n3220 , n3221 );
nand ( n3223 , n3219 , n3222 );
buf ( n3224 , n3223 );
buf ( n3225 , n3224 );
buf ( n3226 , n2649 );
not ( n3227 , n3226 );
buf ( n3228 , n1670 );
not ( n3229 , n3228 );
or ( n3230 , n3227 , n3229 );
buf ( n3231 , n2647 );
xor ( n3232 , n810 , n789 );
buf ( n3233 , n3232 );
nand ( n3234 , n3231 , n3233 );
buf ( n3235 , n3234 );
buf ( n3236 , n3235 );
nand ( n3237 , n3230 , n3236 );
buf ( n3238 , n3237 );
buf ( n3239 , n3238 );
xor ( n3240 , n3225 , n3239 );
buf ( n3241 , n3240 );
buf ( n3242 , n3241 );
xor ( n3243 , n3185 , n3242 );
buf ( n3244 , n2497 );
not ( n3245 , n3244 );
buf ( n3246 , n1965 );
not ( n3247 , n3246 );
or ( n3248 , n3245 , n3247 );
buf ( n3249 , n825 );
buf ( n3250 , n826 );
xnor ( n3251 , n3249 , n3250 );
buf ( n3252 , n3251 );
buf ( n3253 , n3252 );
not ( n3254 , n3253 );
buf ( n3255 , n3254 );
buf ( n3256 , n3255 );
buf ( n3257 , n775 );
buf ( n3258 , n824 );
xor ( n3259 , n3257 , n3258 );
buf ( n3260 , n3259 );
buf ( n3261 , n3260 );
nand ( n3262 , n3256 , n3261 );
buf ( n3263 , n3262 );
buf ( n3264 , n3263 );
nand ( n3265 , n3248 , n3264 );
buf ( n3266 , n3265 );
buf ( n3267 , n2540 );
not ( n3268 , n3267 );
buf ( n3269 , n2526 );
not ( n3270 , n3269 );
or ( n3271 , n3268 , n3270 );
buf ( n3272 , n2010 );
buf ( n3273 , n783 );
buf ( n3274 , n816 );
xor ( n3275 , n3273 , n3274 );
buf ( n3276 , n3275 );
buf ( n3277 , n3276 );
nand ( n3278 , n3272 , n3277 );
buf ( n3279 , n3278 );
buf ( n3280 , n3279 );
nand ( n3281 , n3271 , n3280 );
buf ( n3282 , n3281 );
xor ( n3283 , n3266 , n3282 );
buf ( n3284 , n2626 );
not ( n3285 , n3284 );
buf ( n3286 , n2612 );
not ( n3287 , n3286 );
or ( n3288 , n3285 , n3287 );
buf ( n3289 , n2621 );
buf ( n3290 , n785 );
buf ( n3291 , n814 );
xor ( n3292 , n3290 , n3291 );
buf ( n3293 , n3292 );
buf ( n3294 , n3293 );
nand ( n3295 , n3289 , n3294 );
buf ( n3296 , n3295 );
buf ( n3297 , n3296 );
nand ( n3298 , n3288 , n3297 );
buf ( n3299 , n3298 );
xor ( n3300 , n3283 , n3299 );
buf ( n3301 , n3300 );
xor ( n3302 , n3243 , n3301 );
buf ( n3303 , n3302 );
buf ( n3304 , n3303 );
xor ( n3305 , n3175 , n3304 );
buf ( n3306 , n3305 );
buf ( n3307 , n3306 );
xor ( n3308 , n3146 , n3307 );
xor ( n3309 , n2741 , n3007 );
and ( n3310 , n3309 , n3088 );
and ( n3311 , n2741 , n3007 );
or ( n3312 , n3310 , n3311 );
buf ( n3313 , n3312 );
xor ( n3314 , n3308 , n3313 );
buf ( n3315 , n3314 );
buf ( n3316 , n3315 );
and ( n3317 , n3099 , n3316 );
and ( n3318 , n2561 , n3098 );
or ( n3319 , n3317 , n3318 );
buf ( n3320 , n3319 );
buf ( n3321 , n3320 );
xor ( n3322 , n1214 , n3321 );
buf ( n3323 , n1314 );
not ( n3324 , n3323 );
buf ( n3325 , n2235 );
not ( n3326 , n3325 );
or ( n3327 , n3324 , n3326 );
buf ( n3328 , n790 );
buf ( n3329 , n808 );
xor ( n3330 , n3328 , n3329 );
buf ( n3331 , n3330 );
buf ( n3332 , n3331 );
buf ( n3333 , n1309 );
nand ( n3334 , n3332 , n3333 );
buf ( n3335 , n3334 );
buf ( n3336 , n3335 );
nand ( n3337 , n3327 , n3336 );
buf ( n3338 , n3337 );
buf ( n3339 , n3338 );
buf ( n3340 , n1414 );
not ( n3341 , n3340 );
buf ( n3342 , n1403 );
not ( n3343 , n3342 );
or ( n3344 , n3341 , n3343 );
buf ( n3345 , n2449 );
buf ( n3346 , n792 );
buf ( n3347 , n806 );
xor ( n3348 , n3346 , n3347 );
buf ( n3349 , n3348 );
buf ( n3350 , n3349 );
nand ( n3351 , n3345 , n3350 );
buf ( n3352 , n3351 );
buf ( n3353 , n3352 );
nand ( n3354 , n3344 , n3353 );
buf ( n3355 , n3354 );
buf ( n3356 , n3355 );
xor ( n3357 , n3339 , n3356 );
not ( n3358 , n2672 );
buf ( n3359 , n778 );
buf ( n3360 , n820 );
xor ( n3361 , n3359 , n3360 );
buf ( n3362 , n3361 );
not ( n3363 , n3362 );
or ( n3364 , n3358 , n3363 );
buf ( n3365 , n1344 );
not ( n3366 , n3365 );
buf ( n3367 , n3366 );
or ( n3368 , n2678 , n3367 );
nand ( n3369 , n3364 , n3368 );
buf ( n3370 , n3369 );
xor ( n3371 , n3357 , n3370 );
buf ( n3372 , n3371 );
buf ( n3373 , n3372 );
buf ( n3374 , n3207 );
not ( n3375 , n3374 );
buf ( n3376 , n2916 );
not ( n3377 , n3376 );
or ( n3378 , n3375 , n3377 );
buf ( n3379 , n1693 );
buf ( n3380 , n3379 );
buf ( n3381 , n786 );
buf ( n3382 , n812 );
xor ( n3383 , n3381 , n3382 );
buf ( n3384 , n3383 );
buf ( n3385 , n3384 );
nand ( n3386 , n3380 , n3385 );
buf ( n3387 , n3386 );
buf ( n3388 , n3387 );
nand ( n3389 , n3378 , n3388 );
buf ( n3390 , n3389 );
buf ( n3391 , n3232 );
not ( n3392 , n3391 );
buf ( n3393 , n2641 );
not ( n3394 , n3393 );
or ( n3395 , n3392 , n3394 );
buf ( n3396 , n1676 );
not ( n3397 , n3396 );
buf ( n3398 , n3397 );
buf ( n3399 , n3398 );
buf ( n3400 , n788 );
buf ( n3401 , n810 );
xor ( n3402 , n3400 , n3401 );
buf ( n3403 , n3402 );
buf ( n3404 , n3403 );
nand ( n3405 , n3399 , n3404 );
buf ( n3406 , n3405 );
buf ( n3407 , n3406 );
nand ( n3408 , n3395 , n3407 );
buf ( n3409 , n3408 );
xor ( n3410 , n3390 , n3409 );
buf ( n3411 , n1376 );
not ( n3412 , n3411 );
buf ( n3413 , n1780 );
not ( n3414 , n3413 );
or ( n3415 , n3412 , n3414 );
buf ( n3416 , n1771 );
buf ( n3417 , n772 );
buf ( n3418 , n826 );
xor ( n3419 , n3417 , n3418 );
buf ( n3420 , n3419 );
buf ( n3421 , n3420 );
nand ( n3422 , n3416 , n3421 );
buf ( n3423 , n3422 );
buf ( n3424 , n3423 );
nand ( n3425 , n3415 , n3424 );
buf ( n3426 , n3425 );
xor ( n3427 , n3410 , n3426 );
buf ( n3428 , n3427 );
xor ( n3429 , n3373 , n3428 );
xor ( n3430 , n3158 , n3164 );
and ( n3431 , n3430 , n3171 );
and ( n3432 , n3158 , n3164 );
or ( n3433 , n3431 , n3432 );
buf ( n3434 , n3433 );
buf ( n3435 , n3434 );
xor ( n3436 , n3429 , n3435 );
buf ( n3437 , n3436 );
buf ( n3438 , n3437 );
xor ( n3439 , n3131 , n3136 );
and ( n3440 , n3439 , n3143 );
and ( n3441 , n3131 , n3136 );
or ( n3442 , n3440 , n3441 );
buf ( n3443 , n3442 );
buf ( n3444 , n3443 );
xor ( n3445 , n3438 , n3444 );
xor ( n3446 , n3152 , n3174 );
and ( n3447 , n3446 , n3304 );
and ( n3448 , n3152 , n3174 );
or ( n3449 , n3447 , n3448 );
buf ( n3450 , n3449 );
buf ( n3451 , n3450 );
xor ( n3452 , n3445 , n3451 );
buf ( n3453 , n3452 );
buf ( n3454 , n3453 );
buf ( n3455 , n799 );
buf ( n3456 , n801 );
nand ( n3457 , n3455 , n3456 );
buf ( n3458 , n3457 );
buf ( n3459 , n799 );
buf ( n3460 , n801 );
or ( n3461 , n3459 , n3460 );
buf ( n3462 , n802 );
nand ( n3463 , n3461 , n3462 );
buf ( n3464 , n3463 );
nand ( n3465 , n3458 , n800 , n3464 );
buf ( n3466 , n3465 );
not ( n3467 , n3466 );
buf ( n3468 , n1275 );
not ( n3469 , n3468 );
buf ( n3470 , n1630 );
not ( n3471 , n3470 );
or ( n3472 , n3469 , n3471 );
buf ( n3473 , n768 );
buf ( n3474 , n830 );
xor ( n3475 , n3473 , n3474 );
buf ( n3476 , n3475 );
buf ( n3477 , n3476 );
buf ( n3478 , n831 );
nand ( n3479 , n3477 , n3478 );
buf ( n3480 , n3479 );
buf ( n3481 , n3480 );
nand ( n3482 , n3472 , n3481 );
buf ( n3483 , n3482 );
buf ( n3484 , n3483 );
not ( n3485 , n3484 );
or ( n3486 , n3467 , n3485 );
buf ( n3487 , n3483 );
buf ( n3488 , n3465 );
or ( n3489 , n3487 , n3488 );
nand ( n3490 , n3486 , n3489 );
buf ( n3491 , n3490 );
buf ( n3492 , n3491 );
xor ( n3493 , n1223 , n1261 );
and ( n3494 , n3493 , n1283 );
and ( n3495 , n1223 , n1261 );
or ( n3496 , n3494 , n3495 );
buf ( n3497 , n3496 );
buf ( n3498 , n3497 );
xor ( n3499 , n3492 , n3498 );
not ( n3500 , n3299 );
not ( n3501 , n3266 );
or ( n3502 , n3500 , n3501 );
buf ( n3503 , n3299 );
buf ( n3504 , n3266 );
nor ( n3505 , n3503 , n3504 );
buf ( n3506 , n3505 );
buf ( n3507 , n3282 );
not ( n3508 , n3507 );
buf ( n3509 , n3508 );
or ( n3510 , n3506 , n3509 );
nand ( n3511 , n3502 , n3510 );
buf ( n3512 , n3511 );
xor ( n3513 , n3499 , n3512 );
buf ( n3514 , n3513 );
not ( n3515 , n3198 );
not ( n3516 , n3238 );
or ( n3517 , n3515 , n3516 );
buf ( n3518 , n3198 );
buf ( n3519 , n3238 );
or ( n3520 , n3518 , n3519 );
buf ( n3521 , n3213 );
nand ( n3522 , n3520 , n3521 );
buf ( n3523 , n3522 );
nand ( n3524 , n3517 , n3523 );
not ( n3525 , n3524 );
not ( n3526 , n3525 );
not ( n3527 , n1348 );
not ( n3528 , n1320 );
not ( n3529 , n3528 );
not ( n3530 , n3529 );
or ( n3531 , n3527 , n3530 );
not ( n3532 , n3528 );
not ( n3533 , n1348 );
not ( n3534 , n3533 );
or ( n3535 , n3532 , n3534 );
nand ( n3536 , n3535 , n1382 );
nand ( n3537 , n3531 , n3536 );
not ( n3538 , n3537 );
not ( n3539 , n3538 );
or ( n3540 , n3526 , n3539 );
nand ( n3541 , n3524 , n3537 );
nand ( n3542 , n3540 , n3541 );
not ( n3543 , n1504 );
nand ( n3544 , n1463 , n1421 );
not ( n3545 , n3544 );
or ( n3546 , n3543 , n3545 );
nand ( n3547 , n1460 , n1420 );
nand ( n3548 , n3546 , n3547 );
not ( n3549 , n3548 );
and ( n3550 , n3542 , n3549 );
not ( n3551 , n3542 );
and ( n3552 , n3551 , n3548 );
nor ( n3553 , n3550 , n3552 );
not ( n3554 , n3553 );
xor ( n3555 , n3104 , n3121 );
and ( n3556 , n3555 , n3128 );
and ( n3557 , n3104 , n3121 );
or ( n3558 , n3556 , n3557 );
buf ( n3559 , n3558 );
and ( n3560 , n3554 , n3559 );
not ( n3561 , n3554 );
not ( n3562 , n3559 );
and ( n3563 , n3561 , n3562 );
nor ( n3564 , n3560 , n3563 );
xnor ( n3565 , n3514 , n3564 );
buf ( n3566 , n3565 );
xor ( n3567 , n1286 , n1384 );
and ( n3568 , n3567 , n1510 );
and ( n3569 , n1286 , n1384 );
or ( n3570 , n3568 , n3569 );
buf ( n3571 , n3570 );
buf ( n3572 , n3571 );
xor ( n3573 , n3185 , n3242 );
and ( n3574 , n3573 , n3301 );
and ( n3575 , n3185 , n3242 );
or ( n3576 , n3574 , n3575 );
buf ( n3577 , n3576 );
buf ( n3578 , n3577 );
xor ( n3579 , n3572 , n3578 );
buf ( n3580 , n3114 );
not ( n3581 , n3580 );
buf ( n3582 , n1548 );
not ( n3583 , n3582 );
or ( n3584 , n3581 , n3583 );
buf ( n3585 , n1557 );
buf ( n3586 , n796 );
buf ( n3587 , n802 );
xor ( n3588 , n3586 , n3587 );
buf ( n3589 , n3588 );
buf ( n3590 , n3589 );
nand ( n3591 , n3585 , n3590 );
buf ( n3592 , n3591 );
buf ( n3593 , n3592 );
nand ( n3594 , n3584 , n3593 );
buf ( n3595 , n3594 );
buf ( n3596 , n1454 );
not ( n3597 , n3596 );
buf ( n3598 , n1737 );
not ( n3599 , n3598 );
or ( n3600 , n3597 , n3599 );
buf ( n3601 , n1449 );
buf ( n3602 , n794 );
buf ( n3603 , n804 );
xor ( n3604 , n3602 , n3603 );
buf ( n3605 , n3604 );
buf ( n3606 , n3605 );
nand ( n3607 , n3601 , n3606 );
buf ( n3608 , n3607 );
buf ( n3609 , n3608 );
nand ( n3610 , n3600 , n3609 );
buf ( n3611 , n3610 );
xor ( n3612 , n3595 , n3611 );
buf ( n3613 , n1498 );
not ( n3614 , n3613 );
buf ( n3615 , n1480 );
not ( n3616 , n3615 );
or ( n3617 , n3614 , n3616 );
buf ( n3618 , n1496 );
xor ( n3619 , n818 , n780 );
buf ( n3620 , n3619 );
nand ( n3621 , n3618 , n3620 );
buf ( n3622 , n3621 );
buf ( n3623 , n3622 );
nand ( n3624 , n3617 , n3623 );
buf ( n3625 , n3624 );
xor ( n3626 , n3612 , n3625 );
buf ( n3627 , n3626 );
buf ( n3628 , n3260 );
not ( n3629 , n3628 );
buf ( n3630 , n1965 );
not ( n3631 , n3630 );
or ( n3632 , n3629 , n3631 );
buf ( n3633 , n3255 );
buf ( n3634 , n774 );
buf ( n3635 , n824 );
xor ( n3636 , n3634 , n3635 );
buf ( n3637 , n3636 );
buf ( n3638 , n3637 );
nand ( n3639 , n3633 , n3638 );
buf ( n3640 , n3639 );
buf ( n3641 , n3640 );
nand ( n3642 , n3632 , n3641 );
buf ( n3643 , n3642 );
buf ( n3644 , n3643 );
buf ( n3645 , n799 );
buf ( n3646 , n800 );
xor ( n3647 , n3645 , n3646 );
buf ( n3648 , n3647 );
buf ( n3649 , n3648 );
not ( n3650 , n3649 );
buf ( n3651 , n801 );
buf ( n3652 , n800 );
xnor ( n3653 , n3651 , n3652 );
buf ( n3654 , n3653 );
nor ( n3655 , n3654 , n1218 );
buf ( n3656 , n3655 );
buf ( n3657 , n3656 );
not ( n3658 , n3657 );
or ( n3659 , n3650 , n3658 );
buf ( n3660 , n1218 );
buf ( n3661 , n3660 );
buf ( n3662 , n3661 );
buf ( n3663 , n3662 );
buf ( n3664 , n798 );
buf ( n3665 , n800 );
xor ( n3666 , n3664 , n3665 );
buf ( n3667 , n3666 );
buf ( n3668 , n3667 );
nand ( n3669 , n3663 , n3668 );
buf ( n3670 , n3669 );
buf ( n3671 , n3670 );
nand ( n3672 , n3659 , n3671 );
buf ( n3673 , n3672 );
buf ( n3674 , n3673 );
xor ( n3675 , n3644 , n3674 );
buf ( n3676 , n1254 );
not ( n3677 , n3676 );
buf ( n3678 , n1901 );
buf ( n3679 , n3678 );
buf ( n3680 , n3679 );
buf ( n3681 , n3680 );
not ( n3682 , n3681 );
or ( n3683 , n3677 , n3682 );
buf ( n3684 , n1249 );
buf ( n3685 , n770 );
buf ( n3686 , n828 );
xor ( n3687 , n3685 , n3686 );
buf ( n3688 , n3687 );
buf ( n3689 , n3688 );
nand ( n3690 , n3684 , n3689 );
buf ( n3691 , n3690 );
buf ( n3692 , n3691 );
nand ( n3693 , n3683 , n3692 );
buf ( n3694 , n3693 );
buf ( n3695 , n3694 );
xor ( n3696 , n3675 , n3695 );
buf ( n3697 , n3696 );
buf ( n3698 , n3697 );
xor ( n3699 , n3627 , n3698 );
not ( n3700 , n3293 );
buf ( n3701 , n1931 );
buf ( n3702 , n3701 );
buf ( n3703 , n3702 );
not ( n3704 , n3703 );
or ( n3705 , n3700 , n3704 );
buf ( n3706 , n2621 );
buf ( n3707 , n784 );
buf ( n3708 , n814 );
xor ( n3709 , n3707 , n3708 );
buf ( n3710 , n3709 );
buf ( n3711 , n3710 );
nand ( n3712 , n3706 , n3711 );
buf ( n3713 , n3712 );
nand ( n3714 , n3705 , n3713 );
buf ( n3715 , n3276 );
not ( n3716 , n3715 );
buf ( n3717 , n2004 );
buf ( n3718 , n3717 );
buf ( n3719 , n3718 );
buf ( n3720 , n3719 );
not ( n3721 , n3720 );
or ( n3722 , n3716 , n3721 );
buf ( n3723 , n2535 );
buf ( n3724 , n782 );
buf ( n3725 , n816 );
xor ( n3726 , n3724 , n3725 );
buf ( n3727 , n3726 );
buf ( n3728 , n3727 );
nand ( n3729 , n3723 , n3728 );
buf ( n3730 , n3729 );
buf ( n3731 , n3730 );
nand ( n3732 , n3722 , n3731 );
buf ( n3733 , n3732 );
xor ( n3734 , n3714 , n3733 );
buf ( n3735 , n3192 );
not ( n3736 , n3735 );
buf ( n3737 , n2098 );
buf ( n3738 , n3737 );
buf ( n3739 , n3738 );
buf ( n3740 , n3739 );
not ( n3741 , n3740 );
or ( n3742 , n3736 , n3741 );
buf ( n3743 , n2107 );
buf ( n3744 , n3743 );
buf ( n3745 , n3744 );
buf ( n3746 , n3745 );
buf ( n3747 , n776 );
buf ( n3748 , n822 );
xor ( n3749 , n3747 , n3748 );
buf ( n3750 , n3749 );
buf ( n3751 , n3750 );
nand ( n3752 , n3746 , n3751 );
buf ( n3753 , n3752 );
buf ( n3754 , n3753 );
nand ( n3755 , n3742 , n3754 );
buf ( n3756 , n3755 );
xor ( n3757 , n3734 , n3756 );
buf ( n3758 , n3757 );
xor ( n3759 , n3699 , n3758 );
buf ( n3760 , n3759 );
buf ( n3761 , n3760 );
xor ( n3762 , n3579 , n3761 );
buf ( n3763 , n3762 );
buf ( n3764 , n3763 );
xor ( n3765 , n3566 , n3764 );
xor ( n3766 , n1513 , n2142 );
and ( n3767 , n3766 , n2558 );
and ( n3768 , n1513 , n2142 );
or ( n3769 , n3767 , n3768 );
buf ( n3770 , n3769 );
buf ( n3771 , n3770 );
xor ( n3772 , n3765 , n3771 );
buf ( n3773 , n3772 );
buf ( n3774 , n3773 );
xor ( n3775 , n3454 , n3774 );
xor ( n3776 , n3146 , n3307 );
and ( n3777 , n3776 , n3313 );
and ( n3778 , n3146 , n3307 );
or ( n3779 , n3777 , n3778 );
buf ( n3780 , n3779 );
buf ( n3781 , n3780 );
xor ( n3782 , n3775 , n3781 );
buf ( n3783 , n3782 );
buf ( n3784 , n3783 );
and ( n3785 , n3322 , n3784 );
and ( n3786 , n1214 , n3321 );
or ( n3787 , n3785 , n3786 );
buf ( n3788 , n3787 );
buf ( n3789 , n3788 );
xor ( n3790 , n3454 , n3774 );
and ( n3791 , n3790 , n3781 );
and ( n3792 , n3454 , n3774 );
or ( n3793 , n3791 , n3792 );
buf ( n3794 , n3793 );
buf ( n3795 , n3794 );
not ( n3796 , n3795 );
xor ( n3797 , n3438 , n3444 );
and ( n3798 , n3797 , n3451 );
and ( n3799 , n3438 , n3444 );
or ( n3800 , n3798 , n3799 );
buf ( n3801 , n3800 );
buf ( n3802 , n3801 );
xor ( n3803 , n3566 , n3764 );
and ( n3804 , n3803 , n3771 );
and ( n3805 , n3566 , n3764 );
or ( n3806 , n3804 , n3805 );
buf ( n3807 , n3806 );
buf ( n3808 , n3807 );
xor ( n3809 , n3802 , n3808 );
xor ( n3810 , n3492 , n3498 );
and ( n3811 , n3810 , n3512 );
and ( n3812 , n3492 , n3498 );
or ( n3813 , n3811 , n3812 );
buf ( n3814 , n3813 );
buf ( n3815 , n3814 );
not ( n3816 , n3815 );
buf ( n3817 , n3816 );
buf ( n3818 , n3817 );
buf ( n3819 , n799 );
buf ( n3820 , n800 );
and ( n3821 , n3819 , n3820 );
buf ( n3822 , n3821 );
buf ( n3823 , n3822 );
buf ( n3824 , n3476 );
not ( n3825 , n3824 );
buf ( n3826 , n1161 );
not ( n3827 , n3826 );
or ( n3828 , n3825 , n3827 );
buf ( n3829 , n830 );
buf ( n3830 , n831 );
nand ( n3831 , n3829 , n3830 );
buf ( n3832 , n3831 );
buf ( n3833 , n3832 );
nand ( n3834 , n3828 , n3833 );
buf ( n3835 , n3834 );
buf ( n3836 , n3835 );
xor ( n3837 , n3823 , n3836 );
buf ( n3838 , n3688 );
not ( n3839 , n3838 );
not ( n3840 , n1237 );
xor ( n3841 , n829 , n830 );
nor ( n3842 , n3840 , n3841 );
buf ( n3843 , n3842 );
not ( n3844 , n3843 );
or ( n3845 , n3839 , n3844 );
buf ( n3846 , n1249 );
buf ( n3847 , n769 );
buf ( n3848 , n828 );
xor ( n3849 , n3847 , n3848 );
buf ( n3850 , n3849 );
buf ( n3851 , n3850 );
nand ( n3852 , n3846 , n3851 );
buf ( n3853 , n3852 );
buf ( n3854 , n3853 );
nand ( n3855 , n3845 , n3854 );
buf ( n3856 , n3855 );
buf ( n3857 , n3856 );
xor ( n3858 , n3837 , n3857 );
buf ( n3859 , n3858 );
buf ( n3860 , n3859 );
buf ( n3861 , n3595 );
not ( n3862 , n3861 );
buf ( n3863 , n3611 );
not ( n3864 , n3863 );
or ( n3865 , n3862 , n3864 );
buf ( n3866 , n3611 );
buf ( n3867 , n3595 );
or ( n3868 , n3866 , n3867 );
buf ( n3869 , n3625 );
nand ( n3870 , n3868 , n3869 );
buf ( n3871 , n3870 );
buf ( n3872 , n3871 );
nand ( n3873 , n3865 , n3872 );
buf ( n3874 , n3873 );
buf ( n3875 , n3874 );
xor ( n3876 , n3860 , n3875 );
xor ( n3877 , n3339 , n3356 );
and ( n3878 , n3877 , n3370 );
and ( n3879 , n3339 , n3356 );
or ( n3880 , n3878 , n3879 );
buf ( n3881 , n3880 );
buf ( n3882 , n3881 );
xnor ( n3883 , n3876 , n3882 );
buf ( n3884 , n3883 );
buf ( n3885 , n3884 );
not ( n3886 , n3885 );
buf ( n3887 , n3886 );
buf ( n3888 , n3887 );
xor ( n3889 , n3818 , n3888 );
xor ( n3890 , n3627 , n3698 );
and ( n3891 , n3890 , n3758 );
and ( n3892 , n3627 , n3698 );
or ( n3893 , n3891 , n3892 );
buf ( n3894 , n3893 );
buf ( n3895 , n3894 );
xnor ( n3896 , n3889 , n3895 );
buf ( n3897 , n3896 );
buf ( n3898 , n3897 );
buf ( n3899 , n3750 );
not ( n3900 , n3899 );
buf ( n3901 , n2577 );
not ( n3902 , n3901 );
or ( n3903 , n3900 , n3902 );
buf ( n3904 , n2107 );
buf ( n3905 , n775 );
buf ( n3906 , n822 );
xor ( n3907 , n3905 , n3906 );
buf ( n3908 , n3907 );
buf ( n3909 , n3908 );
nand ( n3910 , n3904 , n3909 );
buf ( n3911 , n3910 );
buf ( n3912 , n3911 );
nand ( n3913 , n3903 , n3912 );
buf ( n3914 , n3913 );
buf ( n3915 , n3914 );
buf ( n3916 , n3710 );
not ( n3917 , n3916 );
not ( n3918 , n814 );
and ( n3919 , n815 , n3918 );
not ( n3920 , n815 );
and ( n3921 , n3920 , n814 );
nor ( n3922 , n3919 , n3921 );
nor ( n3923 , n3922 , n1927 );
buf ( n3924 , n3923 );
not ( n3925 , n3924 );
or ( n3926 , n3917 , n3925 );
buf ( n3927 , n1937 );
buf ( n3928 , n783 );
buf ( n3929 , n814 );
xor ( n3930 , n3928 , n3929 );
buf ( n3931 , n3930 );
buf ( n3932 , n3931 );
nand ( n3933 , n3927 , n3932 );
buf ( n3934 , n3933 );
buf ( n3935 , n3934 );
nand ( n3936 , n3926 , n3935 );
buf ( n3937 , n3936 );
buf ( n3938 , n3937 );
not ( n3939 , n3938 );
buf ( n3940 , n3939 );
buf ( n3941 , n3940 );
and ( n3942 , n3915 , n3941 );
not ( n3943 , n3915 );
buf ( n3944 , n3937 );
and ( n3945 , n3943 , n3944 );
nor ( n3946 , n3942 , n3945 );
buf ( n3947 , n3946 );
buf ( n3948 , n3947 );
buf ( n3949 , n3384 );
not ( n3950 , n3949 );
buf ( n3951 , n2916 );
not ( n3952 , n3951 );
or ( n3953 , n3950 , n3952 );
buf ( n3954 , n1693 );
buf ( n3955 , n785 );
buf ( n3956 , n812 );
xor ( n3957 , n3955 , n3956 );
buf ( n3958 , n3957 );
buf ( n3959 , n3958 );
nand ( n3960 , n3954 , n3959 );
buf ( n3961 , n3960 );
buf ( n3962 , n3961 );
nand ( n3963 , n3953 , n3962 );
buf ( n3964 , n3963 );
buf ( n3965 , n3964 );
and ( n3966 , n3948 , n3965 );
not ( n3967 , n3948 );
buf ( n3968 , n3964 );
not ( n3969 , n3968 );
buf ( n3970 , n3969 );
buf ( n3971 , n3970 );
and ( n3972 , n3967 , n3971 );
nor ( n3973 , n3966 , n3972 );
buf ( n3974 , n3973 );
not ( n3975 , n3362 );
not ( n3976 , n1338 );
or ( n3977 , n3975 , n3976 );
buf ( n3978 , n777 );
buf ( n3979 , n820 );
xor ( n3980 , n3978 , n3979 );
buf ( n3981 , n3980 );
buf ( n3982 , n3981 );
buf ( n3983 , n821 );
buf ( n3984 , n822 );
xor ( n3985 , n3983 , n3984 );
buf ( n3986 , n3985 );
buf ( n3987 , n3986 );
nand ( n3988 , n3982 , n3987 );
buf ( n3989 , n3988 );
nand ( n3990 , n3977 , n3989 );
not ( n3991 , n3990 );
not ( n3992 , n3403 );
not ( n3993 , n2896 );
or ( n3994 , n3992 , n3993 );
buf ( n3995 , n2647 );
buf ( n3996 , n787 );
buf ( n3997 , n810 );
xor ( n3998 , n3996 , n3997 );
buf ( n3999 , n3998 );
buf ( n4000 , n3999 );
nand ( n4001 , n3995 , n4000 );
buf ( n4002 , n4001 );
nand ( n4003 , n3994 , n4002 );
not ( n4004 , n4003 );
or ( n4005 , n3991 , n4004 );
not ( n4006 , n3403 );
not ( n4007 , n2896 );
or ( n4008 , n4006 , n4007 );
nand ( n4009 , n4008 , n4002 );
or ( n4010 , n4009 , n3990 );
nand ( n4011 , n4005 , n4010 );
buf ( n4012 , n1783 );
buf ( n4013 , n3420 );
not ( n4014 , n4013 );
buf ( n4015 , n4014 );
buf ( n4016 , n4015 );
or ( n4017 , n4012 , n4016 );
buf ( n4018 , n1771 );
not ( n4019 , n4018 );
buf ( n4020 , n4019 );
buf ( n4021 , n4020 );
buf ( n4022 , n771 );
buf ( n4023 , n826 );
xor ( n4024 , n4022 , n4023 );
buf ( n4025 , n4024 );
buf ( n4026 , n4025 );
not ( n4027 , n4026 );
buf ( n4028 , n4027 );
buf ( n4029 , n4028 );
or ( n4030 , n4021 , n4029 );
nand ( n4031 , n4017 , n4030 );
buf ( n4032 , n4031 );
and ( n4033 , n4011 , n4032 );
not ( n4034 , n4011 );
buf ( n4035 , n4032 );
not ( n4036 , n4035 );
buf ( n4037 , n4036 );
and ( n4038 , n4034 , n4037 );
nor ( n4039 , n4033 , n4038 );
and ( n4040 , n3974 , n4039 );
not ( n4041 , n3974 );
not ( n4042 , n4039 );
and ( n4043 , n4041 , n4042 );
nor ( n4044 , n4040 , n4043 );
buf ( n4045 , n4044 );
buf ( n4046 , n3331 );
not ( n4047 , n4046 );
buf ( n4048 , n1305 );
not ( n4049 , n4048 );
or ( n4050 , n4047 , n4049 );
buf ( n4051 , n1309 );
buf ( n4052 , n789 );
buf ( n4053 , n808 );
xor ( n4054 , n4052 , n4053 );
buf ( n4055 , n4054 );
buf ( n4056 , n4055 );
nand ( n4057 , n4051 , n4056 );
buf ( n4058 , n4057 );
buf ( n4059 , n4058 );
nand ( n4060 , n4050 , n4059 );
buf ( n4061 , n4060 );
buf ( n4062 , n4061 );
buf ( n4063 , n3349 );
not ( n4064 , n4063 );
buf ( n4065 , n2325 );
not ( n4066 , n4065 );
or ( n4067 , n4064 , n4066 );
buf ( n4068 , n2331 );
buf ( n4069 , n791 );
buf ( n4070 , n806 );
xor ( n4071 , n4069 , n4070 );
buf ( n4072 , n4071 );
buf ( n4073 , n4072 );
nand ( n4074 , n4068 , n4073 );
buf ( n4075 , n4074 );
buf ( n4076 , n4075 );
nand ( n4077 , n4067 , n4076 );
buf ( n4078 , n4077 );
buf ( n4079 , n4078 );
xor ( n4080 , n4062 , n4079 );
buf ( n4081 , n3619 );
not ( n4082 , n4081 );
buf ( n4083 , n1480 );
not ( n4084 , n4083 );
or ( n4085 , n4082 , n4084 );
buf ( n4086 , n1496 );
buf ( n4087 , n779 );
buf ( n4088 , n818 );
xor ( n4089 , n4087 , n4088 );
buf ( n4090 , n4089 );
buf ( n4091 , n4090 );
nand ( n4092 , n4086 , n4091 );
buf ( n4093 , n4092 );
buf ( n4094 , n4093 );
nand ( n4095 , n4085 , n4094 );
buf ( n4096 , n4095 );
buf ( n4097 , n4096 );
xor ( n4098 , n4080 , n4097 );
buf ( n4099 , n4098 );
buf ( n4100 , n4099 );
and ( n4101 , n4045 , n4100 );
not ( n4102 , n4045 );
buf ( n4103 , n4099 );
not ( n4104 , n4103 );
buf ( n4105 , n4104 );
buf ( n4106 , n4105 );
and ( n4107 , n4102 , n4106 );
nor ( n4108 , n4101 , n4107 );
buf ( n4109 , n4108 );
buf ( n4110 , n4109 );
buf ( n4111 , n3756 );
not ( n4112 , n4111 );
buf ( n4113 , n3293 );
not ( n4114 , n4113 );
buf ( n4115 , n3703 );
not ( n4116 , n4115 );
or ( n4117 , n4114 , n4116 );
buf ( n4118 , n3713 );
nand ( n4119 , n4117 , n4118 );
buf ( n4120 , n4119 );
buf ( n4121 , n4120 );
not ( n4122 , n4121 );
or ( n4123 , n4112 , n4122 );
buf ( n4124 , n3756 );
buf ( n4125 , n4120 );
or ( n4126 , n4124 , n4125 );
buf ( n4127 , n3733 );
nand ( n4128 , n4126 , n4127 );
buf ( n4129 , n4128 );
buf ( n4130 , n4129 );
nand ( n4131 , n4123 , n4130 );
buf ( n4132 , n4131 );
buf ( n4133 , n3409 );
not ( n4134 , n4133 );
buf ( n4135 , n3426 );
not ( n4136 , n4135 );
or ( n4137 , n4134 , n4136 );
buf ( n4138 , n3426 );
buf ( n4139 , n3409 );
or ( n4140 , n4138 , n4139 );
buf ( n4141 , n3390 );
nand ( n4142 , n4140 , n4141 );
buf ( n4143 , n4142 );
buf ( n4144 , n4143 );
nand ( n4145 , n4137 , n4144 );
buf ( n4146 , n4145 );
buf ( n4147 , n4146 );
not ( n4148 , n4147 );
buf ( n4149 , n4148 );
xor ( n4150 , n4132 , n4149 );
xor ( n4151 , n3644 , n3674 );
and ( n4152 , n4151 , n3695 );
and ( n4153 , n3644 , n3674 );
or ( n4154 , n4152 , n4153 );
buf ( n4155 , n4154 );
xnor ( n4156 , n4150 , n4155 );
buf ( n4157 , n4156 );
xor ( n4158 , n4110 , n4157 );
xor ( n4159 , n3373 , n3428 );
and ( n4160 , n4159 , n3435 );
and ( n4161 , n3373 , n3428 );
or ( n4162 , n4160 , n4161 );
buf ( n4163 , n4162 );
buf ( n4164 , n4163 );
xor ( n4165 , n4158 , n4164 );
buf ( n4166 , n4165 );
buf ( n4167 , n4166 );
xor ( n4168 , n3898 , n4167 );
buf ( n4169 , n3524 );
not ( n4170 , n4169 );
buf ( n4171 , n3537 );
not ( n4172 , n4171 );
or ( n4173 , n4170 , n4172 );
or ( n4174 , n3524 , n3537 );
nand ( n4175 , n4174 , n3548 );
buf ( n4176 , n4175 );
nand ( n4177 , n4173 , n4176 );
buf ( n4178 , n4177 );
buf ( n4179 , n4178 );
not ( n4180 , n4179 );
buf ( n4181 , n3589 );
not ( n4182 , n4181 );
buf ( n4183 , n1548 );
not ( n4184 , n4183 );
or ( n4185 , n4182 , n4184 );
buf ( n4186 , n1557 );
buf ( n4187 , n795 );
buf ( n4188 , n802 );
xor ( n4189 , n4187 , n4188 );
buf ( n4190 , n4189 );
buf ( n4191 , n4190 );
nand ( n4192 , n4186 , n4191 );
buf ( n4193 , n4192 );
buf ( n4194 , n4193 );
nand ( n4195 , n4185 , n4194 );
buf ( n4196 , n4195 );
buf ( n4197 , n3605 );
not ( n4198 , n4197 );
buf ( n4199 , n1522 );
not ( n4200 , n4199 );
or ( n4201 , n4198 , n4200 );
buf ( n4202 , n1449 );
buf ( n4203 , n793 );
buf ( n4204 , n804 );
xor ( n4205 , n4203 , n4204 );
buf ( n4206 , n4205 );
buf ( n4207 , n4206 );
nand ( n4208 , n4202 , n4207 );
buf ( n4209 , n4208 );
buf ( n4210 , n4209 );
nand ( n4211 , n4201 , n4210 );
buf ( n4212 , n4211 );
xor ( n4213 , n4196 , n4212 );
buf ( n4214 , n3465 );
not ( n4215 , n4214 );
buf ( n4216 , n3483 );
nand ( n4217 , n4215 , n4216 );
buf ( n4218 , n4217 );
and ( n4219 , n4213 , n4218 );
not ( n4220 , n4213 );
buf ( n4221 , n4218 );
not ( n4222 , n4221 );
buf ( n4223 , n4222 );
and ( n4224 , n4220 , n4223 );
nor ( n4225 , n4219 , n4224 );
buf ( n4226 , n4225 );
not ( n4227 , n4226 );
buf ( n4228 , n3667 );
not ( n4229 , n4228 );
buf ( n4230 , n3654 );
buf ( n4231 , n1218 );
nor ( n4232 , n4230 , n4231 );
buf ( n4233 , n4232 );
buf ( n4234 , n4233 );
not ( n4235 , n4234 );
or ( n4236 , n4229 , n4235 );
buf ( n4237 , n1218 );
buf ( n4238 , n797 );
buf ( n4239 , n800 );
xor ( n4240 , n4238 , n4239 );
buf ( n4241 , n4240 );
buf ( n4242 , n4241 );
nand ( n4243 , n4237 , n4242 );
buf ( n4244 , n4243 );
buf ( n4245 , n4244 );
nand ( n4246 , n4236 , n4245 );
buf ( n4247 , n4246 );
buf ( n4248 , n4247 );
buf ( n4249 , n3727 );
not ( n4250 , n4249 );
buf ( n4251 , n2523 );
not ( n4252 , n4251 );
or ( n4253 , n4250 , n4252 );
buf ( n4254 , n2532 );
buf ( n4255 , n781 );
buf ( n4256 , n816 );
xor ( n4257 , n4255 , n4256 );
buf ( n4258 , n4257 );
buf ( n4259 , n4258 );
nand ( n4260 , n4254 , n4259 );
buf ( n4261 , n4260 );
buf ( n4262 , n4261 );
nand ( n4263 , n4253 , n4262 );
buf ( n4264 , n4263 );
buf ( n4265 , n4264 );
xor ( n4266 , n4248 , n4265 );
buf ( n4267 , n3637 );
not ( n4268 , n4267 );
buf ( n4269 , n2790 );
not ( n4270 , n4269 );
or ( n4271 , n4268 , n4270 );
buf ( n4272 , n3255 );
xor ( n4273 , n824 , n773 );
buf ( n4274 , n4273 );
nand ( n4275 , n4272 , n4274 );
buf ( n4276 , n4275 );
buf ( n4277 , n4276 );
nand ( n4278 , n4271 , n4277 );
buf ( n4279 , n4278 );
buf ( n4280 , n4279 );
xor ( n4281 , n4266 , n4280 );
buf ( n4282 , n4281 );
buf ( n4283 , n4282 );
not ( n4284 , n4283 );
and ( n4285 , n4227 , n4284 );
buf ( n4286 , n4225 );
buf ( n4287 , n4282 );
and ( n4288 , n4286 , n4287 );
nor ( n4289 , n4285 , n4288 );
buf ( n4290 , n4289 );
buf ( n4291 , n4290 );
not ( n4292 , n4291 );
or ( n4293 , n4180 , n4292 );
buf ( n4294 , n4290 );
buf ( n4295 , n4178 );
or ( n4296 , n4294 , n4295 );
nand ( n4297 , n4293 , n4296 );
buf ( n4298 , n4297 );
buf ( n4299 , n4298 );
not ( n4300 , n3559 );
not ( n4301 , n3514 );
or ( n4302 , n4300 , n4301 );
buf ( n4303 , n3559 );
buf ( n4304 , n3514 );
or ( n4305 , n4303 , n4304 );
buf ( n4306 , n3553 );
nand ( n4307 , n4305 , n4306 );
buf ( n4308 , n4307 );
nand ( n4309 , n4302 , n4308 );
buf ( n4310 , n4309 );
xor ( n4311 , n4299 , n4310 );
xor ( n4312 , n3572 , n3578 );
and ( n4313 , n4312 , n3761 );
and ( n4314 , n3572 , n3578 );
or ( n4315 , n4313 , n4314 );
buf ( n4316 , n4315 );
buf ( n4317 , n4316 );
xor ( n4318 , n4311 , n4317 );
buf ( n4319 , n4318 );
buf ( n4320 , n4319 );
xor ( n4321 , n4168 , n4320 );
buf ( n4322 , n4321 );
buf ( n4323 , n4322 );
xor ( n4324 , n3809 , n4323 );
buf ( n4325 , n4324 );
buf ( n4326 , n4325 );
not ( n4327 , n4326 );
buf ( n4328 , n4327 );
buf ( n4329 , n4328 );
not ( n4330 , n4329 );
or ( n4331 , n3796 , n4330 );
buf ( n4332 , n4325 );
buf ( n4333 , n3794 );
not ( n4334 , n4333 );
buf ( n4335 , n4334 );
buf ( n4336 , n4335 );
nand ( n4337 , n4332 , n4336 );
buf ( n4338 , n4337 );
buf ( n4339 , n4338 );
nand ( n4340 , n4331 , n4339 );
buf ( n4341 , n4340 );
buf ( n4342 , n4341 );
or ( n4343 , n3789 , n4342 );
buf ( n4344 , n4343 );
buf ( n4345 , n4344 );
buf ( n4346 , n4345 );
buf ( n4347 , n4346 );
buf ( n4348 , n4347 );
nand ( n4349 , n3788 , n4341 );
buf ( n4350 , n4349 );
buf ( n4351 , n4350 );
buf ( n4352 , n4351 );
buf ( n4353 , n4352 );
nand ( n4354 , n4348 , n4353 );
buf ( n4355 , n4354 );
buf ( n4356 , n4355 );
not ( n4357 , n4356 );
xor ( n4358 , n1214 , n3321 );
xor ( n4359 , n4358 , n3784 );
buf ( n4360 , n4359 );
not ( n4361 , n4360 );
buf ( n4362 , n833 );
xor ( n4363 , n2561 , n3098 );
xor ( n4364 , n4363 , n3316 );
buf ( n4365 , n4364 );
buf ( n4366 , n4365 );
xor ( n4367 , n4362 , n4366 );
xor ( n4368 , n2564 , n2568 );
and ( n4369 , n4368 , n3089 );
not ( n4370 , n4368 );
not ( n4371 , n3089 );
and ( n4372 , n4370 , n4371 );
nor ( n4373 , n4369 , n4372 );
not ( n4374 , n4373 );
not ( n4375 , n1790 );
nand ( n4376 , n4375 , n1796 , n1867 );
not ( n4377 , n1867 );
nand ( n4378 , n4377 , n1721 , n1794 );
nand ( n4379 , n1866 , n1790 , n1796 );
nand ( n4380 , n1867 , n1790 , n1721 );
nand ( n4381 , n4376 , n4378 , n4379 , n4380 );
buf ( n4382 , n4381 );
buf ( n4383 , n786 );
buf ( n4384 , n818 );
xor ( n4385 , n4383 , n4384 );
buf ( n4386 , n4385 );
buf ( n4387 , n4386 );
not ( n4388 , n4387 );
buf ( n4389 , n818 );
buf ( n4390 , n819 );
xnor ( n4391 , n4389 , n4390 );
buf ( n4392 , n4391 );
buf ( n4393 , n4392 );
buf ( n4394 , n1478 );
nor ( n4395 , n4393 , n4394 );
buf ( n4396 , n4395 );
buf ( n4397 , n4396 );
not ( n4398 , n4397 );
or ( n4399 , n4388 , n4398 );
buf ( n4400 , n1496 );
buf ( n4401 , n2748 );
nand ( n4402 , n4400 , n4401 );
buf ( n4403 , n4402 );
buf ( n4404 , n4403 );
nand ( n4405 , n4399 , n4404 );
buf ( n4406 , n4405 );
buf ( n4407 , n4406 );
buf ( n4408 , n778 );
buf ( n4409 , n826 );
xor ( n4410 , n4408 , n4409 );
buf ( n4411 , n4410 );
buf ( n4412 , n4411 );
not ( n4413 , n4412 );
buf ( n4414 , n2364 );
not ( n4415 , n4414 );
or ( n4416 , n4413 , n4415 );
buf ( n4417 , n2366 );
buf ( n4418 , n1374 );
nand ( n4419 , n4417 , n4418 );
buf ( n4420 , n4419 );
buf ( n4421 , n4420 );
nand ( n4422 , n4416 , n4421 );
buf ( n4423 , n4422 );
buf ( n4424 , n4423 );
xor ( n4425 , n4407 , n4424 );
not ( n4426 , n2773 );
not ( n4427 , n1249 );
or ( n4428 , n4426 , n4427 );
not ( n4429 , n3841 );
xor ( n4430 , n777 , n828 );
nand ( n4431 , n4429 , n1237 , n4430 );
nand ( n4432 , n4428 , n4431 );
buf ( n4433 , n4432 );
buf ( n4434 , n799 );
buf ( n4435 , n807 );
or ( n4436 , n4434 , n4435 );
buf ( n4437 , n808 );
nand ( n4438 , n4436 , n4437 );
buf ( n4439 , n4438 );
buf ( n4440 , n799 );
buf ( n4441 , n807 );
nand ( n4442 , n4440 , n4441 );
buf ( n4443 , n4442 );
and ( n4444 , n4439 , n4443 , n806 );
buf ( n4445 , n4444 );
and ( n4446 , n4433 , n4445 );
buf ( n4447 , n4446 );
buf ( n4448 , n4447 );
and ( n4449 , n4425 , n4448 );
and ( n4450 , n4407 , n4424 );
or ( n4451 , n4449 , n4450 );
buf ( n4452 , n4451 );
buf ( n4453 , n4452 );
xor ( n4454 , n2055 , n2077 );
xor ( n4455 , n4454 , n2125 );
buf ( n4456 , n4455 );
buf ( n4457 , n4456 );
xor ( n4458 , n4453 , n4457 );
xor ( n4459 , n2761 , n2763 );
xor ( n4460 , n4459 , n2817 );
buf ( n4461 , n4460 );
buf ( n4462 , n4461 );
and ( n4463 , n4458 , n4462 );
and ( n4464 , n4453 , n4457 );
or ( n4465 , n4463 , n4464 );
buf ( n4466 , n4465 );
buf ( n4467 , n4466 );
xor ( n4468 , n4382 , n4467 );
xor ( n4469 , n2889 , n2907 );
xor ( n4470 , n4469 , n2927 );
buf ( n4471 , n4470 );
buf ( n4472 , n4471 );
buf ( n4473 , n799 );
buf ( n4474 , n806 );
xor ( n4475 , n4473 , n4474 );
buf ( n4476 , n4475 );
buf ( n4477 , n4476 );
not ( n4478 , n4477 );
buf ( n4479 , n2325 );
not ( n4480 , n4479 );
or ( n4481 , n4478 , n4480 );
buf ( n4482 , n2331 );
buf ( n4483 , n2976 );
nand ( n4484 , n4482 , n4483 );
buf ( n4485 , n4484 );
buf ( n4486 , n4485 );
nand ( n4487 , n4481 , n4486 );
buf ( n4488 , n4487 );
buf ( n4489 , n4488 );
buf ( n4490 , n779 );
buf ( n4491 , n826 );
xor ( n4492 , n4490 , n4491 );
buf ( n4493 , n4492 );
buf ( n4494 , n4493 );
not ( n4495 , n4494 );
not ( n4496 , n1779 );
buf ( n4497 , n4496 );
not ( n4498 , n4497 );
or ( n4499 , n4495 , n4498 );
buf ( n4500 , n1771 );
buf ( n4501 , n4411 );
nand ( n4502 , n4500 , n4501 );
buf ( n4503 , n4502 );
buf ( n4504 , n4503 );
nand ( n4505 , n4499 , n4504 );
buf ( n4506 , n4505 );
buf ( n4507 , n4506 );
xor ( n4508 , n4489 , n4507 );
buf ( n4509 , n787 );
buf ( n4510 , n818 );
xor ( n4511 , n4509 , n4510 );
buf ( n4512 , n4511 );
buf ( n4513 , n4512 );
not ( n4514 , n4513 );
buf ( n4515 , n1480 );
not ( n4516 , n4515 );
or ( n4517 , n4514 , n4516 );
buf ( n4518 , n1496 );
buf ( n4519 , n4386 );
nand ( n4520 , n4518 , n4519 );
buf ( n4521 , n4520 );
buf ( n4522 , n4521 );
nand ( n4523 , n4517 , n4522 );
buf ( n4524 , n4523 );
buf ( n4525 , n4524 );
and ( n4526 , n4508 , n4525 );
and ( n4527 , n4489 , n4507 );
or ( n4528 , n4526 , n4527 );
buf ( n4529 , n4528 );
buf ( n4530 , n4529 );
xor ( n4531 , n4472 , n4530 );
xor ( n4532 , n2769 , n2786 );
xor ( n4533 , n4532 , n2812 );
buf ( n4534 , n4533 );
buf ( n4535 , n4534 );
and ( n4536 , n4531 , n4535 );
and ( n4537 , n4472 , n4530 );
or ( n4538 , n4536 , n4537 );
buf ( n4539 , n4538 );
buf ( n4540 , n4539 );
not ( n4541 , n2875 );
not ( n4542 , n4541 );
not ( n4543 , n2995 );
not ( n4544 , n2931 );
not ( n4545 , n4544 );
or ( n4546 , n4543 , n4545 );
nand ( n4547 , n2996 , n2931 );
nand ( n4548 , n4546 , n4547 );
not ( n4549 , n4548 );
or ( n4550 , n4542 , n4549 );
or ( n4551 , n4541 , n4548 );
nand ( n4552 , n4550 , n4551 );
buf ( n4553 , n4552 );
or ( n4554 , n4540 , n4553 );
xor ( n4555 , n783 , n822 );
not ( n4556 , n4555 );
not ( n4557 , n2098 );
or ( n4558 , n4556 , n4557 );
buf ( n4559 , n3745 );
buf ( n4560 , n2860 );
nand ( n4561 , n4559 , n4560 );
buf ( n4562 , n4561 );
nand ( n4563 , n4558 , n4562 );
not ( n4564 , n4563 );
xor ( n4565 , n810 , n795 );
buf ( n4566 , n4565 );
not ( n4567 , n4566 );
buf ( n4568 , n1667 );
not ( n4569 , n4568 );
buf ( n4570 , n4569 );
buf ( n4571 , n4570 );
not ( n4572 , n4571 );
or ( n4573 , n4567 , n4572 );
buf ( n4574 , n1679 );
buf ( n4575 , n2890 );
nand ( n4576 , n4574 , n4575 );
buf ( n4577 , n4576 );
buf ( n4578 , n4577 );
nand ( n4579 , n4573 , n4578 );
buf ( n4580 , n4579 );
not ( n4581 , n4580 );
or ( n4582 , n4564 , n4581 );
buf ( n4583 , n4580 );
buf ( n4584 , n4563 );
nor ( n4585 , n4583 , n4584 );
buf ( n4586 , n4585 );
xor ( n4587 , n812 , n793 );
buf ( n4588 , n4587 );
not ( n4589 , n4588 );
buf ( n4590 , n2066 );
not ( n4591 , n4590 );
or ( n4592 , n4589 , n4591 );
buf ( n4593 , n3379 );
buf ( n4594 , n2912 );
nand ( n4595 , n4593 , n4594 );
buf ( n4596 , n4595 );
buf ( n4597 , n4596 );
nand ( n4598 , n4592 , n4597 );
buf ( n4599 , n4598 );
buf ( n4600 , n4599 );
not ( n4601 , n4600 );
buf ( n4602 , n4601 );
or ( n4603 , n4586 , n4602 );
nand ( n4604 , n4582 , n4603 );
buf ( n4605 , n791 );
buf ( n4606 , n814 );
xor ( n4607 , n4605 , n4606 );
buf ( n4608 , n4607 );
buf ( n4609 , n4608 );
not ( n4610 , n4609 );
buf ( n4611 , n2612 );
not ( n4612 , n4611 );
or ( n4613 , n4610 , n4612 );
buf ( n4614 , n1937 );
buf ( n4615 , n2827 );
nand ( n4616 , n4614 , n4615 );
buf ( n4617 , n4616 );
buf ( n4618 , n4617 );
nand ( n4619 , n4613 , n4618 );
buf ( n4620 , n4619 );
buf ( n4621 , n4620 );
not ( n4622 , n4621 );
buf ( n4623 , n781 );
buf ( n4624 , n824 );
xor ( n4625 , n4623 , n4624 );
buf ( n4626 , n4625 );
buf ( n4627 , n4626 );
not ( n4628 , n4627 );
buf ( n4629 , n2790 );
not ( n4630 , n4629 );
or ( n4631 , n4628 , n4630 );
buf ( n4632 , n3255 );
buf ( n4633 , n2798 );
nand ( n4634 , n4632 , n4633 );
buf ( n4635 , n4634 );
buf ( n4636 , n4635 );
nand ( n4637 , n4631 , n4636 );
buf ( n4638 , n4637 );
buf ( n4639 , n4638 );
not ( n4640 , n4639 );
or ( n4641 , n4622 , n4640 );
buf ( n4642 , n4638 );
buf ( n4643 , n4620 );
or ( n4644 , n4642 , n4643 );
buf ( n4645 , n789 );
buf ( n4646 , n816 );
xor ( n4647 , n4645 , n4646 );
buf ( n4648 , n4647 );
buf ( n4649 , n4648 );
not ( n4650 , n4649 );
buf ( n4651 , n2526 );
not ( n4652 , n4651 );
or ( n4653 , n4650 , n4652 );
buf ( n4654 , n2010 );
buf ( n4655 , n2843 );
nand ( n4656 , n4654 , n4655 );
buf ( n4657 , n4656 );
buf ( n4658 , n4657 );
nand ( n4659 , n4653 , n4658 );
buf ( n4660 , n4659 );
buf ( n4661 , n4660 );
nand ( n4662 , n4644 , n4661 );
buf ( n4663 , n4662 );
buf ( n4664 , n4663 );
nand ( n4665 , n4641 , n4664 );
buf ( n4666 , n4665 );
xor ( n4667 , n4604 , n4666 );
buf ( n4668 , n775 );
buf ( n4669 , n830 );
xor ( n4670 , n4668 , n4669 );
buf ( n4671 , n4670 );
buf ( n4672 , n4671 );
not ( n4673 , n4672 );
buf ( n4674 , n1630 );
not ( n4675 , n4674 );
or ( n4676 , n4673 , n4675 );
buf ( n4677 , n2881 );
buf ( n4678 , n831 );
nand ( n4679 , n4677 , n4678 );
buf ( n4680 , n4679 );
buf ( n4681 , n4680 );
nand ( n4682 , n4676 , n4681 );
buf ( n4683 , n4682 );
buf ( n4684 , n4683 );
buf ( n4685 , n797 );
buf ( n4686 , n808 );
xor ( n4687 , n4685 , n4686 );
buf ( n4688 , n4687 );
buf ( n4689 , n4688 );
not ( n4690 , n4689 );
buf ( n4691 , n2235 );
not ( n4692 , n4691 );
or ( n4693 , n4690 , n4692 );
buf ( n4694 , n1309 );
buf ( n4695 , n2936 );
nand ( n4696 , n4694 , n4695 );
buf ( n4697 , n4696 );
buf ( n4698 , n4697 );
nand ( n4699 , n4693 , n4698 );
buf ( n4700 , n4699 );
buf ( n4701 , n4700 );
xor ( n4702 , n4684 , n4701 );
not ( n4703 , n1346 );
not ( n4704 , n2954 );
or ( n4705 , n4703 , n4704 );
buf ( n4706 , n785 );
buf ( n4707 , n820 );
xnor ( n4708 , n4706 , n4707 );
buf ( n4709 , n4708 );
or ( n4710 , n2678 , n4709 );
nand ( n4711 , n4705 , n4710 );
buf ( n4712 , n4711 );
and ( n4713 , n4702 , n4712 );
and ( n4714 , n4684 , n4701 );
or ( n4715 , n4713 , n4714 );
buf ( n4716 , n4715 );
and ( n4717 , n4667 , n4716 );
and ( n4718 , n4604 , n4666 );
or ( n4719 , n4717 , n4718 );
buf ( n4720 , n4719 );
nand ( n4721 , n4554 , n4720 );
buf ( n4722 , n4721 );
buf ( n4723 , n4722 );
buf ( n4724 , n4539 );
buf ( n4725 , n4552 );
nand ( n4726 , n4724 , n4725 );
buf ( n4727 , n4726 );
buf ( n4728 , n4727 );
nand ( n4729 , n4723 , n4728 );
buf ( n4730 , n4729 );
buf ( n4731 , n4730 );
and ( n4732 , n4468 , n4731 );
and ( n4733 , n4382 , n4467 );
or ( n4734 , n4732 , n4733 );
buf ( n4735 , n4734 );
buf ( n4736 , n4735 );
not ( n4737 , n4736 );
buf ( n4738 , n4737 );
not ( n4739 , n4738 );
and ( n4740 , n4374 , n4739 );
buf ( n4741 , n4735 );
not ( n4742 , n4741 );
buf ( n4743 , n4373 );
nand ( n4744 , n4742 , n4743 );
buf ( n4745 , n4744 );
xor ( n4746 , n2744 , n2822 );
xor ( n4747 , n4746 , n3003 );
buf ( n4748 , n4747 );
buf ( n4749 , n4748 );
xor ( n4750 , n4407 , n4424 );
xor ( n4751 , n4750 , n4448 );
buf ( n4752 , n4751 );
not ( n4753 , n4752 );
buf ( n4754 , n4753 );
not ( n4755 , n4754 );
not ( n4756 , n2989 );
not ( n4757 , n4756 );
not ( n4758 , n2966 );
not ( n4759 , n4758 );
or ( n4760 , n4757 , n4759 );
nand ( n4761 , n2989 , n2966 );
nand ( n4762 , n4760 , n4761 );
buf ( n4763 , n2948 );
not ( n4764 , n4763 );
buf ( n4765 , n4764 );
or ( n4766 , n4762 , n4765 );
nand ( n4767 , n4762 , n4765 );
nand ( n4768 , n4766 , n4767 );
buf ( n4769 , n4768 );
not ( n4770 , n4769 );
or ( n4771 , n4755 , n4770 );
xor ( n4772 , n2839 , n2855 );
xor ( n4773 , n4772 , n2872 );
buf ( n4774 , n4773 );
buf ( n4775 , n4774 );
nand ( n4776 , n4771 , n4775 );
buf ( n4777 , n4776 );
buf ( n4778 , n4752 );
not ( n4779 , n4768 );
buf ( n4780 , n4779 );
nand ( n4781 , n4778 , n4780 );
buf ( n4782 , n4781 );
and ( n4783 , n4777 , n4782 );
buf ( n4784 , n4783 );
not ( n4785 , n4784 );
and ( n4786 , n3072 , n3026 );
not ( n4787 , n3072 );
and ( n4788 , n4787 , n3054 );
nor ( n4789 , n4786 , n4788 );
and ( n4790 , n4789 , n3049 );
not ( n4791 , n4789 );
and ( n4792 , n4791 , n3046 );
nor ( n4793 , n4790 , n4792 );
buf ( n4794 , n4793 );
not ( n4795 , n4794 );
or ( n4796 , n4785 , n4795 );
xor ( n4797 , n4453 , n4457 );
xor ( n4798 , n4797 , n4462 );
buf ( n4799 , n4798 );
buf ( n4800 , n4799 );
nand ( n4801 , n4796 , n4800 );
buf ( n4802 , n4801 );
buf ( n4803 , n4802 );
buf ( n4804 , n4793 );
not ( n4805 , n4804 );
buf ( n4806 , n4777 );
buf ( n4807 , n4782 );
nand ( n4808 , n4806 , n4807 );
buf ( n4809 , n4808 );
buf ( n4810 , n4809 );
nand ( n4811 , n4805 , n4810 );
buf ( n4812 , n4811 );
buf ( n4813 , n4812 );
nand ( n4814 , n4803 , n4813 );
buf ( n4815 , n4814 );
buf ( n4816 , n4815 );
xor ( n4817 , n4749 , n4816 );
buf ( n4818 , n3077 );
not ( n4819 , n4818 );
buf ( n4820 , n3018 );
not ( n4821 , n4820 );
or ( n4822 , n4819 , n4821 );
buf ( n4823 , n3077 );
buf ( n4824 , n3018 );
or ( n4825 , n4823 , n4824 );
nand ( n4826 , n4822 , n4825 );
buf ( n4827 , n4826 );
buf ( n4828 , n4827 );
buf ( n4829 , n3011 );
xor ( n4830 , n4828 , n4829 );
buf ( n4831 , n4830 );
buf ( n4832 , n4831 );
and ( n4833 , n4817 , n4832 );
and ( n4834 , n4749 , n4816 );
or ( n4835 , n4833 , n4834 );
buf ( n4836 , n4835 );
buf ( n4837 , n4836 );
and ( n4838 , n4745 , n4837 );
nor ( n4839 , n4740 , n4838 );
buf ( n4840 , n4839 );
not ( n4841 , n4840 );
buf ( n4842 , n4841 );
buf ( n4843 , n4842 );
and ( n4844 , n4367 , n4843 );
and ( n4845 , n4362 , n4366 );
or ( n4846 , n4844 , n4845 );
buf ( n4847 , n4846 );
not ( n4848 , n4847 );
and ( n4849 , n4361 , n4848 );
xor ( n4850 , n4362 , n4366 );
xor ( n4851 , n4850 , n4843 );
buf ( n4852 , n4851 );
buf ( n4853 , n4852 );
buf ( n4854 , n834 );
xor ( n4855 , n4382 , n4467 );
xor ( n4856 , n4855 , n4731 );
buf ( n4857 , n4856 );
buf ( n4858 , n4857 );
xor ( n4859 , n2875 , n4548 );
xnor ( n4860 , n4859 , n4719 );
not ( n4861 , n4539 );
and ( n4862 , n4860 , n4861 );
not ( n4863 , n4860 );
and ( n4864 , n4863 , n4539 );
nor ( n4865 , n4862 , n4864 );
not ( n4866 , n4865 );
xor ( n4867 , n4604 , n4666 );
xor ( n4868 , n4867 , n4716 );
buf ( n4869 , n4868 );
xor ( n4870 , n4472 , n4530 );
xor ( n4871 , n4870 , n4535 );
buf ( n4872 , n4871 );
buf ( n4873 , n4872 );
or ( n4874 , n4869 , n4873 );
and ( n4875 , n4773 , n4752 );
not ( n4876 , n4773 );
and ( n4877 , n4876 , n4753 );
nor ( n4878 , n4875 , n4877 );
buf ( n4879 , n4878 );
buf ( n4880 , n4779 );
and ( n4881 , n4879 , n4880 );
not ( n4882 , n4879 );
not ( n4883 , n4779 );
buf ( n4884 , n4883 );
and ( n4885 , n4882 , n4884 );
nor ( n4886 , n4881 , n4885 );
buf ( n4887 , n4886 );
buf ( n4888 , n4887 );
nand ( n4889 , n4874 , n4888 );
buf ( n4890 , n4889 );
buf ( n4891 , n4872 );
buf ( n4892 , n4868 );
nand ( n4893 , n4891 , n4892 );
buf ( n4894 , n4893 );
nand ( n4895 , n4890 , n4894 );
not ( n4896 , n4895 );
not ( n4897 , n4896 );
not ( n4898 , n4897 );
or ( n4899 , n4866 , n4898 );
or ( n4900 , n4897 , n4865 );
xor ( n4901 , n4563 , n4599 );
xor ( n4902 , n4901 , n4580 );
xor ( n4903 , n4684 , n4701 );
xor ( n4904 , n4903 , n4712 );
buf ( n4905 , n4904 );
xor ( n4906 , n4902 , n4905 );
xnor ( n4907 , n4638 , n4660 );
xnor ( n4908 , n4620 , n4907 );
and ( n4909 , n4906 , n4908 );
and ( n4910 , n4902 , n4905 );
or ( n4911 , n4909 , n4910 );
not ( n4912 , n4911 );
buf ( n4913 , n792 );
buf ( n4914 , n814 );
xor ( n4915 , n4913 , n4914 );
buf ( n4916 , n4915 );
buf ( n4917 , n4916 );
not ( n4918 , n4917 );
buf ( n4919 , n3703 );
not ( n4920 , n4919 );
or ( n4921 , n4918 , n4920 );
buf ( n4922 , n1940 );
buf ( n4923 , n4608 );
nand ( n4924 , n4922 , n4923 );
buf ( n4925 , n4924 );
buf ( n4926 , n4925 );
nand ( n4927 , n4921 , n4926 );
buf ( n4928 , n4927 );
buf ( n4929 , n4928 );
buf ( n4930 , n790 );
buf ( n4931 , n816 );
xor ( n4932 , n4930 , n4931 );
buf ( n4933 , n4932 );
buf ( n4934 , n4933 );
not ( n4935 , n4934 );
buf ( n4936 , n3719 );
not ( n4937 , n4936 );
or ( n4938 , n4935 , n4937 );
buf ( n4939 , n2535 );
buf ( n4940 , n4648 );
nand ( n4941 , n4939 , n4940 );
buf ( n4942 , n4941 );
buf ( n4943 , n4942 );
nand ( n4944 , n4938 , n4943 );
buf ( n4945 , n4944 );
buf ( n4946 , n4945 );
xor ( n4947 , n4929 , n4946 );
xor ( n4948 , n822 , n784 );
buf ( n4949 , n4948 );
not ( n4950 , n4949 );
buf ( n4951 , n2101 );
not ( n4952 , n4951 );
or ( n4953 , n4950 , n4952 );
nand ( n4954 , n2113 , n4555 );
buf ( n4955 , n4954 );
nand ( n4956 , n4953 , n4955 );
buf ( n4957 , n4956 );
buf ( n4958 , n4957 );
and ( n4959 , n4947 , n4958 );
and ( n4960 , n4929 , n4946 );
or ( n4961 , n4959 , n4960 );
buf ( n4962 , n4961 );
buf ( n4963 , n4962 );
not ( n4964 , n4963 );
buf ( n4965 , n4964 );
buf ( n4966 , n4965 );
xor ( n4967 , n830 , n776 );
buf ( n4968 , n4967 );
not ( n4969 , n4968 );
buf ( n4970 , n1161 );
not ( n4971 , n4970 );
or ( n4972 , n4969 , n4971 );
buf ( n4973 , n4671 );
buf ( n4974 , n831 );
nand ( n4975 , n4973 , n4974 );
buf ( n4976 , n4975 );
buf ( n4977 , n4976 );
nand ( n4978 , n4972 , n4977 );
buf ( n4979 , n4978 );
buf ( n4980 , n4979 );
xor ( n4981 , n810 , n796 );
buf ( n4982 , n4981 );
not ( n4983 , n4982 );
buf ( n4984 , n1670 );
not ( n4985 , n4984 );
or ( n4986 , n4983 , n4985 );
buf ( n4987 , n2647 );
buf ( n4988 , n4565 );
nand ( n4989 , n4987 , n4988 );
buf ( n4990 , n4989 );
buf ( n4991 , n4990 );
nand ( n4992 , n4986 , n4991 );
buf ( n4993 , n4992 );
buf ( n4994 , n4993 );
xor ( n4995 , n4980 , n4994 );
buf ( n4996 , n794 );
buf ( n4997 , n812 );
xor ( n4998 , n4996 , n4997 );
buf ( n4999 , n4998 );
buf ( n5000 , n4999 );
not ( n5001 , n5000 );
buf ( n5002 , n2066 );
not ( n5003 , n5002 );
or ( n5004 , n5001 , n5003 );
buf ( n5005 , n1693 );
buf ( n5006 , n4587 );
nand ( n5007 , n5005 , n5006 );
buf ( n5008 , n5007 );
buf ( n5009 , n5008 );
nand ( n5010 , n5004 , n5009 );
buf ( n5011 , n5010 );
buf ( n5012 , n5011 );
and ( n5013 , n4995 , n5012 );
and ( n5014 , n4980 , n4994 );
or ( n5015 , n5013 , n5014 );
buf ( n5016 , n5015 );
xor ( n5017 , n4444 , n4432 );
nor ( n5018 , n5016 , n5017 );
buf ( n5019 , n5018 );
or ( n5020 , n4966 , n5019 );
nand ( n5021 , n5016 , n5017 );
buf ( n5022 , n5021 );
nand ( n5023 , n5020 , n5022 );
buf ( n5024 , n5023 );
not ( n5025 , n5024 );
buf ( n5026 , n1409 );
buf ( n5027 , n799 );
and ( n5028 , n5026 , n5027 );
buf ( n5029 , n5028 );
buf ( n5030 , n5029 );
buf ( n5031 , n778 );
buf ( n5032 , n828 );
xor ( n5033 , n5031 , n5032 );
buf ( n5034 , n5033 );
buf ( n5035 , n5034 );
not ( n5036 , n5035 );
buf ( n5037 , n1239 );
not ( n5038 , n5037 );
or ( n5039 , n5036 , n5038 );
buf ( n5040 , n1249 );
buf ( n5041 , n4430 );
nand ( n5042 , n5040 , n5041 );
buf ( n5043 , n5042 );
buf ( n5044 , n5043 );
nand ( n5045 , n5039 , n5044 );
buf ( n5046 , n5045 );
buf ( n5047 , n5046 );
xor ( n5048 , n5030 , n5047 );
xor ( n5049 , n824 , n782 );
buf ( n5050 , n5049 );
not ( n5051 , n5050 );
buf ( n5052 , n1965 );
not ( n5053 , n5052 );
or ( n5054 , n5051 , n5053 );
buf ( n5055 , n3255 );
buf ( n5056 , n4626 );
nand ( n5057 , n5055 , n5056 );
buf ( n5058 , n5057 );
buf ( n5059 , n5058 );
nand ( n5060 , n5054 , n5059 );
buf ( n5061 , n5060 );
buf ( n5062 , n5061 );
and ( n5063 , n5048 , n5062 );
and ( n5064 , n5030 , n5047 );
or ( n5065 , n5063 , n5064 );
buf ( n5066 , n5065 );
buf ( n5067 , n5066 );
buf ( n5068 , n798 );
buf ( n5069 , n808 );
xor ( n5070 , n5068 , n5069 );
buf ( n5071 , n5070 );
buf ( n5072 , n5071 );
not ( n5073 , n5072 );
buf ( n5074 , n1305 );
not ( n5075 , n5074 );
or ( n5076 , n5073 , n5075 );
buf ( n5077 , n1309 );
buf ( n5078 , n4688 );
nand ( n5079 , n5077 , n5078 );
buf ( n5080 , n5079 );
buf ( n5081 , n5080 );
nand ( n5082 , n5076 , n5081 );
buf ( n5083 , n5082 );
buf ( n5084 , n5083 );
buf ( n5085 , n786 );
buf ( n5086 , n820 );
xor ( n5087 , n5085 , n5086 );
buf ( n5088 , n5087 );
not ( n5089 , n5088 );
not ( n5090 , n1338 );
or ( n5091 , n5089 , n5090 );
not ( n5092 , n4709 );
nand ( n5093 , n5092 , n3986 );
nand ( n5094 , n5091 , n5093 );
buf ( n5095 , n5094 );
xor ( n5096 , n5084 , n5095 );
not ( n5097 , n4493 );
or ( n5098 , n5097 , n2371 );
and ( n5099 , n826 , n780 );
not ( n5100 , n826 );
and ( n5101 , n5100 , n1321 );
nor ( n5102 , n5099 , n5101 );
nand ( n5103 , n5102 , n1356 );
nand ( n5104 , n5098 , n5103 );
buf ( n5105 , n5104 );
and ( n5106 , n5096 , n5105 );
and ( n5107 , n5084 , n5095 );
or ( n5108 , n5106 , n5107 );
buf ( n5109 , n5108 );
buf ( n5110 , n5109 );
xor ( n5111 , n5067 , n5110 );
xor ( n5112 , n4489 , n4507 );
xor ( n5113 , n5112 , n4525 );
buf ( n5114 , n5113 );
buf ( n5115 , n5114 );
and ( n5116 , n5111 , n5115 );
and ( n5117 , n5067 , n5110 );
or ( n5118 , n5116 , n5117 );
buf ( n5119 , n5118 );
not ( n5120 , n5119 );
nand ( n5121 , n5025 , n5120 );
not ( n5122 , n5121 );
or ( n5123 , n4912 , n5122 );
not ( n5124 , n5025 );
nand ( n5125 , n5124 , n5119 );
nand ( n5126 , n5123 , n5125 );
buf ( n5127 , n5126 );
nand ( n5128 , n4900 , n5127 );
nand ( n5129 , n4899 , n5128 );
buf ( n5130 , n5129 );
xor ( n5131 , n4858 , n5130 );
xor ( n5132 , n4749 , n4816 );
xor ( n5133 , n5132 , n4832 );
buf ( n5134 , n5133 );
buf ( n5135 , n5134 );
and ( n5136 , n5131 , n5135 );
and ( n5137 , n4858 , n5130 );
or ( n5138 , n5136 , n5137 );
buf ( n5139 , n5138 );
buf ( n5140 , n5139 );
xor ( n5141 , n4854 , n5140 );
not ( n5142 , n4373 );
buf ( n5143 , n5142 );
not ( n5144 , n5143 );
buf ( n5145 , n4836 );
not ( n5146 , n5145 );
buf ( n5147 , n4738 );
not ( n5148 , n5147 );
and ( n5149 , n5146 , n5148 );
buf ( n5150 , n4836 );
buf ( n5151 , n4738 );
and ( n5152 , n5150 , n5151 );
nor ( n5153 , n5149 , n5152 );
buf ( n5154 , n5153 );
buf ( n5155 , n5154 );
not ( n5156 , n5155 );
or ( n5157 , n5144 , n5156 );
buf ( n5158 , n5154 );
not ( n5159 , n5158 );
buf ( n5160 , n5159 );
buf ( n5161 , n5160 );
not ( n5162 , n5142 );
buf ( n5163 , n5162 );
nand ( n5164 , n5161 , n5163 );
buf ( n5165 , n5164 );
buf ( n5166 , n5165 );
nand ( n5167 , n5157 , n5166 );
buf ( n5168 , n5167 );
buf ( n5169 , n5168 );
and ( n5170 , n5141 , n5169 );
and ( n5171 , n4854 , n5140 );
or ( n5172 , n5170 , n5171 );
buf ( n5173 , n5172 );
buf ( n5174 , n5173 );
nor ( n5175 , n4853 , n5174 );
buf ( n5176 , n5175 );
nor ( n5177 , n4849 , n5176 );
buf ( n5178 , n5177 );
xor ( n5179 , n4854 , n5140 );
xor ( n5180 , n5179 , n5169 );
buf ( n5181 , n5180 );
buf ( n5182 , n5181 );
not ( n5183 , n5182 );
buf ( n5184 , n5183 );
buf ( n5185 , n5184 );
buf ( n5186 , n835 );
buf ( n5187 , n4793 );
not ( n5188 , n5187 );
buf ( n5189 , n5188 );
xor ( n5190 , n4783 , n5189 );
xnor ( n5191 , n5190 , n4799 );
buf ( n5192 , n5191 );
buf ( n5193 , n788 );
buf ( n5194 , n818 );
xor ( n5195 , n5193 , n5194 );
buf ( n5196 , n5195 );
buf ( n5197 , n5196 );
not ( n5198 , n5197 );
buf ( n5199 , n1480 );
not ( n5200 , n5199 );
or ( n5201 , n5198 , n5200 );
buf ( n5202 , n1496 );
buf ( n5203 , n4512 );
nand ( n5204 , n5202 , n5203 );
buf ( n5205 , n5204 );
buf ( n5206 , n5205 );
nand ( n5207 , n5201 , n5206 );
buf ( n5208 , n5207 );
buf ( n5209 , n5208 );
buf ( n5210 , n799 );
buf ( n5211 , n809 );
or ( n5212 , n5210 , n5211 );
buf ( n5213 , n810 );
nand ( n5214 , n5212 , n5213 );
buf ( n5215 , n5214 );
buf ( n5216 , n5215 );
buf ( n5217 , n799 );
buf ( n5218 , n809 );
nand ( n5219 , n5217 , n5218 );
buf ( n5220 , n5219 );
buf ( n5221 , n5220 );
buf ( n5222 , n808 );
and ( n5223 , n5216 , n5221 , n5222 );
buf ( n5224 , n5223 );
buf ( n5225 , n5224 );
buf ( n5226 , n779 );
buf ( n5227 , n828 );
xor ( n5228 , n5226 , n5227 );
buf ( n5229 , n5228 );
buf ( n5230 , n5229 );
not ( n5231 , n5230 );
buf ( n5232 , n1239 );
not ( n5233 , n5232 );
or ( n5234 , n5231 , n5233 );
buf ( n5235 , n1249 );
buf ( n5236 , n5034 );
nand ( n5237 , n5235 , n5236 );
buf ( n5238 , n5237 );
buf ( n5239 , n5238 );
nand ( n5240 , n5234 , n5239 );
buf ( n5241 , n5240 );
buf ( n5242 , n5241 );
and ( n5243 , n5225 , n5242 );
buf ( n5244 , n5243 );
buf ( n5245 , n5244 );
xor ( n5246 , n5209 , n5245 );
buf ( n5247 , n795 );
buf ( n5248 , n812 );
xor ( n5249 , n5247 , n5248 );
buf ( n5250 , n5249 );
buf ( n5251 , n5250 );
not ( n5252 , n5251 );
buf ( n5253 , n1712 );
not ( n5254 , n5253 );
or ( n5255 , n5252 , n5254 );
buf ( n5256 , n1693 );
buf ( n5257 , n4999 );
nand ( n5258 , n5256 , n5257 );
buf ( n5259 , n5258 );
buf ( n5260 , n5259 );
nand ( n5261 , n5255 , n5260 );
buf ( n5262 , n5261 );
buf ( n5263 , n5262 );
xor ( n5264 , n810 , n797 );
buf ( n5265 , n5264 );
not ( n5266 , n5265 );
buf ( n5267 , n2641 );
not ( n5268 , n5267 );
or ( n5269 , n5266 , n5268 );
buf ( n5270 , n1676 );
not ( n5271 , n5270 );
buf ( n5272 , n5271 );
buf ( n5273 , n5272 );
buf ( n5274 , n4981 );
nand ( n5275 , n5273 , n5274 );
buf ( n5276 , n5275 );
buf ( n5277 , n5276 );
nand ( n5278 , n5269 , n5277 );
buf ( n5279 , n5278 );
buf ( n5280 , n5279 );
xor ( n5281 , n5263 , n5280 );
xor ( n5282 , n822 , n785 );
buf ( n5283 , n5282 );
not ( n5284 , n5283 );
buf ( n5285 , n3739 );
not ( n5286 , n5285 );
or ( n5287 , n5284 , n5286 );
buf ( n5288 , n2113 );
buf ( n5289 , n4948 );
nand ( n5290 , n5288 , n5289 );
buf ( n5291 , n5290 );
buf ( n5292 , n5291 );
nand ( n5293 , n5287 , n5292 );
buf ( n5294 , n5293 );
buf ( n5295 , n5294 );
and ( n5296 , n5281 , n5295 );
and ( n5297 , n5263 , n5280 );
or ( n5298 , n5296 , n5297 );
buf ( n5299 , n5298 );
buf ( n5300 , n5299 );
and ( n5301 , n5246 , n5300 );
and ( n5302 , n5209 , n5245 );
or ( n5303 , n5301 , n5302 );
buf ( n5304 , n5303 );
buf ( n5305 , n5304 );
xor ( n5306 , n5067 , n5110 );
xor ( n5307 , n5306 , n5115 );
buf ( n5308 , n5307 );
buf ( n5309 , n5308 );
xor ( n5310 , n5305 , n5309 );
xor ( n5311 , n5030 , n5047 );
xor ( n5312 , n5311 , n5062 );
buf ( n5313 , n5312 );
buf ( n5314 , n5313 );
xor ( n5315 , n4980 , n4994 );
xor ( n5316 , n5315 , n5012 );
buf ( n5317 , n5316 );
buf ( n5318 , n5317 );
xor ( n5319 , n5314 , n5318 );
xor ( n5320 , n4929 , n4946 );
xor ( n5321 , n5320 , n4958 );
buf ( n5322 , n5321 );
buf ( n5323 , n5322 );
and ( n5324 , n5319 , n5323 );
and ( n5325 , n5314 , n5318 );
or ( n5326 , n5324 , n5325 );
buf ( n5327 , n5326 );
buf ( n5328 , n5327 );
and ( n5329 , n5310 , n5328 );
and ( n5330 , n5305 , n5309 );
or ( n5331 , n5329 , n5330 );
buf ( n5332 , n5331 );
buf ( n5333 , n5332 );
not ( n5334 , n831 );
not ( n5335 , n4967 );
or ( n5336 , n5334 , n5335 );
xor ( n5337 , n830 , n777 );
nand ( n5338 , n2207 , n5337 );
nand ( n5339 , n5336 , n5338 );
buf ( n5340 , n799 );
buf ( n5341 , n808 );
xor ( n5342 , n5340 , n5341 );
buf ( n5343 , n5342 );
buf ( n5344 , n5343 );
not ( n5345 , n5344 );
buf ( n5346 , n2235 );
not ( n5347 , n5346 );
or ( n5348 , n5345 , n5347 );
buf ( n5349 , n1309 );
buf ( n5350 , n5071 );
nand ( n5351 , n5349 , n5350 );
buf ( n5352 , n5351 );
buf ( n5353 , n5352 );
nand ( n5354 , n5348 , n5353 );
buf ( n5355 , n5354 );
xor ( n5356 , n5339 , n5355 );
buf ( n5357 , n781 );
buf ( n5358 , n826 );
xor ( n5359 , n5357 , n5358 );
buf ( n5360 , n5359 );
buf ( n5361 , n5360 );
not ( n5362 , n5361 );
buf ( n5363 , n4496 );
not ( n5364 , n5363 );
or ( n5365 , n5362 , n5364 );
buf ( n5366 , n1374 );
buf ( n5367 , n5102 );
nand ( n5368 , n5366 , n5367 );
buf ( n5369 , n5368 );
buf ( n5370 , n5369 );
nand ( n5371 , n5365 , n5370 );
buf ( n5372 , n5371 );
and ( n5373 , n5356 , n5372 );
and ( n5374 , n5339 , n5355 );
or ( n5375 , n5373 , n5374 );
buf ( n5376 , n793 );
buf ( n5377 , n814 );
xor ( n5378 , n5376 , n5377 );
buf ( n5379 , n5378 );
buf ( n5380 , n5379 );
not ( n5381 , n5380 );
buf ( n5382 , n3923 );
not ( n5383 , n5382 );
or ( n5384 , n5381 , n5383 );
buf ( n5385 , n1937 );
buf ( n5386 , n4916 );
nand ( n5387 , n5385 , n5386 );
buf ( n5388 , n5387 );
buf ( n5389 , n5388 );
nand ( n5390 , n5384 , n5389 );
buf ( n5391 , n5390 );
buf ( n5392 , n5391 );
xor ( n5393 , n824 , n783 );
buf ( n5394 , n5393 );
not ( n5395 , n5394 );
buf ( n5396 , n2790 );
not ( n5397 , n5396 );
or ( n5398 , n5395 , n5397 );
buf ( n5399 , n2492 );
buf ( n5400 , n5049 );
nand ( n5401 , n5399 , n5400 );
buf ( n5402 , n5401 );
buf ( n5403 , n5402 );
nand ( n5404 , n5398 , n5403 );
buf ( n5405 , n5404 );
buf ( n5406 , n5405 );
xor ( n5407 , n5392 , n5406 );
buf ( n5408 , n791 );
buf ( n5409 , n816 );
xor ( n5410 , n5408 , n5409 );
buf ( n5411 , n5410 );
buf ( n5412 , n5411 );
not ( n5413 , n5412 );
buf ( n5414 , n3719 );
not ( n5415 , n5414 );
or ( n5416 , n5413 , n5415 );
buf ( n5417 , n2010 );
buf ( n5418 , n4933 );
nand ( n5419 , n5417 , n5418 );
buf ( n5420 , n5419 );
buf ( n5421 , n5420 );
nand ( n5422 , n5416 , n5421 );
buf ( n5423 , n5422 );
buf ( n5424 , n5423 );
and ( n5425 , n5407 , n5424 );
and ( n5426 , n5392 , n5406 );
or ( n5427 , n5425 , n5426 );
buf ( n5428 , n5427 );
xor ( n5429 , n5375 , n5428 );
xor ( n5430 , n5084 , n5095 );
xor ( n5431 , n5430 , n5105 );
buf ( n5432 , n5431 );
and ( n5433 , n5429 , n5432 );
and ( n5434 , n5375 , n5428 );
or ( n5435 , n5433 , n5434 );
not ( n5436 , n5435 );
not ( n5437 , n4962 );
not ( n5438 , n5017 );
and ( n5439 , n5438 , n5016 );
not ( n5440 , n5438 );
not ( n5441 , n5016 );
and ( n5442 , n5440 , n5441 );
nor ( n5443 , n5439 , n5442 );
not ( n5444 , n5443 );
not ( n5445 , n5444 );
or ( n5446 , n5437 , n5445 );
nand ( n5447 , n4965 , n5443 );
nand ( n5448 , n5446 , n5447 );
not ( n5449 , n5448 );
not ( n5450 , n5449 );
or ( n5451 , n5436 , n5450 );
not ( n5452 , n5435 );
not ( n5453 , n5452 );
not ( n5454 , n5448 );
or ( n5455 , n5453 , n5454 );
xor ( n5456 , n4902 , n4905 );
xor ( n5457 , n5456 , n4908 );
nand ( n5458 , n5455 , n5457 );
nand ( n5459 , n5451 , n5458 );
buf ( n5460 , n5459 );
xor ( n5461 , n5333 , n5460 );
not ( n5462 , n5024 );
xor ( n5463 , n5119 , n5462 );
xnor ( n5464 , n5463 , n4911 );
buf ( n5465 , n5464 );
and ( n5466 , n5461 , n5465 );
and ( n5467 , n5333 , n5460 );
or ( n5468 , n5466 , n5467 );
buf ( n5469 , n5468 );
buf ( n5470 , n5469 );
xor ( n5471 , n5192 , n5470 );
not ( n5472 , n4895 );
not ( n5473 , n5472 );
not ( n5474 , n5126 );
or ( n5475 , n5473 , n5474 );
or ( n5476 , n4896 , n5126 );
nand ( n5477 , n5475 , n5476 );
and ( n5478 , n5477 , n4865 );
not ( n5479 , n5477 );
not ( n5480 , n4865 );
and ( n5481 , n5479 , n5480 );
nor ( n5482 , n5478 , n5481 );
buf ( n5483 , n5482 );
and ( n5484 , n5471 , n5483 );
and ( n5485 , n5192 , n5470 );
or ( n5486 , n5484 , n5485 );
buf ( n5487 , n5486 );
buf ( n5488 , n5487 );
xor ( n5489 , n5186 , n5488 );
xor ( n5490 , n4858 , n5130 );
xor ( n5491 , n5490 , n5135 );
buf ( n5492 , n5491 );
buf ( n5493 , n5492 );
and ( n5494 , n5489 , n5493 );
and ( n5495 , n5186 , n5488 );
or ( n5496 , n5494 , n5495 );
buf ( n5497 , n5496 );
buf ( n5498 , n5497 );
not ( n5499 , n5498 );
buf ( n5500 , n5499 );
buf ( n5501 , n5500 );
nand ( n5502 , n5185 , n5501 );
buf ( n5503 , n5502 );
buf ( n5504 , n5503 );
buf ( n5505 , n836 );
buf ( n5506 , n4887 );
buf ( n5507 , n4868 );
not ( n5508 , n5507 );
buf ( n5509 , n5508 );
buf ( n5510 , n5509 );
and ( n5511 , n5506 , n5510 );
not ( n5512 , n5506 );
buf ( n5513 , n4868 );
and ( n5514 , n5512 , n5513 );
nor ( n5515 , n5511 , n5514 );
buf ( n5516 , n5515 );
buf ( n5517 , n5516 );
buf ( n5518 , n4872 );
buf ( n5519 , n5518 );
buf ( n5520 , n5519 );
buf ( n5521 , n5520 );
not ( n5522 , n5521 );
buf ( n5523 , n5522 );
buf ( n5524 , n5523 );
and ( n5525 , n5517 , n5524 );
not ( n5526 , n5517 );
buf ( n5527 , n5520 );
and ( n5528 , n5526 , n5527 );
nor ( n5529 , n5525 , n5528 );
buf ( n5530 , n5529 );
buf ( n5531 , n5530 );
buf ( n5532 , n789 );
buf ( n5533 , n818 );
xor ( n5534 , n5532 , n5533 );
buf ( n5535 , n5534 );
buf ( n5536 , n5535 );
not ( n5537 , n5536 );
buf ( n5538 , n1480 );
not ( n5539 , n5538 );
or ( n5540 , n5537 , n5539 );
buf ( n5541 , n1496 );
buf ( n5542 , n5196 );
nand ( n5543 , n5541 , n5542 );
buf ( n5544 , n5543 );
buf ( n5545 , n5544 );
nand ( n5546 , n5540 , n5545 );
buf ( n5547 , n5546 );
buf ( n5548 , n5547 );
buf ( n5549 , n787 );
buf ( n5550 , n820 );
xor ( n5551 , n5549 , n5550 );
buf ( n5552 , n5551 );
buf ( n5553 , n5552 );
not ( n5554 , n5553 );
buf ( n5555 , n2267 );
not ( n5556 , n5555 );
or ( n5557 , n5554 , n5556 );
buf ( n5558 , n1346 );
buf ( n5559 , n5088 );
nand ( n5560 , n5558 , n5559 );
buf ( n5561 , n5560 );
buf ( n5562 , n5561 );
nand ( n5563 , n5557 , n5562 );
buf ( n5564 , n5563 );
buf ( n5565 , n5564 );
xor ( n5566 , n5548 , n5565 );
xor ( n5567 , n5225 , n5242 );
buf ( n5568 , n5567 );
buf ( n5569 , n5568 );
and ( n5570 , n5566 , n5569 );
and ( n5571 , n5548 , n5565 );
or ( n5572 , n5570 , n5571 );
buf ( n5573 , n5572 );
buf ( n5574 , n5573 );
xor ( n5575 , n824 , n784 );
buf ( n5576 , n5575 );
not ( n5577 , n5576 );
buf ( n5578 , n1965 );
not ( n5579 , n5578 );
or ( n5580 , n5577 , n5579 );
buf ( n5581 , n3255 );
buf ( n5582 , n5393 );
nand ( n5583 , n5581 , n5582 );
buf ( n5584 , n5583 );
buf ( n5585 , n5584 );
nand ( n5586 , n5580 , n5585 );
buf ( n5587 , n5586 );
buf ( n5588 , n5587 );
buf ( n5589 , n1309 );
not ( n5590 , n5589 );
buf ( n5591 , n1156 );
nor ( n5592 , n5590 , n5591 );
buf ( n5593 , n5592 );
buf ( n5594 , n5593 );
or ( n5595 , n5588 , n5594 );
not ( n5596 , n5229 );
not ( n5597 , n1249 );
or ( n5598 , n5596 , n5597 );
buf ( n5599 , n780 );
buf ( n5600 , n828 );
xor ( n5601 , n5599 , n5600 );
buf ( n5602 , n5601 );
nand ( n5603 , n5602 , n3842 );
nand ( n5604 , n5598 , n5603 );
buf ( n5605 , n5604 );
nand ( n5606 , n5595 , n5605 );
buf ( n5607 , n5606 );
buf ( n5608 , n5607 );
buf ( n5609 , n5587 );
buf ( n5610 , n1309 );
buf ( n5611 , n799 );
and ( n5612 , n5610 , n5611 );
buf ( n5613 , n5612 );
buf ( n5614 , n5613 );
nand ( n5615 , n5609 , n5614 );
buf ( n5616 , n5615 );
buf ( n5617 , n5616 );
nand ( n5618 , n5608 , n5617 );
buf ( n5619 , n5618 );
buf ( n5620 , n5619 );
not ( n5621 , n2207 );
buf ( n5622 , n778 );
buf ( n5623 , n830 );
xor ( n5624 , n5622 , n5623 );
buf ( n5625 , n5624 );
not ( n5626 , n5625 );
or ( n5627 , n5621 , n5626 );
nand ( n5628 , n5337 , n831 );
nand ( n5629 , n5627 , n5628 );
buf ( n5630 , n5629 );
buf ( n5631 , n796 );
buf ( n5632 , n812 );
xor ( n5633 , n5631 , n5632 );
buf ( n5634 , n5633 );
buf ( n5635 , n5634 );
not ( n5636 , n5635 );
buf ( n5637 , n1712 );
not ( n5638 , n5637 );
or ( n5639 , n5636 , n5638 );
buf ( n5640 , n1693 );
buf ( n5641 , n5250 );
nand ( n5642 , n5640 , n5641 );
buf ( n5643 , n5642 );
buf ( n5644 , n5643 );
nand ( n5645 , n5639 , n5644 );
buf ( n5646 , n5645 );
buf ( n5647 , n5646 );
xor ( n5648 , n5630 , n5647 );
xor ( n5649 , n810 , n798 );
buf ( n5650 , n5649 );
not ( n5651 , n5650 );
buf ( n5652 , n2641 );
not ( n5653 , n5652 );
or ( n5654 , n5651 , n5653 );
buf ( n5655 , n1679 );
buf ( n5656 , n5264 );
nand ( n5657 , n5655 , n5656 );
buf ( n5658 , n5657 );
buf ( n5659 , n5658 );
nand ( n5660 , n5654 , n5659 );
buf ( n5661 , n5660 );
buf ( n5662 , n5661 );
and ( n5663 , n5648 , n5662 );
and ( n5664 , n5630 , n5647 );
or ( n5665 , n5663 , n5664 );
buf ( n5666 , n5665 );
buf ( n5667 , n5666 );
xor ( n5668 , n5620 , n5667 );
buf ( n5669 , n782 );
buf ( n5670 , n826 );
xor ( n5671 , n5669 , n5670 );
buf ( n5672 , n5671 );
buf ( n5673 , n5672 );
not ( n5674 , n5673 );
buf ( n5675 , n2364 );
not ( n5676 , n5675 );
or ( n5677 , n5674 , n5676 );
buf ( n5678 , n1374 );
buf ( n5679 , n5360 );
nand ( n5680 , n5678 , n5679 );
buf ( n5681 , n5680 );
buf ( n5682 , n5681 );
nand ( n5683 , n5677 , n5682 );
buf ( n5684 , n5683 );
not ( n5685 , n5684 );
buf ( n5686 , n5685 );
not ( n5687 , n5686 );
buf ( n5688 , n788 );
buf ( n5689 , n820 );
xor ( n5690 , n5688 , n5689 );
buf ( n5691 , n5690 );
not ( n5692 , n5691 );
not ( n5693 , n1338 );
or ( n5694 , n5692 , n5693 );
buf ( n5695 , n5552 );
buf ( n5696 , n3986 );
nand ( n5697 , n5695 , n5696 );
buf ( n5698 , n5697 );
nand ( n5699 , n5694 , n5698 );
not ( n5700 , n5699 );
buf ( n5701 , n5700 );
not ( n5702 , n5701 );
or ( n5703 , n5687 , n5702 );
buf ( n5704 , n790 );
buf ( n5705 , n818 );
xor ( n5706 , n5704 , n5705 );
buf ( n5707 , n5706 );
buf ( n5708 , n5707 );
not ( n5709 , n5708 );
buf ( n5710 , n1480 );
not ( n5711 , n5710 );
or ( n5712 , n5709 , n5711 );
buf ( n5713 , n1496 );
buf ( n5714 , n5535 );
nand ( n5715 , n5713 , n5714 );
buf ( n5716 , n5715 );
buf ( n5717 , n5716 );
nand ( n5718 , n5712 , n5717 );
buf ( n5719 , n5718 );
buf ( n5720 , n5719 );
nand ( n5721 , n5703 , n5720 );
buf ( n5722 , n5721 );
buf ( n5723 , n5722 );
buf ( n5724 , n5699 );
buf ( n5725 , n5684 );
nand ( n5726 , n5724 , n5725 );
buf ( n5727 , n5726 );
buf ( n5728 , n5727 );
nand ( n5729 , n5723 , n5728 );
buf ( n5730 , n5729 );
buf ( n5731 , n5730 );
and ( n5732 , n5668 , n5731 );
and ( n5733 , n5620 , n5667 );
or ( n5734 , n5732 , n5733 );
buf ( n5735 , n5734 );
buf ( n5736 , n5735 );
xor ( n5737 , n5574 , n5736 );
xor ( n5738 , n5209 , n5245 );
xor ( n5739 , n5738 , n5300 );
buf ( n5740 , n5739 );
buf ( n5741 , n5740 );
and ( n5742 , n5737 , n5741 );
and ( n5743 , n5574 , n5736 );
or ( n5744 , n5742 , n5743 );
buf ( n5745 , n5744 );
buf ( n5746 , n5745 );
xor ( n5747 , n5305 , n5309 );
xor ( n5748 , n5747 , n5328 );
buf ( n5749 , n5748 );
buf ( n5750 , n5749 );
xor ( n5751 , n5746 , n5750 );
xor ( n5752 , n5314 , n5318 );
xor ( n5753 , n5752 , n5323 );
buf ( n5754 , n5753 );
not ( n5755 , n5754 );
not ( n5756 , n5755 );
not ( n5757 , n5756 );
xor ( n5758 , n5339 , n5355 );
xor ( n5759 , n5758 , n5372 );
buf ( n5760 , n5759 );
buf ( n5761 , n792 );
buf ( n5762 , n816 );
xor ( n5763 , n5761 , n5762 );
buf ( n5764 , n5763 );
buf ( n5765 , n5764 );
not ( n5766 , n5765 );
buf ( n5767 , n2004 );
not ( n5768 , n5767 );
or ( n5769 , n5766 , n5768 );
buf ( n5770 , n2535 );
buf ( n5771 , n5411 );
nand ( n5772 , n5770 , n5771 );
buf ( n5773 , n5772 );
buf ( n5774 , n5773 );
nand ( n5775 , n5769 , n5774 );
buf ( n5776 , n5775 );
buf ( n5777 , n5776 );
not ( n5778 , n5777 );
buf ( n5779 , n5778 );
buf ( n5780 , n5779 );
buf ( n5781 , n5780 );
buf ( n5782 , n5781 );
buf ( n5783 , n5782 );
buf ( n5784 , n794 );
buf ( n5785 , n814 );
xor ( n5786 , n5784 , n5785 );
buf ( n5787 , n5786 );
buf ( n5788 , n5787 );
not ( n5789 , n5788 );
buf ( n5790 , n1931 );
not ( n5791 , n5790 );
or ( n5792 , n5789 , n5791 );
buf ( n5793 , n1937 );
buf ( n5794 , n5379 );
nand ( n5795 , n5793 , n5794 );
buf ( n5796 , n5795 );
buf ( n5797 , n5796 );
nand ( n5798 , n5792 , n5797 );
buf ( n5799 , n5798 );
buf ( n5800 , n5799 );
xor ( n5801 , n822 , n786 );
buf ( n5802 , n5801 );
not ( n5803 , n5802 );
buf ( n5804 , n2098 );
not ( n5805 , n5804 );
or ( n5806 , n5803 , n5805 );
buf ( n5807 , n2113 );
buf ( n5808 , n5282 );
nand ( n5809 , n5807 , n5808 );
buf ( n5810 , n5809 );
buf ( n5811 , n5810 );
nand ( n5812 , n5806 , n5811 );
buf ( n5813 , n5812 );
buf ( n5814 , n5813 );
nor ( n5815 , n5800 , n5814 );
buf ( n5816 , n5815 );
buf ( n5817 , n5816 );
or ( n5818 , n5783 , n5817 );
buf ( n5819 , n5799 );
buf ( n5820 , n5813 );
nand ( n5821 , n5819 , n5820 );
buf ( n5822 , n5821 );
buf ( n5823 , n5822 );
nand ( n5824 , n5818 , n5823 );
buf ( n5825 , n5824 );
buf ( n5826 , n5825 );
xor ( n5827 , n5760 , n5826 );
xor ( n5828 , n5263 , n5280 );
xor ( n5829 , n5828 , n5295 );
buf ( n5830 , n5829 );
buf ( n5831 , n5830 );
and ( n5832 , n5827 , n5831 );
and ( n5833 , n5760 , n5826 );
or ( n5834 , n5832 , n5833 );
buf ( n5835 , n5834 );
not ( n5836 , n5835 );
or ( n5837 , n5757 , n5836 );
not ( n5838 , n5835 );
not ( n5839 , n5838 );
not ( n5840 , n5755 );
or ( n5841 , n5839 , n5840 );
xor ( n5842 , n5375 , n5428 );
xor ( n5843 , n5842 , n5432 );
nand ( n5844 , n5841 , n5843 );
nand ( n5845 , n5837 , n5844 );
buf ( n5846 , n5845 );
and ( n5847 , n5751 , n5846 );
and ( n5848 , n5746 , n5750 );
or ( n5849 , n5847 , n5848 );
buf ( n5850 , n5849 );
buf ( n5851 , n5850 );
xor ( n5852 , n5531 , n5851 );
xor ( n5853 , n5333 , n5460 );
xor ( n5854 , n5853 , n5465 );
buf ( n5855 , n5854 );
buf ( n5856 , n5855 );
and ( n5857 , n5852 , n5856 );
and ( n5858 , n5531 , n5851 );
or ( n5859 , n5857 , n5858 );
buf ( n5860 , n5859 );
buf ( n5861 , n5860 );
xor ( n5862 , n5505 , n5861 );
xor ( n5863 , n5192 , n5470 );
xor ( n5864 , n5863 , n5483 );
buf ( n5865 , n5864 );
buf ( n5866 , n5865 );
and ( n5867 , n5862 , n5866 );
and ( n5868 , n5505 , n5861 );
or ( n5869 , n5867 , n5868 );
buf ( n5870 , n5869 );
not ( n5871 , n5870 );
xor ( n5872 , n5186 , n5488 );
xor ( n5873 , n5872 , n5493 );
buf ( n5874 , n5873 );
buf ( n5875 , n5874 );
not ( n5876 , n5875 );
buf ( n5877 , n5876 );
nand ( n5878 , n5871 , n5877 );
buf ( n5879 , n5878 );
nand ( n5880 , n5504 , n5879 );
buf ( n5881 , n5880 );
buf ( n5882 , n5881 );
not ( n5883 , n5882 );
buf ( n5884 , n5883 );
buf ( n5885 , n5884 );
nand ( n5886 , n5178 , n5885 );
buf ( n5887 , n5886 );
buf ( n5888 , n5887 );
not ( n5889 , n5888 );
buf ( n5890 , n837 );
buf ( n5891 , n5457 );
not ( n5892 , n5891 );
buf ( n5893 , n5892 );
not ( n5894 , n5452 );
not ( n5895 , n5449 );
or ( n5896 , n5894 , n5895 );
nand ( n5897 , n5448 , n5435 );
nand ( n5898 , n5896 , n5897 );
or ( n5899 , n5893 , n5898 );
nand ( n5900 , n5898 , n5893 );
nand ( n5901 , n5899 , n5900 );
buf ( n5902 , n5901 );
xor ( n5903 , n5392 , n5406 );
xor ( n5904 , n5903 , n5424 );
buf ( n5905 , n5904 );
buf ( n5906 , n5905 );
xor ( n5907 , n5548 , n5565 );
xor ( n5908 , n5907 , n5569 );
buf ( n5909 , n5908 );
buf ( n5910 , n5909 );
xor ( n5911 , n5906 , n5910 );
buf ( n5912 , n799 );
buf ( n5913 , n811 );
or ( n5914 , n5912 , n5913 );
buf ( n5915 , n812 );
nand ( n5916 , n5914 , n5915 );
buf ( n5917 , n5916 );
buf ( n5918 , n5917 );
buf ( n5919 , n799 );
buf ( n5920 , n811 );
nand ( n5921 , n5919 , n5920 );
buf ( n5922 , n5921 );
buf ( n5923 , n5922 );
buf ( n5924 , n810 );
and ( n5925 , n5918 , n5923 , n5924 );
buf ( n5926 , n5925 );
buf ( n5927 , n5926 );
xor ( n5928 , n828 , n781 );
buf ( n5929 , n5928 );
not ( n5930 , n5929 );
buf ( n5931 , n1239 );
not ( n5932 , n5931 );
or ( n5933 , n5930 , n5932 );
buf ( n5934 , n1249 );
buf ( n5935 , n5602 );
nand ( n5936 , n5934 , n5935 );
buf ( n5937 , n5936 );
buf ( n5938 , n5937 );
nand ( n5939 , n5933 , n5938 );
buf ( n5940 , n5939 );
buf ( n5941 , n5940 );
and ( n5942 , n5927 , n5941 );
buf ( n5943 , n5942 );
xor ( n5944 , n822 , n787 );
buf ( n5945 , n5944 );
not ( n5946 , n5945 );
buf ( n5947 , n2098 );
not ( n5948 , n5947 );
or ( n5949 , n5946 , n5948 );
buf ( n5950 , n2107 );
buf ( n5951 , n5801 );
nand ( n5952 , n5950 , n5951 );
buf ( n5953 , n5952 );
buf ( n5954 , n5953 );
nand ( n5955 , n5949 , n5954 );
buf ( n5956 , n5955 );
xor ( n5957 , n812 , n797 );
buf ( n5958 , n5957 );
not ( n5959 , n5958 );
buf ( n5960 , n1712 );
not ( n5961 , n5960 );
or ( n5962 , n5959 , n5961 );
buf ( n5963 , n1693 );
buf ( n5964 , n5634 );
nand ( n5965 , n5963 , n5964 );
buf ( n5966 , n5965 );
buf ( n5967 , n5966 );
nand ( n5968 , n5962 , n5967 );
buf ( n5969 , n5968 );
or ( n5970 , n5956 , n5969 );
not ( n5971 , n5970 );
buf ( n5972 , n810 );
not ( n5973 , n5972 );
buf ( n5974 , n799 );
nand ( n5975 , n5973 , n5974 );
buf ( n5976 , n5975 );
buf ( n5977 , n5976 );
not ( n5978 , n5977 );
buf ( n5979 , n799 );
not ( n5980 , n5979 );
buf ( n5981 , n810 );
nand ( n5982 , n5980 , n5981 );
buf ( n5983 , n5982 );
buf ( n5984 , n5983 );
not ( n5985 , n5984 );
or ( n5986 , n5978 , n5985 );
buf ( n5987 , n2641 );
nand ( n5988 , n5986 , n5987 );
buf ( n5989 , n5988 );
buf ( n5990 , n5989 );
buf ( n5991 , n5272 );
buf ( n5992 , n5649 );
nand ( n5993 , n5991 , n5992 );
buf ( n5994 , n5993 );
buf ( n5995 , n5994 );
nand ( n5996 , n5990 , n5995 );
buf ( n5997 , n5996 );
not ( n5998 , n5997 );
or ( n5999 , n5971 , n5998 );
nand ( n6000 , n5969 , n5956 );
nand ( n6001 , n5999 , n6000 );
nand ( n6002 , n5943 , n6001 );
buf ( n6003 , n779 );
buf ( n6004 , n830 );
xor ( n6005 , n6003 , n6004 );
buf ( n6006 , n6005 );
buf ( n6007 , n6006 );
not ( n6008 , n6007 );
buf ( n6009 , n1161 );
not ( n6010 , n6009 );
or ( n6011 , n6008 , n6010 );
buf ( n6012 , n5625 );
buf ( n6013 , n831 );
nand ( n6014 , n6012 , n6013 );
buf ( n6015 , n6014 );
buf ( n6016 , n6015 );
nand ( n6017 , n6011 , n6016 );
buf ( n6018 , n6017 );
buf ( n6019 , n6018 );
buf ( n6020 , n783 );
buf ( n6021 , n826 );
xor ( n6022 , n6020 , n6021 );
buf ( n6023 , n6022 );
buf ( n6024 , n6023 );
not ( n6025 , n6024 );
buf ( n6026 , n4496 );
not ( n6027 , n6026 );
or ( n6028 , n6025 , n6027 );
buf ( n6029 , n1374 );
buf ( n6030 , n5672 );
nand ( n6031 , n6029 , n6030 );
buf ( n6032 , n6031 );
buf ( n6033 , n6032 );
nand ( n6034 , n6028 , n6033 );
buf ( n6035 , n6034 );
buf ( n6036 , n6035 );
xor ( n6037 , n6019 , n6036 );
not ( n6038 , n1346 );
not ( n6039 , n5691 );
or ( n6040 , n6038 , n6039 );
buf ( n6041 , n789 );
buf ( n6042 , n820 );
xor ( n6043 , n6041 , n6042 );
buf ( n6044 , n6043 );
buf ( n6045 , n6044 );
not ( n6046 , n6045 );
buf ( n6047 , n6046 );
or ( n6048 , n2678 , n6047 );
nand ( n6049 , n6040 , n6048 );
buf ( n6050 , n6049 );
and ( n6051 , n6037 , n6050 );
and ( n6052 , n6019 , n6036 );
or ( n6053 , n6051 , n6052 );
buf ( n6054 , n6053 );
nand ( n6055 , n5943 , n6054 );
nand ( n6056 , n6001 , n6054 );
nand ( n6057 , n6002 , n6055 , n6056 );
buf ( n6058 , n6057 );
and ( n6059 , n5911 , n6058 );
and ( n6060 , n5906 , n5910 );
or ( n6061 , n6059 , n6060 );
buf ( n6062 , n6061 );
buf ( n6063 , n6062 );
xor ( n6064 , n5574 , n5736 );
xor ( n6065 , n6064 , n5741 );
buf ( n6066 , n6065 );
buf ( n6067 , n6066 );
xor ( n6068 , n6063 , n6067 );
xor ( n6069 , n5620 , n5667 );
xor ( n6070 , n6069 , n5731 );
buf ( n6071 , n6070 );
buf ( n6072 , n6071 );
buf ( n6073 , n5799 );
buf ( n6074 , n5779 );
and ( n6075 , n6073 , n6074 );
not ( n6076 , n6073 );
buf ( n6077 , n5776 );
and ( n6078 , n6076 , n6077 );
nor ( n6079 , n6075 , n6078 );
buf ( n6080 , n6079 );
not ( n6081 , n6080 );
and ( n6082 , n6081 , n5813 );
not ( n6083 , n6081 );
not ( n6084 , n5813 );
and ( n6085 , n6083 , n6084 );
nor ( n6086 , n6082 , n6085 );
not ( n6087 , n6086 );
buf ( n6088 , n5787 );
not ( n6089 , n6088 );
buf ( n6090 , n1940 );
not ( n6091 , n6090 );
or ( n6092 , n6089 , n6091 );
buf ( n6093 , n3703 );
xor ( n6094 , n814 , n795 );
buf ( n6095 , n6094 );
nand ( n6096 , n6093 , n6095 );
buf ( n6097 , n6096 );
buf ( n6098 , n6097 );
nand ( n6099 , n6092 , n6098 );
buf ( n6100 , n6099 );
not ( n6101 , n6100 );
xor ( n6102 , n824 , n785 );
buf ( n6103 , n6102 );
not ( n6104 , n6103 );
buf ( n6105 , n2483 );
not ( n6106 , n6105 );
or ( n6107 , n6104 , n6106 );
buf ( n6108 , n1859 );
buf ( n6109 , n5575 );
nand ( n6110 , n6108 , n6109 );
buf ( n6111 , n6110 );
buf ( n6112 , n6111 );
nand ( n6113 , n6107 , n6112 );
buf ( n6114 , n6113 );
not ( n6115 , n6114 );
buf ( n6116 , n793 );
buf ( n6117 , n816 );
xor ( n6118 , n6116 , n6117 );
buf ( n6119 , n6118 );
buf ( n6120 , n6119 );
not ( n6121 , n6120 );
xnor ( n6122 , n817 , n816 );
nor ( n6123 , n6122 , n2000 );
buf ( n6124 , n6123 );
not ( n6125 , n6124 );
or ( n6126 , n6121 , n6125 );
buf ( n6127 , n2532 );
buf ( n6128 , n5764 );
nand ( n6129 , n6127 , n6128 );
buf ( n6130 , n6129 );
buf ( n6131 , n6130 );
nand ( n6132 , n6126 , n6131 );
buf ( n6133 , n6132 );
not ( n6134 , n6133 );
nand ( n6135 , n6115 , n6134 );
not ( n6136 , n6135 );
or ( n6137 , n6101 , n6136 );
not ( n6138 , n6134 );
nand ( n6139 , n6138 , n6114 );
nand ( n6140 , n6137 , n6139 );
not ( n6141 , n6140 );
or ( n6142 , n6087 , n6141 );
not ( n6143 , n6140 );
not ( n6144 , n6143 );
not ( n6145 , n6084 );
not ( n6146 , n6080 );
or ( n6147 , n6145 , n6146 );
not ( n6148 , n6081 );
or ( n6149 , n6084 , n6148 );
nand ( n6150 , n6147 , n6149 );
not ( n6151 , n6150 );
or ( n6152 , n6144 , n6151 );
and ( n6153 , n5700 , n5685 );
not ( n6154 , n5700 );
and ( n6155 , n6154 , n5684 );
nor ( n6156 , n6153 , n6155 );
not ( n6157 , n5719 );
xor ( n6158 , n6156 , n6157 );
buf ( n6159 , n6158 );
not ( n6160 , n6159 );
buf ( n6161 , n6160 );
nand ( n6162 , n6152 , n6161 );
nand ( n6163 , n6142 , n6162 );
buf ( n6164 , n6163 );
xor ( n6165 , n6072 , n6164 );
xor ( n6166 , n5760 , n5826 );
xor ( n6167 , n6166 , n5831 );
buf ( n6168 , n6167 );
buf ( n6169 , n6168 );
and ( n6170 , n6165 , n6169 );
and ( n6171 , n6072 , n6164 );
or ( n6172 , n6170 , n6171 );
buf ( n6173 , n6172 );
buf ( n6174 , n6173 );
and ( n6175 , n6068 , n6174 );
and ( n6176 , n6063 , n6067 );
or ( n6177 , n6175 , n6176 );
buf ( n6178 , n6177 );
buf ( n6179 , n6178 );
xor ( n6180 , n5902 , n6179 );
xor ( n6181 , n5746 , n5750 );
xor ( n6182 , n6181 , n5846 );
buf ( n6183 , n6182 );
buf ( n6184 , n6183 );
and ( n6185 , n6180 , n6184 );
and ( n6186 , n5902 , n6179 );
or ( n6187 , n6185 , n6186 );
buf ( n6188 , n6187 );
buf ( n6189 , n6188 );
xor ( n6190 , n5890 , n6189 );
xor ( n6191 , n5531 , n5851 );
xor ( n6192 , n6191 , n5856 );
buf ( n6193 , n6192 );
buf ( n6194 , n6193 );
xor ( n6195 , n6190 , n6194 );
buf ( n6196 , n6195 );
buf ( n6197 , n6196 );
buf ( n6198 , n838 );
xor ( n6199 , n5843 , n5835 );
xor ( n6200 , n6199 , n5756 );
buf ( n6201 , n6200 );
xor ( n6202 , n5604 , n5613 );
xor ( n6203 , n6202 , n5587 );
buf ( n6204 , n6203 );
xor ( n6205 , n5630 , n5647 );
xor ( n6206 , n6205 , n5662 );
buf ( n6207 , n6206 );
buf ( n6208 , n6207 );
xor ( n6209 , n6204 , n6208 );
buf ( n6210 , n791 );
buf ( n6211 , n818 );
xor ( n6212 , n6210 , n6211 );
buf ( n6213 , n6212 );
buf ( n6214 , n6213 );
not ( n6215 , n6214 );
buf ( n6216 , n1480 );
not ( n6217 , n6216 );
or ( n6218 , n6215 , n6217 );
buf ( n6219 , n1496 );
buf ( n6220 , n5707 );
nand ( n6221 , n6219 , n6220 );
buf ( n6222 , n6221 );
buf ( n6223 , n6222 );
nand ( n6224 , n6218 , n6223 );
buf ( n6225 , n6224 );
buf ( n6226 , n6225 );
xor ( n6227 , n5927 , n5941 );
buf ( n6228 , n6227 );
buf ( n6229 , n6228 );
xor ( n6230 , n6226 , n6229 );
xor ( n6231 , n794 , n816 );
not ( n6232 , n6231 );
not ( n6233 , n6123 );
or ( n6234 , n6232 , n6233 );
buf ( n6235 , n2532 );
buf ( n6236 , n6119 );
nand ( n6237 , n6235 , n6236 );
buf ( n6238 , n6237 );
nand ( n6239 , n6234 , n6238 );
buf ( n6240 , n6239 );
buf ( n6241 , n796 );
buf ( n6242 , n814 );
xor ( n6243 , n6241 , n6242 );
buf ( n6244 , n6243 );
buf ( n6245 , n6244 );
not ( n6246 , n6245 );
buf ( n6247 , n3923 );
not ( n6248 , n6247 );
or ( n6249 , n6246 , n6248 );
buf ( n6250 , n1937 );
buf ( n6251 , n6094 );
nand ( n6252 , n6250 , n6251 );
buf ( n6253 , n6252 );
buf ( n6254 , n6253 );
nand ( n6255 , n6249 , n6254 );
buf ( n6256 , n6255 );
buf ( n6257 , n6256 );
xor ( n6258 , n6240 , n6257 );
buf ( n6259 , n782 );
buf ( n6260 , n828 );
xor ( n6261 , n6259 , n6260 );
buf ( n6262 , n6261 );
buf ( n6263 , n6262 );
not ( n6264 , n6263 );
buf ( n6265 , n1901 );
not ( n6266 , n6265 );
or ( n6267 , n6264 , n6266 );
buf ( n6268 , n1249 );
buf ( n6269 , n5928 );
nand ( n6270 , n6268 , n6269 );
buf ( n6271 , n6270 );
buf ( n6272 , n6271 );
nand ( n6273 , n6267 , n6272 );
buf ( n6274 , n6273 );
buf ( n6275 , n6274 );
and ( n6276 , n6258 , n6275 );
and ( n6277 , n6240 , n6257 );
or ( n6278 , n6276 , n6277 );
buf ( n6279 , n6278 );
buf ( n6280 , n6279 );
and ( n6281 , n6230 , n6280 );
and ( n6282 , n6226 , n6229 );
or ( n6283 , n6281 , n6282 );
buf ( n6284 , n6283 );
buf ( n6285 , n6284 );
and ( n6286 , n6209 , n6285 );
and ( n6287 , n6204 , n6208 );
or ( n6288 , n6286 , n6287 );
buf ( n6289 , n6288 );
buf ( n6290 , n6289 );
xor ( n6291 , n5906 , n5910 );
xor ( n6292 , n6291 , n6058 );
buf ( n6293 , n6292 );
buf ( n6294 , n6293 );
xor ( n6295 , n6290 , n6294 );
xor ( n6296 , n6072 , n6164 );
xor ( n6297 , n6296 , n6169 );
buf ( n6298 , n6297 );
buf ( n6299 , n6298 );
and ( n6300 , n6295 , n6299 );
and ( n6301 , n6290 , n6294 );
or ( n6302 , n6300 , n6301 );
buf ( n6303 , n6302 );
buf ( n6304 , n6303 );
xor ( n6305 , n6201 , n6304 );
xor ( n6306 , n6063 , n6067 );
xor ( n6307 , n6306 , n6174 );
buf ( n6308 , n6307 );
buf ( n6309 , n6308 );
and ( n6310 , n6305 , n6309 );
and ( n6311 , n6201 , n6304 );
or ( n6312 , n6310 , n6311 );
buf ( n6313 , n6312 );
buf ( n6314 , n6313 );
xor ( n6315 , n6198 , n6314 );
xor ( n6316 , n5902 , n6179 );
xor ( n6317 , n6316 , n6184 );
buf ( n6318 , n6317 );
buf ( n6319 , n6318 );
and ( n6320 , n6315 , n6319 );
and ( n6321 , n6198 , n6314 );
or ( n6322 , n6320 , n6321 );
buf ( n6323 , n6322 );
buf ( n6324 , n6323 );
nand ( n6325 , n6197 , n6324 );
buf ( n6326 , n6325 );
buf ( n6327 , n6326 );
not ( n6328 , n6327 );
buf ( n6329 , n6328 );
not ( n6330 , n6329 );
xor ( n6331 , n5505 , n5861 );
xor ( n6332 , n6331 , n5866 );
buf ( n6333 , n6332 );
xor ( n6334 , n5890 , n6189 );
and ( n6335 , n6334 , n6194 );
and ( n6336 , n5890 , n6189 );
or ( n6337 , n6335 , n6336 );
buf ( n6338 , n6337 );
nor ( n6339 , n6333 , n6338 );
not ( n6340 , n6339 );
not ( n6341 , n6340 );
or ( n6342 , n6330 , n6341 );
buf ( n6343 , n6333 );
buf ( n6344 , n6343 );
buf ( n6345 , n6344 );
buf ( n6346 , n6345 );
buf ( n6347 , n6338 );
buf ( n6348 , n6347 );
buf ( n6349 , n6348 );
buf ( n6350 , n6349 );
nand ( n6351 , n6346 , n6350 );
buf ( n6352 , n6351 );
nand ( n6353 , n6342 , n6352 );
not ( n6354 , n6353 );
xor ( n6355 , n6198 , n6314 );
xor ( n6356 , n6355 , n6319 );
buf ( n6357 , n6356 );
buf ( n6358 , n6357 );
buf ( n6359 , n839 );
xor ( n6360 , n5943 , n6001 );
xor ( n6361 , n6360 , n6054 );
buf ( n6362 , n6361 );
buf ( n6363 , n1679 );
buf ( n6364 , n799 );
nand ( n6365 , n6363 , n6364 );
buf ( n6366 , n6365 );
buf ( n6367 , n6366 );
not ( n6368 , n6367 );
not ( n6369 , n831 );
not ( n6370 , n6006 );
or ( n6371 , n6369 , n6370 );
nand ( n6372 , n1159 , n830 );
not ( n6373 , n6372 );
and ( n6374 , n830 , n780 );
not ( n6375 , n830 );
and ( n6376 , n6375 , n1321 );
nor ( n6377 , n6374 , n6376 );
nand ( n6378 , n6373 , n6377 );
nand ( n6379 , n6371 , n6378 );
buf ( n6380 , n6379 );
not ( n6381 , n6380 );
buf ( n6382 , n6381 );
buf ( n6383 , n6382 );
not ( n6384 , n6383 );
or ( n6385 , n6368 , n6384 );
buf ( n6386 , n786 );
buf ( n6387 , n824 );
xor ( n6388 , n6386 , n6387 );
buf ( n6389 , n6388 );
buf ( n6390 , n6389 );
not ( n6391 , n6390 );
buf ( n6392 , n1965 );
not ( n6393 , n6392 );
or ( n6394 , n6391 , n6393 );
buf ( n6395 , n3255 );
buf ( n6396 , n6102 );
nand ( n6397 , n6395 , n6396 );
buf ( n6398 , n6397 );
buf ( n6399 , n6398 );
nand ( n6400 , n6394 , n6399 );
buf ( n6401 , n6400 );
buf ( n6402 , n6401 );
nand ( n6403 , n6385 , n6402 );
buf ( n6404 , n6403 );
buf ( n6405 , n6404 );
buf ( n6406 , n6366 );
not ( n6407 , n6406 );
buf ( n6408 , n6379 );
nand ( n6409 , n6407 , n6408 );
buf ( n6410 , n6409 );
buf ( n6411 , n6410 );
nand ( n6412 , n6405 , n6411 );
buf ( n6413 , n6412 );
buf ( n6414 , n6413 );
xor ( n6415 , n6019 , n6036 );
xor ( n6416 , n6415 , n6050 );
buf ( n6417 , n6416 );
buf ( n6418 , n6417 );
xor ( n6419 , n6414 , n6418 );
buf ( n6420 , n788 );
buf ( n6421 , n822 );
xor ( n6422 , n6420 , n6421 );
buf ( n6423 , n6422 );
buf ( n6424 , n6423 );
not ( n6425 , n6424 );
buf ( n6426 , n2098 );
not ( n6427 , n6426 );
or ( n6428 , n6425 , n6427 );
buf ( n6429 , n2107 );
buf ( n6430 , n5944 );
nand ( n6431 , n6429 , n6430 );
buf ( n6432 , n6431 );
buf ( n6433 , n6432 );
nand ( n6434 , n6428 , n6433 );
buf ( n6435 , n6434 );
buf ( n6436 , n6435 );
buf ( n6437 , n798 );
buf ( n6438 , n812 );
xor ( n6439 , n6437 , n6438 );
buf ( n6440 , n6439 );
buf ( n6441 , n6440 );
not ( n6442 , n6441 );
buf ( n6443 , n2916 );
not ( n6444 , n6443 );
or ( n6445 , n6442 , n6444 );
buf ( n6446 , n1693 );
buf ( n6447 , n6446 );
buf ( n6448 , n5957 );
nand ( n6449 , n6447 , n6448 );
buf ( n6450 , n6449 );
buf ( n6451 , n6450 );
nand ( n6452 , n6445 , n6451 );
buf ( n6453 , n6452 );
buf ( n6454 , n6453 );
xor ( n6455 , n6436 , n6454 );
buf ( n6456 , n6023 );
not ( n6457 , n6456 );
buf ( n6458 , n1771 );
not ( n6459 , n6458 );
or ( n6460 , n6457 , n6459 );
buf ( n6461 , n4496 );
not ( n6462 , n6461 );
buf ( n6463 , n6462 );
buf ( n6464 , n6463 );
xor ( n6465 , n826 , n784 );
buf ( n6466 , n6465 );
not ( n6467 , n6466 );
buf ( n6468 , n6467 );
buf ( n6469 , n6468 );
or ( n6470 , n6464 , n6469 );
nand ( n6471 , n6460 , n6470 );
buf ( n6472 , n6471 );
buf ( n6473 , n6472 );
and ( n6474 , n6455 , n6473 );
and ( n6475 , n6436 , n6454 );
or ( n6476 , n6474 , n6475 );
buf ( n6477 , n6476 );
buf ( n6478 , n6477 );
and ( n6479 , n6419 , n6478 );
and ( n6480 , n6414 , n6418 );
or ( n6481 , n6479 , n6480 );
buf ( n6482 , n6481 );
buf ( n6483 , n6482 );
xor ( n6484 , n6362 , n6483 );
xor ( n6485 , n6134 , n6114 );
xor ( n6486 , n6485 , n6100 );
not ( n6487 , n6486 );
not ( n6488 , n6487 );
buf ( n6489 , n5956 );
xor ( n6490 , n5969 , n6489 );
xnor ( n6491 , n6490 , n5997 );
not ( n6492 , n6491 );
not ( n6493 , n6492 );
or ( n6494 , n6488 , n6493 );
not ( n6495 , n6491 );
not ( n6496 , n6486 );
or ( n6497 , n6495 , n6496 );
xor ( n6498 , n820 , n790 );
buf ( n6499 , n6498 );
not ( n6500 , n6499 );
buf ( n6501 , n2410 );
not ( n6502 , n6501 );
or ( n6503 , n6500 , n6502 );
buf ( n6504 , n1346 );
buf ( n6505 , n6044 );
nand ( n6506 , n6504 , n6505 );
buf ( n6507 , n6506 );
buf ( n6508 , n6507 );
nand ( n6509 , n6503 , n6508 );
buf ( n6510 , n6509 );
not ( n6511 , n6510 );
buf ( n6512 , n792 );
buf ( n6513 , n818 );
xor ( n6514 , n6512 , n6513 );
buf ( n6515 , n6514 );
buf ( n6516 , n6515 );
not ( n6517 , n6516 );
buf ( n6518 , n1480 );
not ( n6519 , n6518 );
or ( n6520 , n6517 , n6519 );
buf ( n6521 , n1496 );
buf ( n6522 , n6213 );
nand ( n6523 , n6521 , n6522 );
buf ( n6524 , n6523 );
buf ( n6525 , n6524 );
nand ( n6526 , n6520 , n6525 );
buf ( n6527 , n6526 );
not ( n6528 , n6527 );
or ( n6529 , n6511 , n6528 );
or ( n6530 , n6527 , n6510 );
buf ( n6531 , n799 );
buf ( n6532 , n813 );
or ( n6533 , n6531 , n6532 );
buf ( n6534 , n814 );
nand ( n6535 , n6533 , n6534 );
buf ( n6536 , n6535 );
buf ( n6537 , n799 );
buf ( n6538 , n813 );
nand ( n6539 , n6537 , n6538 );
buf ( n6540 , n6539 );
and ( n6541 , n6536 , n6540 , n812 );
not ( n6542 , n1630 );
buf ( n6543 , n781 );
buf ( n6544 , n830 );
xor ( n6545 , n6543 , n6544 );
buf ( n6546 , n6545 );
not ( n6547 , n6546 );
or ( n6548 , n6542 , n6547 );
buf ( n6549 , n6377 );
buf ( n6550 , n831 );
nand ( n6551 , n6549 , n6550 );
buf ( n6552 , n6551 );
nand ( n6553 , n6548 , n6552 );
and ( n6554 , n6541 , n6553 );
nand ( n6555 , n6530 , n6554 );
nand ( n6556 , n6529 , n6555 );
nand ( n6557 , n6497 , n6556 );
nand ( n6558 , n6494 , n6557 );
buf ( n6559 , n6558 );
and ( n6560 , n6484 , n6559 );
and ( n6561 , n6362 , n6483 );
or ( n6562 , n6560 , n6561 );
buf ( n6563 , n6562 );
buf ( n6564 , n6563 );
and ( n6565 , n6158 , n6143 );
not ( n6566 , n6158 );
and ( n6567 , n6566 , n6140 );
nor ( n6568 , n6565 , n6567 );
buf ( n6569 , n6568 );
buf ( n6570 , n6086 );
and ( n6571 , n6569 , n6570 );
not ( n6572 , n6569 );
buf ( n6573 , n6150 );
buf ( n6574 , n6573 );
and ( n6575 , n6572 , n6574 );
nor ( n6576 , n6571 , n6575 );
buf ( n6577 , n6576 );
buf ( n6578 , n6577 );
xor ( n6579 , n6204 , n6208 );
xor ( n6580 , n6579 , n6285 );
buf ( n6581 , n6580 );
buf ( n6582 , n6581 );
xor ( n6583 , n6578 , n6582 );
xor ( n6584 , n6226 , n6229 );
xor ( n6585 , n6584 , n6280 );
buf ( n6586 , n6585 );
buf ( n6587 , n6586 );
buf ( n6588 , n787 );
buf ( n6589 , n824 );
xor ( n6590 , n6588 , n6589 );
buf ( n6591 , n6590 );
not ( n6592 , n6591 );
not ( n6593 , n1838 );
or ( n6594 , n6592 , n6593 );
not ( n6595 , n3252 );
nand ( n6596 , n6595 , n6389 );
nand ( n6597 , n6594 , n6596 );
buf ( n6598 , n6597 );
not ( n6599 , n6598 );
xor ( n6600 , n814 , n797 );
buf ( n6601 , n6600 );
not ( n6602 , n6601 );
buf ( n6603 , n1931 );
not ( n6604 , n6603 );
or ( n6605 , n6602 , n6604 );
buf ( n6606 , n1937 );
buf ( n6607 , n6244 );
nand ( n6608 , n6606 , n6607 );
buf ( n6609 , n6608 );
buf ( n6610 , n6609 );
nand ( n6611 , n6605 , n6610 );
buf ( n6612 , n6611 );
buf ( n6613 , n6612 );
not ( n6614 , n6613 );
or ( n6615 , n6599 , n6614 );
buf ( n6616 , n6597 );
buf ( n6617 , n6612 );
or ( n6618 , n6616 , n6617 );
xor ( n6619 , n795 , n816 );
not ( n6620 , n6619 );
not ( n6621 , n6123 );
or ( n6622 , n6620 , n6621 );
nand ( n6623 , n2532 , n6231 );
nand ( n6624 , n6622 , n6623 );
buf ( n6625 , n6624 );
nand ( n6626 , n6618 , n6625 );
buf ( n6627 , n6626 );
buf ( n6628 , n6627 );
nand ( n6629 , n6615 , n6628 );
buf ( n6630 , n6629 );
buf ( n6631 , n6630 );
buf ( n6632 , n789 );
buf ( n6633 , n822 );
xor ( n6634 , n6632 , n6633 );
buf ( n6635 , n6634 );
buf ( n6636 , n6635 );
not ( n6637 , n6636 );
buf ( n6638 , n2098 );
not ( n6639 , n6638 );
or ( n6640 , n6637 , n6639 );
buf ( n6641 , n2107 );
buf ( n6642 , n6423 );
nand ( n6643 , n6641 , n6642 );
buf ( n6644 , n6643 );
buf ( n6645 , n6644 );
nand ( n6646 , n6640 , n6645 );
buf ( n6647 , n6646 );
not ( n6648 , n6647 );
buf ( n6649 , n783 );
buf ( n6650 , n828 );
xor ( n6651 , n6649 , n6650 );
buf ( n6652 , n6651 );
buf ( n6653 , n6652 );
not ( n6654 , n6653 );
buf ( n6655 , n1239 );
not ( n6656 , n6655 );
or ( n6657 , n6654 , n6656 );
buf ( n6658 , n1249 );
buf ( n6659 , n6262 );
nand ( n6660 , n6658 , n6659 );
buf ( n6661 , n6660 );
buf ( n6662 , n6661 );
nand ( n6663 , n6657 , n6662 );
buf ( n6664 , n6663 );
not ( n6665 , n6664 );
or ( n6666 , n6648 , n6665 );
buf ( n6667 , n6664 );
buf ( n6668 , n6647 );
nor ( n6669 , n6667 , n6668 );
buf ( n6670 , n6669 );
buf ( n6671 , n799 );
buf ( n6672 , n812 );
xor ( n6673 , n6671 , n6672 );
buf ( n6674 , n6673 );
buf ( n6675 , n6674 );
not ( n6676 , n6675 );
buf ( n6677 , n2916 );
not ( n6678 , n6677 );
or ( n6679 , n6676 , n6678 );
buf ( n6680 , n1693 );
buf ( n6681 , n6440 );
nand ( n6682 , n6680 , n6681 );
buf ( n6683 , n6682 );
buf ( n6684 , n6683 );
nand ( n6685 , n6679 , n6684 );
buf ( n6686 , n6685 );
buf ( n6687 , n6686 );
not ( n6688 , n6687 );
buf ( n6689 , n6688 );
or ( n6690 , n6670 , n6689 );
nand ( n6691 , n6666 , n6690 );
buf ( n6692 , n6691 );
xor ( n6693 , n6631 , n6692 );
xor ( n6694 , n820 , n791 );
not ( n6695 , n6694 );
not ( n6696 , n2410 );
or ( n6697 , n6695 , n6696 );
buf ( n6698 , n2672 );
buf ( n6699 , n6498 );
nand ( n6700 , n6698 , n6699 );
buf ( n6701 , n6700 );
nand ( n6702 , n6697 , n6701 );
not ( n6703 , n6702 );
xor ( n6704 , n818 , n793 );
not ( n6705 , n6704 );
not ( n6706 , n1480 );
or ( n6707 , n6705 , n6706 );
buf ( n6708 , n1496 );
buf ( n6709 , n6515 );
nand ( n6710 , n6708 , n6709 );
buf ( n6711 , n6710 );
nand ( n6712 , n6707 , n6711 );
not ( n6713 , n6712 );
or ( n6714 , n6703 , n6713 );
nor ( n6715 , n6702 , n6712 );
xor ( n6716 , n826 , n785 );
not ( n6717 , n6716 );
not ( n6718 , n2364 );
or ( n6719 , n6717 , n6718 );
buf ( n6720 , n1771 );
buf ( n6721 , n6465 );
nand ( n6722 , n6720 , n6721 );
buf ( n6723 , n6722 );
nand ( n6724 , n6719 , n6723 );
not ( n6725 , n6724 );
or ( n6726 , n6715 , n6725 );
nand ( n6727 , n6714 , n6726 );
buf ( n6728 , n6727 );
and ( n6729 , n6693 , n6728 );
and ( n6730 , n6631 , n6692 );
or ( n6731 , n6729 , n6730 );
buf ( n6732 , n6731 );
buf ( n6733 , n6732 );
xor ( n6734 , n6587 , n6733 );
xor ( n6735 , n6414 , n6418 );
xor ( n6736 , n6735 , n6478 );
buf ( n6737 , n6736 );
buf ( n6738 , n6737 );
and ( n6739 , n6734 , n6738 );
and ( n6740 , n6587 , n6733 );
or ( n6741 , n6739 , n6740 );
buf ( n6742 , n6741 );
buf ( n6743 , n6742 );
and ( n6744 , n6583 , n6743 );
and ( n6745 , n6578 , n6582 );
or ( n6746 , n6744 , n6745 );
buf ( n6747 , n6746 );
buf ( n6748 , n6747 );
xor ( n6749 , n6564 , n6748 );
xor ( n6750 , n6290 , n6294 );
xor ( n6751 , n6750 , n6299 );
buf ( n6752 , n6751 );
buf ( n6753 , n6752 );
and ( n6754 , n6749 , n6753 );
and ( n6755 , n6564 , n6748 );
or ( n6756 , n6754 , n6755 );
buf ( n6757 , n6756 );
buf ( n6758 , n6757 );
xor ( n6759 , n6359 , n6758 );
xor ( n6760 , n6201 , n6304 );
xor ( n6761 , n6760 , n6309 );
buf ( n6762 , n6761 );
buf ( n6763 , n6762 );
and ( n6764 , n6759 , n6763 );
and ( n6765 , n6359 , n6758 );
or ( n6766 , n6764 , n6765 );
buf ( n6767 , n6766 );
buf ( n6768 , n6767 );
nor ( n6769 , n6358 , n6768 );
buf ( n6770 , n6769 );
buf ( n6771 , n6770 );
xor ( n6772 , n6359 , n6758 );
xor ( n6773 , n6772 , n6763 );
buf ( n6774 , n6773 );
buf ( n6775 , n6774 );
buf ( n6776 , n840 );
xor ( n6777 , n6362 , n6483 );
xor ( n6778 , n6777 , n6559 );
buf ( n6779 , n6778 );
buf ( n6780 , n6779 );
xor ( n6781 , n6578 , n6582 );
xor ( n6782 , n6781 , n6743 );
buf ( n6783 , n6782 );
buf ( n6784 , n6783 );
xor ( n6785 , n6780 , n6784 );
buf ( n6786 , n6401 );
not ( n6787 , n6786 );
buf ( n6788 , n6379 );
not ( n6789 , n6788 );
buf ( n6790 , n6366 );
not ( n6791 , n6790 );
and ( n6792 , n6789 , n6791 );
buf ( n6793 , n6379 );
buf ( n6794 , n6366 );
and ( n6795 , n6793 , n6794 );
nor ( n6796 , n6792 , n6795 );
buf ( n6797 , n6796 );
buf ( n6798 , n6797 );
not ( n6799 , n6798 );
or ( n6800 , n6787 , n6799 );
buf ( n6801 , n6797 );
buf ( n6802 , n6401 );
or ( n6803 , n6801 , n6802 );
nand ( n6804 , n6800 , n6803 );
buf ( n6805 , n6804 );
buf ( n6806 , n6805 );
xor ( n6807 , n6240 , n6257 );
xor ( n6808 , n6807 , n6275 );
buf ( n6809 , n6808 );
buf ( n6810 , n6809 );
xor ( n6811 , n6806 , n6810 );
xor ( n6812 , n6436 , n6454 );
xor ( n6813 , n6812 , n6473 );
buf ( n6814 , n6813 );
buf ( n6815 , n6814 );
and ( n6816 , n6811 , n6815 );
and ( n6817 , n6806 , n6810 );
or ( n6818 , n6816 , n6817 );
buf ( n6819 , n6818 );
buf ( n6820 , n6819 );
nand ( n6821 , n6487 , n6556 , n6492 );
not ( n6822 , n6556 );
nand ( n6823 , n6486 , n6822 , n6492 );
nand ( n6824 , n6487 , n6822 , n6491 );
nand ( n6825 , n6491 , n6556 , n6486 );
nand ( n6826 , n6821 , n6823 , n6824 , n6825 );
buf ( n6827 , n6826 );
xor ( n6828 , n6820 , n6827 );
xor ( n6829 , n6587 , n6733 );
xor ( n6830 , n6829 , n6738 );
buf ( n6831 , n6830 );
buf ( n6832 , n6831 );
and ( n6833 , n6828 , n6832 );
and ( n6834 , n6820 , n6827 );
or ( n6835 , n6833 , n6834 );
buf ( n6836 , n6835 );
buf ( n6837 , n6836 );
and ( n6838 , n6785 , n6837 );
and ( n6839 , n6780 , n6784 );
or ( n6840 , n6838 , n6839 );
buf ( n6841 , n6840 );
buf ( n6842 , n6841 );
xor ( n6843 , n6776 , n6842 );
xor ( n6844 , n6564 , n6748 );
xor ( n6845 , n6844 , n6753 );
buf ( n6846 , n6845 );
buf ( n6847 , n6846 );
and ( n6848 , n6843 , n6847 );
and ( n6849 , n6776 , n6842 );
or ( n6850 , n6848 , n6849 );
buf ( n6851 , n6850 );
buf ( n6852 , n6851 );
nor ( n6853 , n6775 , n6852 );
buf ( n6854 , n6853 );
buf ( n6855 , n6854 );
nor ( n6856 , n6771 , n6855 );
buf ( n6857 , n6856 );
buf ( n6858 , n6857 );
buf ( n6859 , n6858 );
buf ( n6860 , n6859 );
buf ( n6861 , n6860 );
not ( n6862 , n6861 );
buf ( n6863 , n6862 );
buf ( n6864 , n6774 );
buf ( n6865 , n6851 );
nand ( n6866 , n6864 , n6865 );
buf ( n6867 , n6866 );
buf ( n6868 , n6867 );
not ( n6869 , n6868 );
buf ( n6870 , n6869 );
not ( n6871 , n6870 );
buf ( n6872 , n6770 );
not ( n6873 , n6872 );
buf ( n6874 , n6873 );
not ( n6875 , n6874 );
or ( n6876 , n6871 , n6875 );
buf ( n6877 , n6357 );
buf ( n6878 , n6877 );
buf ( n6879 , n6878 );
buf ( n6880 , n6879 );
buf ( n6881 , n6767 );
nand ( n6882 , n6880 , n6881 );
buf ( n6883 , n6882 );
nand ( n6884 , n6876 , n6883 );
not ( n6885 , n6884 );
nand ( n6886 , n6354 , n6863 , n6885 );
buf ( n6887 , n6886 );
xor ( n6888 , n6776 , n6842 );
xor ( n6889 , n6888 , n6847 );
buf ( n6890 , n6889 );
buf ( n6891 , n6890 );
buf ( n6892 , n841 );
xor ( n6893 , n6527 , n6510 );
xor ( n6894 , n6893 , n6554 );
buf ( n6895 , n788 );
buf ( n6896 , n824 );
xor ( n6897 , n6895 , n6896 );
buf ( n6898 , n6897 );
not ( n6899 , n6898 );
not ( n6900 , n2790 );
or ( n6901 , n6899 , n6900 );
buf ( n6902 , n3255 );
buf ( n6903 , n6591 );
nand ( n6904 , n6902 , n6903 );
buf ( n6905 , n6904 );
nand ( n6906 , n6901 , n6905 );
not ( n6907 , n6906 );
buf ( n6908 , n1693 );
buf ( n6909 , n799 );
and ( n6910 , n6908 , n6909 );
buf ( n6911 , n6910 );
not ( n6912 , n6911 );
buf ( n6913 , n782 );
buf ( n6914 , n830 );
xor ( n6915 , n6913 , n6914 );
buf ( n6916 , n6915 );
buf ( n6917 , n6916 );
not ( n6918 , n6917 );
buf ( n6919 , n1161 );
not ( n6920 , n6919 );
or ( n6921 , n6918 , n6920 );
buf ( n6922 , n6546 );
buf ( n6923 , n831 );
nand ( n6924 , n6922 , n6923 );
buf ( n6925 , n6924 );
buf ( n6926 , n6925 );
nand ( n6927 , n6921 , n6926 );
buf ( n6928 , n6927 );
not ( n6929 , n6928 );
nand ( n6930 , n6912 , n6929 );
not ( n6931 , n6930 );
or ( n6932 , n6907 , n6931 );
nand ( n6933 , n6928 , n6911 );
nand ( n6934 , n6932 , n6933 );
not ( n6935 , n6934 );
xor ( n6936 , n6541 , n6553 );
not ( n6937 , n6936 );
nand ( n6938 , n6935 , n6937 );
not ( n6939 , n6938 );
buf ( n6940 , n796 );
buf ( n6941 , n816 );
xor ( n6942 , n6940 , n6941 );
buf ( n6943 , n6942 );
buf ( n6944 , n6943 );
not ( n6945 , n6944 );
buf ( n6946 , n2526 );
not ( n6947 , n6946 );
or ( n6948 , n6945 , n6947 );
nand ( n6949 , n6619 , n2010 );
buf ( n6950 , n6949 );
nand ( n6951 , n6948 , n6950 );
buf ( n6952 , n6951 );
buf ( n6953 , n6952 );
not ( n6954 , n6953 );
buf ( n6955 , n6954 );
buf ( n6956 , n6955 );
not ( n6957 , n6956 );
buf ( n6958 , n798 );
buf ( n6959 , n814 );
xor ( n6960 , n6958 , n6959 );
buf ( n6961 , n6960 );
buf ( n6962 , n6961 );
not ( n6963 , n6962 );
buf ( n6964 , n3703 );
not ( n6965 , n6964 );
or ( n6966 , n6963 , n6965 );
buf ( n6967 , n1940 );
buf ( n6968 , n6600 );
nand ( n6969 , n6967 , n6968 );
buf ( n6970 , n6969 );
buf ( n6971 , n6970 );
nand ( n6972 , n6966 , n6971 );
buf ( n6973 , n6972 );
buf ( n6974 , n6973 );
not ( n6975 , n6974 );
buf ( n6976 , n6975 );
buf ( n6977 , n6976 );
not ( n6978 , n6977 );
or ( n6979 , n6957 , n6978 );
buf ( n6980 , n784 );
buf ( n6981 , n828 );
xor ( n6982 , n6980 , n6981 );
buf ( n6983 , n6982 );
buf ( n6984 , n6983 );
not ( n6985 , n6984 );
buf ( n6986 , n3680 );
not ( n6987 , n6986 );
or ( n6988 , n6985 , n6987 );
buf ( n6989 , n1249 );
buf ( n6990 , n6652 );
nand ( n6991 , n6989 , n6990 );
buf ( n6992 , n6991 );
buf ( n6993 , n6992 );
nand ( n6994 , n6988 , n6993 );
buf ( n6995 , n6994 );
buf ( n6996 , n6995 );
nand ( n6997 , n6979 , n6996 );
buf ( n6998 , n6997 );
buf ( n6999 , n6961 );
not ( n7000 , n6999 );
buf ( n7001 , n3703 );
not ( n7002 , n7001 );
or ( n7003 , n7000 , n7002 );
buf ( n7004 , n6970 );
nand ( n7005 , n7003 , n7004 );
buf ( n7006 , n7005 );
buf ( n7007 , n7006 );
buf ( n7008 , n6952 );
nand ( n7009 , n7007 , n7008 );
buf ( n7010 , n7009 );
nand ( n7011 , n6998 , n7010 );
not ( n7012 , n7011 );
or ( n7013 , n6939 , n7012 );
nand ( n7014 , n6936 , n6934 );
nand ( n7015 , n7013 , n7014 );
xor ( n7016 , n6894 , n7015 );
buf ( n7017 , n6597 );
not ( n7018 , n7017 );
buf ( n7019 , n6624 );
not ( n7020 , n7019 );
buf ( n7021 , n7020 );
buf ( n7022 , n7021 );
not ( n7023 , n7022 );
or ( n7024 , n7018 , n7023 );
buf ( n7025 , n7021 );
buf ( n7026 , n6597 );
or ( n7027 , n7025 , n7026 );
nand ( n7028 , n7024 , n7027 );
buf ( n7029 , n7028 );
buf ( n7030 , n7029 );
buf ( n7031 , n6612 );
and ( n7032 , n7030 , n7031 );
not ( n7033 , n7030 );
buf ( n7034 , n6612 );
not ( n7035 , n7034 );
buf ( n7036 , n7035 );
buf ( n7037 , n7036 );
and ( n7038 , n7033 , n7037 );
nor ( n7039 , n7032 , n7038 );
buf ( n7040 , n7039 );
buf ( n7041 , n7040 );
buf ( n7042 , n790 );
buf ( n7043 , n822 );
xor ( n7044 , n7042 , n7043 );
buf ( n7045 , n7044 );
buf ( n7046 , n7045 );
not ( n7047 , n7046 );
buf ( n7048 , n2098 );
not ( n7049 , n7048 );
or ( n7050 , n7047 , n7049 );
buf ( n7051 , n2107 );
buf ( n7052 , n6635 );
nand ( n7053 , n7051 , n7052 );
buf ( n7054 , n7053 );
buf ( n7055 , n7054 );
nand ( n7056 , n7050 , n7055 );
buf ( n7057 , n7056 );
buf ( n7058 , n7057 );
xor ( n7059 , n820 , n792 );
not ( n7060 , n7059 );
not ( n7061 , n2410 );
or ( n7062 , n7060 , n7061 );
nand ( n7063 , n6694 , n1345 );
nand ( n7064 , n7062 , n7063 );
buf ( n7065 , n7064 );
xor ( n7066 , n7058 , n7065 );
buf ( n7067 , n6716 );
not ( n7068 , n7067 );
buf ( n7069 , n1771 );
not ( n7070 , n7069 );
or ( n7071 , n7068 , n7070 );
buf ( n7072 , n1783 );
buf ( n7073 , n786 );
buf ( n7074 , n826 );
xor ( n7075 , n7073 , n7074 );
buf ( n7076 , n7075 );
buf ( n7077 , n7076 );
not ( n7078 , n7077 );
buf ( n7079 , n7078 );
buf ( n7080 , n7079 );
or ( n7081 , n7072 , n7080 );
nand ( n7082 , n7071 , n7081 );
buf ( n7083 , n7082 );
buf ( n7084 , n7083 );
and ( n7085 , n7066 , n7084 );
and ( n7086 , n7058 , n7065 );
or ( n7087 , n7085 , n7086 );
buf ( n7088 , n7087 );
buf ( n7089 , n7088 );
xor ( n7090 , n7041 , n7089 );
xor ( n7091 , n6724 , n6712 );
xor ( n7092 , n7091 , n6702 );
buf ( n7093 , n7092 );
and ( n7094 , n7090 , n7093 );
and ( n7095 , n7041 , n7089 );
or ( n7096 , n7094 , n7095 );
buf ( n7097 , n7096 );
and ( n7098 , n7016 , n7097 );
and ( n7099 , n6894 , n7015 );
or ( n7100 , n7098 , n7099 );
buf ( n7101 , n7100 );
xor ( n7102 , n6631 , n6692 );
xor ( n7103 , n7102 , n6728 );
buf ( n7104 , n7103 );
not ( n7105 , n7104 );
xor ( n7106 , n6806 , n6810 );
xor ( n7107 , n7106 , n6815 );
buf ( n7108 , n7107 );
not ( n7109 , n7108 );
nand ( n7110 , n7105 , n7109 );
not ( n7111 , n7110 );
xor ( n7112 , n6894 , n7015 );
xor ( n7113 , n7112 , n7097 );
not ( n7114 , n7113 );
or ( n7115 , n7111 , n7114 );
not ( n7116 , n7109 );
nand ( n7117 , n7116 , n7104 );
nand ( n7118 , n7115 , n7117 );
buf ( n7119 , n7118 );
xor ( n7120 , n7101 , n7119 );
xor ( n7121 , n6820 , n6827 );
xor ( n7122 , n7121 , n6832 );
buf ( n7123 , n7122 );
buf ( n7124 , n7123 );
and ( n7125 , n7120 , n7124 );
and ( n7126 , n7101 , n7119 );
or ( n7127 , n7125 , n7126 );
buf ( n7128 , n7127 );
buf ( n7129 , n7128 );
xor ( n7130 , n6892 , n7129 );
xor ( n7131 , n6780 , n6784 );
xor ( n7132 , n7131 , n6837 );
buf ( n7133 , n7132 );
buf ( n7134 , n7133 );
and ( n7135 , n7130 , n7134 );
and ( n7136 , n6892 , n7129 );
or ( n7137 , n7135 , n7136 );
buf ( n7138 , n7137 );
buf ( n7139 , n7138 );
nor ( n7140 , n6891 , n7139 );
buf ( n7141 , n7140 );
xor ( n7142 , n6892 , n7129 );
xor ( n7143 , n7142 , n7134 );
buf ( n7144 , n7143 );
buf ( n7145 , n7144 );
buf ( n7146 , n842 );
xor ( n7147 , n6686 , n6664 );
xor ( n7148 , n7147 , n6647 );
buf ( n7149 , n7148 );
xor ( n7150 , n6937 , n6934 );
xnor ( n7151 , n7150 , n7011 );
buf ( n7152 , n7151 );
xor ( n7153 , n7149 , n7152 );
buf ( n7154 , n6704 );
not ( n7155 , n7154 );
buf ( n7156 , n1496 );
not ( n7157 , n7156 );
or ( n7158 , n7155 , n7157 );
buf ( n7159 , n1480 );
buf ( n7160 , n794 );
buf ( n7161 , n818 );
xor ( n7162 , n7160 , n7161 );
buf ( n7163 , n7162 );
buf ( n7164 , n7163 );
nand ( n7165 , n7159 , n7164 );
buf ( n7166 , n7165 );
buf ( n7167 , n7166 );
nand ( n7168 , n7158 , n7167 );
buf ( n7169 , n7168 );
not ( n7170 , n7169 );
buf ( n7171 , n783 );
buf ( n7172 , n830 );
xor ( n7173 , n7171 , n7172 );
buf ( n7174 , n7173 );
buf ( n7175 , n7174 );
not ( n7176 , n7175 );
buf ( n7177 , n1630 );
not ( n7178 , n7177 );
or ( n7179 , n7176 , n7178 );
buf ( n7180 , n6916 );
buf ( n7181 , n831 );
nand ( n7182 , n7180 , n7181 );
buf ( n7183 , n7182 );
buf ( n7184 , n7183 );
nand ( n7185 , n7179 , n7184 );
buf ( n7186 , n7185 );
buf ( n7187 , n799 );
buf ( n7188 , n815 );
or ( n7189 , n7187 , n7188 );
buf ( n7190 , n816 );
nand ( n7191 , n7189 , n7190 );
buf ( n7192 , n7191 );
buf ( n7193 , n7192 );
buf ( n7194 , n799 );
buf ( n7195 , n815 );
nand ( n7196 , n7194 , n7195 );
buf ( n7197 , n7196 );
buf ( n7198 , n7197 );
buf ( n7199 , n814 );
nand ( n7200 , n7193 , n7198 , n7199 );
buf ( n7201 , n7200 );
not ( n7202 , n7201 );
and ( n7203 , n7186 , n7202 );
not ( n7204 , n7203 );
nand ( n7205 , n7170 , n7204 );
buf ( n7206 , n7205 );
not ( n7207 , n7206 );
buf ( n7208 , n3255 );
buf ( n7209 , n6898 );
nand ( n7210 , n7208 , n7209 );
buf ( n7211 , n7210 );
buf ( n7212 , n789 );
buf ( n7213 , n824 );
xor ( n7214 , n7212 , n7213 );
buf ( n7215 , n7214 );
nand ( n7216 , n2790 , n7215 );
and ( n7217 , n7211 , n7216 );
not ( n7218 , n7217 );
buf ( n7219 , n799 );
buf ( n7220 , n814 );
xor ( n7221 , n7219 , n7220 );
buf ( n7222 , n7221 );
not ( n7223 , n7222 );
not ( n7224 , n2612 );
or ( n7225 , n7223 , n7224 );
buf ( n7226 , n1940 );
buf ( n7227 , n6961 );
nand ( n7228 , n7226 , n7227 );
buf ( n7229 , n7228 );
nand ( n7230 , n7225 , n7229 );
or ( n7231 , n7218 , n7230 );
buf ( n7232 , n797 );
buf ( n7233 , n816 );
xor ( n7234 , n7232 , n7233 );
buf ( n7235 , n7234 );
not ( n7236 , n7235 );
not ( n7237 , n2526 );
or ( n7238 , n7236 , n7237 );
buf ( n7239 , n2010 );
buf ( n7240 , n6943 );
nand ( n7241 , n7239 , n7240 );
buf ( n7242 , n7241 );
nand ( n7243 , n7238 , n7242 );
nand ( n7244 , n7231 , n7243 );
nand ( n7245 , n7218 , n7230 );
nand ( n7246 , n7244 , n7245 );
buf ( n7247 , n7246 );
not ( n7248 , n7247 );
or ( n7249 , n7207 , n7248 );
nand ( n7250 , n7169 , n7203 );
buf ( n7251 , n7250 );
nand ( n7252 , n7249 , n7251 );
buf ( n7253 , n7252 );
buf ( n7254 , n7253 );
and ( n7255 , n7153 , n7254 );
and ( n7256 , n7149 , n7152 );
or ( n7257 , n7255 , n7256 );
buf ( n7258 , n7257 );
xor ( n7259 , n7041 , n7089 );
xor ( n7260 , n7259 , n7093 );
buf ( n7261 , n7260 );
xor ( n7262 , n6911 , n6929 );
xnor ( n7263 , n7262 , n6906 );
buf ( n7264 , n791 );
buf ( n7265 , n822 );
xor ( n7266 , n7264 , n7265 );
buf ( n7267 , n7266 );
buf ( n7268 , n7267 );
not ( n7269 , n7268 );
buf ( n7270 , n2101 );
not ( n7271 , n7270 );
or ( n7272 , n7269 , n7271 );
buf ( n7273 , n2107 );
buf ( n7274 , n7045 );
nand ( n7275 , n7273 , n7274 );
buf ( n7276 , n7275 );
buf ( n7277 , n7276 );
nand ( n7278 , n7272 , n7277 );
buf ( n7279 , n7278 );
not ( n7280 , n7279 );
not ( n7281 , n1353 );
not ( n7282 , n1351 );
or ( n7283 , n7281 , n7282 );
nand ( n7284 , n7283 , n1355 );
buf ( n7285 , n7284 );
not ( n7286 , n7285 );
buf ( n7287 , n787 );
buf ( n7288 , n826 );
xnor ( n7289 , n7287 , n7288 );
buf ( n7290 , n7289 );
buf ( n7291 , n7290 );
not ( n7292 , n7291 );
and ( n7293 , n7286 , n7292 );
buf ( n7294 , n1771 );
buf ( n7295 , n7076 );
and ( n7296 , n7294 , n7295 );
nor ( n7297 , n7293 , n7296 );
buf ( n7298 , n7297 );
not ( n7299 , n7298 );
not ( n7300 , n7299 );
or ( n7301 , n7280 , n7300 );
not ( n7302 , n7298 );
buf ( n7303 , n7267 );
not ( n7304 , n7303 );
buf ( n7305 , n2101 );
not ( n7306 , n7305 );
or ( n7307 , n7304 , n7306 );
buf ( n7308 , n7276 );
nand ( n7309 , n7307 , n7308 );
buf ( n7310 , n7309 );
buf ( n7311 , n7310 );
not ( n7312 , n7311 );
buf ( n7313 , n7312 );
not ( n7314 , n7313 );
or ( n7315 , n7302 , n7314 );
buf ( n7316 , n785 );
buf ( n7317 , n828 );
xor ( n7318 , n7316 , n7317 );
buf ( n7319 , n7318 );
buf ( n7320 , n7319 );
not ( n7321 , n7320 );
buf ( n7322 , n3680 );
not ( n7323 , n7322 );
or ( n7324 , n7321 , n7323 );
buf ( n7325 , n1249 );
buf ( n7326 , n6983 );
nand ( n7327 , n7325 , n7326 );
buf ( n7328 , n7327 );
buf ( n7329 , n7328 );
nand ( n7330 , n7324 , n7329 );
buf ( n7331 , n7330 );
nand ( n7332 , n7315 , n7331 );
nand ( n7333 , n7301 , n7332 );
xor ( n7334 , n7263 , n7333 );
xor ( n7335 , n7058 , n7065 );
xor ( n7336 , n7335 , n7084 );
buf ( n7337 , n7336 );
and ( n7338 , n7334 , n7337 );
and ( n7339 , n7263 , n7333 );
or ( n7340 , n7338 , n7339 );
xor ( n7341 , n7261 , n7340 );
buf ( n7342 , n6976 );
not ( n7343 , n7342 );
buf ( n7344 , n6952 );
not ( n7345 , n7344 );
and ( n7346 , n7343 , n7345 );
buf ( n7347 , n6952 );
buf ( n7348 , n6976 );
and ( n7349 , n7347 , n7348 );
nor ( n7350 , n7346 , n7349 );
buf ( n7351 , n7350 );
buf ( n7352 , n7351 );
buf ( n7353 , n6995 );
not ( n7354 , n7353 );
buf ( n7355 , n7354 );
buf ( n7356 , n7355 );
and ( n7357 , n7352 , n7356 );
not ( n7358 , n7352 );
buf ( n7359 , n6995 );
and ( n7360 , n7358 , n7359 );
nor ( n7361 , n7357 , n7360 );
buf ( n7362 , n7361 );
not ( n7363 , n7362 );
xor ( n7364 , n820 , n793 );
buf ( n7365 , n7364 );
not ( n7366 , n7365 );
buf ( n7367 , n2410 );
not ( n7368 , n7367 );
or ( n7369 , n7366 , n7368 );
buf ( n7370 , n2672 );
buf ( n7371 , n7059 );
nand ( n7372 , n7370 , n7371 );
buf ( n7373 , n7372 );
buf ( n7374 , n7373 );
nand ( n7375 , n7369 , n7374 );
buf ( n7376 , n7375 );
buf ( n7377 , n7376 );
not ( n7378 , n7377 );
buf ( n7379 , n7201 );
not ( n7380 , n7379 );
buf ( n7381 , n7186 );
not ( n7382 , n7381 );
or ( n7383 , n7380 , n7382 );
buf ( n7384 , n7186 );
buf ( n7385 , n7201 );
or ( n7386 , n7384 , n7385 );
nand ( n7387 , n7383 , n7386 );
buf ( n7388 , n7387 );
buf ( n7389 , n7388 );
not ( n7390 , n7389 );
or ( n7391 , n7378 , n7390 );
buf ( n7392 , n7388 );
buf ( n7393 , n7376 );
or ( n7394 , n7392 , n7393 );
buf ( n7395 , n795 );
buf ( n7396 , n818 );
xor ( n7397 , n7395 , n7396 );
buf ( n7398 , n7397 );
buf ( n7399 , n7398 );
not ( n7400 , n7399 );
buf ( n7401 , n1480 );
not ( n7402 , n7401 );
or ( n7403 , n7400 , n7402 );
buf ( n7404 , n1496 );
buf ( n7405 , n7163 );
nand ( n7406 , n7404 , n7405 );
buf ( n7407 , n7406 );
buf ( n7408 , n7407 );
nand ( n7409 , n7403 , n7408 );
buf ( n7410 , n7409 );
buf ( n7411 , n7410 );
nand ( n7412 , n7394 , n7411 );
buf ( n7413 , n7412 );
buf ( n7414 , n7413 );
nand ( n7415 , n7391 , n7414 );
buf ( n7416 , n7415 );
not ( n7417 , n7416 );
or ( n7418 , n7363 , n7417 );
buf ( n7419 , n7362 );
buf ( n7420 , n7416 );
nor ( n7421 , n7419 , n7420 );
buf ( n7422 , n7421 );
and ( n7423 , n7204 , n7169 );
not ( n7424 , n7204 );
and ( n7425 , n7424 , n7170 );
nor ( n7426 , n7423 , n7425 );
xor ( n7427 , n7246 , n7426 );
or ( n7428 , n7422 , n7427 );
nand ( n7429 , n7418 , n7428 );
and ( n7430 , n7341 , n7429 );
and ( n7431 , n7261 , n7340 );
or ( n7432 , n7430 , n7431 );
xor ( n7433 , n7258 , n7432 );
not ( n7434 , n7108 );
and ( n7435 , n7104 , n7434 );
not ( n7436 , n7104 );
and ( n7437 , n7436 , n7108 );
nor ( n7438 , n7435 , n7437 );
not ( n7439 , n7113 );
and ( n7440 , n7438 , n7439 );
not ( n7441 , n7438 );
and ( n7442 , n7441 , n7113 );
nor ( n7443 , n7440 , n7442 );
and ( n7444 , n7433 , n7443 );
and ( n7445 , n7258 , n7432 );
or ( n7446 , n7444 , n7445 );
buf ( n7447 , n7446 );
xor ( n7448 , n7146 , n7447 );
xor ( n7449 , n7101 , n7119 );
xor ( n7450 , n7449 , n7124 );
buf ( n7451 , n7450 );
buf ( n7452 , n7451 );
and ( n7453 , n7448 , n7452 );
and ( n7454 , n7146 , n7447 );
or ( n7455 , n7453 , n7454 );
buf ( n7456 , n7455 );
buf ( n7457 , n7456 );
nor ( n7458 , n7145 , n7457 );
buf ( n7459 , n7458 );
nor ( n7460 , n7141 , n7459 );
xor ( n7461 , n7146 , n7447 );
xor ( n7462 , n7461 , n7452 );
buf ( n7463 , n7462 );
buf ( n7464 , n7463 );
buf ( n7465 , n843 );
xor ( n7466 , n7149 , n7152 );
xor ( n7467 , n7466 , n7254 );
buf ( n7468 , n7467 );
buf ( n7469 , n1937 );
buf ( n7470 , n799 );
nand ( n7471 , n7469 , n7470 );
buf ( n7472 , n7471 );
buf ( n7473 , n7472 );
not ( n7474 , n7473 );
not ( n7475 , n831 );
not ( n7476 , n7174 );
or ( n7477 , n7475 , n7476 );
not ( n7478 , n1629 );
buf ( n7479 , n784 );
buf ( n7480 , n830 );
xor ( n7481 , n7479 , n7480 );
buf ( n7482 , n7481 );
nand ( n7483 , n7478 , n7482 );
nand ( n7484 , n7477 , n7483 );
buf ( n7485 , n7484 );
not ( n7486 , n7485 );
buf ( n7487 , n7486 );
buf ( n7488 , n7487 );
not ( n7489 , n7488 );
or ( n7490 , n7474 , n7489 );
buf ( n7491 , n786 );
buf ( n7492 , n828 );
xor ( n7493 , n7491 , n7492 );
buf ( n7494 , n7493 );
buf ( n7495 , n7494 );
not ( n7496 , n7495 );
buf ( n7497 , n1239 );
not ( n7498 , n7497 );
or ( n7499 , n7496 , n7498 );
buf ( n7500 , n1249 );
buf ( n7501 , n7319 );
nand ( n7502 , n7500 , n7501 );
buf ( n7503 , n7502 );
buf ( n7504 , n7503 );
nand ( n7505 , n7499 , n7504 );
buf ( n7506 , n7505 );
buf ( n7507 , n7506 );
nand ( n7508 , n7490 , n7507 );
buf ( n7509 , n7508 );
buf ( n7510 , n7509 );
buf ( n7511 , n7472 );
not ( n7512 , n7511 );
buf ( n7513 , n7484 );
nand ( n7514 , n7512 , n7513 );
buf ( n7515 , n7514 );
buf ( n7516 , n7515 );
nand ( n7517 , n7510 , n7516 );
buf ( n7518 , n7517 );
buf ( n7519 , n7518 );
not ( n7520 , n7519 );
buf ( n7521 , n7520 );
buf ( n7522 , n7521 );
not ( n7523 , n7522 );
buf ( n7524 , n788 );
buf ( n7525 , n826 );
xor ( n7526 , n7524 , n7525 );
buf ( n7527 , n7526 );
buf ( n7528 , n7527 );
not ( n7529 , n7528 );
buf ( n7530 , n7529 );
or ( n7531 , n7530 , n1357 );
or ( n7532 , n4020 , n7290 );
nand ( n7533 , n7531 , n7532 );
buf ( n7534 , n7533 );
not ( n7535 , n7534 );
xor ( n7536 , n820 , n794 );
buf ( n7537 , n7536 );
not ( n7538 , n7537 );
buf ( n7539 , n2410 );
not ( n7540 , n7539 );
or ( n7541 , n7538 , n7540 );
buf ( n7542 , n2672 );
buf ( n7543 , n7364 );
nand ( n7544 , n7542 , n7543 );
buf ( n7545 , n7544 );
buf ( n7546 , n7545 );
nand ( n7547 , n7541 , n7546 );
buf ( n7548 , n7547 );
buf ( n7549 , n7548 );
not ( n7550 , n7549 );
or ( n7551 , n7535 , n7550 );
buf ( n7552 , n7533 );
buf ( n7553 , n7548 );
or ( n7554 , n7552 , n7553 );
buf ( n7555 , n796 );
buf ( n7556 , n818 );
xor ( n7557 , n7555 , n7556 );
buf ( n7558 , n7557 );
buf ( n7559 , n7558 );
not ( n7560 , n7559 );
buf ( n7561 , n1480 );
not ( n7562 , n7561 );
or ( n7563 , n7560 , n7562 );
buf ( n7564 , n1496 );
buf ( n7565 , n7398 );
nand ( n7566 , n7564 , n7565 );
buf ( n7567 , n7566 );
buf ( n7568 , n7567 );
nand ( n7569 , n7563 , n7568 );
buf ( n7570 , n7569 );
buf ( n7571 , n7570 );
nand ( n7572 , n7554 , n7571 );
buf ( n7573 , n7572 );
buf ( n7574 , n7573 );
nand ( n7575 , n7551 , n7574 );
buf ( n7576 , n7575 );
not ( n7577 , n7576 );
buf ( n7578 , n7577 );
not ( n7579 , n7578 );
or ( n7580 , n7523 , n7579 );
buf ( n7581 , n790 );
buf ( n7582 , n824 );
xor ( n7583 , n7581 , n7582 );
buf ( n7584 , n7583 );
buf ( n7585 , n7584 );
not ( n7586 , n7585 );
buf ( n7587 , n2790 );
not ( n7588 , n7587 );
or ( n7589 , n7586 , n7588 );
buf ( n7590 , n2492 );
buf ( n7591 , n7215 );
nand ( n7592 , n7590 , n7591 );
buf ( n7593 , n7592 );
buf ( n7594 , n7593 );
nand ( n7595 , n7589 , n7594 );
buf ( n7596 , n7595 );
not ( n7597 , n7596 );
buf ( n7598 , n3739 );
xor ( n7599 , n822 , n792 );
buf ( n7600 , n7599 );
and ( n7601 , n7598 , n7600 );
buf ( n7602 , n3745 );
buf ( n7603 , n7267 );
and ( n7604 , n7602 , n7603 );
nor ( n7605 , n7601 , n7604 );
buf ( n7606 , n7605 );
buf ( n7607 , n7606 );
not ( n7608 , n7607 );
buf ( n7609 , n7608 );
not ( n7610 , n7609 );
or ( n7611 , n7597 , n7610 );
buf ( n7612 , n7606 );
not ( n7613 , n7612 );
buf ( n7614 , n7596 );
not ( n7615 , n7614 );
buf ( n7616 , n7615 );
buf ( n7617 , n7616 );
not ( n7618 , n7617 );
or ( n7619 , n7613 , n7618 );
buf ( n7620 , n798 );
buf ( n7621 , n816 );
xor ( n7622 , n7620 , n7621 );
buf ( n7623 , n7622 );
buf ( n7624 , n7623 );
not ( n7625 , n7624 );
buf ( n7626 , n2526 );
buf ( n7627 , n7626 );
buf ( n7628 , n7627 );
buf ( n7629 , n7628 );
not ( n7630 , n7629 );
or ( n7631 , n7625 , n7630 );
buf ( n7632 , n2010 );
buf ( n7633 , n7235 );
nand ( n7634 , n7632 , n7633 );
buf ( n7635 , n7634 );
buf ( n7636 , n7635 );
nand ( n7637 , n7631 , n7636 );
buf ( n7638 , n7637 );
buf ( n7639 , n7638 );
nand ( n7640 , n7619 , n7639 );
buf ( n7641 , n7640 );
nand ( n7642 , n7611 , n7641 );
buf ( n7643 , n7642 );
nand ( n7644 , n7580 , n7643 );
buf ( n7645 , n7644 );
buf ( n7646 , n7645 );
buf ( n7647 , n7576 );
buf ( n7648 , n7518 );
nand ( n7649 , n7647 , n7648 );
buf ( n7650 , n7649 );
buf ( n7651 , n7650 );
nand ( n7652 , n7646 , n7651 );
buf ( n7653 , n7652 );
not ( n7654 , n7653 );
xor ( n7655 , n7263 , n7333 );
xor ( n7656 , n7655 , n7337 );
not ( n7657 , n7656 );
or ( n7658 , n7654 , n7657 );
or ( n7659 , n7656 , n7653 );
not ( n7660 , n7243 );
not ( n7661 , n7217 );
or ( n7662 , n7660 , n7661 );
or ( n7663 , n7217 , n7243 );
nand ( n7664 , n7662 , n7663 );
buf ( n7665 , n7664 );
buf ( n7666 , n7230 );
xnor ( n7667 , n7665 , n7666 );
buf ( n7668 , n7667 );
buf ( n7669 , n7668 );
not ( n7670 , n7669 );
buf ( n7671 , n7670 );
buf ( n7672 , n7671 );
not ( n7673 , n7672 );
xor ( n7674 , n7410 , n7376 );
buf ( n7675 , n7674 );
buf ( n7676 , n7388 );
xnor ( n7677 , n7675 , n7676 );
buf ( n7678 , n7677 );
not ( n7679 , n7678 );
buf ( n7680 , n7679 );
not ( n7681 , n7680 );
or ( n7682 , n7673 , n7681 );
buf ( n7683 , n7678 );
not ( n7684 , n7683 );
buf ( n7685 , n7668 );
not ( n7686 , n7685 );
or ( n7687 , n7684 , n7686 );
xor ( n7688 , n7313 , n7331 );
buf ( n7689 , n7688 );
buf ( n7690 , n7298 );
buf ( n7691 , n7690 );
and ( n7692 , n7689 , n7691 );
not ( n7693 , n7689 );
not ( n7694 , n7690 );
buf ( n7695 , n7694 );
and ( n7696 , n7693 , n7695 );
nor ( n7697 , n7692 , n7696 );
buf ( n7698 , n7697 );
buf ( n7699 , n7698 );
nand ( n7700 , n7687 , n7699 );
buf ( n7701 , n7700 );
buf ( n7702 , n7701 );
nand ( n7703 , n7682 , n7702 );
buf ( n7704 , n7703 );
nand ( n7705 , n7659 , n7704 );
nand ( n7706 , n7658 , n7705 );
xor ( n7707 , n7468 , n7706 );
xor ( n7708 , n7261 , n7340 );
xor ( n7709 , n7708 , n7429 );
and ( n7710 , n7707 , n7709 );
and ( n7711 , n7468 , n7706 );
or ( n7712 , n7710 , n7711 );
buf ( n7713 , n7712 );
xor ( n7714 , n7465 , n7713 );
xor ( n7715 , n7258 , n7432 );
xor ( n7716 , n7715 , n7443 );
buf ( n7717 , n7716 );
and ( n7718 , n7714 , n7717 );
and ( n7719 , n7465 , n7713 );
or ( n7720 , n7718 , n7719 );
buf ( n7721 , n7720 );
buf ( n7722 , n7721 );
nor ( n7723 , n7464 , n7722 );
buf ( n7724 , n7723 );
xor ( n7725 , n7465 , n7713 );
xor ( n7726 , n7725 , n7717 );
buf ( n7727 , n7726 );
buf ( n7728 , n844 );
buf ( n7729 , n7427 );
not ( n7730 , n7729 );
xor ( n7731 , n7416 , n7362 );
buf ( n7732 , n7731 );
not ( n7733 , n7732 );
or ( n7734 , n7730 , n7733 );
buf ( n7735 , n7731 );
buf ( n7736 , n7427 );
or ( n7737 , n7735 , n7736 );
nand ( n7738 , n7734 , n7737 );
buf ( n7739 , n7738 );
buf ( n7740 , n7739 );
not ( n7741 , n7740 );
buf ( n7742 , n799 );
buf ( n7743 , n817 );
or ( n7744 , n7742 , n7743 );
buf ( n7745 , n818 );
nand ( n7746 , n7744 , n7745 );
buf ( n7747 , n7746 );
buf ( n7748 , n7747 );
buf ( n7749 , n799 );
buf ( n7750 , n817 );
nand ( n7751 , n7749 , n7750 );
buf ( n7752 , n7751 );
buf ( n7753 , n7752 );
buf ( n7754 , n816 );
and ( n7755 , n7748 , n7753 , n7754 );
buf ( n7756 , n7755 );
buf ( n7757 , n7756 );
buf ( n7758 , n785 );
buf ( n7759 , n830 );
xor ( n7760 , n7758 , n7759 );
buf ( n7761 , n7760 );
buf ( n7762 , n7761 );
not ( n7763 , n7762 );
buf ( n7764 , n1161 );
not ( n7765 , n7764 );
or ( n7766 , n7763 , n7765 );
buf ( n7767 , n7482 );
buf ( n7768 , n831 );
nand ( n7769 , n7767 , n7768 );
buf ( n7770 , n7769 );
buf ( n7771 , n7770 );
nand ( n7772 , n7766 , n7771 );
buf ( n7773 , n7772 );
buf ( n7774 , n7773 );
and ( n7775 , n7757 , n7774 );
buf ( n7776 , n7775 );
buf ( n7777 , n791 );
buf ( n7778 , n824 );
xor ( n7779 , n7777 , n7778 );
buf ( n7780 , n7779 );
buf ( n7781 , n7780 );
not ( n7782 , n7781 );
buf ( n7783 , n2790 );
not ( n7784 , n7783 );
or ( n7785 , n7782 , n7784 );
buf ( n7786 , n2492 );
buf ( n7787 , n7584 );
nand ( n7788 , n7786 , n7787 );
buf ( n7789 , n7788 );
buf ( n7790 , n7789 );
nand ( n7791 , n7785 , n7790 );
buf ( n7792 , n7791 );
not ( n7793 , n7792 );
not ( n7794 , n2010 );
not ( n7795 , n7623 );
or ( n7796 , n7794 , n7795 );
not ( n7797 , n2526 );
buf ( n7798 , n799 );
buf ( n7799 , n816 );
xor ( n7800 , n7798 , n7799 );
buf ( n7801 , n7800 );
not ( n7802 , n7801 );
or ( n7803 , n7797 , n7802 );
nand ( n7804 , n7796 , n7803 );
not ( n7805 , n7804 );
or ( n7806 , n7793 , n7805 );
or ( n7807 , n7804 , n7792 );
buf ( n7808 , n787 );
buf ( n7809 , n828 );
xor ( n7810 , n7808 , n7809 );
buf ( n7811 , n7810 );
buf ( n7812 , n7811 );
not ( n7813 , n7812 );
buf ( n7814 , n1239 );
not ( n7815 , n7814 );
or ( n7816 , n7813 , n7815 );
buf ( n7817 , n1249 );
buf ( n7818 , n7494 );
nand ( n7819 , n7817 , n7818 );
buf ( n7820 , n7819 );
buf ( n7821 , n7820 );
nand ( n7822 , n7816 , n7821 );
buf ( n7823 , n7822 );
nand ( n7824 , n7807 , n7823 );
nand ( n7825 , n7806 , n7824 );
xor ( n7826 , n7776 , n7825 );
buf ( n7827 , n795 );
buf ( n7828 , n820 );
xor ( n7829 , n7827 , n7828 );
buf ( n7830 , n7829 );
buf ( n7831 , n7830 );
not ( n7832 , n7831 );
buf ( n7833 , n2410 );
not ( n7834 , n7833 );
or ( n7835 , n7832 , n7834 );
buf ( n7836 , n7536 );
buf ( n7837 , n1346 );
nand ( n7838 , n7836 , n7837 );
buf ( n7839 , n7838 );
buf ( n7840 , n7839 );
nand ( n7841 , n7835 , n7840 );
buf ( n7842 , n7841 );
buf ( n7843 , n7842 );
not ( n7844 , n2101 );
xor ( n7845 , n822 , n793 );
not ( n7846 , n7845 );
or ( n7847 , n7844 , n7846 );
buf ( n7848 , n2113 );
buf ( n7849 , n7599 );
nand ( n7850 , n7848 , n7849 );
buf ( n7851 , n7850 );
nand ( n7852 , n7847 , n7851 );
buf ( n7853 , n7852 );
or ( n7854 , n7843 , n7853 );
buf ( n7855 , n789 );
buf ( n7856 , n826 );
xor ( n7857 , n7855 , n7856 );
buf ( n7858 , n7857 );
buf ( n7859 , n7858 );
not ( n7860 , n7859 );
buf ( n7861 , n1780 );
not ( n7862 , n7861 );
or ( n7863 , n7860 , n7862 );
buf ( n7864 , n1771 );
buf ( n7865 , n7527 );
nand ( n7866 , n7864 , n7865 );
buf ( n7867 , n7866 );
buf ( n7868 , n7867 );
nand ( n7869 , n7863 , n7868 );
buf ( n7870 , n7869 );
buf ( n7871 , n7870 );
nand ( n7872 , n7854 , n7871 );
buf ( n7873 , n7872 );
buf ( n7874 , n7873 );
buf ( n7875 , n7842 );
buf ( n7876 , n7852 );
nand ( n7877 , n7875 , n7876 );
buf ( n7878 , n7877 );
buf ( n7879 , n7878 );
nand ( n7880 , n7874 , n7879 );
buf ( n7881 , n7880 );
and ( n7882 , n7826 , n7881 );
and ( n7883 , n7776 , n7825 );
or ( n7884 , n7882 , n7883 );
buf ( n7885 , n7884 );
not ( n7886 , n7885 );
not ( n7887 , n7576 );
not ( n7888 , n7518 );
or ( n7889 , n7887 , n7888 );
nand ( n7890 , n7521 , n7577 );
nand ( n7891 , n7889 , n7890 );
xor ( n7892 , n7891 , n7642 );
not ( n7893 , n7892 );
buf ( n7894 , n7893 );
not ( n7895 , n7894 );
or ( n7896 , n7886 , n7895 );
buf ( n7897 , n7892 );
not ( n7898 , n7897 );
buf ( n7899 , n7884 );
not ( n7900 , n7899 );
buf ( n7901 , n7900 );
buf ( n7902 , n7901 );
not ( n7903 , n7902 );
or ( n7904 , n7898 , n7903 );
not ( n7905 , n7472 );
not ( n7906 , n7905 );
not ( n7907 , n7484 );
or ( n7908 , n7906 , n7907 );
or ( n7909 , n7905 , n7484 );
nand ( n7910 , n7908 , n7909 );
xnor ( n7911 , n7506 , n7910 );
buf ( n7912 , n7911 );
not ( n7913 , n7533 );
not ( n7914 , n7913 );
not ( n7915 , n7548 );
not ( n7916 , n7570 );
not ( n7917 , n7916 );
or ( n7918 , n7915 , n7917 );
not ( n7919 , n7548 );
nand ( n7920 , n7919 , n7570 );
nand ( n7921 , n7918 , n7920 );
not ( n7922 , n7921 );
or ( n7923 , n7914 , n7922 );
or ( n7924 , n7921 , n7913 );
nand ( n7925 , n7923 , n7924 );
buf ( n7926 , n7925 );
xor ( n7927 , n7912 , n7926 );
xor ( n7928 , n7616 , n7638 );
xnor ( n7929 , n7928 , n7609 );
buf ( n7930 , n7929 );
and ( n7931 , n7927 , n7930 );
and ( n7932 , n7912 , n7926 );
or ( n7933 , n7931 , n7932 );
buf ( n7934 , n7933 );
buf ( n7935 , n7934 );
nand ( n7936 , n7904 , n7935 );
buf ( n7937 , n7936 );
buf ( n7938 , n7937 );
nand ( n7939 , n7896 , n7938 );
buf ( n7940 , n7939 );
not ( n7941 , n7940 );
or ( n7942 , n7741 , n7941 );
or ( n7943 , n7940 , n7740 );
xor ( n7944 , n7653 , n7656 );
xor ( n7945 , n7944 , n7704 );
nand ( n7946 , n7943 , n7945 );
nand ( n7947 , n7942 , n7946 );
buf ( n7948 , n7947 );
xor ( n7949 , n7728 , n7948 );
xor ( n7950 , n7468 , n7706 );
xor ( n7951 , n7950 , n7709 );
buf ( n7952 , n7951 );
and ( n7953 , n7949 , n7952 );
and ( n7954 , n7728 , n7948 );
or ( n7955 , n7953 , n7954 );
buf ( n7956 , n7955 );
nor ( n7957 , n7727 , n7956 );
nor ( n7958 , n7724 , n7957 );
nand ( n7959 , n7460 , n7958 );
not ( n7960 , n7959 );
buf ( n7961 , n845 );
buf ( n7962 , n7668 );
not ( n7963 , n7962 );
buf ( n7964 , n7698 );
not ( n7965 , n7964 );
and ( n7966 , n7963 , n7965 );
buf ( n7967 , n7668 );
buf ( n7968 , n7698 );
and ( n7969 , n7967 , n7968 );
nor ( n7970 , n7966 , n7969 );
buf ( n7971 , n7970 );
buf ( n7972 , n7971 );
not ( n7973 , n7679 );
buf ( n7974 , n7973 );
and ( n7975 , n7972 , n7974 );
not ( n7976 , n7972 );
buf ( n7977 , n7679 );
and ( n7978 , n7976 , n7977 );
nor ( n7979 , n7975 , n7978 );
buf ( n7980 , n7979 );
buf ( n7981 , n7980 );
buf ( n7982 , n797 );
buf ( n7983 , n818 );
xor ( n7984 , n7982 , n7983 );
buf ( n7985 , n7984 );
buf ( n7986 , n7985 );
not ( n7987 , n7986 );
buf ( n7988 , n2725 );
not ( n7989 , n7988 );
or ( n7990 , n7987 , n7989 );
buf ( n7991 , n1496 );
buf ( n7992 , n7558 );
nand ( n7993 , n7991 , n7992 );
buf ( n7994 , n7993 );
buf ( n7995 , n7994 );
nand ( n7996 , n7990 , n7995 );
buf ( n7997 , n7996 );
buf ( n7998 , n7997 );
xor ( n7999 , n7757 , n7774 );
buf ( n8000 , n7999 );
buf ( n8001 , n8000 );
xor ( n8002 , n7998 , n8001 );
buf ( n8003 , n2010 );
buf ( n8004 , n799 );
and ( n8005 , n8003 , n8004 );
buf ( n8006 , n8005 );
buf ( n8007 , n8006 );
buf ( n8008 , n786 );
buf ( n8009 , n830 );
xor ( n8010 , n8008 , n8009 );
buf ( n8011 , n8010 );
buf ( n8012 , n8011 );
not ( n8013 , n8012 );
buf ( n8014 , n1630 );
not ( n8015 , n8014 );
or ( n8016 , n8013 , n8015 );
buf ( n8017 , n7761 );
buf ( n8018 , n831 );
nand ( n8019 , n8017 , n8018 );
buf ( n8020 , n8019 );
buf ( n8021 , n8020 );
nand ( n8022 , n8016 , n8021 );
buf ( n8023 , n8022 );
buf ( n8024 , n8023 );
xor ( n8025 , n8007 , n8024 );
buf ( n8026 , n788 );
buf ( n8027 , n828 );
xor ( n8028 , n8026 , n8027 );
buf ( n8029 , n8028 );
buf ( n8030 , n8029 );
not ( n8031 , n8030 );
buf ( n8032 , n1901 );
not ( n8033 , n8032 );
or ( n8034 , n8031 , n8033 );
buf ( n8035 , n1249 );
buf ( n8036 , n7811 );
nand ( n8037 , n8035 , n8036 );
buf ( n8038 , n8037 );
buf ( n8039 , n8038 );
nand ( n8040 , n8034 , n8039 );
buf ( n8041 , n8040 );
buf ( n8042 , n8041 );
and ( n8043 , n8025 , n8042 );
and ( n8044 , n8007 , n8024 );
or ( n8045 , n8043 , n8044 );
buf ( n8046 , n8045 );
buf ( n8047 , n8046 );
and ( n8048 , n8002 , n8047 );
and ( n8049 , n7998 , n8001 );
or ( n8050 , n8048 , n8049 );
buf ( n8051 , n8050 );
buf ( n8052 , n8051 );
xor ( n8053 , n7776 , n7825 );
xor ( n8054 , n8053 , n7881 );
buf ( n8055 , n8054 );
xor ( n8056 , n8052 , n8055 );
buf ( n8057 , n794 );
buf ( n8058 , n822 );
xor ( n8059 , n8057 , n8058 );
buf ( n8060 , n8059 );
not ( n8061 , n8060 );
not ( n8062 , n3739 );
or ( n8063 , n8061 , n8062 );
buf ( n8064 , n2113 );
buf ( n8065 , n7845 );
nand ( n8066 , n8064 , n8065 );
buf ( n8067 , n8066 );
nand ( n8068 , n8063 , n8067 );
not ( n8069 , n8068 );
buf ( n8070 , n792 );
buf ( n8071 , n824 );
xor ( n8072 , n8070 , n8071 );
buf ( n8073 , n8072 );
not ( n8074 , n8073 );
not ( n8075 , n2790 );
or ( n8076 , n8074 , n8075 );
buf ( n8077 , n2492 );
buf ( n8078 , n7780 );
nand ( n8079 , n8077 , n8078 );
buf ( n8080 , n8079 );
nand ( n8081 , n8076 , n8080 );
not ( n8082 , n8081 );
or ( n8083 , n8069 , n8082 );
or ( n8084 , n8081 , n8068 );
xor ( n8085 , n826 , n790 );
buf ( n8086 , n8085 );
not ( n8087 , n8086 );
buf ( n8088 , n6463 );
not ( n8089 , n8088 );
buf ( n8090 , n8089 );
buf ( n8091 , n8090 );
not ( n8092 , n8091 );
or ( n8093 , n8087 , n8092 );
buf ( n8094 , n1771 );
buf ( n8095 , n7858 );
nand ( n8096 , n8094 , n8095 );
buf ( n8097 , n8096 );
buf ( n8098 , n8097 );
nand ( n8099 , n8093 , n8098 );
buf ( n8100 , n8099 );
nand ( n8101 , n8084 , n8100 );
nand ( n8102 , n8083 , n8101 );
buf ( n8103 , n8102 );
xor ( n8104 , n7792 , n7823 );
xor ( n8105 , n8104 , n7804 );
buf ( n8106 , n8105 );
xor ( n8107 , n8103 , n8106 );
buf ( n8108 , n7852 );
not ( n8109 , n8108 );
not ( n8110 , n7870 );
xor ( n8111 , n7842 , n8110 );
buf ( n8112 , n8111 );
not ( n8113 , n8112 );
or ( n8114 , n8109 , n8113 );
buf ( n8115 , n8111 );
buf ( n8116 , n7852 );
or ( n8117 , n8115 , n8116 );
nand ( n8118 , n8114 , n8117 );
buf ( n8119 , n8118 );
buf ( n8120 , n8119 );
and ( n8121 , n8107 , n8120 );
and ( n8122 , n8103 , n8106 );
or ( n8123 , n8121 , n8122 );
buf ( n8124 , n8123 );
buf ( n8125 , n8124 );
and ( n8126 , n8056 , n8125 );
and ( n8127 , n8052 , n8055 );
or ( n8128 , n8126 , n8127 );
buf ( n8129 , n8128 );
buf ( n8130 , n8129 );
xor ( n8131 , n7981 , n8130 );
buf ( n8132 , n7893 );
not ( n8133 , n8132 );
buf ( n8134 , n7901 );
not ( n8135 , n8134 );
or ( n8136 , n8133 , n8135 );
buf ( n8137 , n7892 );
buf ( n8138 , n7884 );
nand ( n8139 , n8137 , n8138 );
buf ( n8140 , n8139 );
buf ( n8141 , n8140 );
nand ( n8142 , n8136 , n8141 );
buf ( n8143 , n8142 );
buf ( n8144 , n8143 );
buf ( n8145 , n7934 );
and ( n8146 , n8144 , n8145 );
not ( n8147 , n8144 );
buf ( n8148 , n7934 );
not ( n8149 , n8148 );
buf ( n8150 , n8149 );
buf ( n8151 , n8150 );
and ( n8152 , n8147 , n8151 );
nor ( n8153 , n8146 , n8152 );
buf ( n8154 , n8153 );
buf ( n8155 , n8154 );
and ( n8156 , n8131 , n8155 );
and ( n8157 , n7981 , n8130 );
or ( n8158 , n8156 , n8157 );
buf ( n8159 , n8158 );
buf ( n8160 , n8159 );
xor ( n8161 , n7961 , n8160 );
xor ( n8162 , n7739 , n7940 );
xor ( n8163 , n8162 , n7945 );
buf ( n8164 , n8163 );
xor ( n8165 , n8161 , n8164 );
buf ( n8166 , n8165 );
buf ( n8167 , n8166 );
buf ( n8168 , n846 );
xor ( n8169 , n7912 , n7926 );
xor ( n8170 , n8169 , n7930 );
buf ( n8171 , n8170 );
buf ( n8172 , n8171 );
buf ( n8173 , n787 );
buf ( n8174 , n830 );
xor ( n8175 , n8173 , n8174 );
buf ( n8176 , n8175 );
buf ( n8177 , n8176 );
not ( n8178 , n8177 );
buf ( n8179 , n1161 );
not ( n8180 , n8179 );
or ( n8181 , n8178 , n8180 );
buf ( n8182 , n8011 );
buf ( n8183 , n831 );
nand ( n8184 , n8182 , n8183 );
buf ( n8185 , n8184 );
buf ( n8186 , n8185 );
nand ( n8187 , n8181 , n8186 );
buf ( n8188 , n8187 );
buf ( n8189 , n8188 );
buf ( n8190 , n799 );
buf ( n8191 , n819 );
or ( n8192 , n8190 , n8191 );
buf ( n8193 , n820 );
nand ( n8194 , n8192 , n8193 );
buf ( n8195 , n8194 );
buf ( n8196 , n8195 );
buf ( n8197 , n799 );
buf ( n8198 , n819 );
nand ( n8199 , n8197 , n8198 );
buf ( n8200 , n8199 );
buf ( n8201 , n8200 );
buf ( n8202 , n818 );
nand ( n8203 , n8196 , n8201 , n8202 );
buf ( n8204 , n8203 );
buf ( n8205 , n8204 );
not ( n8206 , n8205 );
buf ( n8207 , n8206 );
buf ( n8208 , n8207 );
and ( n8209 , n8189 , n8208 );
buf ( n8210 , n8209 );
buf ( n8211 , n8210 );
xor ( n8212 , n820 , n796 );
buf ( n8213 , n8212 );
not ( n8214 , n8213 );
buf ( n8215 , n2267 );
not ( n8216 , n8215 );
or ( n8217 , n8214 , n8216 );
buf ( n8218 , n2672 );
buf ( n8219 , n7830 );
nand ( n8220 , n8218 , n8219 );
buf ( n8221 , n8220 );
buf ( n8222 , n8221 );
nand ( n8223 , n8217 , n8222 );
buf ( n8224 , n8223 );
buf ( n8225 , n8224 );
nor ( n8226 , n8211 , n8225 );
buf ( n8227 , n8226 );
buf ( n8228 , n8227 );
buf ( n8229 , n798 );
buf ( n8230 , n818 );
xor ( n8231 , n8229 , n8230 );
buf ( n8232 , n8231 );
buf ( n8233 , n8232 );
not ( n8234 , n8233 );
buf ( n8235 , n1480 );
not ( n8236 , n8235 );
or ( n8237 , n8234 , n8236 );
buf ( n8238 , n1496 );
buf ( n8239 , n7985 );
nand ( n8240 , n8238 , n8239 );
buf ( n8241 , n8240 );
buf ( n8242 , n8241 );
nand ( n8243 , n8237 , n8242 );
buf ( n8244 , n8243 );
buf ( n8245 , n8244 );
not ( n8246 , n8245 );
buf ( n8247 , n8246 );
buf ( n8248 , n8247 );
or ( n8249 , n8228 , n8248 );
buf ( n8250 , n8224 );
buf ( n8251 , n8210 );
nand ( n8252 , n8250 , n8251 );
buf ( n8253 , n8252 );
buf ( n8254 , n8253 );
nand ( n8255 , n8249 , n8254 );
buf ( n8256 , n8255 );
buf ( n8257 , n8256 );
xor ( n8258 , n7998 , n8001 );
xor ( n8259 , n8258 , n8047 );
buf ( n8260 , n8259 );
buf ( n8261 , n8260 );
xor ( n8262 , n8257 , n8261 );
xor ( n8263 , n8007 , n8024 );
xor ( n8264 , n8263 , n8042 );
buf ( n8265 , n8264 );
xor ( n8266 , n826 , n791 );
buf ( n8267 , n8266 );
not ( n8268 , n8267 );
buf ( n8269 , n4496 );
not ( n8270 , n8269 );
or ( n8271 , n8268 , n8270 );
buf ( n8272 , n1771 );
buf ( n8273 , n8085 );
nand ( n8274 , n8272 , n8273 );
buf ( n8275 , n8274 );
buf ( n8276 , n8275 );
nand ( n8277 , n8271 , n8276 );
buf ( n8278 , n8277 );
buf ( n8279 , n8278 );
not ( n8280 , n8279 );
xor ( n8281 , n820 , n797 );
buf ( n8282 , n8281 );
not ( n8283 , n8282 );
buf ( n8284 , n2410 );
not ( n8285 , n8284 );
or ( n8286 , n8283 , n8285 );
buf ( n8287 , n1346 );
buf ( n8288 , n8212 );
nand ( n8289 , n8287 , n8288 );
buf ( n8290 , n8289 );
buf ( n8291 , n8290 );
nand ( n8292 , n8286 , n8291 );
buf ( n8293 , n8292 );
buf ( n8294 , n8293 );
not ( n8295 , n8294 );
or ( n8296 , n8280 , n8295 );
buf ( n8297 , n8293 );
buf ( n8298 , n8278 );
or ( n8299 , n8297 , n8298 );
buf ( n8300 , n799 );
buf ( n8301 , n818 );
xor ( n8302 , n8300 , n8301 );
buf ( n8303 , n8302 );
buf ( n8304 , n8303 );
not ( n8305 , n8304 );
buf ( n8306 , n1480 );
not ( n8307 , n8306 );
or ( n8308 , n8305 , n8307 );
buf ( n8309 , n1496 );
buf ( n8310 , n8232 );
nand ( n8311 , n8309 , n8310 );
buf ( n8312 , n8311 );
buf ( n8313 , n8312 );
nand ( n8314 , n8308 , n8313 );
buf ( n8315 , n8314 );
buf ( n8316 , n8315 );
nand ( n8317 , n8299 , n8316 );
buf ( n8318 , n8317 );
buf ( n8319 , n8318 );
nand ( n8320 , n8296 , n8319 );
buf ( n8321 , n8320 );
and ( n8322 , n8265 , n8321 );
not ( n8323 , n8322 );
not ( n8324 , n8265 );
not ( n8325 , n8324 );
not ( n8326 , n8321 );
not ( n8327 , n8326 );
or ( n8328 , n8325 , n8327 );
xor ( n8329 , n828 , n789 );
buf ( n8330 , n8329 );
not ( n8331 , n8330 );
buf ( n8332 , n3680 );
not ( n8333 , n8332 );
or ( n8334 , n8331 , n8333 );
buf ( n8335 , n1249 );
buf ( n8336 , n8029 );
nand ( n8337 , n8335 , n8336 );
buf ( n8338 , n8337 );
buf ( n8339 , n8338 );
nand ( n8340 , n8334 , n8339 );
buf ( n8341 , n8340 );
not ( n8342 , n8341 );
buf ( n8343 , n793 );
buf ( n8344 , n824 );
xor ( n8345 , n8343 , n8344 );
buf ( n8346 , n8345 );
buf ( n8347 , n8346 );
not ( n8348 , n8347 );
buf ( n8349 , n2790 );
not ( n8350 , n8349 );
or ( n8351 , n8348 , n8350 );
buf ( n8352 , n2489 );
not ( n8353 , n8352 );
buf ( n8354 , n8353 );
buf ( n8355 , n8354 );
buf ( n8356 , n8073 );
nand ( n8357 , n8355 , n8356 );
buf ( n8358 , n8357 );
buf ( n8359 , n8358 );
nand ( n8360 , n8351 , n8359 );
buf ( n8361 , n8360 );
not ( n8362 , n8361 );
nand ( n8363 , n8342 , n8362 );
not ( n8364 , n8363 );
buf ( n8365 , n795 );
buf ( n8366 , n822 );
xor ( n8367 , n8365 , n8366 );
buf ( n8368 , n8367 );
buf ( n8369 , n8368 );
not ( n8370 , n8369 );
buf ( n8371 , n3739 );
not ( n8372 , n8371 );
or ( n8373 , n8370 , n8372 );
buf ( n8374 , n3745 );
buf ( n8375 , n8060 );
nand ( n8376 , n8374 , n8375 );
buf ( n8377 , n8376 );
buf ( n8378 , n8377 );
nand ( n8379 , n8373 , n8378 );
buf ( n8380 , n8379 );
not ( n8381 , n8380 );
or ( n8382 , n8364 , n8381 );
nand ( n8383 , n8361 , n8341 );
nand ( n8384 , n8382 , n8383 );
nand ( n8385 , n8328 , n8384 );
nand ( n8386 , n8323 , n8385 );
buf ( n8387 , n8386 );
and ( n8388 , n8262 , n8387 );
and ( n8389 , n8257 , n8261 );
or ( n8390 , n8388 , n8389 );
buf ( n8391 , n8390 );
buf ( n8392 , n8391 );
xor ( n8393 , n8172 , n8392 );
xor ( n8394 , n8052 , n8055 );
xor ( n8395 , n8394 , n8125 );
buf ( n8396 , n8395 );
buf ( n8397 , n8396 );
and ( n8398 , n8393 , n8397 );
and ( n8399 , n8172 , n8392 );
or ( n8400 , n8398 , n8399 );
buf ( n8401 , n8400 );
buf ( n8402 , n8401 );
xor ( n8403 , n8168 , n8402 );
xor ( n8404 , n7981 , n8130 );
xor ( n8405 , n8404 , n8155 );
buf ( n8406 , n8405 );
buf ( n8407 , n8406 );
and ( n8408 , n8403 , n8407 );
and ( n8409 , n8168 , n8402 );
or ( n8410 , n8408 , n8409 );
buf ( n8411 , n8410 );
buf ( n8412 , n8411 );
nor ( n8413 , n8167 , n8412 );
buf ( n8414 , n8413 );
xor ( n8415 , n7961 , n8160 );
and ( n8416 , n8415 , n8164 );
and ( n8417 , n7961 , n8160 );
or ( n8418 , n8416 , n8417 );
buf ( n8419 , n8418 );
buf ( n8420 , n8419 );
xor ( n8421 , n7728 , n7948 );
xor ( n8422 , n8421 , n7952 );
buf ( n8423 , n8422 );
buf ( n8424 , n8423 );
nor ( n8425 , n8420 , n8424 );
buf ( n8426 , n8425 );
nor ( n8427 , n8414 , n8426 );
not ( n8428 , n8427 );
buf ( n8429 , n848 );
not ( n8430 , n8384 );
not ( n8431 , n8324 );
not ( n8432 , n8321 );
or ( n8433 , n8431 , n8432 );
nand ( n8434 , n8326 , n8265 );
nand ( n8435 , n8433 , n8434 );
nand ( n8436 , n8430 , n8435 );
nand ( n8437 , n8322 , n8384 );
nand ( n8438 , n8384 , n8324 , n8326 );
nand ( n8439 , n8436 , n8437 , n8438 );
buf ( n8440 , n8439 );
xor ( n8441 , n8341 , n8362 );
not ( n8442 , n8380 );
xor ( n8443 , n8441 , n8442 );
xor ( n8444 , n8315 , n8278 );
xor ( n8445 , n8444 , n8293 );
xor ( n8446 , n8443 , n8445 );
buf ( n8447 , n826 );
buf ( n8448 , n792 );
xor ( n8449 , n8447 , n8448 );
buf ( n8450 , n8449 );
buf ( n8451 , n8450 );
not ( n8452 , n8451 );
buf ( n8453 , n1780 );
not ( n8454 , n8453 );
or ( n8455 , n8452 , n8454 );
buf ( n8456 , n1771 );
buf ( n8457 , n8266 );
nand ( n8458 , n8456 , n8457 );
buf ( n8459 , n8458 );
buf ( n8460 , n8459 );
nand ( n8461 , n8455 , n8460 );
buf ( n8462 , n8461 );
buf ( n8463 , n8462 );
buf ( n8464 , n791 );
buf ( n8465 , n828 );
xor ( n8466 , n8464 , n8465 );
buf ( n8467 , n8466 );
buf ( n8468 , n8467 );
not ( n8469 , n8468 );
buf ( n8470 , n3680 );
not ( n8471 , n8470 );
or ( n8472 , n8469 , n8471 );
buf ( n8473 , n1249 );
xor ( n8474 , n828 , n790 );
buf ( n8475 , n8474 );
nand ( n8476 , n8473 , n8475 );
buf ( n8477 , n8476 );
buf ( n8478 , n8477 );
nand ( n8479 , n8472 , n8478 );
buf ( n8480 , n8479 );
buf ( n8481 , n8480 );
not ( n8482 , n8481 );
buf ( n8483 , n799 );
buf ( n8484 , n821 );
or ( n8485 , n8483 , n8484 );
buf ( n8486 , n822 );
nand ( n8487 , n8485 , n8486 );
buf ( n8488 , n8487 );
buf ( n8489 , n8488 );
buf ( n8490 , n799 );
buf ( n8491 , n821 );
nand ( n8492 , n8490 , n8491 );
buf ( n8493 , n8492 );
buf ( n8494 , n8493 );
buf ( n8495 , n820 );
nand ( n8496 , n8489 , n8494 , n8495 );
buf ( n8497 , n8496 );
buf ( n8498 , n8497 );
nor ( n8499 , n8482 , n8498 );
buf ( n8500 , n8499 );
buf ( n8501 , n8500 );
xor ( n8502 , n8463 , n8501 );
buf ( n8503 , n789 );
buf ( n8504 , n830 );
xor ( n8505 , n8503 , n8504 );
buf ( n8506 , n8505 );
buf ( n8507 , n8506 );
not ( n8508 , n8507 );
buf ( n8509 , n1161 );
not ( n8510 , n8509 );
or ( n8511 , n8508 , n8510 );
buf ( n8512 , n788 );
buf ( n8513 , n830 );
xor ( n8514 , n8512 , n8513 );
buf ( n8515 , n8514 );
buf ( n8516 , n8515 );
buf ( n8517 , n831 );
nand ( n8518 , n8516 , n8517 );
buf ( n8519 , n8518 );
buf ( n8520 , n8519 );
nand ( n8521 , n8511 , n8520 );
buf ( n8522 , n8521 );
buf ( n8523 , n8522 );
buf ( n8524 , n795 );
buf ( n8525 , n824 );
xor ( n8526 , n8524 , n8525 );
buf ( n8527 , n8526 );
buf ( n8528 , n8527 );
not ( n8529 , n8528 );
buf ( n8530 , n2790 );
not ( n8531 , n8530 );
or ( n8532 , n8529 , n8531 );
buf ( n8533 , n8354 );
buf ( n8534 , n794 );
buf ( n8535 , n824 );
xor ( n8536 , n8534 , n8535 );
buf ( n8537 , n8536 );
buf ( n8538 , n8537 );
nand ( n8539 , n8533 , n8538 );
buf ( n8540 , n8539 );
buf ( n8541 , n8540 );
nand ( n8542 , n8532 , n8541 );
buf ( n8543 , n8542 );
buf ( n8544 , n8543 );
xor ( n8545 , n8523 , n8544 );
buf ( n8546 , n797 );
buf ( n8547 , n822 );
xor ( n8548 , n8546 , n8547 );
buf ( n8549 , n8548 );
buf ( n8550 , n8549 );
not ( n8551 , n8550 );
buf ( n8552 , n2101 );
not ( n8553 , n8552 );
or ( n8554 , n8551 , n8553 );
buf ( n8555 , n3745 );
buf ( n8556 , n796 );
buf ( n8557 , n822 );
xor ( n8558 , n8556 , n8557 );
buf ( n8559 , n8558 );
buf ( n8560 , n8559 );
nand ( n8561 , n8555 , n8560 );
buf ( n8562 , n8561 );
buf ( n8563 , n8562 );
nand ( n8564 , n8554 , n8563 );
buf ( n8565 , n8564 );
buf ( n8566 , n8565 );
and ( n8567 , n8545 , n8566 );
and ( n8568 , n8523 , n8544 );
or ( n8569 , n8567 , n8568 );
buf ( n8570 , n8569 );
buf ( n8571 , n8570 );
and ( n8572 , n8502 , n8571 );
and ( n8573 , n8463 , n8501 );
or ( n8574 , n8572 , n8573 );
buf ( n8575 , n8574 );
and ( n8576 , n8446 , n8575 );
and ( n8577 , n8443 , n8445 );
or ( n8578 , n8576 , n8577 );
buf ( n8579 , n8578 );
xor ( n8580 , n8440 , n8579 );
xor ( n8581 , n8081 , n8068 );
xor ( n8582 , n8581 , n8100 );
buf ( n8583 , n8582 );
buf ( n8584 , n8227 );
not ( n8585 , n8584 );
buf ( n8586 , n8253 );
nand ( n8587 , n8585 , n8586 );
buf ( n8588 , n8587 );
buf ( n8589 , n8588 );
buf ( n8590 , n8247 );
and ( n8591 , n8589 , n8590 );
not ( n8592 , n8589 );
buf ( n8593 , n8244 );
and ( n8594 , n8592 , n8593 );
nor ( n8595 , n8591 , n8594 );
buf ( n8596 , n8595 );
buf ( n8597 , n8596 );
xor ( n8598 , n8583 , n8597 );
buf ( n8599 , n8188 );
buf ( n8600 , n8207 );
and ( n8601 , n8599 , n8600 );
not ( n8602 , n8599 );
buf ( n8603 , n8204 );
and ( n8604 , n8602 , n8603 );
nor ( n8605 , n8601 , n8604 );
buf ( n8606 , n8605 );
buf ( n8607 , n8606 );
buf ( n8608 , n1496 );
buf ( n8609 , n799 );
and ( n8610 , n8608 , n8609 );
buf ( n8611 , n8610 );
buf ( n8612 , n8611 );
buf ( n8613 , n8537 );
not ( n8614 , n8613 );
buf ( n8615 , n2790 );
not ( n8616 , n8615 );
or ( n8617 , n8614 , n8616 );
buf ( n8618 , n2492 );
buf ( n8619 , n8346 );
nand ( n8620 , n8618 , n8619 );
buf ( n8621 , n8620 );
buf ( n8622 , n8621 );
nand ( n8623 , n8617 , n8622 );
buf ( n8624 , n8623 );
buf ( n8625 , n8624 );
xor ( n8626 , n8612 , n8625 );
buf ( n8627 , n8474 );
not ( n8628 , n8627 );
buf ( n8629 , n3680 );
not ( n8630 , n8629 );
or ( n8631 , n8628 , n8630 );
buf ( n8632 , n1249 );
buf ( n8633 , n8329 );
nand ( n8634 , n8632 , n8633 );
buf ( n8635 , n8634 );
buf ( n8636 , n8635 );
nand ( n8637 , n8631 , n8636 );
buf ( n8638 , n8637 );
buf ( n8639 , n8638 );
and ( n8640 , n8626 , n8639 );
and ( n8641 , n8612 , n8625 );
or ( n8642 , n8640 , n8641 );
buf ( n8643 , n8642 );
buf ( n8644 , n8643 );
xor ( n8645 , n8607 , n8644 );
buf ( n8646 , n8515 );
not ( n8647 , n8646 );
buf ( n8648 , n1161 );
not ( n8649 , n8648 );
or ( n8650 , n8647 , n8649 );
buf ( n8651 , n8176 );
buf ( n8652 , n831 );
nand ( n8653 , n8651 , n8652 );
buf ( n8654 , n8653 );
buf ( n8655 , n8654 );
nand ( n8656 , n8650 , n8655 );
buf ( n8657 , n8656 );
buf ( n8658 , n8657 );
buf ( n8659 , n798 );
buf ( n8660 , n820 );
xor ( n8661 , n8659 , n8660 );
buf ( n8662 , n8661 );
buf ( n8663 , n8662 );
not ( n8664 , n8663 );
buf ( n8665 , n2410 );
not ( n8666 , n8665 );
or ( n8667 , n8664 , n8666 );
buf ( n8668 , n2672 );
buf ( n8669 , n8281 );
nand ( n8670 , n8668 , n8669 );
buf ( n8671 , n8670 );
buf ( n8672 , n8671 );
nand ( n8673 , n8667 , n8672 );
buf ( n8674 , n8673 );
buf ( n8675 , n8674 );
xor ( n8676 , n8658 , n8675 );
buf ( n8677 , n8559 );
not ( n8678 , n8677 );
buf ( n8679 , n3739 );
not ( n8680 , n8679 );
or ( n8681 , n8678 , n8680 );
buf ( n8682 , n3745 );
buf ( n8683 , n8368 );
nand ( n8684 , n8682 , n8683 );
buf ( n8685 , n8684 );
buf ( n8686 , n8685 );
nand ( n8687 , n8681 , n8686 );
buf ( n8688 , n8687 );
buf ( n8689 , n8688 );
and ( n8690 , n8676 , n8689 );
and ( n8691 , n8658 , n8675 );
or ( n8692 , n8690 , n8691 );
buf ( n8693 , n8692 );
buf ( n8694 , n8693 );
and ( n8695 , n8645 , n8694 );
and ( n8696 , n8607 , n8644 );
or ( n8697 , n8695 , n8696 );
buf ( n8698 , n8697 );
buf ( n8699 , n8698 );
xor ( n8700 , n8598 , n8699 );
buf ( n8701 , n8700 );
buf ( n8702 , n8701 );
and ( n8703 , n8580 , n8702 );
and ( n8704 , n8440 , n8579 );
or ( n8705 , n8703 , n8704 );
buf ( n8706 , n8705 );
buf ( n8707 , n8706 );
xor ( n8708 , n8429 , n8707 );
xor ( n8709 , n8103 , n8106 );
xor ( n8710 , n8709 , n8120 );
buf ( n8711 , n8710 );
buf ( n8712 , n8711 );
xor ( n8713 , n8257 , n8261 );
xor ( n8714 , n8713 , n8387 );
buf ( n8715 , n8714 );
buf ( n8716 , n8715 );
xor ( n8717 , n8712 , n8716 );
xor ( n8718 , n8583 , n8597 );
and ( n8719 , n8718 , n8699 );
and ( n8720 , n8583 , n8597 );
or ( n8721 , n8719 , n8720 );
buf ( n8722 , n8721 );
buf ( n8723 , n8722 );
xor ( n8724 , n8717 , n8723 );
buf ( n8725 , n8724 );
buf ( n8726 , n8725 );
and ( n8727 , n8708 , n8726 );
and ( n8728 , n8429 , n8707 );
or ( n8729 , n8727 , n8728 );
buf ( n8730 , n8729 );
buf ( n8731 , n8730 );
buf ( n8732 , n847 );
xor ( n8733 , n8712 , n8716 );
and ( n8734 , n8733 , n8723 );
and ( n8735 , n8712 , n8716 );
or ( n8736 , n8734 , n8735 );
buf ( n8737 , n8736 );
buf ( n8738 , n8737 );
xor ( n8739 , n8732 , n8738 );
xor ( n8740 , n8172 , n8392 );
xor ( n8741 , n8740 , n8397 );
buf ( n8742 , n8741 );
buf ( n8743 , n8742 );
xor ( n8744 , n8739 , n8743 );
buf ( n8745 , n8744 );
buf ( n8746 , n8745 );
nand ( n8747 , n8731 , n8746 );
buf ( n8748 , n8747 );
buf ( n8749 , n8748 );
not ( n8750 , n8749 );
xor ( n8751 , n8168 , n8402 );
xor ( n8752 , n8751 , n8407 );
buf ( n8753 , n8752 );
buf ( n8754 , n8753 );
xor ( n8755 , n8732 , n8738 );
and ( n8756 , n8755 , n8743 );
and ( n8757 , n8732 , n8738 );
or ( n8758 , n8756 , n8757 );
buf ( n8759 , n8758 );
buf ( n8760 , n8759 );
nand ( n8761 , n8754 , n8760 );
buf ( n8762 , n8761 );
buf ( n8763 , n8762 );
not ( n8764 , n8763 );
or ( n8765 , n8750 , n8764 );
or ( n8766 , n8753 , n8759 );
buf ( n8767 , n8766 );
nand ( n8768 , n8765 , n8767 );
buf ( n8769 , n8768 );
buf ( n8770 , n8769 );
not ( n8771 , n8770 );
buf ( n8772 , n8771 );
not ( n8773 , n8772 );
or ( n8774 , n8428 , n8773 );
buf ( n8775 , n8426 );
not ( n8776 , n8775 );
buf ( n8777 , n8776 );
buf ( n8778 , n8777 );
buf ( n8779 , n8166 );
not ( n8780 , n8779 );
buf ( n8781 , n8780 );
buf ( n8782 , n8781 );
buf ( n8783 , n8411 );
not ( n8784 , n8783 );
buf ( n8785 , n8784 );
buf ( n8786 , n8785 );
nor ( n8787 , n8782 , n8786 );
buf ( n8788 , n8787 );
buf ( n8789 , n8788 );
and ( n8790 , n8778 , n8789 );
buf ( n8791 , n8423 );
buf ( n8792 , n8419 );
and ( n8793 , n8791 , n8792 );
buf ( n8794 , n8793 );
buf ( n8795 , n8794 );
nor ( n8796 , n8790 , n8795 );
buf ( n8797 , n8796 );
nand ( n8798 , n8774 , n8797 );
nand ( n8799 , n7960 , n8798 );
not ( n8800 , n6890 );
not ( n8801 , n7138 );
and ( n8802 , n8800 , n8801 );
buf ( n8803 , n7456 );
buf ( n8804 , n7144 );
nor ( n8805 , n8803 , n8804 );
buf ( n8806 , n8805 );
nor ( n8807 , n8802 , n8806 );
buf ( n8808 , n8807 );
not ( n8809 , n8808 );
buf ( n8810 , n7727 );
buf ( n8811 , n7956 );
and ( n8812 , n8810 , n8811 );
buf ( n8813 , n8812 );
buf ( n8814 , n8813 );
not ( n8815 , n8814 );
not ( n8816 , n7721 );
buf ( n8817 , n7463 );
not ( n8818 , n8817 );
buf ( n8819 , n8818 );
nand ( n8820 , n8816 , n8819 );
buf ( n8821 , n8820 );
not ( n8822 , n8821 );
or ( n8823 , n8815 , n8822 );
not ( n8824 , n8819 );
nand ( n8825 , n8824 , n7721 );
buf ( n8826 , n8825 );
nand ( n8827 , n8823 , n8826 );
buf ( n8828 , n8827 );
buf ( n8829 , n8828 );
not ( n8830 , n8829 );
or ( n8831 , n8809 , n8830 );
buf ( n8832 , n7141 );
not ( n8833 , n8832 );
buf ( n8834 , n8833 );
buf ( n8835 , n8834 );
buf ( n8836 , n7144 );
buf ( n8837 , n7456 );
nand ( n8838 , n8836 , n8837 );
buf ( n8839 , n8838 );
buf ( n8840 , n8839 );
not ( n8841 , n8840 );
buf ( n8842 , n8841 );
buf ( n8843 , n8842 );
and ( n8844 , n8835 , n8843 );
buf ( n8845 , n7138 );
buf ( n8846 , n6890 );
and ( n8847 , n8845 , n8846 );
buf ( n8848 , n8847 );
buf ( n8849 , n8848 );
nor ( n8850 , n8844 , n8849 );
buf ( n8851 , n8850 );
buf ( n8852 , n8851 );
nand ( n8853 , n8831 , n8852 );
buf ( n8854 , n8853 );
nor ( n8855 , n6884 , n8854 );
nand ( n8856 , n6354 , n8799 , n8855 );
buf ( n8857 , n8856 );
buf ( n8858 , n6196 );
buf ( n8859 , n6323 );
nor ( n8860 , n8858 , n8859 );
buf ( n8861 , n8860 );
nor ( n8862 , n6339 , n8861 );
buf ( n8863 , n8862 );
buf ( n8864 , n8863 );
buf ( n8865 , n8864 );
not ( n8866 , n8865 );
nand ( n8867 , n8866 , n6354 );
buf ( n8868 , n8867 );
nand ( n8869 , n5889 , n6887 , n8857 , n8868 );
buf ( n8870 , n8869 );
buf ( n8871 , n8870 );
buf ( n8872 , n8781 );
buf ( n8873 , n8785 );
nand ( n8874 , n8872 , n8873 );
buf ( n8875 , n8874 );
buf ( n8876 , n8875 );
not ( n8877 , n8753 );
not ( n8878 , n8759 );
and ( n8879 , n8877 , n8878 );
buf ( n8880 , n8730 );
buf ( n8881 , n8745 );
nor ( n8882 , n8880 , n8881 );
buf ( n8883 , n8882 );
nor ( n8884 , n8879 , n8883 );
buf ( n8885 , n8884 );
buf ( n8886 , n8777 );
and ( n8887 , n8876 , n8885 , n8886 );
buf ( n8888 , n8887 );
buf ( n8889 , n8888 );
not ( n8890 , n8889 );
buf ( n8891 , n8890 );
buf ( n8892 , n8891 );
not ( n8893 , n8892 );
buf ( n8894 , n8893 );
not ( n8895 , n7959 );
and ( n8896 , n5884 , n8894 , n6860 , n8895 );
buf ( n8897 , n8896 );
buf ( n8898 , n5177 );
buf ( n8899 , n8865 );
xor ( n8900 , n8429 , n8707 );
xor ( n8901 , n8900 , n8726 );
buf ( n8902 , n8901 );
buf ( n8903 , n8902 );
buf ( n8904 , n849 );
xor ( n8905 , n8607 , n8644 );
xor ( n8906 , n8905 , n8694 );
buf ( n8907 , n8906 );
buf ( n8908 , n8907 );
xor ( n8909 , n8612 , n8625 );
xor ( n8910 , n8909 , n8639 );
buf ( n8911 , n8910 );
buf ( n8912 , n8911 );
xor ( n8913 , n8658 , n8675 );
xor ( n8914 , n8913 , n8689 );
buf ( n8915 , n8914 );
buf ( n8916 , n8915 );
xor ( n8917 , n8912 , n8916 );
buf ( n8918 , n799 );
buf ( n8919 , n820 );
xor ( n8920 , n8918 , n8919 );
buf ( n8921 , n8920 );
buf ( n8922 , n8921 );
not ( n8923 , n8922 );
buf ( n8924 , n2410 );
not ( n8925 , n8924 );
or ( n8926 , n8923 , n8925 );
buf ( n8927 , n2672 );
buf ( n8928 , n8662 );
nand ( n8929 , n8927 , n8928 );
buf ( n8930 , n8929 );
buf ( n8931 , n8930 );
nand ( n8932 , n8926 , n8931 );
buf ( n8933 , n8932 );
buf ( n8934 , n8933 );
xor ( n8935 , n826 , n793 );
buf ( n8936 , n8935 );
not ( n8937 , n8936 );
buf ( n8938 , n8090 );
not ( n8939 , n8938 );
or ( n8940 , n8937 , n8939 );
buf ( n8941 , n1771 );
buf ( n8942 , n8450 );
nand ( n8943 , n8941 , n8942 );
buf ( n8944 , n8943 );
buf ( n8945 , n8944 );
nand ( n8946 , n8940 , n8945 );
buf ( n8947 , n8946 );
buf ( n8948 , n8947 );
xor ( n8949 , n8934 , n8948 );
buf ( n8950 , n8497 );
not ( n8951 , n8950 );
buf ( n8952 , n8480 );
not ( n8953 , n8952 );
or ( n8954 , n8951 , n8953 );
buf ( n8955 , n8480 );
buf ( n8956 , n8497 );
or ( n8957 , n8955 , n8956 );
nand ( n8958 , n8954 , n8957 );
buf ( n8959 , n8958 );
buf ( n8960 , n8959 );
and ( n8961 , n8949 , n8960 );
and ( n8962 , n8934 , n8948 );
or ( n8963 , n8961 , n8962 );
buf ( n8964 , n8963 );
buf ( n8965 , n8964 );
and ( n8966 , n8917 , n8965 );
and ( n8967 , n8912 , n8916 );
or ( n8968 , n8966 , n8967 );
buf ( n8969 , n8968 );
buf ( n8970 , n8969 );
xor ( n8971 , n8908 , n8970 );
xor ( n8972 , n8443 , n8445 );
xor ( n8973 , n8972 , n8575 );
buf ( n8974 , n8973 );
and ( n8975 , n8971 , n8974 );
and ( n8976 , n8908 , n8970 );
or ( n8977 , n8975 , n8976 );
buf ( n8978 , n8977 );
buf ( n8979 , n8978 );
xor ( n8980 , n8904 , n8979 );
xor ( n8981 , n8440 , n8579 );
xor ( n8982 , n8981 , n8702 );
buf ( n8983 , n8982 );
buf ( n8984 , n8983 );
and ( n8985 , n8980 , n8984 );
and ( n8986 , n8904 , n8979 );
or ( n8987 , n8985 , n8986 );
buf ( n8988 , n8987 );
buf ( n8989 , n8988 );
nor ( n8990 , n8903 , n8989 );
buf ( n8991 , n8990 );
buf ( n8992 , n8991 );
xor ( n8993 , n8904 , n8979 );
xor ( n8994 , n8993 , n8984 );
buf ( n8995 , n8994 );
buf ( n8996 , n8995 );
buf ( n8997 , n850 );
xor ( n8998 , n8463 , n8501 );
xor ( n8999 , n8998 , n8571 );
buf ( n9000 , n8999 );
buf ( n9001 , n9000 );
buf ( n9002 , n1346 );
buf ( n9003 , n799 );
and ( n9004 , n9002 , n9003 );
buf ( n9005 , n9004 );
buf ( n9006 , n9005 );
buf ( n9007 , n792 );
buf ( n9008 , n828 );
xor ( n9009 , n9007 , n9008 );
buf ( n9010 , n9009 );
buf ( n9011 , n9010 );
not ( n9012 , n9011 );
buf ( n9013 , n3680 );
not ( n9014 , n9013 );
or ( n9015 , n9012 , n9014 );
buf ( n9016 , n1249 );
buf ( n9017 , n8467 );
nand ( n9018 , n9016 , n9017 );
buf ( n9019 , n9018 );
buf ( n9020 , n9019 );
nand ( n9021 , n9015 , n9020 );
buf ( n9022 , n9021 );
buf ( n9023 , n9022 );
xor ( n9024 , n9006 , n9023 );
buf ( n9025 , n796 );
buf ( n9026 , n824 );
xor ( n9027 , n9025 , n9026 );
buf ( n9028 , n9027 );
buf ( n9029 , n9028 );
not ( n9030 , n9029 );
buf ( n9031 , n2790 );
not ( n9032 , n9031 );
or ( n9033 , n9030 , n9032 );
buf ( n9034 , n8354 );
buf ( n9035 , n8527 );
nand ( n9036 , n9034 , n9035 );
buf ( n9037 , n9036 );
buf ( n9038 , n9037 );
nand ( n9039 , n9033 , n9038 );
buf ( n9040 , n9039 );
buf ( n9041 , n9040 );
and ( n9042 , n9024 , n9041 );
and ( n9043 , n9006 , n9023 );
or ( n9044 , n9042 , n9043 );
buf ( n9045 , n9044 );
buf ( n9046 , n9045 );
buf ( n9047 , n790 );
buf ( n9048 , n830 );
xor ( n9049 , n9047 , n9048 );
buf ( n9050 , n9049 );
buf ( n9051 , n9050 );
not ( n9052 , n9051 );
buf ( n9053 , n1161 );
not ( n9054 , n9053 );
or ( n9055 , n9052 , n9054 );
buf ( n9056 , n8506 );
buf ( n9057 , n831 );
nand ( n9058 , n9056 , n9057 );
buf ( n9059 , n9058 );
buf ( n9060 , n9059 );
nand ( n9061 , n9055 , n9060 );
buf ( n9062 , n9061 );
buf ( n9063 , n9062 );
buf ( n9064 , n798 );
buf ( n9065 , n822 );
xor ( n9066 , n9064 , n9065 );
buf ( n9067 , n9066 );
buf ( n9068 , n9067 );
not ( n9069 , n9068 );
buf ( n9070 , n3739 );
not ( n9071 , n9070 );
or ( n9072 , n9069 , n9071 );
buf ( n9073 , n3745 );
buf ( n9074 , n8549 );
nand ( n9075 , n9073 , n9074 );
buf ( n9076 , n9075 );
buf ( n9077 , n9076 );
nand ( n9078 , n9072 , n9077 );
buf ( n9079 , n9078 );
buf ( n9080 , n9079 );
xor ( n9081 , n9063 , n9080 );
buf ( n9082 , n8935 );
not ( n9083 , n9082 );
buf ( n9084 , n1771 );
not ( n9085 , n9084 );
or ( n9086 , n9083 , n9085 );
buf ( n9087 , n1783 );
buf ( n9088 , n794 );
buf ( n9089 , n826 );
xor ( n9090 , n9088 , n9089 );
buf ( n9091 , n9090 );
buf ( n9092 , n9091 );
not ( n9093 , n9092 );
buf ( n9094 , n9093 );
buf ( n9095 , n9094 );
or ( n9096 , n9087 , n9095 );
nand ( n9097 , n9086 , n9096 );
buf ( n9098 , n9097 );
buf ( n9099 , n9098 );
and ( n9100 , n9081 , n9099 );
and ( n9101 , n9063 , n9080 );
or ( n9102 , n9100 , n9101 );
buf ( n9103 , n9102 );
buf ( n9104 , n9103 );
xor ( n9105 , n9046 , n9104 );
xor ( n9106 , n8523 , n8544 );
xor ( n9107 , n9106 , n8566 );
buf ( n9108 , n9107 );
buf ( n9109 , n9108 );
and ( n9110 , n9105 , n9109 );
and ( n9111 , n9046 , n9104 );
or ( n9112 , n9110 , n9111 );
buf ( n9113 , n9112 );
buf ( n9114 , n9113 );
xor ( n9115 , n9001 , n9114 );
xor ( n9116 , n8912 , n8916 );
xor ( n9117 , n9116 , n8965 );
buf ( n9118 , n9117 );
buf ( n9119 , n9118 );
and ( n9120 , n9115 , n9119 );
and ( n9121 , n9001 , n9114 );
or ( n9122 , n9120 , n9121 );
buf ( n9123 , n9122 );
buf ( n9124 , n9123 );
xor ( n9125 , n8997 , n9124 );
xor ( n9126 , n8908 , n8970 );
xor ( n9127 , n9126 , n8974 );
buf ( n9128 , n9127 );
buf ( n9129 , n9128 );
and ( n9130 , n9125 , n9129 );
and ( n9131 , n8997 , n9124 );
or ( n9132 , n9130 , n9131 );
buf ( n9133 , n9132 );
buf ( n9134 , n9133 );
nor ( n9135 , n8996 , n9134 );
buf ( n9136 , n9135 );
buf ( n9137 , n9136 );
nor ( n9138 , n8992 , n9137 );
buf ( n9139 , n9138 );
buf ( n9140 , n9139 );
xor ( n9141 , n8997 , n9124 );
xor ( n9142 , n9141 , n9129 );
buf ( n9143 , n9142 );
not ( n9144 , n9143 );
buf ( n9145 , n851 );
xor ( n9146 , n8934 , n8948 );
xor ( n9147 , n9146 , n8960 );
buf ( n9148 , n9147 );
buf ( n9149 , n9148 );
buf ( n9150 , n793 );
buf ( n9151 , n828 );
xor ( n9152 , n9150 , n9151 );
buf ( n9153 , n9152 );
buf ( n9154 , n9153 );
not ( n9155 , n9154 );
buf ( n9156 , n3680 );
not ( n9157 , n9156 );
or ( n9158 , n9155 , n9157 );
buf ( n9159 , n1249 );
buf ( n9160 , n9010 );
nand ( n9161 , n9159 , n9160 );
buf ( n9162 , n9161 );
buf ( n9163 , n9162 );
nand ( n9164 , n9158 , n9163 );
buf ( n9165 , n9164 );
buf ( n9166 , n9165 );
not ( n9167 , n9166 );
buf ( n9168 , n799 );
buf ( n9169 , n823 );
or ( n9170 , n9168 , n9169 );
buf ( n9171 , n824 );
nand ( n9172 , n9170 , n9171 );
buf ( n9173 , n9172 );
buf ( n9174 , n9173 );
buf ( n9175 , n799 );
buf ( n9176 , n823 );
nand ( n9177 , n9175 , n9176 );
buf ( n9178 , n9177 );
buf ( n9179 , n9178 );
buf ( n9180 , n822 );
nand ( n9181 , n9174 , n9179 , n9180 );
buf ( n9182 , n9181 );
buf ( n9183 , n9182 );
nor ( n9184 , n9167 , n9183 );
buf ( n9185 , n9184 );
buf ( n9186 , n9185 );
xor ( n9187 , n9006 , n9023 );
xor ( n9188 , n9187 , n9041 );
buf ( n9189 , n9188 );
buf ( n9190 , n9189 );
xor ( n9191 , n9186 , n9190 );
buf ( n9192 , n791 );
buf ( n9193 , n830 );
xor ( n9194 , n9192 , n9193 );
buf ( n9195 , n9194 );
buf ( n9196 , n9195 );
not ( n9197 , n9196 );
buf ( n9198 , n1161 );
not ( n9199 , n9198 );
or ( n9200 , n9197 , n9199 );
buf ( n9201 , n9050 );
buf ( n9202 , n831 );
nand ( n9203 , n9201 , n9202 );
buf ( n9204 , n9203 );
buf ( n9205 , n9204 );
nand ( n9206 , n9200 , n9205 );
buf ( n9207 , n9206 );
xor ( n9208 , n824 , n797 );
buf ( n9209 , n9208 );
not ( n9210 , n9209 );
buf ( n9211 , n2790 );
not ( n9212 , n9211 );
or ( n9213 , n9210 , n9212 );
buf ( n9214 , n1859 );
buf ( n9215 , n9028 );
nand ( n9216 , n9214 , n9215 );
buf ( n9217 , n9216 );
buf ( n9218 , n9217 );
nand ( n9219 , n9213 , n9218 );
buf ( n9220 , n9219 );
xor ( n9221 , n9207 , n9220 );
xor ( n9222 , n822 , n799 );
not ( n9223 , n9222 );
not ( n9224 , n3739 );
or ( n9225 , n9223 , n9224 );
buf ( n9226 , n3745 );
buf ( n9227 , n9067 );
nand ( n9228 , n9226 , n9227 );
buf ( n9229 , n9228 );
nand ( n9230 , n9225 , n9229 );
and ( n9231 , n9221 , n9230 );
and ( n9232 , n9207 , n9220 );
or ( n9233 , n9231 , n9232 );
buf ( n9234 , n9233 );
and ( n9235 , n9191 , n9234 );
and ( n9236 , n9186 , n9190 );
or ( n9237 , n9235 , n9236 );
buf ( n9238 , n9237 );
buf ( n9239 , n9238 );
xor ( n9240 , n9149 , n9239 );
xor ( n9241 , n9046 , n9104 );
xor ( n9242 , n9241 , n9109 );
buf ( n9243 , n9242 );
buf ( n9244 , n9243 );
and ( n9245 , n9240 , n9244 );
and ( n9246 , n9149 , n9239 );
or ( n9247 , n9245 , n9246 );
buf ( n9248 , n9247 );
buf ( n9249 , n9248 );
xor ( n9250 , n9145 , n9249 );
xor ( n9251 , n9001 , n9114 );
xor ( n9252 , n9251 , n9119 );
buf ( n9253 , n9252 );
buf ( n9254 , n9253 );
and ( n9255 , n9250 , n9254 );
and ( n9256 , n9145 , n9249 );
or ( n9257 , n9255 , n9256 );
buf ( n9258 , n9257 );
not ( n9259 , n9258 );
and ( n9260 , n9144 , n9259 );
xor ( n9261 , n9145 , n9249 );
xor ( n9262 , n9261 , n9254 );
buf ( n9263 , n9262 );
buf ( n9264 , n9263 );
buf ( n9265 , n852 );
xor ( n9266 , n9063 , n9080 );
xor ( n9267 , n9266 , n9099 );
buf ( n9268 , n9267 );
buf ( n9269 , n9268 );
buf ( n9270 , n795 );
buf ( n9271 , n826 );
xor ( n9272 , n9270 , n9271 );
buf ( n9273 , n9272 );
buf ( n9274 , n9273 );
not ( n9275 , n9274 );
buf ( n9276 , n8090 );
not ( n9277 , n9276 );
or ( n9278 , n9275 , n9277 );
buf ( n9279 , n1771 );
buf ( n9280 , n9091 );
nand ( n9281 , n9279 , n9280 );
buf ( n9282 , n9281 );
buf ( n9283 , n9282 );
nand ( n9284 , n9278 , n9283 );
buf ( n9285 , n9284 );
buf ( n9286 , n9285 );
buf ( n9287 , n2107 );
buf ( n9288 , n799 );
and ( n9289 , n9287 , n9288 );
buf ( n9290 , n9289 );
buf ( n9291 , n9290 );
buf ( n9292 , n792 );
buf ( n9293 , n830 );
xor ( n9294 , n9292 , n9293 );
buf ( n9295 , n9294 );
buf ( n9296 , n9295 );
not ( n9297 , n9296 );
buf ( n9298 , n1161 );
not ( n9299 , n9298 );
or ( n9300 , n9297 , n9299 );
buf ( n9301 , n9195 );
buf ( n9302 , n831 );
nand ( n9303 , n9301 , n9302 );
buf ( n9304 , n9303 );
buf ( n9305 , n9304 );
nand ( n9306 , n9300 , n9305 );
buf ( n9307 , n9306 );
buf ( n9308 , n9307 );
xor ( n9309 , n9291 , n9308 );
xor ( n9310 , n824 , n798 );
buf ( n9311 , n9310 );
not ( n9312 , n9311 );
buf ( n9313 , n2790 );
not ( n9314 , n9313 );
or ( n9315 , n9312 , n9314 );
buf ( n9316 , n8354 );
buf ( n9317 , n9208 );
nand ( n9318 , n9316 , n9317 );
buf ( n9319 , n9318 );
buf ( n9320 , n9319 );
nand ( n9321 , n9315 , n9320 );
buf ( n9322 , n9321 );
buf ( n9323 , n9322 );
and ( n9324 , n9309 , n9323 );
and ( n9325 , n9291 , n9308 );
or ( n9326 , n9324 , n9325 );
buf ( n9327 , n9326 );
buf ( n9328 , n9327 );
xor ( n9329 , n9286 , n9328 );
buf ( n9330 , n9182 );
not ( n9331 , n9330 );
buf ( n9332 , n9165 );
not ( n9333 , n9332 );
or ( n9334 , n9331 , n9333 );
buf ( n9335 , n9165 );
buf ( n9336 , n9182 );
or ( n9337 , n9335 , n9336 );
nand ( n9338 , n9334 , n9337 );
buf ( n9339 , n9338 );
buf ( n9340 , n9339 );
and ( n9341 , n9329 , n9340 );
and ( n9342 , n9286 , n9328 );
or ( n9343 , n9341 , n9342 );
buf ( n9344 , n9343 );
buf ( n9345 , n9344 );
xor ( n9346 , n9269 , n9345 );
xor ( n9347 , n9186 , n9190 );
xor ( n9348 , n9347 , n9234 );
buf ( n9349 , n9348 );
buf ( n9350 , n9349 );
and ( n9351 , n9346 , n9350 );
and ( n9352 , n9269 , n9345 );
or ( n9353 , n9351 , n9352 );
buf ( n9354 , n9353 );
buf ( n9355 , n9354 );
xor ( n9356 , n9265 , n9355 );
xor ( n9357 , n9149 , n9239 );
xor ( n9358 , n9357 , n9244 );
buf ( n9359 , n9358 );
buf ( n9360 , n9359 );
and ( n9361 , n9356 , n9360 );
and ( n9362 , n9265 , n9355 );
or ( n9363 , n9361 , n9362 );
buf ( n9364 , n9363 );
buf ( n9365 , n9364 );
nor ( n9366 , n9264 , n9365 );
buf ( n9367 , n9366 );
nor ( n9368 , n9260 , n9367 );
buf ( n9369 , n9368 );
and ( n9370 , n9140 , n9369 );
buf ( n9371 , n9370 );
buf ( n9372 , n9371 );
not ( n9373 , n9372 );
xor ( n9374 , n9265 , n9355 );
xor ( n9375 , n9374 , n9360 );
buf ( n9376 , n9375 );
buf ( n9377 , n9376 );
not ( n9378 , n9377 );
buf ( n9379 , n9378 );
buf ( n9380 , n9379 );
buf ( n9381 , n793 );
buf ( n9382 , n830 );
xor ( n9383 , n9381 , n9382 );
buf ( n9384 , n9383 );
buf ( n9385 , n9384 );
not ( n9386 , n9385 );
buf ( n9387 , n1161 );
not ( n9388 , n9387 );
or ( n9389 , n9386 , n9388 );
buf ( n9390 , n9295 );
buf ( n9391 , n831 );
nand ( n9392 , n9390 , n9391 );
buf ( n9393 , n9392 );
buf ( n9394 , n9393 );
nand ( n9395 , n9389 , n9394 );
buf ( n9396 , n9395 );
buf ( n9397 , n9396 );
buf ( n9398 , n799 );
buf ( n9399 , n825 );
or ( n9400 , n9398 , n9399 );
buf ( n9401 , n826 );
nand ( n9402 , n9400 , n9401 );
buf ( n9403 , n9402 );
buf ( n9404 , n9403 );
buf ( n9405 , n799 );
buf ( n9406 , n825 );
nand ( n9407 , n9405 , n9406 );
buf ( n9408 , n9407 );
buf ( n9409 , n9408 );
buf ( n9410 , n824 );
nand ( n9411 , n9404 , n9409 , n9410 );
buf ( n9412 , n9411 );
buf ( n9413 , n9412 );
not ( n9414 , n9413 );
buf ( n9415 , n9414 );
buf ( n9416 , n9415 );
nand ( n9417 , n9397 , n9416 );
buf ( n9418 , n9417 );
buf ( n9419 , n9418 );
not ( n9420 , n9419 );
buf ( n9421 , n796 );
buf ( n9422 , n826 );
xor ( n9423 , n9421 , n9422 );
buf ( n9424 , n9423 );
buf ( n9425 , n9424 );
not ( n9426 , n9425 );
buf ( n9427 , n1780 );
not ( n9428 , n9427 );
or ( n9429 , n9426 , n9428 );
buf ( n9430 , n1771 );
buf ( n9431 , n9273 );
nand ( n9432 , n9430 , n9431 );
buf ( n9433 , n9432 );
buf ( n9434 , n9433 );
nand ( n9435 , n9429 , n9434 );
buf ( n9436 , n9435 );
buf ( n9437 , n9436 );
not ( n9438 , n9437 );
buf ( n9439 , n9438 );
buf ( n9440 , n9439 );
not ( n9441 , n9440 );
or ( n9442 , n9420 , n9441 );
buf ( n9443 , n794 );
buf ( n9444 , n828 );
xor ( n9445 , n9443 , n9444 );
buf ( n9446 , n9445 );
buf ( n9447 , n9446 );
not ( n9448 , n9447 );
buf ( n9449 , n3680 );
not ( n9450 , n9449 );
or ( n9451 , n9448 , n9450 );
buf ( n9452 , n1249 );
not ( n9453 , n9452 );
buf ( n9454 , n9453 );
buf ( n9455 , n9454 );
not ( n9456 , n9455 );
buf ( n9457 , n9456 );
buf ( n9458 , n9457 );
buf ( n9459 , n9153 );
nand ( n9460 , n9458 , n9459 );
buf ( n9461 , n9460 );
buf ( n9462 , n9461 );
nand ( n9463 , n9451 , n9462 );
buf ( n9464 , n9463 );
buf ( n9465 , n9464 );
nand ( n9466 , n9442 , n9465 );
buf ( n9467 , n9466 );
buf ( n9468 , n9467 );
buf ( n9469 , n9418 );
not ( n9470 , n9469 );
buf ( n9471 , n9436 );
nand ( n9472 , n9470 , n9471 );
buf ( n9473 , n9472 );
buf ( n9474 , n9473 );
nand ( n9475 , n9468 , n9474 );
buf ( n9476 , n9475 );
buf ( n9477 , n9476 );
xor ( n9478 , n9207 , n9220 );
xor ( n9479 , n9478 , n9230 );
buf ( n9480 , n9479 );
xor ( n9481 , n9477 , n9480 );
xor ( n9482 , n9286 , n9328 );
xor ( n9483 , n9482 , n9340 );
buf ( n9484 , n9483 );
buf ( n9485 , n9484 );
and ( n9486 , n9481 , n9485 );
and ( n9487 , n9477 , n9480 );
or ( n9488 , n9486 , n9487 );
buf ( n9489 , n9488 );
buf ( n9490 , n9489 );
buf ( n9491 , n9490 );
buf ( n9492 , n9491 );
buf ( n9493 , n9492 );
not ( n9494 , n9493 );
xor ( n9495 , n9269 , n9345 );
xor ( n9496 , n9495 , n9350 );
buf ( n9497 , n9496 );
buf ( n9498 , n9497 );
buf ( n9499 , n9498 );
not ( n9500 , n9499 );
or ( n9501 , n9494 , n9500 );
buf ( n9502 , n9498 );
buf ( n9503 , n9492 );
or ( n9504 , n9502 , n9503 );
buf ( n9505 , n853 );
nand ( n9506 , n9504 , n9505 );
buf ( n9507 , n9506 );
buf ( n9508 , n9507 );
nand ( n9509 , n9501 , n9508 );
buf ( n9510 , n9509 );
buf ( n9511 , n9510 );
not ( n9512 , n9511 );
buf ( n9513 , n9512 );
buf ( n9514 , n9513 );
nand ( n9515 , n9380 , n9514 );
buf ( n9516 , n9515 );
buf ( n9517 , n9489 );
not ( n9518 , n9517 );
buf ( n9519 , n9518 );
and ( n9520 , n853 , n9519 );
not ( n9521 , n853 );
and ( n9522 , n9521 , n9489 );
or ( n9523 , n9520 , n9522 );
buf ( n9524 , n9523 );
buf ( n9525 , n9498 );
and ( n9526 , n9524 , n9525 );
not ( n9527 , n9524 );
buf ( n9528 , n9498 );
not ( n9529 , n9528 );
buf ( n9530 , n9529 );
buf ( n9531 , n9530 );
and ( n9532 , n9527 , n9531 );
nor ( n9533 , n9526 , n9532 );
buf ( n9534 , n9533 );
buf ( n9535 , n9534 );
not ( n9536 , n9535 );
buf ( n9537 , n9536 );
buf ( n9538 , n9537 );
buf ( n9539 , n854 );
xor ( n9540 , n9291 , n9308 );
xor ( n9541 , n9540 , n9323 );
buf ( n9542 , n9541 );
buf ( n9543 , n9542 );
buf ( n9544 , n797 );
buf ( n9545 , n826 );
xor ( n9546 , n9544 , n9545 );
buf ( n9547 , n9546 );
buf ( n9548 , n9547 );
not ( n9549 , n9548 );
buf ( n9550 , n1780 );
not ( n9551 , n9550 );
or ( n9552 , n9549 , n9551 );
buf ( n9553 , n1771 );
buf ( n9554 , n9424 );
nand ( n9555 , n9553 , n9554 );
buf ( n9556 , n9555 );
buf ( n9557 , n9556 );
nand ( n9558 , n9552 , n9557 );
buf ( n9559 , n9558 );
buf ( n9560 , n9559 );
xor ( n9561 , n824 , n799 );
buf ( n9562 , n9561 );
not ( n9563 , n9562 );
buf ( n9564 , n2790 );
not ( n9565 , n9564 );
or ( n9566 , n9563 , n9565 );
buf ( n9567 , n2492 );
buf ( n9568 , n9310 );
nand ( n9569 , n9567 , n9568 );
buf ( n9570 , n9569 );
buf ( n9571 , n9570 );
nand ( n9572 , n9566 , n9571 );
buf ( n9573 , n9572 );
buf ( n9574 , n9573 );
or ( n9575 , n9560 , n9574 );
buf ( n9576 , n795 );
buf ( n9577 , n828 );
xor ( n9578 , n9576 , n9577 );
buf ( n9579 , n9578 );
buf ( n9580 , n9579 );
not ( n9581 , n9580 );
buf ( n9582 , n3680 );
not ( n9583 , n9582 );
or ( n9584 , n9581 , n9583 );
buf ( n9585 , n9457 );
buf ( n9586 , n9446 );
nand ( n9587 , n9585 , n9586 );
buf ( n9588 , n9587 );
buf ( n9589 , n9588 );
nand ( n9590 , n9584 , n9589 );
buf ( n9591 , n9590 );
buf ( n9592 , n9591 );
nand ( n9593 , n9575 , n9592 );
buf ( n9594 , n9593 );
buf ( n9595 , n9594 );
buf ( n9596 , n9559 );
buf ( n9597 , n9573 );
nand ( n9598 , n9596 , n9597 );
buf ( n9599 , n9598 );
buf ( n9600 , n9599 );
nand ( n9601 , n9595 , n9600 );
buf ( n9602 , n9601 );
buf ( n9603 , n9602 );
xor ( n9604 , n9543 , n9603 );
xor ( n9605 , n9418 , n9436 );
buf ( n9606 , n9605 );
buf ( n9607 , n9464 );
xnor ( n9608 , n9606 , n9607 );
buf ( n9609 , n9608 );
buf ( n9610 , n9609 );
and ( n9611 , n9604 , n9610 );
and ( n9612 , n9543 , n9603 );
or ( n9613 , n9611 , n9612 );
buf ( n9614 , n9613 );
buf ( n9615 , n9614 );
xor ( n9616 , n9539 , n9615 );
xor ( n9617 , n9477 , n9480 );
xor ( n9618 , n9617 , n9485 );
buf ( n9619 , n9618 );
buf ( n9620 , n9619 );
and ( n9621 , n9616 , n9620 );
and ( n9622 , n9539 , n9615 );
or ( n9623 , n9621 , n9622 );
buf ( n9624 , n9623 );
buf ( n9625 , n9624 );
not ( n9626 , n9625 );
buf ( n9627 , n9626 );
buf ( n9628 , n9627 );
nand ( n9629 , n9538 , n9628 );
buf ( n9630 , n9629 );
buf ( n9631 , n855 );
buf ( n9632 , n9396 );
buf ( n9633 , n9415 );
and ( n9634 , n9632 , n9633 );
not ( n9635 , n9632 );
buf ( n9636 , n9412 );
and ( n9637 , n9635 , n9636 );
nor ( n9638 , n9634 , n9637 );
buf ( n9639 , n9638 );
buf ( n9640 , n9639 );
not ( n9641 , n9640 );
buf ( n9642 , n9641 );
buf ( n9643 , n8354 );
buf ( n9644 , n799 );
nand ( n9645 , n9643 , n9644 );
buf ( n9646 , n9645 );
buf ( n9647 , n9646 );
not ( n9648 , n9647 );
buf ( n9649 , n9648 );
buf ( n9650 , n9649 );
not ( n9651 , n9650 );
buf ( n9652 , n794 );
buf ( n9653 , n830 );
xor ( n9654 , n9652 , n9653 );
buf ( n9655 , n9654 );
buf ( n9656 , n9655 );
not ( n9657 , n9656 );
buf ( n9658 , n1161 );
not ( n9659 , n9658 );
or ( n9660 , n9657 , n9659 );
buf ( n9661 , n9384 );
buf ( n9662 , n831 );
nand ( n9663 , n9661 , n9662 );
buf ( n9664 , n9663 );
buf ( n9665 , n9664 );
nand ( n9666 , n9660 , n9665 );
buf ( n9667 , n9666 );
buf ( n9668 , n9667 );
not ( n9669 , n9668 );
or ( n9670 , n9651 , n9669 );
buf ( n9671 , n9646 );
not ( n9672 , n9671 );
buf ( n9673 , n9667 );
not ( n9674 , n9673 );
buf ( n9675 , n9674 );
buf ( n9676 , n9675 );
not ( n9677 , n9676 );
or ( n9678 , n9672 , n9677 );
buf ( n9679 , n796 );
buf ( n9680 , n828 );
xor ( n9681 , n9679 , n9680 );
buf ( n9682 , n9681 );
buf ( n9683 , n9682 );
not ( n9684 , n9683 );
buf ( n9685 , n3680 );
not ( n9686 , n9685 );
or ( n9687 , n9684 , n9686 );
buf ( n9688 , n9579 );
buf ( n9689 , n1249 );
nand ( n9690 , n9688 , n9689 );
buf ( n9691 , n9690 );
buf ( n9692 , n9691 );
nand ( n9693 , n9687 , n9692 );
buf ( n9694 , n9693 );
buf ( n9695 , n9694 );
nand ( n9696 , n9678 , n9695 );
buf ( n9697 , n9696 );
buf ( n9698 , n9697 );
nand ( n9699 , n9670 , n9698 );
buf ( n9700 , n9699 );
not ( n9701 , n9700 );
and ( n9702 , n9642 , n9701 );
not ( n9703 , n9702 );
buf ( n9704 , n9703 );
not ( n9705 , n9704 );
xor ( n9706 , n9559 , n9573 );
xnor ( n9707 , n9706 , n9591 );
buf ( n9708 , n9707 );
not ( n9709 , n9708 );
buf ( n9710 , n9709 );
buf ( n9711 , n9710 );
not ( n9712 , n9711 );
or ( n9713 , n9705 , n9712 );
buf ( n9714 , n9700 );
buf ( n9715 , n9639 );
nand ( n9716 , n9714 , n9715 );
buf ( n9717 , n9716 );
buf ( n9718 , n9717 );
nand ( n9719 , n9713 , n9718 );
buf ( n9720 , n9719 );
buf ( n9721 , n9720 );
xor ( n9722 , n9631 , n9721 );
xor ( n9723 , n9543 , n9603 );
xor ( n9724 , n9723 , n9610 );
buf ( n9725 , n9724 );
buf ( n9726 , n9725 );
and ( n9727 , n9722 , n9726 );
and ( n9728 , n9631 , n9721 );
or ( n9729 , n9727 , n9728 );
buf ( n9730 , n9729 );
buf ( n9731 , n9730 );
xor ( n9732 , n9539 , n9615 );
xor ( n9733 , n9732 , n9620 );
buf ( n9734 , n9733 );
buf ( n9735 , n9734 );
nor ( n9736 , n9731 , n9735 );
buf ( n9737 , n9736 );
buf ( n9738 , n9737 );
xor ( n9739 , n9631 , n9721 );
xor ( n9740 , n9739 , n9726 );
buf ( n9741 , n9740 );
buf ( n9742 , n9741 );
buf ( n9743 , n799 );
buf ( n9744 , n827 );
or ( n9745 , n9743 , n9744 );
buf ( n9746 , n828 );
nand ( n9747 , n9745 , n9746 );
buf ( n9748 , n9747 );
buf ( n9749 , n9748 );
buf ( n9750 , n799 );
buf ( n9751 , n827 );
nand ( n9752 , n9750 , n9751 );
buf ( n9753 , n9752 );
buf ( n9754 , n9753 );
buf ( n9755 , n826 );
and ( n9756 , n9749 , n9754 , n9755 );
buf ( n9757 , n9756 );
buf ( n9758 , n9757 );
buf ( n9759 , n795 );
buf ( n9760 , n830 );
xor ( n9761 , n9759 , n9760 );
buf ( n9762 , n9761 );
buf ( n9763 , n9762 );
not ( n9764 , n9763 );
buf ( n9765 , n1161 );
not ( n9766 , n9765 );
or ( n9767 , n9764 , n9766 );
buf ( n9768 , n9655 );
buf ( n9769 , n831 );
nand ( n9770 , n9768 , n9769 );
buf ( n9771 , n9770 );
buf ( n9772 , n9771 );
nand ( n9773 , n9767 , n9772 );
buf ( n9774 , n9773 );
buf ( n9775 , n9774 );
and ( n9776 , n9758 , n9775 );
buf ( n9777 , n9776 );
buf ( n9778 , n798 );
buf ( n9779 , n826 );
xor ( n9780 , n9778 , n9779 );
buf ( n9781 , n9780 );
buf ( n9782 , n9781 );
not ( n9783 , n9782 );
buf ( n9784 , n8090 );
not ( n9785 , n9784 );
or ( n9786 , n9783 , n9785 );
buf ( n9787 , n1771 );
buf ( n9788 , n9547 );
nand ( n9789 , n9787 , n9788 );
buf ( n9790 , n9789 );
buf ( n9791 , n9790 );
nand ( n9792 , n9786 , n9791 );
buf ( n9793 , n9792 );
xor ( n9794 , n9777 , n9793 );
xor ( n9795 , n9646 , n9667 );
xnor ( n9796 , n9795 , n9694 );
and ( n9797 , n9794 , n9796 );
and ( n9798 , n9777 , n9793 );
or ( n9799 , n9797 , n9798 );
buf ( n9800 , n9799 );
buf ( n9801 , n9800 );
buf ( n9802 , n9801 );
buf ( n9803 , n9802 );
not ( n9804 , n9803 );
not ( n9805 , n9700 );
xor ( n9806 , n9642 , n9805 );
buf ( n9807 , n9806 );
not ( n9808 , n9807 );
buf ( n9809 , n9808 );
buf ( n9810 , n9809 );
not ( n9811 , n9810 );
buf ( n9812 , n9710 );
not ( n9813 , n9812 );
or ( n9814 , n9811 , n9813 );
buf ( n9815 , n9806 );
buf ( n9816 , n9707 );
nand ( n9817 , n9815 , n9816 );
buf ( n9818 , n9817 );
buf ( n9819 , n9818 );
nand ( n9820 , n9814 , n9819 );
buf ( n9821 , n9820 );
buf ( n9822 , n9821 );
buf ( n9823 , n9822 );
buf ( n9824 , n9823 );
buf ( n9825 , n9824 );
buf ( n9826 , n9825 );
not ( n9827 , n9826 );
or ( n9828 , n9804 , n9827 );
buf ( n9829 , n9825 );
buf ( n9830 , n9802 );
or ( n9831 , n9829 , n9830 );
buf ( n9832 , n856 );
nand ( n9833 , n9831 , n9832 );
buf ( n9834 , n9833 );
buf ( n9835 , n9834 );
nand ( n9836 , n9828 , n9835 );
buf ( n9837 , n9836 );
buf ( n9838 , n9837 );
nor ( n9839 , n9742 , n9838 );
buf ( n9840 , n9839 );
buf ( n9841 , n9840 );
nor ( n9842 , n9738 , n9841 );
buf ( n9843 , n9842 );
and ( n9844 , n9516 , n9630 , n9843 );
buf ( n9845 , n856 );
not ( n9846 , n9845 );
buf ( n9847 , n9799 );
not ( n9848 , n9847 );
buf ( n9849 , n9848 );
buf ( n9850 , n9849 );
not ( n9851 , n9850 );
or ( n9852 , n9846 , n9851 );
not ( n9853 , n856 );
nand ( n9854 , n9853 , n9799 );
buf ( n9855 , n9854 );
nand ( n9856 , n9852 , n9855 );
buf ( n9857 , n9856 );
buf ( n9858 , n9857 );
buf ( n9859 , n9822 );
and ( n9860 , n9858 , n9859 );
not ( n9861 , n9858 );
buf ( n9862 , n9822 );
not ( n9863 , n9862 );
buf ( n9864 , n9863 );
buf ( n9865 , n9864 );
and ( n9866 , n9861 , n9865 );
nor ( n9867 , n9860 , n9866 );
buf ( n9868 , n9867 );
buf ( n9869 , n9868 );
buf ( n9870 , n857 );
buf ( n9871 , n797 );
buf ( n9872 , n828 );
xor ( n9873 , n9871 , n9872 );
buf ( n9874 , n9873 );
buf ( n9875 , n9874 );
not ( n9876 , n9875 );
buf ( n9877 , n3680 );
not ( n9878 , n9877 );
or ( n9879 , n9876 , n9878 );
buf ( n9880 , n1249 );
buf ( n9881 , n9682 );
nand ( n9882 , n9880 , n9881 );
buf ( n9883 , n9882 );
buf ( n9884 , n9883 );
nand ( n9885 , n9879 , n9884 );
buf ( n9886 , n9885 );
buf ( n9887 , n9886 );
xor ( n9888 , n9758 , n9775 );
buf ( n9889 , n9888 );
buf ( n9890 , n9889 );
xor ( n9891 , n9887 , n9890 );
buf ( n9892 , n826 );
buf ( n9893 , n799 );
xor ( n9894 , n9892 , n9893 );
buf ( n9895 , n9894 );
buf ( n9896 , n9895 );
not ( n9897 , n9896 );
buf ( n9898 , n8090 );
not ( n9899 , n9898 );
or ( n9900 , n9897 , n9899 );
buf ( n9901 , n1771 );
buf ( n9902 , n9781 );
nand ( n9903 , n9901 , n9902 );
buf ( n9904 , n9903 );
buf ( n9905 , n9904 );
nand ( n9906 , n9900 , n9905 );
buf ( n9907 , n9906 );
buf ( n9908 , n9907 );
and ( n9909 , n9891 , n9908 );
and ( n9910 , n9887 , n9890 );
or ( n9911 , n9909 , n9910 );
buf ( n9912 , n9911 );
buf ( n9913 , n9912 );
xor ( n9914 , n9870 , n9913 );
xor ( n9915 , n9777 , n9793 );
xor ( n9916 , n9915 , n9796 );
buf ( n9917 , n9916 );
and ( n9918 , n9914 , n9917 );
and ( n9919 , n9870 , n9913 );
or ( n9920 , n9918 , n9919 );
buf ( n9921 , n9920 );
buf ( n9922 , n9921 );
or ( n9923 , n9869 , n9922 );
buf ( n9924 , n9923 );
buf ( n9925 , n9924 );
xor ( n9926 , n9870 , n9913 );
xor ( n9927 , n9926 , n9917 );
buf ( n9928 , n9927 );
buf ( n9929 , n9928 );
buf ( n9930 , n858 );
buf ( n9931 , n796 );
buf ( n9932 , n830 );
xor ( n9933 , n9931 , n9932 );
buf ( n9934 , n9933 );
buf ( n9935 , n9934 );
not ( n9936 , n9935 );
buf ( n9937 , n1161 );
not ( n9938 , n9937 );
or ( n9939 , n9936 , n9938 );
buf ( n9940 , n9762 );
buf ( n9941 , n831 );
nand ( n9942 , n9940 , n9941 );
buf ( n9943 , n9942 );
buf ( n9944 , n9943 );
nand ( n9945 , n9939 , n9944 );
buf ( n9946 , n9945 );
not ( n9947 , n9946 );
buf ( n9948 , n799 );
buf ( n9949 , n1771 );
nand ( n9950 , n9948 , n9949 );
buf ( n9951 , n9950 );
buf ( n9952 , n9951 );
not ( n9953 , n9952 );
buf ( n9954 , n9953 );
not ( n9955 , n9954 );
or ( n9956 , n9947 , n9955 );
buf ( n9957 , n9951 );
not ( n9958 , n9957 );
buf ( n9959 , n9946 );
not ( n9960 , n9959 );
buf ( n9961 , n9960 );
buf ( n9962 , n9961 );
not ( n9963 , n9962 );
or ( n9964 , n9958 , n9963 );
buf ( n9965 , n798 );
buf ( n9966 , n828 );
xor ( n9967 , n9965 , n9966 );
buf ( n9968 , n9967 );
buf ( n9969 , n9968 );
not ( n9970 , n9969 );
buf ( n9971 , n3680 );
not ( n9972 , n9971 );
or ( n9973 , n9970 , n9972 );
buf ( n9974 , n1249 );
buf ( n9975 , n9874 );
nand ( n9976 , n9974 , n9975 );
buf ( n9977 , n9976 );
buf ( n9978 , n9977 );
nand ( n9979 , n9973 , n9978 );
buf ( n9980 , n9979 );
buf ( n9981 , n9980 );
nand ( n9982 , n9964 , n9981 );
buf ( n9983 , n9982 );
nand ( n9984 , n9956 , n9983 );
buf ( n9985 , n9984 );
xor ( n9986 , n9930 , n9985 );
xor ( n9987 , n9887 , n9890 );
xor ( n9988 , n9987 , n9908 );
buf ( n9989 , n9988 );
buf ( n9990 , n9989 );
and ( n9991 , n9986 , n9990 );
and ( n9992 , n9930 , n9985 );
or ( n9993 , n9991 , n9992 );
buf ( n9994 , n9993 );
buf ( n9995 , n9994 );
nand ( n9996 , n9929 , n9995 );
buf ( n9997 , n9996 );
buf ( n9998 , n9997 );
not ( n9999 , n9998 );
buf ( n10000 , n9999 );
buf ( n10001 , n10000 );
and ( n10002 , n9925 , n10001 );
buf ( n10003 , n9868 );
buf ( n10004 , n9921 );
and ( n10005 , n10003 , n10004 );
buf ( n10006 , n10005 );
buf ( n10007 , n10006 );
nor ( n10008 , n10002 , n10007 );
buf ( n10009 , n10008 );
buf ( n10010 , n10009 );
buf ( n10011 , n9924 );
buf ( n10012 , n859 );
buf ( n10013 , n1161 );
not ( n10014 , n10013 );
buf ( n10015 , n797 );
buf ( n10016 , n830 );
xor ( n10017 , n10015 , n10016 );
buf ( n10018 , n10017 );
buf ( n10019 , n10018 );
not ( n10020 , n10019 );
or ( n10021 , n10014 , n10020 );
buf ( n10022 , n9934 );
buf ( n10023 , n831 );
nand ( n10024 , n10022 , n10023 );
buf ( n10025 , n10024 );
buf ( n10026 , n10025 );
nand ( n10027 , n10021 , n10026 );
buf ( n10028 , n10027 );
buf ( n10029 , n10028 );
buf ( n10030 , n799 );
buf ( n10031 , n829 );
or ( n10032 , n10030 , n10031 );
buf ( n10033 , n830 );
nand ( n10034 , n10032 , n10033 );
buf ( n10035 , n10034 );
buf ( n10036 , n10035 );
buf ( n10037 , n799 );
buf ( n10038 , n829 );
nand ( n10039 , n10037 , n10038 );
buf ( n10040 , n10039 );
buf ( n10041 , n10040 );
buf ( n10042 , n828 );
nand ( n10043 , n10036 , n10041 , n10042 );
buf ( n10044 , n10043 );
buf ( n10045 , n10044 );
not ( n10046 , n10045 );
buf ( n10047 , n10046 );
buf ( n10048 , n10047 );
and ( n10049 , n10029 , n10048 );
buf ( n10050 , n10049 );
buf ( n10051 , n10050 );
xor ( n10052 , n10012 , n10051 );
xor ( n10053 , n9954 , n9961 );
xnor ( n10054 , n10053 , n9980 );
buf ( n10055 , n10054 );
and ( n10056 , n10052 , n10055 );
and ( n10057 , n10012 , n10051 );
or ( n10058 , n10056 , n10057 );
buf ( n10059 , n10058 );
buf ( n10060 , n10059 );
xor ( n10061 , n9930 , n9985 );
xor ( n10062 , n10061 , n9990 );
buf ( n10063 , n10062 );
buf ( n10064 , n10063 );
nor ( n10065 , n10060 , n10064 );
buf ( n10066 , n10065 );
buf ( n10067 , n10066 );
xor ( n10068 , n10012 , n10051 );
xor ( n10069 , n10068 , n10055 );
buf ( n10070 , n10069 );
buf ( n10071 , n10070 );
buf ( n10072 , n860 );
buf ( n10073 , n799 );
buf ( n10074 , n828 );
xor ( n10075 , n10073 , n10074 );
buf ( n10076 , n10075 );
buf ( n10077 , n10076 );
not ( n10078 , n10077 );
buf ( n10079 , n3680 );
not ( n10080 , n10079 );
or ( n10081 , n10078 , n10080 );
buf ( n10082 , n1249 );
buf ( n10083 , n9968 );
nand ( n10084 , n10082 , n10083 );
buf ( n10085 , n10084 );
buf ( n10086 , n10085 );
nand ( n10087 , n10081 , n10086 );
buf ( n10088 , n10087 );
buf ( n10089 , n10088 );
xor ( n10090 , n10072 , n10089 );
buf ( n10091 , n10044 );
not ( n10092 , n10091 );
buf ( n10093 , n10028 );
not ( n10094 , n10093 );
or ( n10095 , n10092 , n10094 );
buf ( n10096 , n6372 );
buf ( n10097 , n10096 );
buf ( n10098 , n10018 );
not ( n10099 , n10098 );
buf ( n10100 , n10099 );
buf ( n10101 , n10100 );
or ( n10102 , n10097 , n10101 );
not ( n10103 , n831 );
buf ( n10104 , n10103 );
buf ( n10105 , n9934 );
not ( n10106 , n10105 );
buf ( n10107 , n10106 );
buf ( n10108 , n10107 );
or ( n10109 , n10104 , n10108 );
buf ( n10110 , n10047 );
nand ( n10111 , n10102 , n10109 , n10110 );
buf ( n10112 , n10111 );
buf ( n10113 , n10112 );
nand ( n10114 , n10095 , n10113 );
buf ( n10115 , n10114 );
buf ( n10116 , n10115 );
and ( n10117 , n10090 , n10116 );
and ( n10118 , n10072 , n10089 );
or ( n10119 , n10117 , n10118 );
buf ( n10120 , n10119 );
buf ( n10121 , n10120 );
nand ( n10122 , n10071 , n10121 );
buf ( n10123 , n10122 );
buf ( n10124 , n10123 );
or ( n10125 , n10067 , n10124 );
buf ( n10126 , n10063 );
buf ( n10127 , n10126 );
buf ( n10128 , n10127 );
buf ( n10129 , n10128 );
buf ( n10130 , n10059 );
nand ( n10131 , n10129 , n10130 );
buf ( n10132 , n10131 );
buf ( n10133 , n10132 );
nand ( n10134 , n10125 , n10133 );
buf ( n10135 , n10134 );
buf ( n10136 , n10135 );
buf ( n10137 , n9928 );
buf ( n10138 , n9994 );
nor ( n10139 , n10137 , n10138 );
buf ( n10140 , n10139 );
buf ( n10141 , n10140 );
not ( n10142 , n10141 );
buf ( n10143 , n10142 );
buf ( n10144 , n10143 );
nand ( n10145 , n10011 , n10136 , n10144 );
buf ( n10146 , n10145 );
buf ( n10147 , n10146 );
buf ( n10148 , n9924 );
buf ( n10149 , n10063 );
buf ( n10150 , n10059 );
nor ( n10151 , n10149 , n10150 );
buf ( n10152 , n10151 );
buf ( n10153 , n10152 );
buf ( n10154 , n10070 );
buf ( n10155 , n10120 );
nor ( n10156 , n10154 , n10155 );
buf ( n10157 , n10156 );
buf ( n10158 , n10157 );
nor ( n10159 , n10153 , n10158 );
buf ( n10160 , n10159 );
buf ( n10161 , n10160 );
buf ( n10162 , n861 );
buf ( n10163 , n1168 );
not ( n10164 , n10163 );
buf ( n10165 , n1161 );
not ( n10166 , n10165 );
or ( n10167 , n10164 , n10166 );
buf ( n10168 , n831 );
buf ( n10169 , n10018 );
nand ( n10170 , n10168 , n10169 );
buf ( n10171 , n10170 );
buf ( n10172 , n10171 );
nand ( n10173 , n10167 , n10172 );
buf ( n10174 , n10173 );
buf ( n10175 , n10174 );
xor ( n10176 , n10162 , n10175 );
buf ( n10177 , n9457 );
buf ( n10178 , n799 );
and ( n10179 , n10177 , n10178 );
buf ( n10180 , n10179 );
buf ( n10181 , n10180 );
xor ( n10182 , n10176 , n10181 );
buf ( n10183 , n10182 );
buf ( n10184 , n10183 );
and ( n10185 , n1202 , n1203 );
buf ( n10186 , n10185 );
buf ( n10187 , n10186 );
nor ( n10188 , n10184 , n10187 );
buf ( n10189 , n10188 );
buf ( n10190 , n10189 );
buf ( n10191 , n1175 );
not ( n10192 , n10191 );
buf ( n10193 , n1208 );
nand ( n10194 , n10192 , n10193 );
buf ( n10195 , n10194 );
buf ( n10196 , n1201 );
not ( n10197 , n10196 );
buf ( n10198 , n10197 );
and ( n10199 , n10195 , n10198 );
and ( n10200 , n1175 , n1205 );
nor ( n10201 , n10199 , n10200 );
buf ( n10202 , n10201 );
nor ( n10203 , n10190 , n10202 );
buf ( n10204 , n10203 );
buf ( n10205 , n10204 );
not ( n10206 , n10205 );
buf ( n10207 , n10183 );
buf ( n10208 , n10186 );
nand ( n10209 , n10207 , n10208 );
buf ( n10210 , n10209 );
buf ( n10211 , n10210 );
nand ( n10212 , n10206 , n10211 );
buf ( n10213 , n10212 );
not ( n10214 , n10213 );
xor ( n10215 , n10072 , n10089 );
xor ( n10216 , n10215 , n10116 );
buf ( n10217 , n10216 );
buf ( n10218 , n10217 );
xor ( n10219 , n10162 , n10175 );
and ( n10220 , n10219 , n10181 );
and ( n10221 , n10162 , n10175 );
or ( n10222 , n10220 , n10221 );
buf ( n10223 , n10222 );
buf ( n10224 , n10223 );
nor ( n10225 , n10218 , n10224 );
buf ( n10226 , n10225 );
buf ( n10227 , n10226 );
not ( n10228 , n10227 );
buf ( n10229 , n10228 );
not ( n10230 , n10229 );
or ( n10231 , n10214 , n10230 );
buf ( n10232 , n10217 );
buf ( n10233 , n10232 );
buf ( n10234 , n10233 );
buf ( n10235 , n10234 );
buf ( n10236 , n10223 );
nand ( n10237 , n10235 , n10236 );
buf ( n10238 , n10237 );
nand ( n10239 , n10231 , n10238 );
buf ( n10240 , n10239 );
and ( n10241 , n10161 , n10240 );
buf ( n10242 , n10241 );
buf ( n10243 , n10242 );
buf ( n10244 , n10143 );
nand ( n10245 , n10148 , n10243 , n10244 );
buf ( n10246 , n10245 );
buf ( n10247 , n10246 );
nand ( n10248 , n10010 , n10147 , n10247 );
buf ( n10249 , n10248 );
buf ( n10250 , n10249 );
not ( n10251 , n10250 );
buf ( n10252 , n10251 );
buf ( n10253 , n10252 );
not ( n10254 , n10253 );
buf ( n10255 , n10254 );
nand ( n10256 , n9844 , n10255 );
buf ( n10257 , n9737 );
buf ( n10258 , n9741 );
buf ( n10259 , n9837 );
nand ( n10260 , n10258 , n10259 );
buf ( n10261 , n10260 );
buf ( n10262 , n10261 );
or ( n10263 , n10257 , n10262 );
buf ( n10264 , n9734 );
buf ( n10265 , n9730 );
nand ( n10266 , n10264 , n10265 );
buf ( n10267 , n10266 );
buf ( n10268 , n10267 );
nand ( n10269 , n10263 , n10268 );
buf ( n10270 , n10269 );
buf ( n10271 , n10270 );
not ( n10272 , n10271 );
not ( n10273 , n9376 );
not ( n10274 , n9510 );
and ( n10275 , n10273 , n10274 );
buf ( n10276 , n9534 );
buf ( n10277 , n9624 );
nor ( n10278 , n10276 , n10277 );
buf ( n10279 , n10278 );
nor ( n10280 , n10275 , n10279 );
buf ( n10281 , n10280 );
not ( n10282 , n10281 );
or ( n10283 , n10272 , n10282 );
buf ( n10284 , n9516 );
buf ( n10285 , n9534 );
buf ( n10286 , n9624 );
nand ( n10287 , n10285 , n10286 );
buf ( n10288 , n10287 );
buf ( n10289 , n10288 );
not ( n10290 , n10289 );
buf ( n10291 , n10290 );
buf ( n10292 , n10291 );
and ( n10293 , n10284 , n10292 );
buf ( n10294 , n9379 );
buf ( n10295 , n9513 );
nor ( n10296 , n10294 , n10295 );
buf ( n10297 , n10296 );
buf ( n10298 , n10297 );
nor ( n10299 , n10293 , n10298 );
buf ( n10300 , n10299 );
buf ( n10301 , n10300 );
nand ( n10302 , n10283 , n10301 );
buf ( n10303 , n10302 );
buf ( n10304 , n10303 );
not ( n10305 , n10304 );
buf ( n10306 , n10305 );
nand ( n10307 , n10256 , n10306 );
buf ( n10308 , n10307 );
not ( n10309 , n10308 );
or ( n10310 , n9373 , n10309 );
buf ( n10311 , n9143 );
buf ( n10312 , n9258 );
nor ( n10313 , n10311 , n10312 );
buf ( n10314 , n10313 );
buf ( n10315 , n10314 );
buf ( n10316 , n9263 );
buf ( n10317 , n9364 );
nand ( n10318 , n10316 , n10317 );
buf ( n10319 , n10318 );
buf ( n10320 , n10319 );
or ( n10321 , n10315 , n10320 );
buf ( n10322 , n9143 );
buf ( n10323 , n9258 );
nand ( n10324 , n10322 , n10323 );
buf ( n10325 , n10324 );
buf ( n10326 , n10325 );
nand ( n10327 , n10321 , n10326 );
buf ( n10328 , n10327 );
not ( n10329 , n10328 );
not ( n10330 , n9139 );
or ( n10331 , n10329 , n10330 );
buf ( n10332 , n8995 );
buf ( n10333 , n9133 );
and ( n10334 , n10332 , n10333 );
buf ( n10335 , n10334 );
buf ( n10336 , n10335 );
buf ( n10337 , n8988 );
not ( n10338 , n10337 );
buf ( n10339 , n8902 );
not ( n10340 , n10339 );
buf ( n10341 , n10340 );
buf ( n10342 , n10341 );
nand ( n10343 , n10338 , n10342 );
buf ( n10344 , n10343 );
buf ( n10345 , n10344 );
and ( n10346 , n10336 , n10345 );
buf ( n10347 , n8988 );
not ( n10348 , n10347 );
buf ( n10349 , n10341 );
nor ( n10350 , n10348 , n10349 );
buf ( n10351 , n10350 );
buf ( n10352 , n10351 );
nor ( n10353 , n10346 , n10352 );
buf ( n10354 , n10353 );
nand ( n10355 , n10331 , n10354 );
not ( n10356 , n10355 );
buf ( n10357 , n10356 );
nand ( n10358 , n10310 , n10357 );
buf ( n10359 , n10358 );
buf ( n10360 , n10359 );
and ( n10361 , n8898 , n8899 , n10360 );
buf ( n10362 , n10361 );
buf ( n10363 , n10362 );
and ( n10364 , n8897 , n10363 );
buf ( n10365 , n5870 );
not ( n10366 , n10365 );
buf ( n10367 , n5877 );
nor ( n10368 , n10366 , n10367 );
buf ( n10369 , n10368 );
buf ( n10370 , n10369 );
not ( n10371 , n10370 );
buf ( n10372 , n5503 );
not ( n10373 , n10372 );
or ( n10374 , n10371 , n10373 );
buf ( n10375 , n5497 );
buf ( n10376 , n5181 );
nand ( n10377 , n10375 , n10376 );
buf ( n10378 , n10377 );
buf ( n10379 , n10378 );
nand ( n10380 , n10374 , n10379 );
buf ( n10381 , n10380 );
buf ( n10382 , n10381 );
not ( n10383 , n10382 );
buf ( n10384 , n5177 );
not ( n10385 , n10384 );
or ( n10386 , n10383 , n10385 );
not ( n10387 , n4847 );
not ( n10388 , n4360 );
nand ( n10389 , n10387 , n10388 );
buf ( n10390 , n4852 );
buf ( n10391 , n5173 );
nand ( n10392 , n10390 , n10391 );
buf ( n10393 , n10392 );
buf ( n10394 , n10393 );
not ( n10395 , n10394 );
buf ( n10396 , n10395 );
and ( n10397 , n10389 , n10396 );
buf ( n10398 , n4360 );
buf ( n10399 , n4847 );
nand ( n10400 , n10398 , n10399 );
buf ( n10401 , n10400 );
buf ( n10402 , n10401 );
not ( n10403 , n10402 );
buf ( n10404 , n10403 );
nor ( n10405 , n10397 , n10404 );
buf ( n10406 , n10405 );
nand ( n10407 , n10386 , n10406 );
buf ( n10408 , n10407 );
buf ( n10409 , n10408 );
nor ( n10410 , n10364 , n10409 );
buf ( n10411 , n10410 );
buf ( n10412 , n10411 );
nand ( n10413 , n8871 , n10412 );
buf ( n10414 , n10413 );
buf ( n10415 , n10414 );
buf ( n10416 , n10415 );
buf ( n10417 , n10416 );
buf ( n10418 , n10417 );
not ( n10419 , n10418 );
or ( n10420 , n4357 , n10419 );
buf ( n10421 , n8870 );
buf ( n10422 , n10411 );
nand ( n10423 , n10421 , n10422 );
buf ( n10424 , n10423 );
buf ( n10425 , n10424 );
buf ( n10426 , n10425 );
buf ( n10427 , n10426 );
buf ( n10428 , n10427 );
buf ( n10429 , n10428 );
buf ( n10430 , n10429 );
buf ( n10431 , n10430 );
buf ( n10432 , n4355 );
or ( n10433 , n10431 , n10432 );
nand ( n10434 , n10420 , n10433 );
buf ( n10435 , n10434 );
buf ( n10436 , n10435 );
buf ( n10437 , n795 );
buf ( n10438 , n800 );
and ( n10439 , n10437 , n10438 );
buf ( n10440 , n10439 );
buf ( n10441 , n10440 );
buf ( n10442 , n794 );
buf ( n10443 , n800 );
xor ( n10444 , n10442 , n10443 );
buf ( n10445 , n10444 );
buf ( n10446 , n10445 );
not ( n10447 , n10446 );
buf ( n10448 , n3656 );
not ( n10449 , n10448 );
or ( n10450 , n10447 , n10449 );
buf ( n10451 , n3662 );
xor ( n10452 , n800 , n793 );
buf ( n10453 , n10452 );
nand ( n10454 , n10451 , n10453 );
buf ( n10455 , n10454 );
buf ( n10456 , n10455 );
nand ( n10457 , n10450 , n10456 );
buf ( n10458 , n10457 );
buf ( n10459 , n10458 );
xor ( n10460 , n10441 , n10459 );
buf ( n10461 , n768 );
buf ( n10462 , n826 );
xor ( n10463 , n10461 , n10462 );
buf ( n10464 , n10463 );
buf ( n10465 , n10464 );
not ( n10466 , n10465 );
buf ( n10467 , n4496 );
not ( n10468 , n10467 );
or ( n10469 , n10466 , n10468 );
buf ( n10470 , n1771 );
buf ( n10471 , n826 );
nand ( n10472 , n10470 , n10471 );
buf ( n10473 , n10472 );
buf ( n10474 , n10473 );
nand ( n10475 , n10469 , n10474 );
buf ( n10476 , n10475 );
buf ( n10477 , n10476 );
not ( n10478 , n10477 );
buf ( n10479 , n10478 );
buf ( n10480 , n10479 );
xor ( n10481 , n10460 , n10480 );
buf ( n10482 , n10481 );
buf ( n10483 , n10482 );
buf ( n10484 , n768 );
buf ( n10485 , n828 );
xor ( n10486 , n10484 , n10485 );
buf ( n10487 , n10486 );
buf ( n10488 , n10487 );
not ( n10489 , n10488 );
buf ( n10490 , n3680 );
not ( n10491 , n10490 );
or ( n10492 , n10489 , n10491 );
buf ( n10493 , n828 );
buf ( n10494 , n1249 );
nand ( n10495 , n10493 , n10494 );
buf ( n10496 , n10495 );
buf ( n10497 , n10496 );
nand ( n10498 , n10492 , n10497 );
buf ( n10499 , n10498 );
buf ( n10500 , n10499 );
buf ( n10501 , n795 );
buf ( n10502 , n800 );
xor ( n10503 , n10501 , n10502 );
buf ( n10504 , n10503 );
buf ( n10505 , n10504 );
not ( n10506 , n10505 );
buf ( n10507 , n3656 );
buf ( n10508 , n10507 );
buf ( n10509 , n10508 );
buf ( n10510 , n10509 );
not ( n10511 , n10510 );
or ( n10512 , n10506 , n10511 );
buf ( n10513 , n3662 );
buf ( n10514 , n10445 );
nand ( n10515 , n10513 , n10514 );
buf ( n10516 , n10515 );
buf ( n10517 , n10516 );
nand ( n10518 , n10512 , n10517 );
buf ( n10519 , n10518 );
buf ( n10520 , n10519 );
xor ( n10521 , n10500 , n10520 );
buf ( n10522 , n797 );
buf ( n10523 , n800 );
and ( n10524 , n10522 , n10523 );
buf ( n10525 , n10524 );
buf ( n10526 , n10525 );
buf ( n10527 , n774 );
buf ( n10528 , n822 );
xor ( n10529 , n10527 , n10528 );
buf ( n10530 , n10529 );
buf ( n10531 , n10530 );
not ( n10532 , n10531 );
buf ( n10533 , n2577 );
not ( n10534 , n10533 );
or ( n10535 , n10532 , n10534 );
buf ( n10536 , n2107 );
buf ( n10537 , n773 );
buf ( n10538 , n822 );
xor ( n10539 , n10537 , n10538 );
buf ( n10540 , n10539 );
buf ( n10541 , n10540 );
nand ( n10542 , n10536 , n10541 );
buf ( n10543 , n10542 );
buf ( n10544 , n10543 );
nand ( n10545 , n10535 , n10544 );
buf ( n10546 , n10545 );
buf ( n10547 , n10546 );
xor ( n10548 , n10526 , n10547 );
buf ( n10549 , n770 );
buf ( n10550 , n826 );
xor ( n10551 , n10549 , n10550 );
buf ( n10552 , n10551 );
buf ( n10553 , n10552 );
not ( n10554 , n10553 );
buf ( n10555 , n1780 );
not ( n10556 , n10555 );
or ( n10557 , n10554 , n10556 );
buf ( n10558 , n1374 );
buf ( n10559 , n769 );
buf ( n10560 , n826 );
xor ( n10561 , n10559 , n10560 );
buf ( n10562 , n10561 );
buf ( n10563 , n10562 );
nand ( n10564 , n10558 , n10563 );
buf ( n10565 , n10564 );
buf ( n10566 , n10565 );
nand ( n10567 , n10557 , n10566 );
buf ( n10568 , n10567 );
buf ( n10569 , n10568 );
and ( n10570 , n10548 , n10569 );
and ( n10571 , n10526 , n10547 );
or ( n10572 , n10570 , n10571 );
buf ( n10573 , n10572 );
buf ( n10574 , n10573 );
and ( n10575 , n10521 , n10574 );
and ( n10576 , n10500 , n10520 );
or ( n10577 , n10575 , n10576 );
buf ( n10578 , n10577 );
buf ( n10579 , n10578 );
xor ( n10580 , n10483 , n10579 );
buf ( n10581 , n782 );
buf ( n10582 , n814 );
xor ( n10583 , n10581 , n10582 );
buf ( n10584 , n10583 );
buf ( n10585 , n10584 );
not ( n10586 , n10585 );
buf ( n10587 , n1931 );
not ( n10588 , n10587 );
or ( n10589 , n10586 , n10588 );
buf ( n10590 , n2621 );
buf ( n10591 , n781 );
buf ( n10592 , n814 );
xor ( n10593 , n10591 , n10592 );
buf ( n10594 , n10593 );
buf ( n10595 , n10594 );
nand ( n10596 , n10590 , n10595 );
buf ( n10597 , n10596 );
buf ( n10598 , n10597 );
nand ( n10599 , n10589 , n10598 );
buf ( n10600 , n10599 );
buf ( n10601 , n10600 );
not ( n10602 , n10601 );
not ( n10603 , n1346 );
xor ( n10604 , n820 , n775 );
not ( n10605 , n10604 );
or ( n10606 , n10603 , n10605 );
buf ( n10607 , n776 );
buf ( n10608 , n820 );
xnor ( n10609 , n10607 , n10608 );
buf ( n10610 , n10609 );
or ( n10611 , n2678 , n10610 );
nand ( n10612 , n10606 , n10611 );
buf ( n10613 , n10612 );
not ( n10614 , n10613 );
or ( n10615 , n10602 , n10614 );
buf ( n10616 , n10600 );
buf ( n10617 , n10612 );
or ( n10618 , n10616 , n10617 );
buf ( n10619 , n784 );
buf ( n10620 , n812 );
xor ( n10621 , n10619 , n10620 );
buf ( n10622 , n10621 );
buf ( n10623 , n10622 );
not ( n10624 , n10623 );
buf ( n10625 , n1712 );
not ( n10626 , n10625 );
or ( n10627 , n10624 , n10626 );
buf ( n10628 , n1693 );
buf ( n10629 , n783 );
buf ( n10630 , n812 );
xor ( n10631 , n10629 , n10630 );
buf ( n10632 , n10631 );
buf ( n10633 , n10632 );
nand ( n10634 , n10628 , n10633 );
buf ( n10635 , n10634 );
buf ( n10636 , n10635 );
nand ( n10637 , n10627 , n10636 );
buf ( n10638 , n10637 );
buf ( n10639 , n10638 );
nand ( n10640 , n10618 , n10639 );
buf ( n10641 , n10640 );
buf ( n10642 , n10641 );
nand ( n10643 , n10615 , n10642 );
buf ( n10644 , n10643 );
buf ( n10645 , n10644 );
buf ( n10646 , n772 );
buf ( n10647 , n824 );
xor ( n10648 , n10646 , n10647 );
buf ( n10649 , n10648 );
buf ( n10650 , n10649 );
not ( n10651 , n10650 );
buf ( n10652 , n1844 );
not ( n10653 , n10652 );
or ( n10654 , n10651 , n10653 );
buf ( n10655 , n3255 );
buf ( n10656 , n771 );
buf ( n10657 , n824 );
xor ( n10658 , n10656 , n10657 );
buf ( n10659 , n10658 );
buf ( n10660 , n10659 );
nand ( n10661 , n10655 , n10660 );
buf ( n10662 , n10661 );
buf ( n10663 , n10662 );
nand ( n10664 , n10654 , n10663 );
buf ( n10665 , n10664 );
buf ( n10666 , n788 );
buf ( n10667 , n808 );
xor ( n10668 , n10666 , n10667 );
buf ( n10669 , n10668 );
buf ( n10670 , n10669 );
not ( n10671 , n10670 );
buf ( n10672 , n2232 );
not ( n10673 , n10672 );
buf ( n10674 , n10673 );
buf ( n10675 , n10674 );
not ( n10676 , n10675 );
or ( n10677 , n10671 , n10676 );
buf ( n10678 , n1309 );
buf ( n10679 , n787 );
buf ( n10680 , n808 );
xor ( n10681 , n10679 , n10680 );
buf ( n10682 , n10681 );
buf ( n10683 , n10682 );
nand ( n10684 , n10678 , n10683 );
buf ( n10685 , n10684 );
buf ( n10686 , n10685 );
nand ( n10687 , n10677 , n10686 );
buf ( n10688 , n10687 );
or ( n10689 , n10665 , n10688 );
buf ( n10690 , n786 );
buf ( n10691 , n810 );
xor ( n10692 , n10690 , n10691 );
buf ( n10693 , n10692 );
buf ( n10694 , n10693 );
not ( n10695 , n10694 );
buf ( n10696 , n2896 );
not ( n10697 , n10696 );
or ( n10698 , n10695 , n10697 );
buf ( n10699 , n2647 );
buf ( n10700 , n785 );
buf ( n10701 , n810 );
xor ( n10702 , n10700 , n10701 );
buf ( n10703 , n10702 );
buf ( n10704 , n10703 );
nand ( n10705 , n10699 , n10704 );
buf ( n10706 , n10705 );
buf ( n10707 , n10706 );
nand ( n10708 , n10698 , n10707 );
buf ( n10709 , n10708 );
nand ( n10710 , n10689 , n10709 );
buf ( n10711 , n10665 );
buf ( n10712 , n10688 );
nand ( n10713 , n10711 , n10712 );
buf ( n10714 , n10713 );
nand ( n10715 , n10710 , n10714 );
buf ( n10716 , n10715 );
or ( n10717 , n10645 , n10716 );
buf ( n10718 , n790 );
buf ( n10719 , n806 );
xor ( n10720 , n10718 , n10719 );
buf ( n10721 , n10720 );
buf ( n10722 , n10721 );
not ( n10723 , n10722 );
buf ( n10724 , n2325 );
not ( n10725 , n10724 );
or ( n10726 , n10723 , n10725 );
buf ( n10727 , n2331 );
buf ( n10728 , n789 );
buf ( n10729 , n806 );
xor ( n10730 , n10728 , n10729 );
buf ( n10731 , n10730 );
buf ( n10732 , n10731 );
nand ( n10733 , n10727 , n10732 );
buf ( n10734 , n10733 );
buf ( n10735 , n10734 );
nand ( n10736 , n10726 , n10735 );
buf ( n10737 , n10736 );
buf ( n10738 , n10737 );
buf ( n10739 , n792 );
buf ( n10740 , n804 );
xor ( n10741 , n10739 , n10740 );
buf ( n10742 , n10741 );
buf ( n10743 , n10742 );
not ( n10744 , n10743 );
buf ( n10745 , n1522 );
not ( n10746 , n10745 );
or ( n10747 , n10744 , n10746 );
buf ( n10748 , n1449 );
buf ( n10749 , n791 );
buf ( n10750 , n804 );
xor ( n10751 , n10749 , n10750 );
buf ( n10752 , n10751 );
buf ( n10753 , n10752 );
nand ( n10754 , n10748 , n10753 );
buf ( n10755 , n10754 );
buf ( n10756 , n10755 );
nand ( n10757 , n10747 , n10756 );
buf ( n10758 , n10757 );
buf ( n10759 , n10758 );
xor ( n10760 , n10738 , n10759 );
buf ( n10761 , n778 );
buf ( n10762 , n818 );
xor ( n10763 , n10761 , n10762 );
buf ( n10764 , n10763 );
buf ( n10765 , n10764 );
not ( n10766 , n10765 );
buf ( n10767 , n1480 );
not ( n10768 , n10767 );
or ( n10769 , n10766 , n10768 );
buf ( n10770 , n1496 );
xor ( n10771 , n777 , n818 );
buf ( n10772 , n10771 );
nand ( n10773 , n10770 , n10772 );
buf ( n10774 , n10773 );
buf ( n10775 , n10774 );
nand ( n10776 , n10769 , n10775 );
buf ( n10777 , n10776 );
buf ( n10778 , n10777 );
and ( n10779 , n10760 , n10778 );
and ( n10780 , n10738 , n10759 );
or ( n10781 , n10779 , n10780 );
buf ( n10782 , n10781 );
buf ( n10783 , n10782 );
nand ( n10784 , n10717 , n10783 );
buf ( n10785 , n10784 );
buf ( n10786 , n10785 );
buf ( n10787 , n10644 );
buf ( n10788 , n10715 );
nand ( n10789 , n10787 , n10788 );
buf ( n10790 , n10789 );
buf ( n10791 , n10790 );
nand ( n10792 , n10786 , n10791 );
buf ( n10793 , n10792 );
buf ( n10794 , n10793 );
and ( n10795 , n10580 , n10794 );
and ( n10796 , n10483 , n10579 );
or ( n10797 , n10795 , n10796 );
buf ( n10798 , n10797 );
buf ( n10799 , n10798 );
buf ( n10800 , n796 );
buf ( n10801 , n800 );
and ( n10802 , n10800 , n10801 );
buf ( n10803 , n10802 );
buf ( n10804 , n10803 );
buf ( n10805 , n10632 );
not ( n10806 , n10805 );
buf ( n10807 , n1712 );
not ( n10808 , n10807 );
or ( n10809 , n10806 , n10808 );
buf ( n10810 , n1693 );
buf ( n10811 , n782 );
buf ( n10812 , n812 );
xor ( n10813 , n10811 , n10812 );
buf ( n10814 , n10813 );
buf ( n10815 , n10814 );
nand ( n10816 , n10810 , n10815 );
buf ( n10817 , n10816 );
buf ( n10818 , n10817 );
nand ( n10819 , n10809 , n10818 );
buf ( n10820 , n10819 );
buf ( n10821 , n10820 );
xor ( n10822 , n10804 , n10821 );
buf ( n10823 , n10594 );
not ( n10824 , n10823 );
buf ( n10825 , n1931 );
not ( n10826 , n10825 );
or ( n10827 , n10824 , n10826 );
buf ( n10828 , n1937 );
buf ( n10829 , n780 );
buf ( n10830 , n814 );
xor ( n10831 , n10829 , n10830 );
buf ( n10832 , n10831 );
buf ( n10833 , n10832 );
nand ( n10834 , n10828 , n10833 );
buf ( n10835 , n10834 );
buf ( n10836 , n10835 );
nand ( n10837 , n10827 , n10836 );
buf ( n10838 , n10837 );
buf ( n10839 , n10838 );
xnor ( n10840 , n10822 , n10839 );
buf ( n10841 , n10840 );
buf ( n10842 , n10841 );
not ( n10843 , n10842 );
buf ( n10844 , n829 );
buf ( n10845 , n830 );
xnor ( n10846 , n10844 , n10845 );
buf ( n10847 , n10846 );
buf ( n10848 , n10847 );
buf ( n10849 , n1237 );
nand ( n10850 , n10848 , n10849 );
buf ( n10851 , n10850 );
buf ( n10852 , n10851 );
not ( n10853 , n10852 );
buf ( n10854 , n9454 );
not ( n10855 , n10854 );
or ( n10856 , n10853 , n10855 );
buf ( n10857 , n828 );
nand ( n10858 , n10856 , n10857 );
buf ( n10859 , n10858 );
buf ( n10860 , n10859 );
not ( n10861 , n10860 );
buf ( n10862 , n10861 );
buf ( n10863 , n10562 );
not ( n10864 , n10863 );
buf ( n10865 , n2364 );
not ( n10866 , n10865 );
or ( n10867 , n10864 , n10866 );
buf ( n10868 , n10464 );
buf ( n10869 , n1771 );
nand ( n10870 , n10868 , n10869 );
buf ( n10871 , n10870 );
buf ( n10872 , n10871 );
nand ( n10873 , n10867 , n10872 );
buf ( n10874 , n10873 );
xor ( n10875 , n10862 , n10874 );
buf ( n10876 , n10540 );
not ( n10877 , n10876 );
buf ( n10878 , n2098 );
not ( n10879 , n10878 );
or ( n10880 , n10877 , n10879 );
buf ( n10881 , n2107 );
buf ( n10882 , n772 );
buf ( n10883 , n822 );
xor ( n10884 , n10882 , n10883 );
buf ( n10885 , n10884 );
buf ( n10886 , n10885 );
nand ( n10887 , n10881 , n10886 );
buf ( n10888 , n10887 );
buf ( n10889 , n10888 );
nand ( n10890 , n10880 , n10889 );
buf ( n10891 , n10890 );
and ( n10892 , n10875 , n10891 );
not ( n10893 , n10875 );
buf ( n10894 , n10891 );
not ( n10895 , n10894 );
buf ( n10896 , n10895 );
and ( n10897 , n10893 , n10896 );
nor ( n10898 , n10892 , n10897 );
buf ( n10899 , n10898 );
not ( n10900 , n10899 );
or ( n10901 , n10843 , n10900 );
buf ( n10902 , n794 );
buf ( n10903 , n802 );
xor ( n10904 , n10902 , n10903 );
buf ( n10905 , n10904 );
buf ( n10906 , n10905 );
not ( n10907 , n10906 );
buf ( n10908 , n802 );
not ( n10909 , n10908 );
buf ( n10910 , n803 );
not ( n10911 , n10910 );
and ( n10912 , n10909 , n10911 );
buf ( n10913 , n802 );
buf ( n10914 , n803 );
and ( n10915 , n10913 , n10914 );
nor ( n10916 , n10912 , n10915 );
buf ( n10917 , n10916 );
buf ( n10918 , n10917 );
not ( n10919 , n10918 );
buf ( n10920 , n1547 );
nor ( n10921 , n10919 , n10920 );
buf ( n10922 , n10921 );
buf ( n10923 , n10922 );
not ( n10924 , n10923 );
or ( n10925 , n10907 , n10924 );
buf ( n10926 , n1557 );
buf ( n10927 , n793 );
buf ( n10928 , n802 );
xor ( n10929 , n10927 , n10928 );
buf ( n10930 , n10929 );
buf ( n10931 , n10930 );
nand ( n10932 , n10926 , n10931 );
buf ( n10933 , n10932 );
buf ( n10934 , n10933 );
nand ( n10935 , n10925 , n10934 );
buf ( n10936 , n10935 );
buf ( n10937 , n10936 );
buf ( n10938 , n796 );
buf ( n10939 , n800 );
xor ( n10940 , n10938 , n10939 );
buf ( n10941 , n10940 );
buf ( n10942 , n10941 );
not ( n10943 , n10942 );
buf ( n10944 , n3656 );
not ( n10945 , n10944 );
or ( n10946 , n10943 , n10945 );
buf ( n10947 , n3662 );
buf ( n10948 , n10504 );
nand ( n10949 , n10947 , n10948 );
buf ( n10950 , n10949 );
buf ( n10951 , n10950 );
nand ( n10952 , n10946 , n10951 );
buf ( n10953 , n10952 );
buf ( n10954 , n10953 );
xor ( n10955 , n10937 , n10954 );
buf ( n10956 , n780 );
buf ( n10957 , n816 );
xor ( n10958 , n10956 , n10957 );
buf ( n10959 , n10958 );
buf ( n10960 , n10959 );
not ( n10961 , n10960 );
buf ( n10962 , n2526 );
not ( n10963 , n10962 );
or ( n10964 , n10961 , n10963 );
buf ( n10965 , n779 );
buf ( n10966 , n816 );
xor ( n10967 , n10965 , n10966 );
buf ( n10968 , n10967 );
buf ( n10969 , n10968 );
buf ( n10970 , n2010 );
nand ( n10971 , n10969 , n10970 );
buf ( n10972 , n10971 );
buf ( n10973 , n10972 );
nand ( n10974 , n10964 , n10973 );
buf ( n10975 , n10974 );
buf ( n10976 , n10975 );
and ( n10977 , n10955 , n10976 );
and ( n10978 , n10937 , n10954 );
or ( n10979 , n10977 , n10978 );
buf ( n10980 , n10979 );
buf ( n10981 , n10980 );
nand ( n10982 , n10901 , n10981 );
buf ( n10983 , n10982 );
buf ( n10984 , n10983 );
buf ( n10985 , n10803 );
buf ( n10986 , n10820 );
xor ( n10987 , n10985 , n10986 );
buf ( n10988 , n10838 );
xnor ( n10989 , n10987 , n10988 );
buf ( n10990 , n10989 );
buf ( n10991 , n10990 );
not ( n10992 , n10991 );
buf ( n10993 , n10898 );
not ( n10994 , n10993 );
buf ( n10995 , n10994 );
buf ( n10996 , n10995 );
nand ( n10997 , n10992 , n10996 );
buf ( n10998 , n10997 );
buf ( n10999 , n10998 );
nand ( n11000 , n10984 , n10999 );
buf ( n11001 , n11000 );
buf ( n11002 , n11001 );
not ( n11003 , n10838 );
not ( n11004 , n10803 );
or ( n11005 , n11003 , n11004 );
buf ( n11006 , n10838 );
buf ( n11007 , n10803 );
nor ( n11008 , n11006 , n11007 );
buf ( n11009 , n11008 );
buf ( n11010 , n10820 );
not ( n11011 , n11010 );
buf ( n11012 , n11011 );
or ( n11013 , n11009 , n11012 );
nand ( n11014 , n11005 , n11013 );
buf ( n11015 , n11014 );
buf ( n11016 , n10874 );
buf ( n11017 , n10891 );
nor ( n11018 , n11016 , n11017 );
buf ( n11019 , n11018 );
buf ( n11020 , n11019 );
buf ( n11021 , n10862 );
or ( n11022 , n11020 , n11021 );
buf ( n11023 , n10874 );
buf ( n11024 , n10891 );
nand ( n11025 , n11023 , n11024 );
buf ( n11026 , n11025 );
buf ( n11027 , n11026 );
nand ( n11028 , n11022 , n11027 );
buf ( n11029 , n11028 );
buf ( n11030 , n11029 );
xor ( n11031 , n11015 , n11030 );
buf ( n11032 , n10682 );
not ( n11033 , n11032 );
buf ( n11034 , n10674 );
not ( n11035 , n11034 );
or ( n11036 , n11033 , n11035 );
buf ( n11037 , n1309 );
xor ( n11038 , n808 , n786 );
buf ( n11039 , n11038 );
nand ( n11040 , n11037 , n11039 );
buf ( n11041 , n11040 );
buf ( n11042 , n11041 );
nand ( n11043 , n11036 , n11042 );
buf ( n11044 , n11043 );
buf ( n11045 , n11044 );
buf ( n11046 , n10703 );
not ( n11047 , n11046 );
buf ( n11048 , n1667 );
not ( n11049 , n11048 );
buf ( n11050 , n11049 );
buf ( n11051 , n11050 );
not ( n11052 , n11051 );
or ( n11053 , n11047 , n11052 );
buf ( n11054 , n3398 );
xor ( n11055 , n810 , n784 );
buf ( n11056 , n11055 );
nand ( n11057 , n11054 , n11056 );
buf ( n11058 , n11057 );
buf ( n11059 , n11058 );
nand ( n11060 , n11053 , n11059 );
buf ( n11061 , n11060 );
buf ( n11062 , n11061 );
xor ( n11063 , n11045 , n11062 );
not ( n11064 , n2672 );
xor ( n11065 , n820 , n774 );
not ( n11066 , n11065 );
or ( n11067 , n11064 , n11066 );
buf ( n11068 , n10604 );
not ( n11069 , n11068 );
buf ( n11070 , n11069 );
or ( n11071 , n2681 , n11070 );
nand ( n11072 , n11067 , n11071 );
buf ( n11073 , n11072 );
and ( n11074 , n11063 , n11073 );
and ( n11075 , n11045 , n11062 );
or ( n11076 , n11074 , n11075 );
buf ( n11077 , n11076 );
buf ( n11078 , n11077 );
xor ( n11079 , n11031 , n11078 );
buf ( n11080 , n11079 );
buf ( n11081 , n11080 );
xor ( n11082 , n11002 , n11081 );
buf ( n11083 , n10659 );
not ( n11084 , n11083 );
buf ( n11085 , n1965 );
not ( n11086 , n11085 );
or ( n11087 , n11084 , n11086 );
buf ( n11088 , n3255 );
buf ( n11089 , n770 );
buf ( n11090 , n824 );
xor ( n11091 , n11089 , n11090 );
buf ( n11092 , n11091 );
buf ( n11093 , n11092 );
nand ( n11094 , n11088 , n11093 );
buf ( n11095 , n11094 );
buf ( n11096 , n11095 );
nand ( n11097 , n11087 , n11096 );
buf ( n11098 , n11097 );
buf ( n11099 , n11098 );
not ( n11100 , n1496 );
xor ( n11101 , n818 , n776 );
not ( n11102 , n11101 );
or ( n11103 , n11100 , n11102 );
not ( n11104 , n1474 );
not ( n11105 , n1478 );
nand ( n11106 , n11104 , n11105 , n10771 );
nand ( n11107 , n11103 , n11106 );
buf ( n11108 , n11107 );
xor ( n11109 , n11099 , n11108 );
buf ( n11110 , n10731 );
not ( n11111 , n11110 );
buf ( n11112 , n1403 );
not ( n11113 , n11112 );
or ( n11114 , n11111 , n11113 );
buf ( n11115 , n2331 );
buf ( n11116 , n788 );
buf ( n11117 , n806 );
xor ( n11118 , n11116 , n11117 );
buf ( n11119 , n11118 );
buf ( n11120 , n11119 );
nand ( n11121 , n11115 , n11120 );
buf ( n11122 , n11121 );
buf ( n11123 , n11122 );
nand ( n11124 , n11114 , n11123 );
buf ( n11125 , n11124 );
buf ( n11126 , n11125 );
and ( n11127 , n11109 , n11126 );
and ( n11128 , n11099 , n11108 );
or ( n11129 , n11127 , n11128 );
buf ( n11130 , n11129 );
buf ( n11131 , n11130 );
not ( n11132 , n10752 );
not ( n11133 , n1440 );
or ( n11134 , n11132 , n11133 );
buf ( n11135 , n1449 );
buf ( n11136 , n11135 );
buf ( n11137 , n11136 );
buf ( n11138 , n11137 );
xor ( n11139 , n804 , n790 );
buf ( n11140 , n11139 );
nand ( n11141 , n11138 , n11140 );
buf ( n11142 , n11141 );
nand ( n11143 , n11134 , n11142 );
buf ( n11144 , n10930 );
not ( n11145 , n11144 );
buf ( n11146 , n1551 );
not ( n11147 , n11146 );
or ( n11148 , n11145 , n11147 );
buf ( n11149 , n1560 );
buf ( n11150 , n792 );
buf ( n11151 , n802 );
xor ( n11152 , n11150 , n11151 );
buf ( n11153 , n11152 );
buf ( n11154 , n11153 );
nand ( n11155 , n11149 , n11154 );
buf ( n11156 , n11155 );
buf ( n11157 , n11156 );
nand ( n11158 , n11148 , n11157 );
buf ( n11159 , n11158 );
or ( n11160 , n11143 , n11159 );
not ( n11161 , n10968 );
not ( n11162 , n2526 );
or ( n11163 , n11161 , n11162 );
buf ( n11164 , n2535 );
buf ( n11165 , n778 );
buf ( n11166 , n816 );
xor ( n11167 , n11165 , n11166 );
buf ( n11168 , n11167 );
buf ( n11169 , n11168 );
nand ( n11170 , n11164 , n11169 );
buf ( n11171 , n11170 );
nand ( n11172 , n11163 , n11171 );
nand ( n11173 , n11160 , n11172 );
buf ( n11174 , n11173 );
buf ( n11175 , n11143 );
buf ( n11176 , n11159 );
nand ( n11177 , n11175 , n11176 );
buf ( n11178 , n11177 );
buf ( n11179 , n11178 );
nand ( n11180 , n11174 , n11179 );
buf ( n11181 , n11180 );
buf ( n11182 , n11181 );
xor ( n11183 , n11131 , n11182 );
buf ( n11184 , n11092 );
not ( n11185 , n11184 );
buf ( n11186 , n2483 );
not ( n11187 , n11186 );
or ( n11188 , n11185 , n11187 );
buf ( n11189 , n8354 );
buf ( n11190 , n769 );
not ( n11191 , n11190 );
buf ( n11192 , n11191 );
and ( n11193 , n824 , n11192 );
not ( n11194 , n824 );
and ( n11195 , n11194 , n769 );
or ( n11196 , n11193 , n11195 );
buf ( n11197 , n11196 );
nand ( n11198 , n11189 , n11197 );
buf ( n11199 , n11198 );
buf ( n11200 , n11199 );
nand ( n11201 , n11188 , n11200 );
buf ( n11202 , n11201 );
buf ( n11203 , n11202 );
buf ( n11204 , n10814 );
not ( n11205 , n11204 );
buf ( n11206 , n2066 );
not ( n11207 , n11206 );
or ( n11208 , n11205 , n11207 );
buf ( n11209 , n3379 );
xor ( n11210 , n812 , n781 );
buf ( n11211 , n11210 );
nand ( n11212 , n11209 , n11211 );
buf ( n11213 , n11212 );
buf ( n11214 , n11213 );
nand ( n11215 , n11208 , n11214 );
buf ( n11216 , n11215 );
buf ( n11217 , n11216 );
xor ( n11218 , n11203 , n11217 );
buf ( n11219 , n11065 );
not ( n11220 , n11219 );
buf ( n11221 , n2410 );
not ( n11222 , n11221 );
or ( n11223 , n11220 , n11222 );
buf ( n11224 , n2672 );
buf ( n11225 , n773 );
buf ( n11226 , n820 );
xor ( n11227 , n11225 , n11226 );
buf ( n11228 , n11227 );
buf ( n11229 , n11228 );
nand ( n11230 , n11224 , n11229 );
buf ( n11231 , n11230 );
buf ( n11232 , n11231 );
nand ( n11233 , n11223 , n11232 );
buf ( n11234 , n11233 );
buf ( n11235 , n11234 );
xor ( n11236 , n11218 , n11235 );
buf ( n11237 , n11236 );
buf ( n11238 , n11237 );
xor ( n11239 , n11183 , n11238 );
buf ( n11240 , n11239 );
buf ( n11241 , n11240 );
and ( n11242 , n11082 , n11241 );
and ( n11243 , n11002 , n11081 );
or ( n11244 , n11242 , n11243 );
buf ( n11245 , n11244 );
buf ( n11246 , n11245 );
xor ( n11247 , n10799 , n11246 );
buf ( n11248 , n10476 );
buf ( n11249 , n11101 );
not ( n11250 , n11249 );
buf ( n11251 , n4396 );
not ( n11252 , n11251 );
or ( n11253 , n11250 , n11252 );
buf ( n11254 , n1493 );
buf ( n11255 , n775 );
buf ( n11256 , n818 );
xor ( n11257 , n11255 , n11256 );
buf ( n11258 , n11257 );
buf ( n11259 , n11258 );
nand ( n11260 , n11254 , n11259 );
buf ( n11261 , n11260 );
buf ( n11262 , n11261 );
nand ( n11263 , n11253 , n11262 );
buf ( n11264 , n11263 );
buf ( n11265 , n11264 );
not ( n11266 , n1305 );
not ( n11267 , n11038 );
or ( n11268 , n11266 , n11267 );
buf ( n11269 , n1309 );
xor ( n11270 , n808 , n785 );
buf ( n11271 , n11270 );
nand ( n11272 , n11269 , n11271 );
buf ( n11273 , n11272 );
nand ( n11274 , n11268 , n11273 );
buf ( n11275 , n11274 );
xor ( n11276 , n11265 , n11275 );
buf ( n11277 , n11055 );
not ( n11278 , n11277 );
buf ( n11279 , n4570 );
not ( n11280 , n11279 );
or ( n11281 , n11278 , n11280 );
buf ( n11282 , n5272 );
xor ( n11283 , n810 , n783 );
buf ( n11284 , n11283 );
nand ( n11285 , n11282 , n11284 );
buf ( n11286 , n11285 );
buf ( n11287 , n11286 );
nand ( n11288 , n11281 , n11287 );
buf ( n11289 , n11288 );
buf ( n11290 , n11289 );
and ( n11291 , n11276 , n11290 );
and ( n11292 , n11265 , n11275 );
or ( n11293 , n11291 , n11292 );
buf ( n11294 , n11293 );
buf ( n11295 , n11294 );
xor ( n11296 , n11248 , n11295 );
xor ( n11297 , n11203 , n11217 );
and ( n11298 , n11297 , n11235 );
and ( n11299 , n11203 , n11217 );
or ( n11300 , n11298 , n11299 );
buf ( n11301 , n11300 );
buf ( n11302 , n11301 );
xor ( n11303 , n11296 , n11302 );
buf ( n11304 , n11303 );
xor ( n11305 , n11131 , n11182 );
and ( n11306 , n11305 , n11238 );
and ( n11307 , n11131 , n11182 );
or ( n11308 , n11306 , n11307 );
buf ( n11309 , n11308 );
xor ( n11310 , n11304 , n11309 );
buf ( n11311 , n11139 );
not ( n11312 , n11311 );
buf ( n11313 , n1737 );
not ( n11314 , n11313 );
or ( n11315 , n11312 , n11314 );
buf ( n11316 , n1433 );
buf ( n11317 , n789 );
buf ( n11318 , n804 );
xor ( n11319 , n11317 , n11318 );
buf ( n11320 , n11319 );
buf ( n11321 , n11320 );
nand ( n11322 , n11316 , n11321 );
buf ( n11323 , n11322 );
buf ( n11324 , n11323 );
nand ( n11325 , n11315 , n11324 );
buf ( n11326 , n11325 );
not ( n11327 , n11326 );
buf ( n11328 , n10832 );
not ( n11329 , n11328 );
buf ( n11330 , n1931 );
not ( n11331 , n11330 );
or ( n11332 , n11329 , n11331 );
buf ( n11333 , n2621 );
buf ( n11334 , n779 );
buf ( n11335 , n814 );
xor ( n11336 , n11334 , n11335 );
buf ( n11337 , n11336 );
buf ( n11338 , n11337 );
nand ( n11339 , n11333 , n11338 );
buf ( n11340 , n11339 );
buf ( n11341 , n11340 );
nand ( n11342 , n11332 , n11341 );
buf ( n11343 , n11342 );
not ( n11344 , n11343 );
or ( n11345 , n11327 , n11344 );
or ( n11346 , n11326 , n11343 );
not ( n11347 , n11153 );
not ( n11348 , n10922 );
or ( n11349 , n11347 , n11348 );
buf ( n11350 , n1557 );
buf ( n11351 , n791 );
buf ( n11352 , n802 );
xor ( n11353 , n11351 , n11352 );
buf ( n11354 , n11353 );
buf ( n11355 , n11354 );
nand ( n11356 , n11350 , n11355 );
buf ( n11357 , n11356 );
nand ( n11358 , n11349 , n11357 );
nand ( n11359 , n11346 , n11358 );
nand ( n11360 , n11345 , n11359 );
buf ( n11361 , n11360 );
buf ( n11362 , n11119 );
not ( n11363 , n11362 );
buf ( n11364 , n1403 );
not ( n11365 , n11364 );
or ( n11366 , n11363 , n11365 );
buf ( n11367 , n2331 );
buf ( n11368 , n787 );
buf ( n11369 , n806 );
xor ( n11370 , n11368 , n11369 );
buf ( n11371 , n11370 );
buf ( n11372 , n11371 );
nand ( n11373 , n11367 , n11372 );
buf ( n11374 , n11373 );
buf ( n11375 , n11374 );
nand ( n11376 , n11366 , n11375 );
buf ( n11377 , n11376 );
buf ( n11378 , n11377 );
not ( n11379 , n11378 );
buf ( n11380 , n10885 );
not ( n11381 , n11380 );
buf ( n11382 , n2101 );
not ( n11383 , n11382 );
or ( n11384 , n11381 , n11383 );
buf ( n11385 , n2107 );
xor ( n11386 , n822 , n771 );
buf ( n11387 , n11386 );
nand ( n11388 , n11385 , n11387 );
buf ( n11389 , n11388 );
buf ( n11390 , n11389 );
nand ( n11391 , n11384 , n11390 );
buf ( n11392 , n11391 );
buf ( n11393 , n11392 );
not ( n11394 , n11393 );
or ( n11395 , n11379 , n11394 );
buf ( n11396 , n11392 );
buf ( n11397 , n11377 );
or ( n11398 , n11396 , n11397 );
buf ( n11399 , n11168 );
not ( n11400 , n11399 );
buf ( n11401 , n2526 );
not ( n11402 , n11401 );
or ( n11403 , n11400 , n11402 );
buf ( n11404 , n2010 );
buf ( n11405 , n777 );
buf ( n11406 , n816 );
xor ( n11407 , n11405 , n11406 );
buf ( n11408 , n11407 );
buf ( n11409 , n11408 );
nand ( n11410 , n11404 , n11409 );
buf ( n11411 , n11410 );
buf ( n11412 , n11411 );
nand ( n11413 , n11403 , n11412 );
buf ( n11414 , n11413 );
buf ( n11415 , n11414 );
nand ( n11416 , n11398 , n11415 );
buf ( n11417 , n11416 );
buf ( n11418 , n11417 );
nand ( n11419 , n11395 , n11418 );
buf ( n11420 , n11419 );
buf ( n11421 , n11420 );
xor ( n11422 , n11361 , n11421 );
buf ( n11423 , n11258 );
not ( n11424 , n11423 );
buf ( n11425 , n1480 );
not ( n11426 , n11425 );
or ( n11427 , n11424 , n11426 );
buf ( n11428 , n1496 );
buf ( n11429 , n774 );
buf ( n11430 , n818 );
xor ( n11431 , n11429 , n11430 );
buf ( n11432 , n11431 );
buf ( n11433 , n11432 );
nand ( n11434 , n11428 , n11433 );
buf ( n11435 , n11434 );
buf ( n11436 , n11435 );
nand ( n11437 , n11427 , n11436 );
buf ( n11438 , n11437 );
buf ( n11439 , n11438 );
buf ( n11440 , n11283 );
not ( n11441 , n11440 );
buf ( n11442 , n4570 );
not ( n11443 , n11442 );
or ( n11444 , n11441 , n11443 );
buf ( n11445 , n3398 );
buf ( n11446 , n782 );
buf ( n11447 , n810 );
xor ( n11448 , n11446 , n11447 );
buf ( n11449 , n11448 );
buf ( n11450 , n11449 );
nand ( n11451 , n11445 , n11450 );
buf ( n11452 , n11451 );
buf ( n11453 , n11452 );
nand ( n11454 , n11444 , n11453 );
buf ( n11455 , n11454 );
buf ( n11456 , n11455 );
xor ( n11457 , n11439 , n11456 );
buf ( n11458 , n11210 );
not ( n11459 , n11458 );
buf ( n11460 , n2066 );
not ( n11461 , n11460 );
or ( n11462 , n11459 , n11461 );
buf ( n11463 , n1694 );
buf ( n11464 , n780 );
buf ( n11465 , n812 );
xor ( n11466 , n11464 , n11465 );
buf ( n11467 , n11466 );
buf ( n11468 , n11467 );
nand ( n11469 , n11463 , n11468 );
buf ( n11470 , n11469 );
buf ( n11471 , n11470 );
nand ( n11472 , n11462 , n11471 );
buf ( n11473 , n11472 );
buf ( n11474 , n11473 );
xor ( n11475 , n11457 , n11474 );
buf ( n11476 , n11475 );
buf ( n11477 , n11476 );
xor ( n11478 , n11422 , n11477 );
buf ( n11479 , n11478 );
xor ( n11480 , n11310 , n11479 );
buf ( n11481 , n11480 );
xor ( n11482 , n11247 , n11481 );
buf ( n11483 , n11482 );
buf ( n11484 , n11483 );
xor ( n11485 , n11099 , n11108 );
xor ( n11486 , n11485 , n11126 );
buf ( n11487 , n11486 );
buf ( n11488 , n11487 );
xor ( n11489 , n11045 , n11062 );
xor ( n11490 , n11489 , n11073 );
buf ( n11491 , n11490 );
buf ( n11492 , n11491 );
xor ( n11493 , n11488 , n11492 );
not ( n11494 , n11159 );
not ( n11495 , n11172 );
not ( n11496 , n11143 );
or ( n11497 , n11495 , n11496 );
or ( n11498 , n11143 , n11172 );
nand ( n11499 , n11497 , n11498 );
not ( n11500 , n11499 );
or ( n11501 , n11494 , n11500 );
or ( n11502 , n11499 , n11159 );
nand ( n11503 , n11501 , n11502 );
buf ( n11504 , n11503 );
and ( n11505 , n11493 , n11504 );
and ( n11506 , n11488 , n11492 );
or ( n11507 , n11505 , n11506 );
buf ( n11508 , n11507 );
buf ( n11509 , n11508 );
xor ( n11510 , n11358 , n11326 );
buf ( n11511 , n11510 );
buf ( n11512 , n11343 );
buf ( n11513 , n11512 );
buf ( n11514 , n11513 );
buf ( n11515 , n11514 );
xnor ( n11516 , n11511 , n11515 );
buf ( n11517 , n11516 );
not ( n11518 , n11517 );
xor ( n11519 , n11265 , n11275 );
xor ( n11520 , n11519 , n11290 );
buf ( n11521 , n11520 );
not ( n11522 , n11521 );
and ( n11523 , n11518 , n11522 );
and ( n11524 , n11517 , n11521 );
nor ( n11525 , n11523 , n11524 );
xor ( n11526 , n11414 , n11392 );
buf ( n11527 , n11526 );
buf ( n11528 , n11377 );
and ( n11529 , n11527 , n11528 );
not ( n11530 , n11527 );
buf ( n11531 , n11377 );
not ( n11532 , n11531 );
buf ( n11533 , n11532 );
buf ( n11534 , n11533 );
and ( n11535 , n11530 , n11534 );
nor ( n11536 , n11529 , n11535 );
buf ( n11537 , n11536 );
and ( n11538 , n11525 , n11537 );
not ( n11539 , n11525 );
buf ( n11540 , n11537 );
not ( n11541 , n11540 );
buf ( n11542 , n11541 );
and ( n11543 , n11539 , n11542 );
nor ( n11544 , n11538 , n11543 );
buf ( n11545 , n11544 );
not ( n11546 , n11545 );
buf ( n11547 , n11546 );
buf ( n11548 , n11547 );
or ( n11549 , n11509 , n11548 );
buf ( n11550 , n10499 );
buf ( n11551 , n830 );
nand ( n11552 , n11550 , n11551 );
buf ( n11553 , n11552 );
buf ( n11554 , n11553 );
not ( n11555 , n11554 );
buf ( n11556 , n798 );
buf ( n11557 , n800 );
and ( n11558 , n11556 , n11557 );
buf ( n11559 , n11558 );
buf ( n11560 , n11559 );
buf ( n11561 , n4241 );
not ( n11562 , n11561 );
buf ( n11563 , n3656 );
not ( n11564 , n11563 );
or ( n11565 , n11562 , n11564 );
buf ( n11566 , n3662 );
buf ( n11567 , n10941 );
nand ( n11568 , n11566 , n11567 );
buf ( n11569 , n11568 );
buf ( n11570 , n11569 );
nand ( n11571 , n11565 , n11570 );
buf ( n11572 , n11571 );
buf ( n11573 , n11572 );
xor ( n11574 , n11560 , n11573 );
buf ( n11575 , n4258 );
not ( n11576 , n11575 );
buf ( n11577 , n2526 );
not ( n11578 , n11577 );
or ( n11579 , n11576 , n11578 );
buf ( n11580 , n2010 );
buf ( n11581 , n10959 );
nand ( n11582 , n11580 , n11581 );
buf ( n11583 , n11582 );
buf ( n11584 , n11583 );
nand ( n11585 , n11579 , n11584 );
buf ( n11586 , n11585 );
buf ( n11587 , n11586 );
and ( n11588 , n11574 , n11587 );
and ( n11589 , n11560 , n11573 );
or ( n11590 , n11588 , n11589 );
buf ( n11591 , n11590 );
buf ( n11592 , n11591 );
not ( n11593 , n11592 );
or ( n11594 , n11555 , n11593 );
buf ( n11595 , n10499 );
not ( n11596 , n11595 );
buf ( n11597 , n830 );
not ( n11598 , n11597 );
buf ( n11599 , n11598 );
buf ( n11600 , n11599 );
nand ( n11601 , n11596 , n11600 );
buf ( n11602 , n11601 );
buf ( n11603 , n11602 );
nand ( n11604 , n11594 , n11603 );
buf ( n11605 , n11604 );
buf ( n11606 , n11605 );
xor ( n11607 , n10500 , n10520 );
xor ( n11608 , n11607 , n10574 );
buf ( n11609 , n11608 );
buf ( n11610 , n11609 );
xor ( n11611 , n11606 , n11610 );
buf ( n11612 , n3999 );
not ( n11613 , n11612 );
buf ( n11614 , n4570 );
not ( n11615 , n11614 );
or ( n11616 , n11613 , n11615 );
buf ( n11617 , n2647 );
buf ( n11618 , n10693 );
nand ( n11619 , n11617 , n11618 );
buf ( n11620 , n11619 );
buf ( n11621 , n11620 );
nand ( n11622 , n11616 , n11621 );
buf ( n11623 , n11622 );
buf ( n11624 , n11623 );
buf ( n11625 , n3908 );
not ( n11626 , n11625 );
buf ( n11627 , n2098 );
not ( n11628 , n11627 );
or ( n11629 , n11626 , n11628 );
buf ( n11630 , n2107 );
buf ( n11631 , n10530 );
nand ( n11632 , n11630 , n11631 );
buf ( n11633 , n11632 );
buf ( n11634 , n11633 );
nand ( n11635 , n11629 , n11634 );
buf ( n11636 , n11635 );
buf ( n11637 , n11636 );
or ( n11638 , n11624 , n11637 );
buf ( n11639 , n3958 );
not ( n11640 , n11639 );
buf ( n11641 , n2066 );
not ( n11642 , n11641 );
or ( n11643 , n11640 , n11642 );
buf ( n11644 , n1693 );
buf ( n11645 , n10622 );
nand ( n11646 , n11644 , n11645 );
buf ( n11647 , n11646 );
buf ( n11648 , n11647 );
nand ( n11649 , n11643 , n11648 );
buf ( n11650 , n11649 );
buf ( n11651 , n11650 );
nand ( n11652 , n11638 , n11651 );
buf ( n11653 , n11652 );
buf ( n11654 , n11636 );
buf ( n11655 , n11623 );
nand ( n11656 , n11654 , n11655 );
buf ( n11657 , n11656 );
nand ( n11658 , n11653 , n11657 );
buf ( n11659 , n11658 );
buf ( n11660 , n3931 );
not ( n11661 , n11660 );
buf ( n11662 , n3923 );
not ( n11663 , n11662 );
or ( n11664 , n11661 , n11663 );
buf ( n11665 , n1937 );
buf ( n11666 , n10584 );
nand ( n11667 , n11665 , n11666 );
buf ( n11668 , n11667 );
buf ( n11669 , n11668 );
nand ( n11670 , n11664 , n11669 );
buf ( n11671 , n11670 );
not ( n11672 , n11671 );
buf ( n11673 , n4273 );
not ( n11674 , n11673 );
buf ( n11675 , n2790 );
not ( n11676 , n11675 );
or ( n11677 , n11674 , n11676 );
buf ( n11678 , n2492 );
buf ( n11679 , n10649 );
nand ( n11680 , n11678 , n11679 );
buf ( n11681 , n11680 );
buf ( n11682 , n11681 );
nand ( n11683 , n11677 , n11682 );
buf ( n11684 , n11683 );
not ( n11685 , n11684 );
or ( n11686 , n11672 , n11685 );
or ( n11687 , n11671 , n11684 );
buf ( n11688 , n3850 );
not ( n11689 , n11688 );
buf ( n11690 , n3842 );
not ( n11691 , n11690 );
or ( n11692 , n11689 , n11691 );
buf ( n11693 , n1249 );
buf ( n11694 , n10487 );
nand ( n11695 , n11693 , n11694 );
buf ( n11696 , n11695 );
buf ( n11697 , n11696 );
nand ( n11698 , n11692 , n11697 );
buf ( n11699 , n11698 );
nand ( n11700 , n11687 , n11699 );
nand ( n11701 , n11686 , n11700 );
buf ( n11702 , n11701 );
or ( n11703 , n11659 , n11702 );
buf ( n11704 , n3981 );
not ( n11705 , n11704 );
buf ( n11706 , n1338 );
not ( n11707 , n11706 );
or ( n11708 , n11705 , n11707 );
buf ( n11709 , n10610 );
not ( n11710 , n11709 );
buf ( n11711 , n3986 );
nand ( n11712 , n11710 , n11711 );
buf ( n11713 , n11712 );
buf ( n11714 , n11713 );
nand ( n11715 , n11708 , n11714 );
buf ( n11716 , n11715 );
buf ( n11717 , n11716 );
buf ( n11718 , n4055 );
not ( n11719 , n11718 );
buf ( n11720 , n2235 );
not ( n11721 , n11720 );
or ( n11722 , n11719 , n11721 );
buf ( n11723 , n1309 );
buf ( n11724 , n10669 );
nand ( n11725 , n11723 , n11724 );
buf ( n11726 , n11725 );
buf ( n11727 , n11726 );
nand ( n11728 , n11722 , n11727 );
buf ( n11729 , n11728 );
buf ( n11730 , n11729 );
xor ( n11731 , n11717 , n11730 );
buf ( n11732 , n4025 );
not ( n11733 , n11732 );
buf ( n11734 , n4496 );
not ( n11735 , n11734 );
or ( n11736 , n11733 , n11735 );
buf ( n11737 , n1374 );
buf ( n11738 , n10552 );
nand ( n11739 , n11737 , n11738 );
buf ( n11740 , n11739 );
buf ( n11741 , n11740 );
nand ( n11742 , n11736 , n11741 );
buf ( n11743 , n11742 );
buf ( n11744 , n11743 );
and ( n11745 , n11731 , n11744 );
and ( n11746 , n11717 , n11730 );
or ( n11747 , n11745 , n11746 );
buf ( n11748 , n11747 );
buf ( n11749 , n11748 );
nand ( n11750 , n11703 , n11749 );
buf ( n11751 , n11750 );
buf ( n11752 , n11751 );
buf ( n11753 , n11658 );
buf ( n11754 , n11701 );
nand ( n11755 , n11753 , n11754 );
buf ( n11756 , n11755 );
buf ( n11757 , n11756 );
nand ( n11758 , n11752 , n11757 );
buf ( n11759 , n11758 );
buf ( n11760 , n11759 );
and ( n11761 , n11611 , n11760 );
and ( n11762 , n11606 , n11610 );
or ( n11763 , n11761 , n11762 );
buf ( n11764 , n11763 );
buf ( n11765 , n11764 );
nand ( n11766 , n11549 , n11765 );
buf ( n11767 , n11766 );
buf ( n11768 , n11767 );
buf ( n11769 , n11547 );
buf ( n11770 , n11508 );
nand ( n11771 , n11769 , n11770 );
buf ( n11772 , n11771 );
buf ( n11773 , n11772 );
nand ( n11774 , n11768 , n11773 );
buf ( n11775 , n11774 );
buf ( n11776 , n11775 );
not ( n11777 , n11521 );
nand ( n11778 , n11777 , n11517 );
not ( n11779 , n11778 );
not ( n11780 , n11537 );
or ( n11781 , n11779 , n11780 );
buf ( n11782 , n11517 );
not ( n11783 , n11782 );
buf ( n11784 , n11521 );
nand ( n11785 , n11783 , n11784 );
buf ( n11786 , n11785 );
nand ( n11787 , n11781 , n11786 );
buf ( n11788 , n11787 );
not ( n11789 , n11354 );
not ( n11790 , n10922 );
or ( n11791 , n11789 , n11790 );
buf ( n11792 , n1557 );
buf ( n11793 , n790 );
buf ( n11794 , n802 );
xor ( n11795 , n11793 , n11794 );
buf ( n11796 , n11795 );
buf ( n11797 , n11796 );
nand ( n11798 , n11792 , n11797 );
buf ( n11799 , n11798 );
nand ( n11800 , n11791 , n11799 );
buf ( n11801 , n1737 );
not ( n11802 , n11801 );
buf ( n11803 , n11802 );
buf ( n11804 , n11803 );
not ( n11805 , n11804 );
buf ( n11806 , n11320 );
not ( n11807 , n11806 );
buf ( n11808 , n11807 );
buf ( n11809 , n11808 );
not ( n11810 , n11809 );
and ( n11811 , n11805 , n11810 );
buf ( n11812 , n1433 );
xor ( n11813 , n804 , n788 );
buf ( n11814 , n11813 );
and ( n11815 , n11812 , n11814 );
buf ( n11816 , n11815 );
buf ( n11817 , n11816 );
nor ( n11818 , n11811 , n11817 );
buf ( n11819 , n11818 );
not ( n11820 , n11819 );
xor ( n11821 , n11800 , n11820 );
buf ( n11822 , n11408 );
not ( n11823 , n11822 );
buf ( n11824 , n2526 );
not ( n11825 , n11824 );
or ( n11826 , n11823 , n11825 );
buf ( n11827 , n2010 );
buf ( n11828 , n776 );
buf ( n11829 , n816 );
xor ( n11830 , n11828 , n11829 );
buf ( n11831 , n11830 );
buf ( n11832 , n11831 );
nand ( n11833 , n11827 , n11832 );
buf ( n11834 , n11833 );
buf ( n11835 , n11834 );
nand ( n11836 , n11826 , n11835 );
buf ( n11837 , n11836 );
xnor ( n11838 , n11821 , n11837 );
not ( n11839 , n10452 );
not ( n11840 , n3656 );
or ( n11841 , n11839 , n11840 );
buf ( n11842 , n3662 );
xor ( n11843 , n800 , n792 );
buf ( n11844 , n11843 );
nand ( n11845 , n11842 , n11844 );
buf ( n11846 , n11845 );
nand ( n11847 , n11841 , n11846 );
buf ( n11848 , n794 );
buf ( n11849 , n800 );
and ( n11850 , n11848 , n11849 );
buf ( n11851 , n11850 );
or ( n11852 , n11847 , n11851 );
buf ( n11853 , n11847 );
buf ( n11854 , n11851 );
nand ( n11855 , n11853 , n11854 );
buf ( n11856 , n11855 );
nand ( n11857 , n11852 , n11856 );
buf ( n11858 , n11337 );
not ( n11859 , n11858 );
buf ( n11860 , n3703 );
not ( n11861 , n11860 );
or ( n11862 , n11859 , n11861 );
buf ( n11863 , n1940 );
buf ( n11864 , n778 );
buf ( n11865 , n814 );
xor ( n11866 , n11864 , n11865 );
buf ( n11867 , n11866 );
buf ( n11868 , n11867 );
nand ( n11869 , n11863 , n11868 );
buf ( n11870 , n11869 );
buf ( n11871 , n11870 );
nand ( n11872 , n11862 , n11871 );
buf ( n11873 , n11872 );
xor ( n11874 , n11857 , n11873 );
xor ( n11875 , n11838 , n11874 );
buf ( n11876 , n2361 );
not ( n11877 , n11876 );
buf ( n11878 , n2371 );
not ( n11879 , n11878 );
or ( n11880 , n11877 , n11879 );
buf ( n11881 , n826 );
nand ( n11882 , n11880 , n11881 );
buf ( n11883 , n11882 );
buf ( n11884 , n11228 );
not ( n11885 , n11884 );
buf ( n11886 , n2267 );
not ( n11887 , n11886 );
or ( n11888 , n11885 , n11887 );
buf ( n11889 , n1346 );
buf ( n11890 , n772 );
buf ( n11891 , n820 );
xor ( n11892 , n11890 , n11891 );
buf ( n11893 , n11892 );
buf ( n11894 , n11893 );
nand ( n11895 , n11889 , n11894 );
buf ( n11896 , n11895 );
buf ( n11897 , n11896 );
nand ( n11898 , n11888 , n11897 );
buf ( n11899 , n11898 );
xnor ( n11900 , n11883 , n11899 );
buf ( n11901 , n11900 );
buf ( n11902 , n11196 );
not ( n11903 , n11902 );
buf ( n11904 , n2790 );
not ( n11905 , n11904 );
or ( n11906 , n11903 , n11905 );
buf ( n11907 , n8354 );
buf ( n11908 , n768 );
buf ( n11909 , n824 );
xor ( n11910 , n11908 , n11909 );
buf ( n11911 , n11910 );
buf ( n11912 , n11911 );
nand ( n11913 , n11907 , n11912 );
buf ( n11914 , n11913 );
buf ( n11915 , n11914 );
nand ( n11916 , n11906 , n11915 );
buf ( n11917 , n11916 );
buf ( n11918 , n11917 );
and ( n11919 , n11901 , n11918 );
not ( n11920 , n11901 );
buf ( n11921 , n11917 );
not ( n11922 , n11921 );
buf ( n11923 , n11922 );
buf ( n11924 , n11923 );
and ( n11925 , n11920 , n11924 );
or ( n11926 , n11919 , n11925 );
buf ( n11927 , n11926 );
xor ( n11928 , n11875 , n11927 );
buf ( n11929 , n11928 );
xor ( n11930 , n11788 , n11929 );
xor ( n11931 , n10441 , n10459 );
and ( n11932 , n11931 , n10480 );
and ( n11933 , n10441 , n10459 );
or ( n11934 , n11932 , n11933 );
buf ( n11935 , n11934 );
buf ( n11936 , n11935 );
buf ( n11937 , n11270 );
not ( n11938 , n11937 );
buf ( n11939 , n2235 );
not ( n11940 , n11939 );
or ( n11941 , n11938 , n11940 );
buf ( n11942 , n1309 );
buf ( n11943 , n784 );
buf ( n11944 , n808 );
xor ( n11945 , n11943 , n11944 );
buf ( n11946 , n11945 );
buf ( n11947 , n11946 );
nand ( n11948 , n11942 , n11947 );
buf ( n11949 , n11948 );
buf ( n11950 , n11949 );
nand ( n11951 , n11941 , n11950 );
buf ( n11952 , n11951 );
buf ( n11953 , n11386 );
not ( n11954 , n11953 );
buf ( n11955 , n2098 );
not ( n11956 , n11955 );
or ( n11957 , n11954 , n11956 );
buf ( n11958 , n2107 );
xor ( n11959 , n822 , n770 );
buf ( n11960 , n11959 );
nand ( n11961 , n11958 , n11960 );
buf ( n11962 , n11961 );
buf ( n11963 , n11962 );
nand ( n11964 , n11957 , n11963 );
buf ( n11965 , n11964 );
xor ( n11966 , n11952 , n11965 );
buf ( n11967 , n11371 );
not ( n11968 , n11967 );
buf ( n11969 , n1403 );
not ( n11970 , n11969 );
or ( n11971 , n11968 , n11970 );
buf ( n11972 , n2331 );
xor ( n11973 , n806 , n786 );
buf ( n11974 , n11973 );
nand ( n11975 , n11972 , n11974 );
buf ( n11976 , n11975 );
buf ( n11977 , n11976 );
nand ( n11978 , n11971 , n11977 );
buf ( n11979 , n11978 );
xor ( n11980 , n11966 , n11979 );
buf ( n11981 , n11980 );
xor ( n11982 , n11936 , n11981 );
xor ( n11983 , n11015 , n11030 );
and ( n11984 , n11983 , n11078 );
and ( n11985 , n11015 , n11030 );
or ( n11986 , n11984 , n11985 );
buf ( n11987 , n11986 );
buf ( n11988 , n11987 );
xor ( n11989 , n11982 , n11988 );
buf ( n11990 , n11989 );
buf ( n11991 , n11990 );
xor ( n11992 , n11930 , n11991 );
buf ( n11993 , n11992 );
buf ( n11994 , n11993 );
xor ( n11995 , n11776 , n11994 );
xor ( n11996 , n10483 , n10579 );
xor ( n11997 , n11996 , n10794 );
buf ( n11998 , n11997 );
buf ( n11999 , n11998 );
xor ( n12000 , n11002 , n11081 );
xor ( n12001 , n12000 , n11241 );
buf ( n12002 , n12001 );
buf ( n12003 , n12002 );
or ( n12004 , n11999 , n12003 );
buf ( n12005 , n4072 );
not ( n12006 , n12005 );
buf ( n12007 , n2325 );
not ( n12008 , n12007 );
or ( n12009 , n12006 , n12008 );
buf ( n12010 , n2982 );
buf ( n12011 , n10721 );
nand ( n12012 , n12010 , n12011 );
buf ( n12013 , n12012 );
buf ( n12014 , n12013 );
nand ( n12015 , n12009 , n12014 );
buf ( n12016 , n12015 );
buf ( n12017 , n12016 );
buf ( n12018 , n4090 );
not ( n12019 , n12018 );
buf ( n12020 , n1480 );
not ( n12021 , n12020 );
or ( n12022 , n12019 , n12021 );
buf ( n12023 , n1496 );
buf ( n12024 , n10764 );
nand ( n12025 , n12023 , n12024 );
buf ( n12026 , n12025 );
buf ( n12027 , n12026 );
nand ( n12028 , n12022 , n12027 );
buf ( n12029 , n12028 );
buf ( n12030 , n12029 );
xor ( n12031 , n12017 , n12030 );
buf ( n12032 , n4206 );
not ( n12033 , n12032 );
buf ( n12034 , n1440 );
not ( n12035 , n12034 );
or ( n12036 , n12033 , n12035 );
buf ( n12037 , n1528 );
buf ( n12038 , n10742 );
nand ( n12039 , n12037 , n12038 );
buf ( n12040 , n12039 );
buf ( n12041 , n12040 );
nand ( n12042 , n12036 , n12041 );
buf ( n12043 , n12042 );
buf ( n12044 , n12043 );
and ( n12045 , n12031 , n12044 );
and ( n12046 , n12017 , n12030 );
or ( n12047 , n12045 , n12046 );
buf ( n12048 , n12047 );
buf ( n12049 , n12048 );
xor ( n12050 , n10937 , n10954 );
xor ( n12051 , n12050 , n10976 );
buf ( n12052 , n12051 );
buf ( n12053 , n12052 );
xor ( n12054 , n12049 , n12053 );
xor ( n12055 , n10612 , n10600 );
xor ( n12056 , n12055 , n10638 );
buf ( n12057 , n12056 );
and ( n12058 , n12054 , n12057 );
and ( n12059 , n12049 , n12053 );
or ( n12060 , n12058 , n12059 );
buf ( n12061 , n12060 );
not ( n12062 , n12061 );
buf ( n12063 , n12062 );
not ( n12064 , n12063 );
buf ( n12065 , n10644 );
buf ( n12066 , n10715 );
and ( n12067 , n12065 , n12066 );
not ( n12068 , n12065 );
buf ( n12069 , n10715 );
not ( n12070 , n12069 );
buf ( n12071 , n12070 );
buf ( n12072 , n12071 );
and ( n12073 , n12068 , n12072 );
nor ( n12074 , n12067 , n12073 );
buf ( n12075 , n12074 );
buf ( n12076 , n12075 );
buf ( n12077 , n10782 );
not ( n12078 , n12077 );
buf ( n12079 , n12078 );
buf ( n12080 , n12079 );
and ( n12081 , n12076 , n12080 );
not ( n12082 , n12076 );
buf ( n12083 , n10782 );
and ( n12084 , n12082 , n12083 );
nor ( n12085 , n12081 , n12084 );
buf ( n12086 , n12085 );
buf ( n12087 , n12086 );
not ( n12088 , n12087 );
or ( n12089 , n12064 , n12088 );
xor ( n12090 , n10526 , n10547 );
xor ( n12091 , n12090 , n10569 );
buf ( n12092 , n12091 );
buf ( n12093 , n12092 );
xor ( n12094 , n10738 , n10759 );
xor ( n12095 , n12094 , n10778 );
buf ( n12096 , n12095 );
buf ( n12097 , n12096 );
xor ( n12098 , n12093 , n12097 );
buf ( n12099 , n10709 );
not ( n12100 , n12099 );
buf ( n12101 , n12100 );
xor ( n12102 , n10688 , n12101 );
xnor ( n12103 , n12102 , n10665 );
buf ( n12104 , n12103 );
and ( n12105 , n12098 , n12104 );
and ( n12106 , n12093 , n12097 );
or ( n12107 , n12105 , n12106 );
buf ( n12108 , n12107 );
buf ( n12109 , n12108 );
nand ( n12110 , n12089 , n12109 );
buf ( n12111 , n12110 );
buf ( n12112 , n12111 );
buf ( n12113 , n12086 );
not ( n12114 , n12113 );
buf ( n12115 , n12061 );
nand ( n12116 , n12114 , n12115 );
buf ( n12117 , n12116 );
buf ( n12118 , n12117 );
nand ( n12119 , n12112 , n12118 );
buf ( n12120 , n12119 );
buf ( n12121 , n12120 );
nand ( n12122 , n12004 , n12121 );
buf ( n12123 , n12122 );
buf ( n12124 , n12123 );
buf ( n12125 , n12002 );
buf ( n12126 , n11998 );
nand ( n12127 , n12125 , n12126 );
buf ( n12128 , n12127 );
buf ( n12129 , n12128 );
nand ( n12130 , n12124 , n12129 );
buf ( n12131 , n12130 );
buf ( n12132 , n12131 );
xor ( n12133 , n11995 , n12132 );
buf ( n12134 , n12133 );
buf ( n12135 , n12134 );
xor ( n12136 , n11484 , n12135 );
buf ( n12137 , n10980 );
not ( n12138 , n12137 );
buf ( n12139 , n10841 );
not ( n12140 , n12139 );
and ( n12141 , n12138 , n12140 );
buf ( n12142 , n10980 );
buf ( n12143 , n10990 );
and ( n12144 , n12142 , n12143 );
nor ( n12145 , n12141 , n12144 );
buf ( n12146 , n12145 );
buf ( n12147 , n12146 );
buf ( n12148 , n10995 );
buf ( n12149 , n12148 );
buf ( n12150 , n12149 );
buf ( n12151 , n12150 );
xnor ( n12152 , n12147 , n12151 );
buf ( n12153 , n12152 );
buf ( n12154 , n12153 );
xor ( n12155 , n11488 , n11492 );
xor ( n12156 , n12155 , n11504 );
buf ( n12157 , n12156 );
buf ( n12158 , n12157 );
xor ( n12159 , n12154 , n12158 );
xor ( n12160 , n11606 , n11610 );
xor ( n12161 , n12160 , n11760 );
buf ( n12162 , n12161 );
buf ( n12163 , n12162 );
and ( n12164 , n12159 , n12163 );
and ( n12165 , n12154 , n12158 );
or ( n12166 , n12164 , n12165 );
buf ( n12167 , n12166 );
buf ( n12168 , n12167 );
xor ( n12169 , n11508 , n11544 );
xnor ( n12170 , n12169 , n11764 );
buf ( n12171 , n12170 );
xor ( n12172 , n12168 , n12171 );
buf ( n12173 , n11591 );
not ( n12174 , n12173 );
buf ( n12175 , n10499 );
not ( n12176 , n12175 );
buf ( n12177 , n11599 );
not ( n12178 , n12177 );
and ( n12179 , n12176 , n12178 );
buf ( n12180 , n10499 );
buf ( n12181 , n11599 );
and ( n12182 , n12180 , n12181 );
nor ( n12183 , n12179 , n12182 );
buf ( n12184 , n12183 );
buf ( n12185 , n12184 );
not ( n12186 , n12185 );
and ( n12187 , n12174 , n12186 );
buf ( n12188 , n11591 );
buf ( n12189 , n12184 );
and ( n12190 , n12188 , n12189 );
nor ( n12191 , n12187 , n12190 );
buf ( n12192 , n12191 );
buf ( n12193 , n12192 );
not ( n12194 , n12193 );
buf ( n12195 , n12194 );
buf ( n12196 , n12195 );
not ( n12197 , n12196 );
xor ( n12198 , n11717 , n11730 );
xor ( n12199 , n12198 , n11744 );
buf ( n12200 , n12199 );
buf ( n12201 , n12200 );
buf ( n12202 , n12201 );
buf ( n12203 , n11636 );
not ( n12204 , n12203 );
buf ( n12205 , n11650 );
not ( n12206 , n12205 );
buf ( n12207 , n12206 );
buf ( n12208 , n12207 );
not ( n12209 , n12208 );
or ( n12210 , n12204 , n12209 );
buf ( n12211 , n12207 );
buf ( n12212 , n11636 );
or ( n12213 , n12211 , n12212 );
nand ( n12214 , n12210 , n12213 );
buf ( n12215 , n12214 );
xor ( n12216 , n12215 , n11623 );
buf ( n12217 , n12216 );
or ( n12218 , n12202 , n12217 );
xnor ( n12219 , n11671 , n11699 );
not ( n12220 , n11684 );
and ( n12221 , n12219 , n12220 );
not ( n12222 , n12219 );
and ( n12223 , n12222 , n11684 );
nor ( n12224 , n12221 , n12223 );
buf ( n12225 , n12224 );
nand ( n12226 , n12218 , n12225 );
buf ( n12227 , n12226 );
buf ( n12228 , n12227 );
buf ( n12229 , n12216 );
buf ( n12230 , n12201 );
nand ( n12231 , n12229 , n12230 );
buf ( n12232 , n12231 );
buf ( n12233 , n12232 );
nand ( n12234 , n12228 , n12233 );
buf ( n12235 , n12234 );
buf ( n12236 , n12235 );
not ( n12237 , n12236 );
or ( n12238 , n12197 , n12237 );
buf ( n12239 , n12192 );
not ( n12240 , n12239 );
buf ( n12241 , n12235 );
not ( n12242 , n12241 );
buf ( n12243 , n12242 );
buf ( n12244 , n12243 );
not ( n12245 , n12244 );
or ( n12246 , n12240 , n12245 );
or ( n12247 , n4003 , n3990 );
not ( n12248 , n12247 );
not ( n12249 , n4032 );
or ( n12250 , n12248 , n12249 );
nand ( n12251 , n4009 , n3990 );
nand ( n12252 , n12250 , n12251 );
buf ( n12253 , n12252 );
not ( n12254 , n12253 );
xor ( n12255 , n12017 , n12030 );
xor ( n12256 , n12255 , n12044 );
buf ( n12257 , n12256 );
buf ( n12258 , n12257 );
not ( n12259 , n12258 );
or ( n12260 , n12254 , n12259 );
buf ( n12261 , n12252 );
buf ( n12262 , n12257 );
or ( n12263 , n12261 , n12262 );
xor ( n12264 , n11560 , n11573 );
xor ( n12265 , n12264 , n11587 );
buf ( n12266 , n12265 );
buf ( n12267 , n12266 );
nand ( n12268 , n12263 , n12267 );
buf ( n12269 , n12268 );
buf ( n12270 , n12269 );
nand ( n12271 , n12260 , n12270 );
buf ( n12272 , n12271 );
buf ( n12273 , n12272 );
nand ( n12274 , n12246 , n12273 );
buf ( n12275 , n12274 );
buf ( n12276 , n12275 );
nand ( n12277 , n12238 , n12276 );
buf ( n12278 , n12277 );
not ( n12279 , n12278 );
buf ( n12280 , n11599 );
not ( n12281 , n12280 );
buf ( n12282 , n4190 );
not ( n12283 , n12282 );
buf ( n12284 , n1551 );
not ( n12285 , n12284 );
or ( n12286 , n12283 , n12285 );
buf ( n12287 , n1560 );
buf ( n12288 , n10905 );
nand ( n12289 , n12287 , n12288 );
buf ( n12290 , n12289 );
buf ( n12291 , n12290 );
nand ( n12292 , n12286 , n12291 );
buf ( n12293 , n12292 );
buf ( n12294 , n12293 );
not ( n12295 , n12294 );
buf ( n12296 , n12295 );
buf ( n12297 , n12296 );
not ( n12298 , n12297 );
or ( n12299 , n12281 , n12298 );
xor ( n12300 , n3823 , n3836 );
and ( n12301 , n12300 , n3857 );
and ( n12302 , n3823 , n3836 );
or ( n12303 , n12301 , n12302 );
buf ( n12304 , n12303 );
buf ( n12305 , n12304 );
nand ( n12306 , n12299 , n12305 );
buf ( n12307 , n12306 );
buf ( n12308 , n12307 );
buf ( n12309 , n12293 );
buf ( n12310 , n830 );
nand ( n12311 , n12309 , n12310 );
buf ( n12312 , n12311 );
buf ( n12313 , n12312 );
nand ( n12314 , n12308 , n12313 );
buf ( n12315 , n12314 );
buf ( n12316 , n12315 );
xor ( n12317 , n4248 , n4265 );
and ( n12318 , n12317 , n4280 );
and ( n12319 , n4248 , n4265 );
or ( n12320 , n12318 , n12319 );
buf ( n12321 , n12320 );
buf ( n12322 , n12321 );
xor ( n12323 , n4062 , n4079 );
and ( n12324 , n12323 , n4097 );
and ( n12325 , n4062 , n4079 );
or ( n12326 , n12324 , n12325 );
buf ( n12327 , n12326 );
buf ( n12328 , n12327 );
xor ( n12329 , n12322 , n12328 );
buf ( n12330 , n3940 );
not ( n12331 , n12330 );
buf ( n12332 , n3914 );
not ( n12333 , n12332 );
buf ( n12334 , n12333 );
buf ( n12335 , n12334 );
not ( n12336 , n12335 );
or ( n12337 , n12331 , n12336 );
buf ( n12338 , n3964 );
nand ( n12339 , n12337 , n12338 );
buf ( n12340 , n12339 );
buf ( n12341 , n12340 );
buf ( n12342 , n3914 );
buf ( n12343 , n3937 );
nand ( n12344 , n12342 , n12343 );
buf ( n12345 , n12344 );
buf ( n12346 , n12345 );
nand ( n12347 , n12341 , n12346 );
buf ( n12348 , n12347 );
buf ( n12349 , n12348 );
and ( n12350 , n12329 , n12349 );
and ( n12351 , n12322 , n12328 );
or ( n12352 , n12350 , n12351 );
buf ( n12353 , n12352 );
buf ( n12354 , n12353 );
xor ( n12355 , n12316 , n12354 );
xor ( n12356 , n11701 , n11658 );
xor ( n12357 , n12356 , n11748 );
buf ( n12358 , n12357 );
and ( n12359 , n12355 , n12358 );
and ( n12360 , n12316 , n12354 );
or ( n12361 , n12359 , n12360 );
buf ( n12362 , n12361 );
not ( n12363 , n12362 );
or ( n12364 , n12279 , n12363 );
buf ( n12365 , n12086 );
not ( n12366 , n12365 );
buf ( n12367 , n12108 );
not ( n12368 , n12367 );
or ( n12369 , n12366 , n12368 );
buf ( n12370 , n12108 );
buf ( n12371 , n12086 );
or ( n12372 , n12370 , n12371 );
nand ( n12373 , n12369 , n12372 );
buf ( n12374 , n12373 );
buf ( n12375 , n12374 );
buf ( n12376 , n12061 );
buf ( n12377 , n12376 );
and ( n12378 , n12375 , n12377 );
not ( n12379 , n12375 );
not ( n12380 , n12376 );
buf ( n12381 , n12380 );
and ( n12382 , n12379 , n12381 );
nor ( n12383 , n12378 , n12382 );
buf ( n12384 , n12383 );
not ( n12385 , n12384 );
nor ( n12386 , n12278 , n12362 );
or ( n12387 , n12385 , n12386 );
nand ( n12388 , n12364 , n12387 );
buf ( n12389 , n12388 );
and ( n12390 , n12172 , n12389 );
and ( n12391 , n12168 , n12171 );
or ( n12392 , n12390 , n12391 );
buf ( n12393 , n12392 );
buf ( n12394 , n12393 );
xor ( n12395 , n12136 , n12394 );
buf ( n12396 , n12395 );
buf ( n12397 , n11998 );
not ( n12398 , n12397 );
buf ( n12399 , n12398 );
buf ( n12400 , n12399 );
not ( n12401 , n12400 );
buf ( n12402 , n12120 );
not ( n12403 , n12402 );
and ( n12404 , n12401 , n12403 );
buf ( n12405 , n12120 );
buf ( n12406 , n12399 );
and ( n12407 , n12405 , n12406 );
nor ( n12408 , n12404 , n12407 );
buf ( n12409 , n12408 );
not ( n12410 , n12409 );
xor ( n12411 , n12002 , n12410 );
buf ( n12412 , n12411 );
xor ( n12413 , n12049 , n12053 );
xor ( n12414 , n12413 , n12057 );
buf ( n12415 , n12414 );
xor ( n12416 , n12093 , n12097 );
xor ( n12417 , n12416 , n12104 );
buf ( n12418 , n12417 );
xor ( n12419 , n12415 , n12418 );
buf ( n12420 , n3974 );
not ( n12421 , n12420 );
buf ( n12422 , n4039 );
not ( n12423 , n12422 );
or ( n12424 , n12421 , n12423 );
buf ( n12425 , n4099 );
nand ( n12426 , n12424 , n12425 );
buf ( n12427 , n12426 );
buf ( n12428 , n12427 );
buf ( n12429 , n3974 );
not ( n12430 , n12429 );
buf ( n12431 , n4042 );
nand ( n12432 , n12430 , n12431 );
buf ( n12433 , n12432 );
buf ( n12434 , n12433 );
nand ( n12435 , n12428 , n12434 );
buf ( n12436 , n12435 );
buf ( n12437 , n12436 );
buf ( n12438 , n12293 );
not ( n12439 , n12438 );
buf ( n12440 , n11599 );
not ( n12441 , n12440 );
and ( n12442 , n12439 , n12441 );
buf ( n12443 , n12293 );
buf ( n12444 , n11599 );
and ( n12445 , n12443 , n12444 );
nor ( n12446 , n12442 , n12445 );
buf ( n12447 , n12446 );
xnor ( n12448 , n12304 , n12447 );
buf ( n12449 , n12448 );
or ( n12450 , n12437 , n12449 );
xor ( n12451 , n12322 , n12328 );
xor ( n12452 , n12451 , n12349 );
buf ( n12453 , n12452 );
buf ( n12454 , n12453 );
nand ( n12455 , n12450 , n12454 );
buf ( n12456 , n12455 );
buf ( n12457 , n12456 );
buf ( n12458 , n12436 );
buf ( n12459 , n12448 );
nand ( n12460 , n12458 , n12459 );
buf ( n12461 , n12460 );
buf ( n12462 , n12461 );
nand ( n12463 , n12457 , n12462 );
buf ( n12464 , n12463 );
and ( n12465 , n12419 , n12464 );
and ( n12466 , n12415 , n12418 );
or ( n12467 , n12465 , n12466 );
xor ( n12468 , n12154 , n12158 );
xor ( n12469 , n12468 , n12163 );
buf ( n12470 , n12469 );
xor ( n12471 , n12467 , n12470 );
xor ( n12472 , n12316 , n12354 );
xor ( n12473 , n12472 , n12358 );
buf ( n12474 , n12473 );
not ( n12475 , n12474 );
buf ( n12476 , n4212 );
not ( n12477 , n12476 );
buf ( n12478 , n12477 );
buf ( n12479 , n12478 );
not ( n12480 , n12479 );
buf ( n12481 , n4218 );
not ( n12482 , n12481 );
or ( n12483 , n12480 , n12482 );
buf ( n12484 , n4196 );
nand ( n12485 , n12483 , n12484 );
buf ( n12486 , n12485 );
buf ( n12487 , n12486 );
buf ( n12488 , n4223 );
buf ( n12489 , n4212 );
nand ( n12490 , n12488 , n12489 );
buf ( n12491 , n12490 );
buf ( n12492 , n12491 );
nand ( n12493 , n12487 , n12492 );
buf ( n12494 , n12493 );
not ( n12495 , n12494 );
buf ( n12496 , n3859 );
not ( n12497 , n12496 );
buf ( n12498 , n3874 );
not ( n12499 , n12498 );
or ( n12500 , n12497 , n12499 );
buf ( n12501 , n3874 );
buf ( n12502 , n3859 );
or ( n12503 , n12501 , n12502 );
buf ( n12504 , n12503 );
buf ( n12505 , n12504 );
buf ( n12506 , n3881 );
nand ( n12507 , n12505 , n12506 );
buf ( n12508 , n12507 );
buf ( n12509 , n12508 );
nand ( n12510 , n12500 , n12509 );
buf ( n12511 , n12510 );
not ( n12512 , n12511 );
or ( n12513 , n12495 , n12512 );
not ( n12514 , n12494 );
not ( n12515 , n12514 );
not ( n12516 , n12511 );
not ( n12517 , n12516 );
or ( n12518 , n12515 , n12517 );
buf ( n12519 , n4132 );
not ( n12520 , n12519 );
buf ( n12521 , n12520 );
buf ( n12522 , n12521 );
not ( n12523 , n12522 );
buf ( n12524 , n4149 );
not ( n12525 , n12524 );
or ( n12526 , n12523 , n12525 );
buf ( n12527 , n4155 );
nand ( n12528 , n12526 , n12527 );
buf ( n12529 , n12528 );
buf ( n12530 , n12529 );
buf ( n12531 , n4132 );
buf ( n12532 , n4146 );
nand ( n12533 , n12531 , n12532 );
buf ( n12534 , n12533 );
buf ( n12535 , n12534 );
nand ( n12536 , n12530 , n12535 );
buf ( n12537 , n12536 );
nand ( n12538 , n12518 , n12537 );
nand ( n12539 , n12513 , n12538 );
not ( n12540 , n12539 );
or ( n12541 , n12475 , n12540 );
nor ( n12542 , n12474 , n12539 );
buf ( n12543 , n12192 );
not ( n12544 , n12543 );
buf ( n12545 , n12272 );
not ( n12546 , n12545 );
or ( n12547 , n12544 , n12546 );
buf ( n12548 , n12272 );
buf ( n12549 , n12192 );
or ( n12550 , n12548 , n12549 );
nand ( n12551 , n12547 , n12550 );
buf ( n12552 , n12551 );
buf ( n12553 , n12552 );
buf ( n12554 , n12235 );
buf ( n12555 , n12554 );
buf ( n12556 , n12555 );
buf ( n12557 , n12556 );
xnor ( n12558 , n12553 , n12557 );
buf ( n12559 , n12558 );
or ( n12560 , n12542 , n12559 );
nand ( n12561 , n12541 , n12560 );
and ( n12562 , n12471 , n12561 );
and ( n12563 , n12467 , n12470 );
or ( n12564 , n12562 , n12563 );
buf ( n12565 , n12564 );
xor ( n12566 , n12412 , n12565 );
xor ( n12567 , n12168 , n12171 );
xor ( n12568 , n12567 , n12389 );
buf ( n12569 , n12568 );
buf ( n12570 , n12569 );
and ( n12571 , n12566 , n12570 );
and ( n12572 , n12412 , n12565 );
or ( n12573 , n12571 , n12572 );
buf ( n12574 , n12573 );
xor ( n12575 , n12396 , n12574 );
not ( n12576 , n12575 );
xor ( n12577 , n12514 , n12511 );
not ( n12578 , n12537 );
xnor ( n12579 , n12577 , n12578 );
not ( n12580 , n12579 );
buf ( n12581 , n3817 );
not ( n12582 , n12581 );
buf ( n12583 , n3884 );
not ( n12584 , n12583 );
or ( n12585 , n12582 , n12584 );
buf ( n12586 , n3894 );
nand ( n12587 , n12585 , n12586 );
buf ( n12588 , n12587 );
buf ( n12589 , n3887 );
buf ( n12590 , n3814 );
nand ( n12591 , n12589 , n12590 );
buf ( n12592 , n12591 );
nand ( n12593 , n12588 , n12592 );
not ( n12594 , n12593 );
not ( n12595 , n12594 );
or ( n12596 , n12580 , n12595 );
xor ( n12597 , n12453 , n12448 );
xor ( n12598 , n12597 , n12436 );
nand ( n12599 , n12596 , n12598 );
buf ( n12600 , n12599 );
not ( n12601 , n12579 );
nand ( n12602 , n12593 , n12601 );
buf ( n12603 , n12602 );
nand ( n12604 , n12600 , n12603 );
buf ( n12605 , n12604 );
buf ( n12606 , n12605 );
not ( n12607 , n12606 );
xor ( n12608 , n12415 , n12418 );
xor ( n12609 , n12608 , n12464 );
buf ( n12610 , n12609 );
buf ( n12611 , n12610 );
not ( n12612 , n12611 );
buf ( n12613 , n12612 );
buf ( n12614 , n12613 );
not ( n12615 , n12220 );
not ( n12616 , n12219 );
and ( n12617 , n12615 , n12616 );
and ( n12618 , n12220 , n12219 );
nor ( n12619 , n12617 , n12618 );
not ( n12620 , n12619 );
not ( n12621 , n12200 );
not ( n12622 , n12621 );
or ( n12623 , n12620 , n12622 );
or ( n12624 , n12619 , n12621 );
nand ( n12625 , n12623 , n12624 );
buf ( n12626 , n12625 );
buf ( n12627 , n12216 );
not ( n12628 , n12627 );
buf ( n12629 , n12628 );
buf ( n12630 , n12629 );
and ( n12631 , n12626 , n12630 );
not ( n12632 , n12626 );
buf ( n12633 , n12216 );
and ( n12634 , n12632 , n12633 );
nor ( n12635 , n12631 , n12634 );
buf ( n12636 , n12635 );
buf ( n12637 , n12636 );
not ( n12638 , n12637 );
buf ( n12639 , n12638 );
not ( n12640 , n12639 );
xor ( n12641 , n12252 , n12266 );
xnor ( n12642 , n12641 , n12257 );
buf ( n12643 , n12642 );
not ( n12644 , n12643 );
buf ( n12645 , n12644 );
not ( n12646 , n12645 );
or ( n12647 , n12640 , n12646 );
not ( n12648 , n12642 );
not ( n12649 , n12636 );
or ( n12650 , n12648 , n12649 );
buf ( n12651 , n4178 );
not ( n12652 , n12651 );
buf ( n12653 , n4282 );
not ( n12654 , n12653 );
buf ( n12655 , n4225 );
nand ( n12656 , n12654 , n12655 );
buf ( n12657 , n12656 );
buf ( n12658 , n12657 );
not ( n12659 , n12658 );
or ( n12660 , n12652 , n12659 );
buf ( n12661 , n4225 );
not ( n12662 , n12661 );
buf ( n12663 , n4282 );
nand ( n12664 , n12662 , n12663 );
buf ( n12665 , n12664 );
buf ( n12666 , n12665 );
nand ( n12667 , n12660 , n12666 );
buf ( n12668 , n12667 );
nand ( n12669 , n12650 , n12668 );
nand ( n12670 , n12647 , n12669 );
buf ( n12671 , n12670 );
not ( n12672 , n12671 );
buf ( n12673 , n12672 );
buf ( n12674 , n12673 );
nand ( n12675 , n12614 , n12674 );
buf ( n12676 , n12675 );
buf ( n12677 , n12676 );
not ( n12678 , n12677 );
or ( n12679 , n12607 , n12678 );
buf ( n12680 , n12610 );
buf ( n12681 , n12670 );
nand ( n12682 , n12680 , n12681 );
buf ( n12683 , n12682 );
buf ( n12684 , n12683 );
nand ( n12685 , n12679 , n12684 );
buf ( n12686 , n12685 );
not ( n12687 , n12686 );
xor ( n12688 , n12467 , n12470 );
xor ( n12689 , n12688 , n12561 );
not ( n12690 , n12689 );
and ( n12691 , n12687 , n12690 );
xor ( n12692 , n12278 , n12362 );
and ( n12693 , n12692 , n12384 );
not ( n12694 , n12692 );
and ( n12695 , n12694 , n12385 );
or ( n12696 , n12693 , n12695 );
nor ( n12697 , n12691 , n12696 );
nor ( n12698 , n12687 , n12690 );
nor ( n12699 , n12697 , n12698 );
not ( n12700 , n12699 );
buf ( n12701 , n12700 );
xor ( n12702 , n12412 , n12565 );
xor ( n12703 , n12702 , n12570 );
buf ( n12704 , n12703 );
buf ( n12705 , n12704 );
and ( n12706 , n12701 , n12705 );
buf ( n12707 , n12706 );
not ( n12708 , n12707 );
and ( n12709 , n12576 , n12708 );
and ( n12710 , n12696 , n12686 );
not ( n12711 , n12696 );
not ( n12712 , n12686 );
and ( n12713 , n12711 , n12712 );
nor ( n12714 , n12710 , n12713 );
xor ( n12715 , n12690 , n12714 );
buf ( n12716 , n12715 );
xor ( n12717 , n12539 , n12474 );
buf ( n12718 , n12717 );
buf ( n12719 , n12559 );
not ( n12720 , n12719 );
buf ( n12721 , n12720 );
buf ( n12722 , n12721 );
and ( n12723 , n12718 , n12722 );
not ( n12724 , n12718 );
buf ( n12725 , n12559 );
and ( n12726 , n12724 , n12725 );
nor ( n12727 , n12723 , n12726 );
buf ( n12728 , n12727 );
buf ( n12729 , n12728 );
not ( n12730 , n12729 );
xor ( n12731 , n4110 , n4157 );
and ( n12732 , n12731 , n4164 );
and ( n12733 , n4110 , n4157 );
or ( n12734 , n12732 , n12733 );
buf ( n12735 , n12734 );
buf ( n12736 , n12735 );
buf ( n12737 , n12642 );
buf ( n12738 , n12737 );
buf ( n12739 , n12738 );
buf ( n12740 , n12739 );
buf ( n12741 , n12668 );
not ( n12742 , n12741 );
buf ( n12743 , n12636 );
not ( n12744 , n12743 );
and ( n12745 , n12742 , n12744 );
buf ( n12746 , n12668 );
buf ( n12747 , n12636 );
and ( n12748 , n12746 , n12747 );
nor ( n12749 , n12745 , n12748 );
buf ( n12750 , n12749 );
buf ( n12751 , n12750 );
xor ( n12752 , n12740 , n12751 );
buf ( n12753 , n12752 );
buf ( n12754 , n12753 );
xor ( n12755 , n12736 , n12754 );
xor ( n12756 , n4299 , n4310 );
and ( n12757 , n12756 , n4317 );
and ( n12758 , n4299 , n4310 );
or ( n12759 , n12757 , n12758 );
buf ( n12760 , n12759 );
buf ( n12761 , n12760 );
and ( n12762 , n12755 , n12761 );
and ( n12763 , n12736 , n12754 );
or ( n12764 , n12762 , n12763 );
buf ( n12765 , n12764 );
buf ( n12766 , n12765 );
not ( n12767 , n12766 );
or ( n12768 , n12730 , n12767 );
buf ( n12769 , n12728 );
not ( n12770 , n12769 );
buf ( n12771 , n12770 );
buf ( n12772 , n12771 );
not ( n12773 , n12772 );
buf ( n12774 , n12765 );
not ( n12775 , n12774 );
buf ( n12776 , n12775 );
buf ( n12777 , n12776 );
not ( n12778 , n12777 );
or ( n12779 , n12773 , n12778 );
not ( n12780 , n12670 );
not ( n12781 , n12609 );
not ( n12782 , n12781 );
or ( n12783 , n12780 , n12782 );
nand ( n12784 , n12609 , n12673 );
nand ( n12785 , n12783 , n12784 );
buf ( n12786 , n12785 );
buf ( n12787 , n12599 );
buf ( n12788 , n12602 );
and ( n12789 , n12787 , n12788 );
buf ( n12790 , n12789 );
buf ( n12791 , n12790 );
xor ( n12792 , n12786 , n12791 );
buf ( n12793 , n12792 );
buf ( n12794 , n12793 );
not ( n12795 , n12794 );
buf ( n12796 , n12795 );
buf ( n12797 , n12796 );
nand ( n12798 , n12779 , n12797 );
buf ( n12799 , n12798 );
buf ( n12800 , n12799 );
nand ( n12801 , n12768 , n12800 );
buf ( n12802 , n12801 );
buf ( n12803 , n12802 );
and ( n12804 , n12716 , n12803 );
buf ( n12805 , n12804 );
xor ( n12806 , n12701 , n12705 );
buf ( n12807 , n12806 );
nor ( n12808 , n12805 , n12807 );
nor ( n12809 , n12709 , n12808 );
buf ( n12810 , n12809 );
xor ( n12811 , n11484 , n12135 );
and ( n12812 , n12811 , n12394 );
and ( n12813 , n11484 , n12135 );
or ( n12814 , n12812 , n12813 );
buf ( n12815 , n12814 );
buf ( n12816 , n12815 );
not ( n12817 , n12816 );
buf ( n12818 , n11874 );
not ( n12819 , n12818 );
buf ( n12820 , n11838 );
not ( n12821 , n12820 );
or ( n12822 , n12819 , n12821 );
buf ( n12823 , n11927 );
nand ( n12824 , n12822 , n12823 );
buf ( n12825 , n12824 );
buf ( n12826 , n12825 );
buf ( n12827 , n11874 );
not ( n12828 , n12827 );
not ( n12829 , n11838 );
buf ( n12830 , n12829 );
nand ( n12831 , n12828 , n12830 );
buf ( n12832 , n12831 );
buf ( n12833 , n12832 );
nand ( n12834 , n12826 , n12833 );
buf ( n12835 , n12834 );
buf ( n12836 , n12835 );
not ( n12837 , n11873 );
not ( n12838 , n11851 );
or ( n12839 , n12837 , n12838 );
buf ( n12840 , n11873 );
buf ( n12841 , n11851 );
nor ( n12842 , n12840 , n12841 );
buf ( n12843 , n12842 );
buf ( n12844 , n11847 );
not ( n12845 , n12844 );
buf ( n12846 , n12845 );
or ( n12847 , n12843 , n12846 );
nand ( n12848 , n12839 , n12847 );
buf ( n12849 , n12848 );
buf ( n12850 , n11946 );
not ( n12851 , n12850 );
buf ( n12852 , n1305 );
not ( n12853 , n12852 );
or ( n12854 , n12851 , n12853 );
buf ( n12855 , n1309 );
buf ( n12856 , n783 );
buf ( n12857 , n808 );
xor ( n12858 , n12856 , n12857 );
buf ( n12859 , n12858 );
buf ( n12860 , n12859 );
nand ( n12861 , n12855 , n12860 );
buf ( n12862 , n12861 );
buf ( n12863 , n12862 );
nand ( n12864 , n12854 , n12863 );
buf ( n12865 , n12864 );
buf ( n12866 , n12865 );
buf ( n12867 , n11432 );
not ( n12868 , n12867 );
buf ( n12869 , n1480 );
not ( n12870 , n12869 );
or ( n12871 , n12868 , n12870 );
buf ( n12872 , n1496 );
buf ( n12873 , n773 );
buf ( n12874 , n818 );
xor ( n12875 , n12873 , n12874 );
buf ( n12876 , n12875 );
buf ( n12877 , n12876 );
nand ( n12878 , n12872 , n12877 );
buf ( n12879 , n12878 );
buf ( n12880 , n12879 );
nand ( n12881 , n12871 , n12880 );
buf ( n12882 , n12881 );
buf ( n12883 , n12882 );
xor ( n12884 , n12866 , n12883 );
buf ( n12885 , n11449 );
not ( n12886 , n12885 );
buf ( n12887 , n1667 );
not ( n12888 , n12887 );
buf ( n12889 , n12888 );
buf ( n12890 , n12889 );
not ( n12891 , n12890 );
or ( n12892 , n12886 , n12891 );
buf ( n12893 , n3398 );
buf ( n12894 , n781 );
buf ( n12895 , n810 );
xor ( n12896 , n12894 , n12895 );
buf ( n12897 , n12896 );
buf ( n12898 , n12897 );
nand ( n12899 , n12893 , n12898 );
buf ( n12900 , n12899 );
buf ( n12901 , n12900 );
nand ( n12902 , n12892 , n12901 );
buf ( n12903 , n12902 );
buf ( n12904 , n12903 );
xor ( n12905 , n12884 , n12904 );
buf ( n12906 , n12905 );
buf ( n12907 , n12906 );
xor ( n12908 , n12849 , n12907 );
buf ( n12909 , n793 );
buf ( n12910 , n800 );
and ( n12911 , n12909 , n12910 );
buf ( n12912 , n12911 );
buf ( n12913 , n12912 );
buf ( n12914 , n11843 );
not ( n12915 , n12914 );
buf ( n12916 , n3656 );
not ( n12917 , n12916 );
or ( n12918 , n12915 , n12917 );
buf ( n12919 , n3662 );
buf ( n12920 , n791 );
buf ( n12921 , n800 );
xor ( n12922 , n12920 , n12921 );
buf ( n12923 , n12922 );
buf ( n12924 , n12923 );
nand ( n12925 , n12919 , n12924 );
buf ( n12926 , n12925 );
buf ( n12927 , n12926 );
nand ( n12928 , n12918 , n12927 );
buf ( n12929 , n12928 );
buf ( n12930 , n12929 );
xor ( n12931 , n12913 , n12930 );
buf ( n12932 , n11893 );
not ( n12933 , n12932 );
buf ( n12934 , n2410 );
not ( n12935 , n12934 );
or ( n12936 , n12933 , n12935 );
buf ( n12937 , n771 );
buf ( n12938 , n820 );
xnor ( n12939 , n12937 , n12938 );
buf ( n12940 , n12939 );
buf ( n12941 , n12940 );
not ( n12942 , n12941 );
buf ( n12943 , n1346 );
nand ( n12944 , n12942 , n12943 );
buf ( n12945 , n12944 );
buf ( n12946 , n12945 );
nand ( n12947 , n12936 , n12946 );
buf ( n12948 , n12947 );
buf ( n12949 , n12948 );
xor ( n12950 , n12931 , n12949 );
buf ( n12951 , n12950 );
buf ( n12952 , n12951 );
xor ( n12953 , n12908 , n12952 );
buf ( n12954 , n12953 );
buf ( n12955 , n12954 );
xor ( n12956 , n12836 , n12955 );
xor ( n12957 , n11936 , n11981 );
and ( n12958 , n12957 , n11988 );
and ( n12959 , n11936 , n11981 );
or ( n12960 , n12958 , n12959 );
buf ( n12961 , n12960 );
buf ( n12962 , n12961 );
xor ( n12963 , n12956 , n12962 );
buf ( n12964 , n12963 );
buf ( n12965 , n12964 );
xor ( n12966 , n11788 , n11929 );
and ( n12967 , n12966 , n11991 );
and ( n12968 , n11788 , n11929 );
or ( n12969 , n12967 , n12968 );
buf ( n12970 , n12969 );
buf ( n12971 , n12970 );
xor ( n12972 , n12965 , n12971 );
not ( n12973 , n11911 );
not ( n12974 , n1965 );
or ( n12975 , n12973 , n12974 );
buf ( n12976 , n1859 );
buf ( n12977 , n824 );
nand ( n12978 , n12976 , n12977 );
buf ( n12979 , n12978 );
nand ( n12980 , n12975 , n12979 );
not ( n12981 , n11867 );
not ( n12982 , n3923 );
or ( n12983 , n12981 , n12982 );
buf ( n12984 , n777 );
buf ( n12985 , n814 );
xor ( n12986 , n12984 , n12985 );
buf ( n12987 , n12986 );
nand ( n12988 , n12987 , n1940 );
nand ( n12989 , n12983 , n12988 );
xor ( n12990 , n12980 , n12989 );
buf ( n12991 , n11796 );
not ( n12992 , n12991 );
buf ( n12993 , n10922 );
not ( n12994 , n12993 );
or ( n12995 , n12992 , n12994 );
buf ( n12996 , n1557 );
buf ( n12997 , n789 );
buf ( n12998 , n802 );
xor ( n12999 , n12997 , n12998 );
buf ( n13000 , n12999 );
buf ( n13001 , n13000 );
nand ( n13002 , n12996 , n13001 );
buf ( n13003 , n13002 );
buf ( n13004 , n13003 );
nand ( n13005 , n12995 , n13004 );
buf ( n13006 , n13005 );
xor ( n13007 , n12990 , n13006 );
buf ( n13008 , n13007 );
buf ( n13009 , n11973 );
not ( n13010 , n13009 );
buf ( n13011 , n1403 );
not ( n13012 , n13011 );
or ( n13013 , n13010 , n13012 );
buf ( n13014 , n2982 );
buf ( n13015 , n785 );
buf ( n13016 , n806 );
xor ( n13017 , n13015 , n13016 );
buf ( n13018 , n13017 );
buf ( n13019 , n13018 );
nand ( n13020 , n13014 , n13019 );
buf ( n13021 , n13020 );
buf ( n13022 , n13021 );
nand ( n13023 , n13013 , n13022 );
buf ( n13024 , n13023 );
not ( n13025 , n11831 );
not ( n13026 , n2004 );
or ( n13027 , n13025 , n13026 );
buf ( n13028 , n775 );
buf ( n13029 , n816 );
xor ( n13030 , n13028 , n13029 );
buf ( n13031 , n13030 );
nand ( n13032 , n2535 , n13031 );
nand ( n13033 , n13027 , n13032 );
xor ( n13034 , n13024 , n13033 );
buf ( n13035 , n11813 );
not ( n13036 , n13035 );
buf ( n13037 , n1522 );
not ( n13038 , n13037 );
or ( n13039 , n13036 , n13038 );
buf ( n13040 , n1449 );
xor ( n13041 , n804 , n787 );
buf ( n13042 , n13041 );
nand ( n13043 , n13040 , n13042 );
buf ( n13044 , n13043 );
buf ( n13045 , n13044 );
nand ( n13046 , n13039 , n13045 );
buf ( n13047 , n13046 );
xor ( n13048 , n13034 , n13047 );
buf ( n13049 , n13048 );
xor ( n13050 , n13008 , n13049 );
buf ( n13051 , n11467 );
not ( n13052 , n13051 );
buf ( n13053 , n2066 );
not ( n13054 , n13053 );
or ( n13055 , n13052 , n13054 );
buf ( n13056 , n6446 );
buf ( n13057 , n779 );
buf ( n13058 , n812 );
xor ( n13059 , n13057 , n13058 );
buf ( n13060 , n13059 );
buf ( n13061 , n13060 );
nand ( n13062 , n13056 , n13061 );
buf ( n13063 , n13062 );
buf ( n13064 , n13063 );
nand ( n13065 , n13055 , n13064 );
buf ( n13066 , n13065 );
buf ( n13067 , n13066 );
buf ( n13068 , n11959 );
not ( n13069 , n13068 );
buf ( n13070 , n2101 );
not ( n13071 , n13070 );
or ( n13072 , n13069 , n13071 );
buf ( n13073 , n3745 );
buf ( n13074 , n769 );
buf ( n13075 , n822 );
xor ( n13076 , n13074 , n13075 );
buf ( n13077 , n13076 );
buf ( n13078 , n13077 );
nand ( n13079 , n13073 , n13078 );
buf ( n13080 , n13079 );
buf ( n13081 , n13080 );
nand ( n13082 , n13072 , n13081 );
buf ( n13083 , n13082 );
buf ( n13084 , n13083 );
not ( n13085 , n13084 );
buf ( n13086 , n13085 );
buf ( n13087 , n13086 );
xor ( n13088 , n13067 , n13087 );
buf ( n13089 , n11800 );
not ( n13090 , n13089 );
buf ( n13091 , n13090 );
buf ( n13092 , n13091 );
not ( n13093 , n13092 );
buf ( n13094 , n11819 );
not ( n13095 , n13094 );
or ( n13096 , n13093 , n13095 );
buf ( n13097 , n11837 );
nand ( n13098 , n13096 , n13097 );
buf ( n13099 , n13098 );
buf ( n13100 , n13099 );
nand ( n13101 , n11820 , n11800 );
buf ( n13102 , n13101 );
nand ( n13103 , n13100 , n13102 );
buf ( n13104 , n13103 );
buf ( n13105 , n13104 );
xor ( n13106 , n13088 , n13105 );
buf ( n13107 , n13106 );
buf ( n13108 , n13107 );
xor ( n13109 , n13050 , n13108 );
buf ( n13110 , n13109 );
buf ( n13111 , n13110 );
buf ( n13112 , n11479 );
not ( n13113 , n13112 );
buf ( n13114 , n11304 );
not ( n13115 , n13114 );
or ( n13116 , n13113 , n13115 );
buf ( n13117 , n11304 );
buf ( n13118 , n11479 );
or ( n13119 , n13117 , n13118 );
buf ( n13120 , n11309 );
nand ( n13121 , n13119 , n13120 );
buf ( n13122 , n13121 );
buf ( n13123 , n13122 );
nand ( n13124 , n13116 , n13123 );
buf ( n13125 , n13124 );
buf ( n13126 , n13125 );
xor ( n13127 , n13111 , n13126 );
xor ( n13128 , n11248 , n11295 );
and ( n13129 , n13128 , n11302 );
and ( n13130 , n11248 , n11295 );
or ( n13131 , n13129 , n13130 );
buf ( n13132 , n13131 );
buf ( n13133 , n13132 );
xor ( n13134 , n11361 , n11421 );
and ( n13135 , n13134 , n11477 );
and ( n13136 , n11361 , n11421 );
or ( n13137 , n13135 , n13136 );
buf ( n13138 , n13137 );
buf ( n13139 , n13138 );
xor ( n13140 , n13133 , n13139 );
buf ( n13141 , n11952 );
buf ( n13142 , n11965 );
nand ( n13143 , n13141 , n13142 );
buf ( n13144 , n13143 );
buf ( n13145 , n13144 );
buf ( n13146 , n11952 );
buf ( n13147 , n11965 );
or ( n13148 , n13146 , n13147 );
buf ( n13149 , n11979 );
nand ( n13150 , n13148 , n13149 );
buf ( n13151 , n13150 );
buf ( n13152 , n13151 );
nand ( n13153 , n13145 , n13152 );
buf ( n13154 , n13153 );
buf ( n13155 , n13154 );
buf ( n13156 , n11917 );
not ( n13157 , n13156 );
buf ( n13158 , n11899 );
not ( n13159 , n13158 );
or ( n13160 , n13157 , n13159 );
buf ( n13161 , n11923 );
not ( n13162 , n13161 );
buf ( n13163 , n11899 );
not ( n13164 , n13163 );
buf ( n13165 , n13164 );
buf ( n13166 , n13165 );
not ( n13167 , n13166 );
or ( n13168 , n13162 , n13167 );
buf ( n13169 , n11883 );
nand ( n13170 , n13168 , n13169 );
buf ( n13171 , n13170 );
buf ( n13172 , n13171 );
nand ( n13173 , n13160 , n13172 );
buf ( n13174 , n13173 );
buf ( n13175 , n13174 );
xor ( n13176 , n13155 , n13175 );
xor ( n13177 , n11439 , n11456 );
and ( n13178 , n13177 , n11474 );
and ( n13179 , n11439 , n11456 );
or ( n13180 , n13178 , n13179 );
buf ( n13181 , n13180 );
buf ( n13182 , n13181 );
xor ( n13183 , n13176 , n13182 );
buf ( n13184 , n13183 );
buf ( n13185 , n13184 );
xor ( n13186 , n13140 , n13185 );
buf ( n13187 , n13186 );
buf ( n13188 , n13187 );
xor ( n13189 , n13127 , n13188 );
buf ( n13190 , n13189 );
buf ( n13191 , n13190 );
xor ( n13192 , n12972 , n13191 );
buf ( n13193 , n13192 );
buf ( n13194 , n13193 );
xor ( n13195 , n10799 , n11246 );
and ( n13196 , n13195 , n11481 );
and ( n13197 , n10799 , n11246 );
or ( n13198 , n13196 , n13197 );
buf ( n13199 , n13198 );
buf ( n13200 , n13199 );
not ( n13201 , n13200 );
buf ( n13202 , n13201 );
buf ( n13203 , n13202 );
and ( n13204 , n13194 , n13203 );
not ( n13205 , n13194 );
buf ( n13206 , n13199 );
and ( n13207 , n13205 , n13206 );
nor ( n13208 , n13204 , n13207 );
buf ( n13209 , n13208 );
buf ( n13210 , n13209 );
xor ( n13211 , n11776 , n11994 );
and ( n13212 , n13211 , n12132 );
and ( n13213 , n11776 , n11994 );
or ( n13214 , n13212 , n13213 );
buf ( n13215 , n13214 );
buf ( n13216 , n13215 );
buf ( n13217 , n13216 );
buf ( n13218 , n13217 );
buf ( n13219 , n13218 );
and ( n13220 , n13210 , n13219 );
not ( n13221 , n13210 );
buf ( n13222 , n13218 );
not ( n13223 , n13222 );
buf ( n13224 , n13223 );
buf ( n13225 , n13224 );
and ( n13226 , n13221 , n13225 );
nor ( n13227 , n13220 , n13226 );
buf ( n13228 , n13227 );
not ( n13229 , n13228 );
not ( n13230 , n13229 );
buf ( n13231 , n13230 );
not ( n13232 , n13231 );
or ( n13233 , n12817 , n13232 );
buf ( n13234 , n12815 );
not ( n13235 , n13234 );
buf ( n13236 , n13235 );
buf ( n13237 , n13236 );
buf ( n13238 , n13229 );
nand ( n13239 , n13237 , n13238 );
buf ( n13240 , n13239 );
buf ( n13241 , n13240 );
nand ( n13242 , n13233 , n13241 );
buf ( n13243 , n13242 );
buf ( n13244 , n13243 );
buf ( n13245 , n12396 );
buf ( n13246 , n12574 );
and ( n13247 , n13245 , n13246 );
buf ( n13248 , n13247 );
buf ( n13249 , n13248 );
nor ( n13250 , n13244 , n13249 );
buf ( n13251 , n13250 );
buf ( n13252 , n13251 );
and ( n13253 , n13229 , n12815 );
buf ( n13254 , n13253 );
buf ( n13255 , n13199 );
not ( n13256 , n13255 );
buf ( n13257 , n13215 );
not ( n13258 , n13257 );
or ( n13259 , n13256 , n13258 );
buf ( n13260 , n13202 );
not ( n13261 , n13260 );
buf ( n13262 , n13215 );
not ( n13263 , n13262 );
buf ( n13264 , n13263 );
buf ( n13265 , n13264 );
not ( n13266 , n13265 );
or ( n13267 , n13261 , n13266 );
buf ( n13268 , n13193 );
buf ( n13269 , n13268 );
buf ( n13270 , n13269 );
buf ( n13271 , n13270 );
nand ( n13272 , n13267 , n13271 );
buf ( n13273 , n13272 );
buf ( n13274 , n13273 );
nand ( n13275 , n13259 , n13274 );
buf ( n13276 , n13275 );
not ( n13277 , n13276 );
not ( n13278 , n13277 );
buf ( n13279 , n13278 );
not ( n13280 , n13279 );
xor ( n13281 , n13111 , n13126 );
and ( n13282 , n13281 , n13188 );
and ( n13283 , n13111 , n13126 );
or ( n13284 , n13282 , n13283 );
buf ( n13285 , n13284 );
buf ( n13286 , n13285 );
xor ( n13287 , n12965 , n12971 );
and ( n13288 , n13287 , n13191 );
and ( n13289 , n12965 , n12971 );
or ( n13290 , n13288 , n13289 );
buf ( n13291 , n13290 );
buf ( n13292 , n13291 );
xor ( n13293 , n13286 , n13292 );
xor ( n13294 , n12836 , n12955 );
and ( n13295 , n13294 , n12962 );
and ( n13296 , n12836 , n12955 );
or ( n13297 , n13295 , n13296 );
buf ( n13298 , n13297 );
xor ( n13299 , n12849 , n12907 );
and ( n13300 , n13299 , n12952 );
and ( n13301 , n12849 , n12907 );
or ( n13302 , n13300 , n13301 );
buf ( n13303 , n13302 );
xor ( n13304 , n12913 , n12930 );
and ( n13305 , n13304 , n12949 );
and ( n13306 , n12913 , n12930 );
or ( n13307 , n13305 , n13306 );
buf ( n13308 , n13307 );
buf ( n13309 , n13308 );
buf ( n13310 , n12859 );
not ( n13311 , n13310 );
buf ( n13312 , n2235 );
not ( n13313 , n13312 );
or ( n13314 , n13311 , n13313 );
buf ( n13315 , n1309 );
buf ( n13316 , n782 );
buf ( n13317 , n808 );
xor ( n13318 , n13316 , n13317 );
buf ( n13319 , n13318 );
buf ( n13320 , n13319 );
nand ( n13321 , n13315 , n13320 );
buf ( n13322 , n13321 );
buf ( n13323 , n13322 );
nand ( n13324 , n13314 , n13323 );
buf ( n13325 , n13324 );
buf ( n13326 , n13325 );
buf ( n13327 , n12897 );
not ( n13328 , n13327 );
buf ( n13329 , n2641 );
not ( n13330 , n13329 );
or ( n13331 , n13328 , n13330 );
buf ( n13332 , n1679 );
buf ( n13333 , n780 );
buf ( n13334 , n810 );
xor ( n13335 , n13333 , n13334 );
buf ( n13336 , n13335 );
buf ( n13337 , n13336 );
nand ( n13338 , n13332 , n13337 );
buf ( n13339 , n13338 );
buf ( n13340 , n13339 );
nand ( n13341 , n13331 , n13340 );
buf ( n13342 , n13341 );
buf ( n13343 , n13342 );
xor ( n13344 , n13326 , n13343 );
buf ( n13345 , n7797 );
buf ( n13346 , n13031 );
not ( n13347 , n13346 );
buf ( n13348 , n13347 );
buf ( n13349 , n13348 );
or ( n13350 , n13345 , n13349 );
buf ( n13351 , n2535 );
not ( n13352 , n13351 );
buf ( n13353 , n13352 );
buf ( n13354 , n13353 );
buf ( n13355 , n774 );
buf ( n13356 , n816 );
xor ( n13357 , n13355 , n13356 );
buf ( n13358 , n13357 );
buf ( n13359 , n13358 );
not ( n13360 , n13359 );
buf ( n13361 , n13360 );
buf ( n13362 , n13361 );
or ( n13363 , n13354 , n13362 );
nand ( n13364 , n13350 , n13363 );
buf ( n13365 , n13364 );
buf ( n13366 , n13365 );
xor ( n13367 , n13344 , n13366 );
buf ( n13368 , n13367 );
buf ( n13369 , n13368 );
xor ( n13370 , n13309 , n13369 );
buf ( n13371 , n12876 );
not ( n13372 , n13371 );
buf ( n13373 , n4396 );
not ( n13374 , n13373 );
or ( n13375 , n13372 , n13374 );
buf ( n13376 , n1496 );
buf ( n13377 , n772 );
buf ( n13378 , n818 );
xor ( n13379 , n13377 , n13378 );
buf ( n13380 , n13379 );
buf ( n13381 , n13380 );
nand ( n13382 , n13376 , n13381 );
buf ( n13383 , n13382 );
buf ( n13384 , n13383 );
nand ( n13385 , n13375 , n13384 );
buf ( n13386 , n13385 );
not ( n13387 , n13386 );
buf ( n13388 , n13077 );
not ( n13389 , n13388 );
buf ( n13390 , n2101 );
not ( n13391 , n13390 );
or ( n13392 , n13389 , n13391 );
buf ( n13393 , n3745 );
buf ( n13394 , n768 );
buf ( n13395 , n822 );
xor ( n13396 , n13394 , n13395 );
buf ( n13397 , n13396 );
buf ( n13398 , n13397 );
nand ( n13399 , n13393 , n13398 );
buf ( n13400 , n13399 );
buf ( n13401 , n13400 );
nand ( n13402 , n13392 , n13401 );
buf ( n13403 , n13402 );
not ( n13404 , n13403 );
buf ( n13405 , n3252 );
not ( n13406 , n13405 );
buf ( n13407 , n1841 );
not ( n13408 , n13407 );
or ( n13409 , n13406 , n13408 );
buf ( n13410 , n824 );
nand ( n13411 , n13409 , n13410 );
buf ( n13412 , n13411 );
nand ( n13413 , n13387 , n13404 , n13412 );
not ( n13414 , n13386 );
nor ( n13415 , n13414 , n13412 );
nand ( n13416 , n13404 , n13415 );
nor ( n13417 , n13412 , n13386 );
nand ( n13418 , n13403 , n13417 );
nand ( n13419 , n13412 , n13386 );
not ( n13420 , n13419 );
nand ( n13421 , n13420 , n13403 );
nand ( n13422 , n13413 , n13416 , n13418 , n13421 );
buf ( n13423 , n13422 );
xor ( n13424 , n13370 , n13423 );
buf ( n13425 , n13424 );
xor ( n13426 , n13303 , n13425 );
buf ( n13427 , n12987 );
not ( n13428 , n13427 );
buf ( n13429 , n1931 );
not ( n13430 , n13429 );
or ( n13431 , n13428 , n13430 );
buf ( n13432 , n1940 );
buf ( n13433 , n776 );
buf ( n13434 , n814 );
xor ( n13435 , n13433 , n13434 );
buf ( n13436 , n13435 );
buf ( n13437 , n13436 );
nand ( n13438 , n13432 , n13437 );
buf ( n13439 , n13438 );
buf ( n13440 , n13439 );
nand ( n13441 , n13431 , n13440 );
buf ( n13442 , n13441 );
buf ( n13443 , n13442 );
not ( n13444 , n13443 );
buf ( n13445 , n13444 );
buf ( n13446 , n13445 );
not ( n13447 , n13446 );
buf ( n13448 , n13000 );
not ( n13449 , n13448 );
buf ( n13450 , n1548 );
buf ( n13451 , n13450 );
not ( n13452 , n13451 );
or ( n13453 , n13449 , n13452 );
buf ( n13454 , n1557 );
buf ( n13455 , n788 );
buf ( n13456 , n802 );
xor ( n13457 , n13455 , n13456 );
buf ( n13458 , n13457 );
buf ( n13459 , n13458 );
nand ( n13460 , n13454 , n13459 );
buf ( n13461 , n13460 );
buf ( n13462 , n13461 );
nand ( n13463 , n13453 , n13462 );
buf ( n13464 , n13463 );
buf ( n13465 , n13464 );
not ( n13466 , n13465 );
and ( n13467 , n13447 , n13466 );
buf ( n13468 , n13464 );
buf ( n13469 , n13445 );
and ( n13470 , n13468 , n13469 );
nor ( n13471 , n13467 , n13470 );
buf ( n13472 , n13471 );
buf ( n13473 , n12923 );
not ( n13474 , n13473 );
buf ( n13475 , n3656 );
not ( n13476 , n13475 );
or ( n13477 , n13474 , n13476 );
buf ( n13478 , n3662 );
buf ( n13479 , n790 );
buf ( n13480 , n800 );
xor ( n13481 , n13479 , n13480 );
buf ( n13482 , n13481 );
buf ( n13483 , n13482 );
nand ( n13484 , n13478 , n13483 );
buf ( n13485 , n13484 );
buf ( n13486 , n13485 );
nand ( n13487 , n13477 , n13486 );
buf ( n13488 , n13487 );
and ( n13489 , n13472 , n13488 );
not ( n13490 , n13472 );
buf ( n13491 , n13488 );
not ( n13492 , n13491 );
buf ( n13493 , n13492 );
and ( n13494 , n13490 , n13493 );
nor ( n13495 , n13489 , n13494 );
buf ( n13496 , n13018 );
not ( n13497 , n13496 );
buf ( n13498 , n2325 );
not ( n13499 , n13498 );
or ( n13500 , n13497 , n13499 );
buf ( n13501 , n2331 );
buf ( n13502 , n784 );
buf ( n13503 , n806 );
xor ( n13504 , n13502 , n13503 );
buf ( n13505 , n13504 );
buf ( n13506 , n13505 );
nand ( n13507 , n13501 , n13506 );
buf ( n13508 , n13507 );
buf ( n13509 , n13508 );
nand ( n13510 , n13500 , n13509 );
buf ( n13511 , n13510 );
buf ( n13512 , n13511 );
not ( n13513 , n2410 );
not ( n13514 , n12940 );
not ( n13515 , n13514 );
or ( n13516 , n13513 , n13515 );
buf ( n13517 , n1345 );
xor ( n13518 , n820 , n770 );
buf ( n13519 , n13518 );
nand ( n13520 , n13517 , n13519 );
buf ( n13521 , n13520 );
nand ( n13522 , n13516 , n13521 );
buf ( n13523 , n13522 );
xor ( n13524 , n13512 , n13523 );
buf ( n13525 , n13041 );
not ( n13526 , n13525 );
buf ( n13527 , n1522 );
not ( n13528 , n13527 );
or ( n13529 , n13526 , n13528 );
buf ( n13530 , n11137 );
buf ( n13531 , n786 );
buf ( n13532 , n804 );
xor ( n13533 , n13531 , n13532 );
buf ( n13534 , n13533 );
buf ( n13535 , n13534 );
nand ( n13536 , n13530 , n13535 );
buf ( n13537 , n13536 );
buf ( n13538 , n13537 );
nand ( n13539 , n13529 , n13538 );
buf ( n13540 , n13539 );
buf ( n13541 , n13540 );
xor ( n13542 , n13524 , n13541 );
buf ( n13543 , n13542 );
not ( n13544 , n13543 );
and ( n13545 , n13495 , n13544 );
not ( n13546 , n13495 );
and ( n13547 , n13546 , n13543 );
nor ( n13548 , n13545 , n13547 );
buf ( n13549 , n13548 );
buf ( n13550 , n792 );
buf ( n13551 , n800 );
and ( n13552 , n13550 , n13551 );
buf ( n13553 , n13552 );
buf ( n13554 , n13553 );
buf ( n13555 , n13083 );
xor ( n13556 , n13554 , n13555 );
buf ( n13557 , n13060 );
not ( n13558 , n13557 );
buf ( n13559 , n2066 );
not ( n13560 , n13559 );
or ( n13561 , n13558 , n13560 );
buf ( n13562 , n1694 );
buf ( n13563 , n778 );
buf ( n13564 , n812 );
xor ( n13565 , n13563 , n13564 );
buf ( n13566 , n13565 );
buf ( n13567 , n13566 );
nand ( n13568 , n13562 , n13567 );
buf ( n13569 , n13568 );
buf ( n13570 , n13569 );
nand ( n13571 , n13561 , n13570 );
buf ( n13572 , n13571 );
buf ( n13573 , n13572 );
xor ( n13574 , n13556 , n13573 );
buf ( n13575 , n13574 );
buf ( n13576 , n13575 );
and ( n13577 , n13549 , n13576 );
not ( n13578 , n13549 );
buf ( n13579 , n13575 );
not ( n13580 , n13579 );
buf ( n13581 , n13580 );
buf ( n13582 , n13581 );
and ( n13583 , n13578 , n13582 );
nor ( n13584 , n13577 , n13583 );
buf ( n13585 , n13584 );
xor ( n13586 , n13426 , n13585 );
xor ( n13587 , n13298 , n13586 );
xor ( n13588 , n13008 , n13049 );
and ( n13589 , n13588 , n13108 );
and ( n13590 , n13008 , n13049 );
or ( n13591 , n13589 , n13590 );
buf ( n13592 , n13591 );
buf ( n13593 , n13592 );
xor ( n13594 , n13067 , n13087 );
and ( n13595 , n13594 , n13105 );
and ( n13596 , n13067 , n13087 );
or ( n13597 , n13595 , n13596 );
buf ( n13598 , n13597 );
buf ( n13599 , n13598 );
buf ( n13600 , n12980 );
not ( n13601 , n13600 );
buf ( n13602 , n12989 );
not ( n13603 , n13602 );
or ( n13604 , n13601 , n13603 );
or ( n13605 , n12989 , n12980 );
nand ( n13606 , n13605 , n13006 );
buf ( n13607 , n13606 );
nand ( n13608 , n13604 , n13607 );
buf ( n13609 , n13608 );
buf ( n13610 , n13609 );
buf ( n13611 , n13047 );
not ( n13612 , n13611 );
buf ( n13613 , n13024 );
not ( n13614 , n13613 );
or ( n13615 , n13612 , n13614 );
buf ( n13616 , n13047 );
buf ( n13617 , n13024 );
or ( n13618 , n13616 , n13617 );
buf ( n13619 , n13033 );
nand ( n13620 , n13618 , n13619 );
buf ( n13621 , n13620 );
buf ( n13622 , n13621 );
nand ( n13623 , n13615 , n13622 );
buf ( n13624 , n13623 );
buf ( n13625 , n13624 );
xor ( n13626 , n13610 , n13625 );
xor ( n13627 , n12866 , n12883 );
and ( n13628 , n13627 , n12904 );
and ( n13629 , n12866 , n12883 );
or ( n13630 , n13628 , n13629 );
buf ( n13631 , n13630 );
buf ( n13632 , n13631 );
xor ( n13633 , n13626 , n13632 );
buf ( n13634 , n13633 );
buf ( n13635 , n13634 );
xor ( n13636 , n13599 , n13635 );
xor ( n13637 , n13155 , n13175 );
and ( n13638 , n13637 , n13182 );
and ( n13639 , n13155 , n13175 );
or ( n13640 , n13638 , n13639 );
buf ( n13641 , n13640 );
buf ( n13642 , n13641 );
xor ( n13643 , n13636 , n13642 );
buf ( n13644 , n13643 );
buf ( n13645 , n13644 );
xor ( n13646 , n13593 , n13645 );
xor ( n13647 , n13133 , n13139 );
and ( n13648 , n13647 , n13185 );
and ( n13649 , n13133 , n13139 );
or ( n13650 , n13648 , n13649 );
buf ( n13651 , n13650 );
buf ( n13652 , n13651 );
xor ( n13653 , n13646 , n13652 );
buf ( n13654 , n13653 );
xor ( n13655 , n13587 , n13654 );
buf ( n13656 , n13655 );
xor ( n13657 , n13293 , n13656 );
buf ( n13658 , n13657 );
buf ( n13659 , n13658 );
not ( n13660 , n13659 );
buf ( n13661 , n13660 );
buf ( n13662 , n13661 );
not ( n13663 , n13662 );
or ( n13664 , n13280 , n13663 );
buf ( n13665 , n13658 );
buf ( n13666 , n13277 );
nand ( n13667 , n13665 , n13666 );
buf ( n13668 , n13667 );
buf ( n13669 , n13668 );
nand ( n13670 , n13664 , n13669 );
buf ( n13671 , n13670 );
buf ( n13672 , n13671 );
nor ( n13673 , n13254 , n13672 );
buf ( n13674 , n13673 );
buf ( n13675 , n13674 );
nor ( n13676 , n13252 , n13675 );
buf ( n13677 , n13676 );
buf ( n13678 , n13677 );
nand ( n13679 , n12810 , n13678 );
buf ( n13680 , n13679 );
buf ( n13681 , n13680 );
not ( n13682 , n13681 );
xor ( n13683 , n12793 , n12728 );
and ( n13684 , n13683 , n12765 );
not ( n13685 , n13683 );
and ( n13686 , n13685 , n12776 );
nor ( n13687 , n13684 , n13686 );
not ( n13688 , n13687 );
xor ( n13689 , n12593 , n12579 );
not ( n13690 , n12598 );
and ( n13691 , n13689 , n13690 );
not ( n13692 , n13689 );
and ( n13693 , n13692 , n12598 );
nor ( n13694 , n13691 , n13693 );
xor ( n13695 , n3898 , n4167 );
and ( n13696 , n13695 , n4320 );
and ( n13697 , n3898 , n4167 );
or ( n13698 , n13696 , n13697 );
buf ( n13699 , n13698 );
xor ( n13700 , n13694 , n13699 );
xor ( n13701 , n12736 , n12754 );
xor ( n13702 , n13701 , n12761 );
buf ( n13703 , n13702 );
and ( n13704 , n13700 , n13703 );
and ( n13705 , n13694 , n13699 );
or ( n13706 , n13704 , n13705 );
and ( n13707 , n13688 , n13706 );
not ( n13708 , n13688 );
not ( n13709 , n13706 );
and ( n13710 , n13708 , n13709 );
nor ( n13711 , n13707 , n13710 );
xor ( n13712 , n13694 , n13699 );
xor ( n13713 , n13712 , n13703 );
buf ( n13714 , n13713 );
xor ( n13715 , n3802 , n3808 );
and ( n13716 , n13715 , n4323 );
and ( n13717 , n3802 , n3808 );
or ( n13718 , n13716 , n13717 );
buf ( n13719 , n13718 );
buf ( n13720 , n13719 );
and ( n13721 , n13714 , n13720 );
buf ( n13722 , n13721 );
nor ( n13723 , n13711 , n13722 );
buf ( n13724 , n13688 );
buf ( n13725 , n13706 );
and ( n13726 , n13724 , n13725 );
buf ( n13727 , n13726 );
buf ( n13728 , n13727 );
xor ( n13729 , n12715 , n12802 );
buf ( n13730 , n13729 );
nor ( n13731 , n13728 , n13730 );
buf ( n13732 , n13731 );
nor ( n13733 , n13723 , n13732 );
buf ( n13734 , n13733 );
not ( n13735 , n13734 );
buf ( n13736 , n4344 );
buf ( n13737 , n13719 );
not ( n13738 , n13737 );
not ( n13739 , n13713 );
buf ( n13740 , n13739 );
not ( n13741 , n13740 );
or ( n13742 , n13738 , n13741 );
buf ( n13743 , n13713 );
buf ( n13744 , n13719 );
not ( n13745 , n13744 );
buf ( n13746 , n13745 );
buf ( n13747 , n13746 );
nand ( n13748 , n13743 , n13747 );
buf ( n13749 , n13748 );
buf ( n13750 , n13749 );
nand ( n13751 , n13742 , n13750 );
buf ( n13752 , n13751 );
not ( n13753 , n13752 );
and ( n13754 , n4325 , n3794 );
not ( n13755 , n13754 );
nand ( n13756 , n13753 , n13755 );
buf ( n13757 , n13756 );
nand ( n13758 , n13736 , n13757 );
buf ( n13759 , n13758 );
buf ( n13760 , n13759 );
nor ( n13761 , n13735 , n13760 );
buf ( n13762 , n13761 );
buf ( n13763 , n13762 );
nand ( n13764 , n13682 , n13763 );
buf ( n13765 , n13764 );
buf ( n13766 , n13765 );
not ( n13767 , n13766 );
buf ( n13768 , n13767 );
buf ( n13769 , n13768 );
not ( n13770 , n13769 );
buf ( n13771 , n13770 );
buf ( n13772 , n13771 );
not ( n13773 , n3662 );
buf ( n13774 , n789 );
buf ( n13775 , n800 );
xor ( n13776 , n13774 , n13775 );
buf ( n13777 , n13776 );
not ( n13778 , n13777 );
or ( n13779 , n13773 , n13778 );
nand ( n13780 , n3656 , n13482 );
nand ( n13781 , n13779 , n13780 );
buf ( n13782 , n13781 );
buf ( n13783 , n13397 );
not ( n13784 , n13783 );
buf ( n13785 , n2098 );
not ( n13786 , n13785 );
or ( n13787 , n13784 , n13786 );
buf ( n13788 , n822 );
buf ( n13789 , n3745 );
nand ( n13790 , n13788 , n13789 );
buf ( n13791 , n13790 );
buf ( n13792 , n13791 );
nand ( n13793 , n13787 , n13792 );
buf ( n13794 , n13793 );
buf ( n13795 , n13794 );
xor ( n13796 , n13782 , n13795 );
buf ( n13797 , n13566 );
not ( n13798 , n13797 );
buf ( n13799 , n2066 );
not ( n13800 , n13799 );
or ( n13801 , n13798 , n13800 );
buf ( n13802 , n6446 );
buf ( n13803 , n777 );
buf ( n13804 , n812 );
xor ( n13805 , n13803 , n13804 );
buf ( n13806 , n13805 );
buf ( n13807 , n13806 );
nand ( n13808 , n13802 , n13807 );
buf ( n13809 , n13808 );
buf ( n13810 , n13809 );
nand ( n13811 , n13801 , n13810 );
buf ( n13812 , n13811 );
buf ( n13813 , n13812 );
xor ( n13814 , n13796 , n13813 );
buf ( n13815 , n13814 );
buf ( n13816 , n13815 );
buf ( n13817 , n13505 );
not ( n13818 , n13817 );
buf ( n13819 , n1403 );
not ( n13820 , n13819 );
or ( n13821 , n13818 , n13820 );
buf ( n13822 , n2982 );
buf ( n13823 , n783 );
buf ( n13824 , n806 );
xor ( n13825 , n13823 , n13824 );
buf ( n13826 , n13825 );
buf ( n13827 , n13826 );
nand ( n13828 , n13822 , n13827 );
buf ( n13829 , n13828 );
buf ( n13830 , n13829 );
nand ( n13831 , n13821 , n13830 );
buf ( n13832 , n13831 );
buf ( n13833 , n13832 );
not ( n13834 , n13833 );
buf ( n13835 , n13834 );
buf ( n13836 , n13835 );
not ( n13837 , n13836 );
buf ( n13838 , n13319 );
not ( n13839 , n13838 );
buf ( n13840 , n10674 );
not ( n13841 , n13840 );
or ( n13842 , n13839 , n13841 );
buf ( n13843 , n1309 );
buf ( n13844 , n781 );
buf ( n13845 , n808 );
xor ( n13846 , n13844 , n13845 );
buf ( n13847 , n13846 );
buf ( n13848 , n13847 );
nand ( n13849 , n13843 , n13848 );
buf ( n13850 , n13849 );
buf ( n13851 , n13850 );
nand ( n13852 , n13842 , n13851 );
buf ( n13853 , n13852 );
buf ( n13854 , n13358 );
not ( n13855 , n13854 );
buf ( n13856 , n2004 );
not ( n13857 , n13856 );
or ( n13858 , n13855 , n13857 );
buf ( n13859 , n2010 );
buf ( n13860 , n773 );
buf ( n13861 , n816 );
xor ( n13862 , n13860 , n13861 );
buf ( n13863 , n13862 );
buf ( n13864 , n13863 );
nand ( n13865 , n13859 , n13864 );
buf ( n13866 , n13865 );
buf ( n13867 , n13866 );
nand ( n13868 , n13858 , n13867 );
buf ( n13869 , n13868 );
xor ( n13870 , n13853 , n13869 );
buf ( n13871 , n13870 );
not ( n13872 , n13871 );
or ( n13873 , n13837 , n13872 );
buf ( n13874 , n13870 );
buf ( n13875 , n13835 );
or ( n13876 , n13874 , n13875 );
nand ( n13877 , n13873 , n13876 );
buf ( n13878 , n13877 );
buf ( n13879 , n13878 );
xor ( n13880 , n13816 , n13879 );
buf ( n13881 , n13436 );
not ( n13882 , n13881 );
buf ( n13883 , n1931 );
not ( n13884 , n13883 );
or ( n13885 , n13882 , n13884 );
buf ( n13886 , n2621 );
buf ( n13887 , n775 );
buf ( n13888 , n814 );
xor ( n13889 , n13887 , n13888 );
buf ( n13890 , n13889 );
buf ( n13891 , n13890 );
nand ( n13892 , n13886 , n13891 );
buf ( n13893 , n13892 );
buf ( n13894 , n13893 );
nand ( n13895 , n13885 , n13894 );
buf ( n13896 , n13895 );
buf ( n13897 , n13534 );
not ( n13898 , n13897 );
buf ( n13899 , n1440 );
not ( n13900 , n13899 );
or ( n13901 , n13898 , n13900 );
buf ( n13902 , n1449 );
xor ( n13903 , n804 , n785 );
buf ( n13904 , n13903 );
nand ( n13905 , n13902 , n13904 );
buf ( n13906 , n13905 );
buf ( n13907 , n13906 );
nand ( n13908 , n13901 , n13907 );
buf ( n13909 , n13908 );
buf ( n13910 , n13909 );
not ( n13911 , n13910 );
buf ( n13912 , n13911 );
xor ( n13913 , n13896 , n13912 );
buf ( n13914 , n13458 );
not ( n13915 , n13914 );
buf ( n13916 , n1551 );
not ( n13917 , n13916 );
or ( n13918 , n13915 , n13917 );
buf ( n13919 , n1560 );
xor ( n13920 , n802 , n787 );
buf ( n13921 , n13920 );
nand ( n13922 , n13919 , n13921 );
buf ( n13923 , n13922 );
buf ( n13924 , n13923 );
nand ( n13925 , n13918 , n13924 );
buf ( n13926 , n13925 );
xnor ( n13927 , n13913 , n13926 );
buf ( n13928 , n13927 );
xor ( n13929 , n13880 , n13928 );
buf ( n13930 , n13929 );
buf ( n13931 , n13930 );
xor ( n13932 , n13599 , n13635 );
and ( n13933 , n13932 , n13642 );
and ( n13934 , n13599 , n13635 );
or ( n13935 , n13933 , n13934 );
buf ( n13936 , n13935 );
buf ( n13937 , n13936 );
xor ( n13938 , n13931 , n13937 );
xor ( n13939 , n13554 , n13555 );
and ( n13940 , n13939 , n13573 );
and ( n13941 , n13554 , n13555 );
or ( n13942 , n13940 , n13941 );
buf ( n13943 , n13942 );
buf ( n13944 , n13943 );
xor ( n13945 , n13610 , n13625 );
and ( n13946 , n13945 , n13632 );
and ( n13947 , n13610 , n13625 );
or ( n13948 , n13946 , n13947 );
buf ( n13949 , n13948 );
buf ( n13950 , n13949 );
xor ( n13951 , n13944 , n13950 );
buf ( n13952 , n13518 );
not ( n13953 , n13952 );
buf ( n13954 , n2267 );
not ( n13955 , n13954 );
or ( n13956 , n13953 , n13955 );
buf ( n13957 , n1346 );
buf ( n13958 , n769 );
buf ( n13959 , n820 );
xor ( n13960 , n13958 , n13959 );
buf ( n13961 , n13960 );
buf ( n13962 , n13961 );
nand ( n13963 , n13957 , n13962 );
buf ( n13964 , n13963 );
buf ( n13965 , n13964 );
nand ( n13966 , n13956 , n13965 );
buf ( n13967 , n13966 );
buf ( n13968 , n13967 );
not ( n13969 , n13968 );
buf ( n13970 , n13969 );
buf ( n13971 , n13970 );
xor ( n13972 , n13326 , n13343 );
and ( n13973 , n13972 , n13366 );
and ( n13974 , n13326 , n13343 );
or ( n13975 , n13973 , n13974 );
buf ( n13976 , n13975 );
buf ( n13977 , n13976 );
xor ( n13978 , n13971 , n13977 );
xor ( n13979 , n13512 , n13523 );
and ( n13980 , n13979 , n13541 );
and ( n13981 , n13512 , n13523 );
or ( n13982 , n13980 , n13981 );
buf ( n13983 , n13982 );
buf ( n13984 , n13983 );
xor ( n13985 , n13978 , n13984 );
buf ( n13986 , n13985 );
buf ( n13987 , n13986 );
xor ( n13988 , n13951 , n13987 );
buf ( n13989 , n13988 );
buf ( n13990 , n13989 );
xor ( n13991 , n13938 , n13990 );
buf ( n13992 , n13991 );
buf ( n13993 , n13992 );
buf ( n13994 , n13488 );
not ( n13995 , n13994 );
buf ( n13996 , n13442 );
not ( n13997 , n13996 );
or ( n13998 , n13995 , n13997 );
buf ( n13999 , n13442 );
buf ( n14000 , n13488 );
or ( n14001 , n13999 , n14000 );
buf ( n14002 , n13464 );
nand ( n14003 , n14001 , n14002 );
buf ( n14004 , n14003 );
buf ( n14005 , n14004 );
nand ( n14006 , n13998 , n14005 );
buf ( n14007 , n14006 );
not ( n14008 , n13412 );
nand ( n14009 , n14008 , n13414 );
not ( n14010 , n14009 );
not ( n14011 , n13403 );
or ( n14012 , n14010 , n14011 );
nand ( n14013 , n14012 , n13419 );
and ( n14014 , n14007 , n14013 );
not ( n14015 , n14007 );
and ( n14016 , n13403 , n14009 );
nor ( n14017 , n14016 , n13420 );
and ( n14018 , n14015 , n14017 );
nor ( n14019 , n14014 , n14018 );
buf ( n14020 , n14019 );
buf ( n14021 , n791 );
buf ( n14022 , n800 );
nand ( n14023 , n14021 , n14022 );
buf ( n14024 , n14023 );
buf ( n14025 , n14024 );
not ( n14026 , n14025 );
buf ( n14027 , n14026 );
buf ( n14028 , n14027 );
buf ( n14029 , n13380 );
not ( n14030 , n14029 );
buf ( n14031 , n4396 );
not ( n14032 , n14031 );
or ( n14033 , n14030 , n14032 );
buf ( n14034 , n1496 );
buf ( n14035 , n771 );
buf ( n14036 , n818 );
xor ( n14037 , n14035 , n14036 );
buf ( n14038 , n14037 );
buf ( n14039 , n14038 );
nand ( n14040 , n14034 , n14039 );
buf ( n14041 , n14040 );
buf ( n14042 , n14041 );
nand ( n14043 , n14033 , n14042 );
buf ( n14044 , n14043 );
buf ( n14045 , n14044 );
xor ( n14046 , n14028 , n14045 );
buf ( n14047 , n13336 );
not ( n14048 , n14047 );
buf ( n14049 , n11050 );
not ( n14050 , n14049 );
or ( n14051 , n14048 , n14050 );
buf ( n14052 , n5272 );
buf ( n14053 , n779 );
buf ( n14054 , n810 );
xor ( n14055 , n14053 , n14054 );
buf ( n14056 , n14055 );
buf ( n14057 , n14056 );
nand ( n14058 , n14052 , n14057 );
buf ( n14059 , n14058 );
buf ( n14060 , n14059 );
nand ( n14061 , n14051 , n14060 );
buf ( n14062 , n14061 );
buf ( n14063 , n14062 );
xnor ( n14064 , n14046 , n14063 );
buf ( n14065 , n14064 );
buf ( n14066 , n14065 );
not ( n14067 , n14066 );
buf ( n14068 , n14067 );
buf ( n14069 , n14068 );
and ( n14070 , n14020 , n14069 );
not ( n14071 , n14020 );
buf ( n14072 , n14065 );
and ( n14073 , n14071 , n14072 );
nor ( n14074 , n14070 , n14073 );
buf ( n14075 , n14074 );
buf ( n14076 , n14075 );
buf ( n14077 , n13543 );
buf ( n14078 , n13575 );
or ( n14079 , n14077 , n14078 );
not ( n14080 , n13495 );
buf ( n14081 , n14080 );
nand ( n14082 , n14079 , n14081 );
buf ( n14083 , n14082 );
buf ( n14084 , n14083 );
buf ( n14085 , n13543 );
buf ( n14086 , n13575 );
nand ( n14087 , n14085 , n14086 );
buf ( n14088 , n14087 );
buf ( n14089 , n14088 );
nand ( n14090 , n14084 , n14089 );
buf ( n14091 , n14090 );
buf ( n14092 , n14091 );
xor ( n14093 , n14076 , n14092 );
xor ( n14094 , n13309 , n13369 );
and ( n14095 , n14094 , n13423 );
and ( n14096 , n13309 , n13369 );
or ( n14097 , n14095 , n14096 );
buf ( n14098 , n14097 );
buf ( n14099 , n14098 );
xor ( n14100 , n14093 , n14099 );
buf ( n14101 , n14100 );
xor ( n14102 , n13303 , n13425 );
and ( n14103 , n14102 , n13585 );
and ( n14104 , n13303 , n13425 );
or ( n14105 , n14103 , n14104 );
xor ( n14106 , n14101 , n14105 );
xor ( n14107 , n13593 , n13645 );
and ( n14108 , n14107 , n13652 );
and ( n14109 , n13593 , n13645 );
or ( n14110 , n14108 , n14109 );
buf ( n14111 , n14110 );
xor ( n14112 , n14106 , n14111 );
buf ( n14113 , n14112 );
xor ( n14114 , n13993 , n14113 );
xor ( n14115 , n13298 , n13586 );
and ( n14116 , n14115 , n13654 );
and ( n14117 , n13298 , n13586 );
or ( n14118 , n14116 , n14117 );
buf ( n14119 , n14118 );
xor ( n14120 , n14114 , n14119 );
buf ( n14121 , n14120 );
xor ( n14122 , n13286 , n13292 );
and ( n14123 , n14122 , n13656 );
and ( n14124 , n13286 , n13292 );
or ( n14125 , n14123 , n14124 );
buf ( n14126 , n14125 );
and ( n14127 , n14121 , n14126 );
not ( n14128 , n14127 );
xor ( n14129 , n13944 , n13950 );
and ( n14130 , n14129 , n13987 );
and ( n14131 , n13944 , n13950 );
or ( n14132 , n14130 , n14131 );
buf ( n14133 , n14132 );
buf ( n14134 , n14133 );
not ( n14135 , n14134 );
buf ( n14136 , n13903 );
not ( n14137 , n14136 );
buf ( n14138 , n1737 );
not ( n14139 , n14138 );
or ( n14140 , n14137 , n14139 );
buf ( n14141 , n1449 );
xor ( n14142 , n804 , n784 );
buf ( n14143 , n14142 );
nand ( n14144 , n14141 , n14143 );
buf ( n14145 , n14144 );
buf ( n14146 , n14145 );
nand ( n14147 , n14140 , n14146 );
buf ( n14148 , n14147 );
buf ( n14149 , n13920 );
not ( n14150 , n14149 );
buf ( n14151 , n10922 );
not ( n14152 , n14151 );
or ( n14153 , n14150 , n14152 );
buf ( n14154 , n1557 );
xor ( n14155 , n802 , n786 );
buf ( n14156 , n14155 );
nand ( n14157 , n14154 , n14156 );
buf ( n14158 , n14157 );
buf ( n14159 , n14158 );
nand ( n14160 , n14153 , n14159 );
buf ( n14161 , n14160 );
xor ( n14162 , n14148 , n14161 );
buf ( n14163 , n14038 );
not ( n14164 , n14163 );
buf ( n14165 , n1480 );
not ( n14166 , n14165 );
or ( n14167 , n14164 , n14166 );
buf ( n14168 , n1496 );
buf ( n14169 , n770 );
buf ( n14170 , n818 );
xor ( n14171 , n14169 , n14170 );
buf ( n14172 , n14171 );
buf ( n14173 , n14172 );
nand ( n14174 , n14168 , n14173 );
buf ( n14175 , n14174 );
buf ( n14176 , n14175 );
nand ( n14177 , n14167 , n14176 );
buf ( n14178 , n14177 );
not ( n14179 , n14178 );
xor ( n14180 , n14162 , n14179 );
buf ( n14181 , n13961 );
not ( n14182 , n14181 );
buf ( n14183 , n2410 );
not ( n14184 , n14183 );
or ( n14185 , n14182 , n14184 );
buf ( n14186 , n768 );
buf ( n14187 , n820 );
xor ( n14188 , n14186 , n14187 );
buf ( n14189 , n14188 );
buf ( n14190 , n14189 );
buf ( n14191 , n1346 );
nand ( n14192 , n14190 , n14191 );
buf ( n14193 , n14192 );
buf ( n14194 , n14193 );
nand ( n14195 , n14185 , n14194 );
buf ( n14196 , n14195 );
buf ( n14197 , n2110 );
not ( n14198 , n14197 );
buf ( n14199 , n2577 );
not ( n14200 , n14199 );
buf ( n14201 , n14200 );
buf ( n14202 , n14201 );
not ( n14203 , n14202 );
or ( n14204 , n14198 , n14203 );
buf ( n14205 , n822 );
nand ( n14206 , n14204 , n14205 );
buf ( n14207 , n14206 );
xor ( n14208 , n14196 , n14207 );
buf ( n14209 , n13863 );
not ( n14210 , n14209 );
buf ( n14211 , n2526 );
not ( n14212 , n14211 );
or ( n14213 , n14210 , n14212 );
buf ( n14214 , n2010 );
buf ( n14215 , n772 );
buf ( n14216 , n816 );
xor ( n14217 , n14215 , n14216 );
buf ( n14218 , n14217 );
buf ( n14219 , n14218 );
nand ( n14220 , n14214 , n14219 );
buf ( n14221 , n14220 );
buf ( n14222 , n14221 );
nand ( n14223 , n14213 , n14222 );
buf ( n14224 , n14223 );
xor ( n14225 , n14208 , n14224 );
xor ( n14226 , n14180 , n14225 );
buf ( n14227 , n13847 );
not ( n14228 , n14227 );
buf ( n14229 , n10674 );
not ( n14230 , n14229 );
or ( n14231 , n14228 , n14230 );
buf ( n14232 , n1309 );
buf ( n14233 , n780 );
buf ( n14234 , n808 );
xor ( n14235 , n14233 , n14234 );
buf ( n14236 , n14235 );
buf ( n14237 , n14236 );
nand ( n14238 , n14232 , n14237 );
buf ( n14239 , n14238 );
buf ( n14240 , n14239 );
nand ( n14241 , n14231 , n14240 );
buf ( n14242 , n14241 );
buf ( n14243 , n14242 );
not ( n14244 , n14243 );
buf ( n14245 , n14244 );
buf ( n14246 , n14245 );
buf ( n14247 , n13890 );
not ( n14248 , n14247 );
buf ( n14249 , n2612 );
not ( n14250 , n14249 );
or ( n14251 , n14248 , n14250 );
buf ( n14252 , n1940 );
buf ( n14253 , n774 );
buf ( n14254 , n814 );
xor ( n14255 , n14253 , n14254 );
buf ( n14256 , n14255 );
buf ( n14257 , n14256 );
nand ( n14258 , n14252 , n14257 );
buf ( n14259 , n14258 );
buf ( n14260 , n14259 );
nand ( n14261 , n14251 , n14260 );
buf ( n14262 , n14261 );
buf ( n14263 , n14262 );
and ( n14264 , n14246 , n14263 );
not ( n14265 , n14246 );
buf ( n14266 , n14262 );
not ( n14267 , n14266 );
buf ( n14268 , n14267 );
buf ( n14269 , n14268 );
and ( n14270 , n14265 , n14269 );
or ( n14271 , n14264 , n14270 );
buf ( n14272 , n14271 );
buf ( n14273 , n14272 );
buf ( n14274 , n13826 );
not ( n14275 , n14274 );
buf ( n14276 , n1403 );
buf ( n14277 , n14276 );
buf ( n14278 , n14277 );
buf ( n14279 , n14278 );
not ( n14280 , n14279 );
or ( n14281 , n14275 , n14280 );
buf ( n14282 , n2982 );
buf ( n14283 , n14282 );
buf ( n14284 , n14283 );
buf ( n14285 , n14284 );
buf ( n14286 , n782 );
buf ( n14287 , n806 );
xor ( n14288 , n14286 , n14287 );
buf ( n14289 , n14288 );
buf ( n14290 , n14289 );
nand ( n14291 , n14285 , n14290 );
buf ( n14292 , n14291 );
buf ( n14293 , n14292 );
nand ( n14294 , n14281 , n14293 );
buf ( n14295 , n14294 );
buf ( n14296 , n14295 );
xnor ( n14297 , n14273 , n14296 );
buf ( n14298 , n14297 );
xnor ( n14299 , n14226 , n14298 );
buf ( n14300 , n14299 );
not ( n14301 , n14300 );
and ( n14302 , n14135 , n14301 );
buf ( n14303 , n14133 );
buf ( n14304 , n14299 );
and ( n14305 , n14303 , n14304 );
nor ( n14306 , n14302 , n14305 );
buf ( n14307 , n14306 );
buf ( n14308 , n14307 );
buf ( n14309 , n790 );
buf ( n14310 , n800 );
and ( n14311 , n14309 , n14310 );
buf ( n14312 , n14311 );
buf ( n14313 , n14312 );
buf ( n14314 , n13777 );
not ( n14315 , n14314 );
buf ( n14316 , n3656 );
not ( n14317 , n14316 );
or ( n14318 , n14315 , n14317 );
xor ( n14319 , n800 , n788 );
nand ( n14320 , n3662 , n14319 );
buf ( n14321 , n14320 );
nand ( n14322 , n14318 , n14321 );
buf ( n14323 , n14322 );
buf ( n14324 , n14323 );
xor ( n14325 , n14313 , n14324 );
buf ( n14326 , n13806 );
not ( n14327 , n14326 );
buf ( n14328 , n2066 );
not ( n14329 , n14328 );
or ( n14330 , n14327 , n14329 );
buf ( n14331 , n1693 );
buf ( n14332 , n14331 );
buf ( n14333 , n776 );
buf ( n14334 , n812 );
xor ( n14335 , n14333 , n14334 );
buf ( n14336 , n14335 );
buf ( n14337 , n14336 );
nand ( n14338 , n14332 , n14337 );
buf ( n14339 , n14338 );
buf ( n14340 , n14339 );
nand ( n14341 , n14330 , n14340 );
buf ( n14342 , n14341 );
buf ( n14343 , n14342 );
xor ( n14344 , n14325 , n14343 );
buf ( n14345 , n14344 );
buf ( n14346 , n13909 );
not ( n14347 , n14346 );
buf ( n14348 , n13896 );
not ( n14349 , n14348 );
or ( n14350 , n14347 , n14349 );
buf ( n14351 , n13912 );
not ( n14352 , n14351 );
buf ( n14353 , n13896 );
not ( n14354 , n14353 );
buf ( n14355 , n14354 );
buf ( n14356 , n14355 );
not ( n14357 , n14356 );
or ( n14358 , n14352 , n14357 );
buf ( n14359 , n13926 );
nand ( n14360 , n14358 , n14359 );
buf ( n14361 , n14360 );
buf ( n14362 , n14361 );
nand ( n14363 , n14350 , n14362 );
buf ( n14364 , n14363 );
buf ( n14365 , n14364 );
not ( n14366 , n14365 );
buf ( n14367 , n13967 );
not ( n14368 , n14367 );
buf ( n14369 , n14056 );
not ( n14370 , n14369 );
buf ( n14371 , n2641 );
not ( n14372 , n14371 );
or ( n14373 , n14370 , n14372 );
buf ( n14374 , n3398 );
buf ( n14375 , n778 );
buf ( n14376 , n810 );
xor ( n14377 , n14375 , n14376 );
buf ( n14378 , n14377 );
buf ( n14379 , n14378 );
nand ( n14380 , n14374 , n14379 );
buf ( n14381 , n14380 );
buf ( n14382 , n14381 );
nand ( n14383 , n14373 , n14382 );
buf ( n14384 , n14383 );
buf ( n14385 , n14384 );
not ( n14386 , n14385 );
buf ( n14387 , n14386 );
buf ( n14388 , n14387 );
not ( n14389 , n14388 );
and ( n14390 , n14368 , n14389 );
buf ( n14391 , n13967 );
buf ( n14392 , n14387 );
and ( n14393 , n14391 , n14392 );
nor ( n14394 , n14390 , n14393 );
buf ( n14395 , n14394 );
buf ( n14396 , n14395 );
not ( n14397 , n14396 );
and ( n14398 , n14366 , n14397 );
buf ( n14399 , n14364 );
buf ( n14400 , n14395 );
and ( n14401 , n14399 , n14400 );
nor ( n14402 , n14398 , n14401 );
buf ( n14403 , n14402 );
xor ( n14404 , n14345 , n14403 );
xor ( n14405 , n13971 , n13977 );
and ( n14406 , n14405 , n13984 );
and ( n14407 , n13971 , n13977 );
or ( n14408 , n14406 , n14407 );
buf ( n14409 , n14408 );
xor ( n14410 , n14404 , n14409 );
not ( n14411 , n14410 );
buf ( n14412 , n14411 );
not ( n14413 , n14412 );
buf ( n14414 , n14413 );
and ( n14415 , n14308 , n14414 );
not ( n14416 , n14308 );
buf ( n14417 , n14412 );
and ( n14418 , n14416 , n14417 );
nor ( n14419 , n14415 , n14418 );
buf ( n14420 , n14419 );
buf ( n14421 , n14420 );
not ( n14422 , n14068 );
not ( n14423 , n14013 );
or ( n14424 , n14422 , n14423 );
not ( n14425 , n14065 );
not ( n14426 , n14017 );
or ( n14427 , n14425 , n14426 );
nand ( n14428 , n14427 , n14007 );
nand ( n14429 , n14424 , n14428 );
buf ( n14430 , n14429 );
not ( n14431 , n14044 );
nand ( n14432 , n14431 , n14024 );
not ( n14433 , n14432 );
not ( n14434 , n14062 );
or ( n14435 , n14433 , n14434 );
buf ( n14436 , n14044 );
buf ( n14437 , n14027 );
nand ( n14438 , n14436 , n14437 );
buf ( n14439 , n14438 );
nand ( n14440 , n14435 , n14439 );
buf ( n14441 , n14440 );
buf ( n14442 , n13853 );
buf ( n14443 , n13832 );
or ( n14444 , n14442 , n14443 );
buf ( n14445 , n13869 );
nand ( n14446 , n14444 , n14445 );
buf ( n14447 , n14446 );
buf ( n14448 , n14447 );
buf ( n14449 , n13853 );
buf ( n14450 , n13832 );
nand ( n14451 , n14449 , n14450 );
buf ( n14452 , n14451 );
buf ( n14453 , n14452 );
nand ( n14454 , n14448 , n14453 );
buf ( n14455 , n14454 );
buf ( n14456 , n14455 );
xor ( n14457 , n14441 , n14456 );
xor ( n14458 , n13782 , n13795 );
and ( n14459 , n14458 , n13813 );
and ( n14460 , n13782 , n13795 );
or ( n14461 , n14459 , n14460 );
buf ( n14462 , n14461 );
buf ( n14463 , n14462 );
xor ( n14464 , n14457 , n14463 );
buf ( n14465 , n14464 );
buf ( n14466 , n14465 );
xor ( n14467 , n14430 , n14466 );
xor ( n14468 , n13816 , n13879 );
and ( n14469 , n14468 , n13928 );
and ( n14470 , n13816 , n13879 );
or ( n14471 , n14469 , n14470 );
buf ( n14472 , n14471 );
buf ( n14473 , n14472 );
xor ( n14474 , n14467 , n14473 );
buf ( n14475 , n14474 );
buf ( n14476 , n14475 );
xor ( n14477 , n14076 , n14092 );
and ( n14478 , n14477 , n14099 );
and ( n14479 , n14076 , n14092 );
or ( n14480 , n14478 , n14479 );
buf ( n14481 , n14480 );
buf ( n14482 , n14481 );
xor ( n14483 , n14476 , n14482 );
xor ( n14484 , n13931 , n13937 );
and ( n14485 , n14484 , n13990 );
and ( n14486 , n13931 , n13937 );
or ( n14487 , n14485 , n14486 );
buf ( n14488 , n14487 );
buf ( n14489 , n14488 );
xor ( n14490 , n14483 , n14489 );
buf ( n14491 , n14490 );
buf ( n14492 , n14491 );
xor ( n14493 , n14421 , n14492 );
xor ( n14494 , n14101 , n14105 );
and ( n14495 , n14494 , n14111 );
and ( n14496 , n14101 , n14105 );
or ( n14497 , n14495 , n14496 );
buf ( n14498 , n14497 );
xor ( n14499 , n14493 , n14498 );
buf ( n14500 , n14499 );
buf ( n14501 , n14500 );
not ( n14502 , n14501 );
buf ( n14503 , n14502 );
buf ( n14504 , n14503 );
not ( n14505 , n14504 );
xor ( n14506 , n13993 , n14113 );
and ( n14507 , n14506 , n14119 );
and ( n14508 , n13993 , n14113 );
or ( n14509 , n14507 , n14508 );
buf ( n14510 , n14509 );
buf ( n14511 , n14510 );
not ( n14512 , n14511 );
or ( n14513 , n14505 , n14512 );
buf ( n14514 , n14510 );
not ( n14515 , n14514 );
buf ( n14516 , n14515 );
buf ( n14517 , n14516 );
buf ( n14518 , n14500 );
nand ( n14519 , n14517 , n14518 );
buf ( n14520 , n14519 );
buf ( n14521 , n14520 );
nand ( n14522 , n14513 , n14521 );
buf ( n14523 , n14522 );
not ( n14524 , n14523 );
and ( n14525 , n14128 , n14524 );
buf ( n14526 , n14126 );
not ( n14527 , n14526 );
not ( n14528 , n14121 );
buf ( n14529 , n14528 );
not ( n14530 , n14529 );
or ( n14531 , n14527 , n14530 );
buf ( n14532 , n14126 );
not ( n14533 , n14532 );
buf ( n14534 , n14533 );
buf ( n14535 , n14534 );
buf ( n14536 , n14121 );
nand ( n14537 , n14535 , n14536 );
buf ( n14538 , n14537 );
buf ( n14539 , n14538 );
nand ( n14540 , n14531 , n14539 );
buf ( n14541 , n14540 );
buf ( n14542 , n14541 );
buf ( n14543 , n13658 );
buf ( n14544 , n13278 );
and ( n14545 , n14543 , n14544 );
buf ( n14546 , n14545 );
buf ( n14547 , n14546 );
nor ( n14548 , n14542 , n14547 );
buf ( n14549 , n14548 );
nor ( n14550 , n14525 , n14549 );
buf ( n14551 , n14550 );
buf ( n14552 , n14155 );
not ( n14553 , n14552 );
buf ( n14554 , n1551 );
not ( n14555 , n14554 );
or ( n14556 , n14553 , n14555 );
buf ( n14557 , n1560 );
buf ( n14558 , n785 );
buf ( n14559 , n802 );
xor ( n14560 , n14558 , n14559 );
buf ( n14561 , n14560 );
buf ( n14562 , n14561 );
nand ( n14563 , n14557 , n14562 );
buf ( n14564 , n14563 );
buf ( n14565 , n14564 );
nand ( n14566 , n14556 , n14565 );
buf ( n14567 , n14566 );
buf ( n14568 , n14567 );
not ( n14569 , n14319 );
not ( n14570 , n10509 );
or ( n14571 , n14569 , n14570 );
buf ( n14572 , n3662 );
buf ( n14573 , n787 );
buf ( n14574 , n800 );
xor ( n14575 , n14573 , n14574 );
buf ( n14576 , n14575 );
buf ( n14577 , n14576 );
nand ( n14578 , n14572 , n14577 );
buf ( n14579 , n14578 );
nand ( n14580 , n14571 , n14579 );
buf ( n14581 , n14580 );
xor ( n14582 , n14568 , n14581 );
buf ( n14583 , n14336 );
not ( n14584 , n14583 );
buf ( n14585 , n2066 );
not ( n14586 , n14585 );
or ( n14587 , n14584 , n14586 );
not ( n14588 , n1694 );
not ( n14589 , n14588 );
buf ( n14590 , n14589 );
buf ( n14591 , n775 );
buf ( n14592 , n812 );
xor ( n14593 , n14591 , n14592 );
buf ( n14594 , n14593 );
buf ( n14595 , n14594 );
nand ( n14596 , n14590 , n14595 );
buf ( n14597 , n14596 );
buf ( n14598 , n14597 );
nand ( n14599 , n14587 , n14598 );
buf ( n14600 , n14599 );
buf ( n14601 , n14600 );
xor ( n14602 , n14582 , n14601 );
buf ( n14603 , n14602 );
buf ( n14604 , n14603 );
buf ( n14605 , n14236 );
not ( n14606 , n14605 );
buf ( n14607 , n10674 );
not ( n14608 , n14607 );
or ( n14609 , n14606 , n14608 );
buf ( n14610 , n1309 );
buf ( n14611 , n779 );
buf ( n14612 , n808 );
xor ( n14613 , n14611 , n14612 );
buf ( n14614 , n14613 );
buf ( n14615 , n14614 );
nand ( n14616 , n14610 , n14615 );
buf ( n14617 , n14616 );
buf ( n14618 , n14617 );
nand ( n14619 , n14609 , n14618 );
buf ( n14620 , n14619 );
buf ( n14621 , n14620 );
buf ( n14622 , n14378 );
not ( n14623 , n14622 );
buf ( n14624 , n12889 );
not ( n14625 , n14624 );
or ( n14626 , n14623 , n14625 );
buf ( n14627 , n5272 );
buf ( n14628 , n777 );
buf ( n14629 , n810 );
xor ( n14630 , n14628 , n14629 );
buf ( n14631 , n14630 );
buf ( n14632 , n14631 );
nand ( n14633 , n14627 , n14632 );
buf ( n14634 , n14633 );
buf ( n14635 , n14634 );
nand ( n14636 , n14626 , n14635 );
buf ( n14637 , n14636 );
buf ( n14638 , n14637 );
xor ( n14639 , n14621 , n14638 );
buf ( n14640 , n14172 );
not ( n14641 , n14640 );
buf ( n14642 , n1480 );
not ( n14643 , n14642 );
or ( n14644 , n14641 , n14643 );
buf ( n14645 , n1496 );
buf ( n14646 , n769 );
buf ( n14647 , n818 );
xor ( n14648 , n14646 , n14647 );
buf ( n14649 , n14648 );
buf ( n14650 , n14649 );
nand ( n14651 , n14645 , n14650 );
buf ( n14652 , n14651 );
buf ( n14653 , n14652 );
nand ( n14654 , n14644 , n14653 );
buf ( n14655 , n14654 );
buf ( n14656 , n14655 );
not ( n14657 , n14656 );
buf ( n14658 , n14657 );
buf ( n14659 , n14658 );
xor ( n14660 , n14639 , n14659 );
buf ( n14661 , n14660 );
buf ( n14662 , n14661 );
xor ( n14663 , n14604 , n14662 );
xor ( n14664 , n14441 , n14456 );
and ( n14665 , n14664 , n14463 );
and ( n14666 , n14441 , n14456 );
or ( n14667 , n14665 , n14666 );
buf ( n14668 , n14667 );
buf ( n14669 , n14668 );
xor ( n14670 , n14663 , n14669 );
buf ( n14671 , n14670 );
buf ( n14672 , n14671 );
buf ( n14673 , n14672 );
buf ( n14674 , n14673 );
buf ( n14675 , n14674 );
not ( n14676 , n14675 );
buf ( n14677 , n14345 );
not ( n14678 , n14677 );
buf ( n14679 , n14403 );
not ( n14680 , n14679 );
buf ( n14681 , n14680 );
buf ( n14682 , n14681 );
not ( n14683 , n14682 );
or ( n14684 , n14678 , n14683 );
buf ( n14685 , n14345 );
not ( n14686 , n14685 );
buf ( n14687 , n14686 );
buf ( n14688 , n14687 );
not ( n14689 , n14688 );
buf ( n14690 , n14403 );
not ( n14691 , n14690 );
or ( n14692 , n14689 , n14691 );
buf ( n14693 , n14409 );
nand ( n14694 , n14692 , n14693 );
buf ( n14695 , n14694 );
buf ( n14696 , n14695 );
nand ( n14697 , n14684 , n14696 );
buf ( n14698 , n14697 );
buf ( n14699 , n14698 );
not ( n14700 , n14699 );
not ( n14701 , n14242 );
not ( n14702 , n14262 );
or ( n14703 , n14701 , n14702 );
buf ( n14704 , n14245 );
not ( n14705 , n14704 );
buf ( n14706 , n14268 );
not ( n14707 , n14706 );
or ( n14708 , n14705 , n14707 );
buf ( n14709 , n14295 );
nand ( n14710 , n14708 , n14709 );
buf ( n14711 , n14710 );
nand ( n14712 , n14703 , n14711 );
not ( n14713 , n14712 );
buf ( n14714 , n789 );
buf ( n14715 , n800 );
and ( n14716 , n14714 , n14715 );
buf ( n14717 , n14716 );
buf ( n14718 , n14717 );
buf ( n14719 , n14218 );
not ( n14720 , n14719 );
buf ( n14721 , n2526 );
not ( n14722 , n14721 );
or ( n14723 , n14720 , n14722 );
buf ( n14724 , n2010 );
buf ( n14725 , n771 );
buf ( n14726 , n816 );
xor ( n14727 , n14725 , n14726 );
buf ( n14728 , n14727 );
buf ( n14729 , n14728 );
nand ( n14730 , n14724 , n14729 );
buf ( n14731 , n14730 );
buf ( n14732 , n14731 );
nand ( n14733 , n14723 , n14732 );
buf ( n14734 , n14733 );
buf ( n14735 , n14734 );
xor ( n14736 , n14718 , n14735 );
buf ( n14737 , n14189 );
not ( n14738 , n14737 );
buf ( n14739 , n2410 );
not ( n14740 , n14739 );
or ( n14741 , n14738 , n14740 );
buf ( n14742 , n820 );
buf ( n14743 , n2672 );
nand ( n14744 , n14742 , n14743 );
buf ( n14745 , n14744 );
buf ( n14746 , n14745 );
nand ( n14747 , n14741 , n14746 );
buf ( n14748 , n14747 );
buf ( n14749 , n14748 );
xor ( n14750 , n14736 , n14749 );
buf ( n14751 , n14750 );
buf ( n14752 , n14751 );
not ( n14753 , n14752 );
buf ( n14754 , n14753 );
not ( n14755 , n14754 );
or ( n14756 , n14713 , n14755 );
not ( n14757 , n14712 );
nand ( n14758 , n14757 , n14751 );
nand ( n14759 , n14756 , n14758 );
not ( n14760 , n14142 );
not ( n14761 , n1522 );
or ( n14762 , n14760 , n14761 );
buf ( n14763 , n1528 );
buf ( n14764 , n783 );
buf ( n14765 , n804 );
xor ( n14766 , n14764 , n14765 );
buf ( n14767 , n14766 );
buf ( n14768 , n14767 );
nand ( n14769 , n14763 , n14768 );
buf ( n14770 , n14769 );
nand ( n14771 , n14762 , n14770 );
buf ( n14772 , n14289 );
not ( n14773 , n14772 );
buf ( n14774 , n1403 );
not ( n14775 , n14774 );
or ( n14776 , n14773 , n14775 );
buf ( n14777 , n2982 );
buf ( n14778 , n781 );
buf ( n14779 , n806 );
xor ( n14780 , n14778 , n14779 );
buf ( n14781 , n14780 );
buf ( n14782 , n14781 );
nand ( n14783 , n14777 , n14782 );
buf ( n14784 , n14783 );
buf ( n14785 , n14784 );
nand ( n14786 , n14776 , n14785 );
buf ( n14787 , n14786 );
xor ( n14788 , n14771 , n14787 );
buf ( n14789 , n14256 );
not ( n14790 , n14789 );
buf ( n14791 , n3703 );
not ( n14792 , n14791 );
or ( n14793 , n14790 , n14792 );
buf ( n14794 , n1940 );
buf ( n14795 , n773 );
buf ( n14796 , n814 );
xor ( n14797 , n14795 , n14796 );
buf ( n14798 , n14797 );
buf ( n14799 , n14798 );
nand ( n14800 , n14794 , n14799 );
buf ( n14801 , n14800 );
buf ( n14802 , n14801 );
nand ( n14803 , n14793 , n14802 );
buf ( n14804 , n14803 );
not ( n14805 , n14804 );
xor ( n14806 , n14788 , n14805 );
and ( n14807 , n14759 , n14806 );
not ( n14808 , n14759 );
not ( n14809 , n14806 );
and ( n14810 , n14808 , n14809 );
nor ( n14811 , n14807 , n14810 );
buf ( n14812 , n14811 );
not ( n14813 , n14812 );
and ( n14814 , n14700 , n14813 );
buf ( n14815 , n14698 );
buf ( n14816 , n14811 );
and ( n14817 , n14815 , n14816 );
nor ( n14818 , n14814 , n14817 );
buf ( n14819 , n14818 );
buf ( n14820 , n14819 );
not ( n14821 , n14820 );
or ( n14822 , n14676 , n14821 );
buf ( n14823 , n14819 );
buf ( n14824 , n14674 );
or ( n14825 , n14823 , n14824 );
nand ( n14826 , n14822 , n14825 );
buf ( n14827 , n14826 );
buf ( n14828 , n14827 );
xor ( n14829 , n14476 , n14482 );
and ( n14830 , n14829 , n14489 );
and ( n14831 , n14476 , n14482 );
or ( n14832 , n14830 , n14831 );
buf ( n14833 , n14832 );
buf ( n14834 , n14833 );
xor ( n14835 , n14828 , n14834 );
xor ( n14836 , n14430 , n14466 );
and ( n14837 , n14836 , n14473 );
and ( n14838 , n14430 , n14466 );
or ( n14839 , n14837 , n14838 );
buf ( n14840 , n14839 );
buf ( n14841 , n14840 );
buf ( n14842 , n13970 );
buf ( n14843 , n14387 );
nand ( n14844 , n14842 , n14843 );
buf ( n14845 , n14844 );
buf ( n14846 , n14845 );
not ( n14847 , n14846 );
buf ( n14848 , n14364 );
not ( n14849 , n14848 );
or ( n14850 , n14847 , n14849 );
buf ( n14851 , n14384 );
buf ( n14852 , n13967 );
nand ( n14853 , n14851 , n14852 );
buf ( n14854 , n14853 );
buf ( n14855 , n14854 );
nand ( n14856 , n14850 , n14855 );
buf ( n14857 , n14856 );
buf ( n14858 , n14857 );
not ( n14859 , n14178 );
buf ( n14860 , n14148 );
buf ( n14861 , n14161 );
or ( n14862 , n14860 , n14861 );
buf ( n14863 , n14862 );
not ( n14864 , n14863 );
or ( n14865 , n14859 , n14864 );
buf ( n14866 , n14148 );
buf ( n14867 , n14161 );
nand ( n14868 , n14866 , n14867 );
buf ( n14869 , n14868 );
nand ( n14870 , n14865 , n14869 );
buf ( n14871 , n14870 );
buf ( n14872 , n14207 );
not ( n14873 , n14872 );
buf ( n14874 , n14196 );
not ( n14875 , n14874 );
or ( n14876 , n14873 , n14875 );
buf ( n14877 , n14196 );
buf ( n14878 , n14207 );
or ( n14879 , n14877 , n14878 );
buf ( n14880 , n14224 );
nand ( n14881 , n14879 , n14880 );
buf ( n14882 , n14881 );
buf ( n14883 , n14882 );
nand ( n14884 , n14876 , n14883 );
buf ( n14885 , n14884 );
buf ( n14886 , n14885 );
xor ( n14887 , n14871 , n14886 );
xor ( n14888 , n14313 , n14324 );
and ( n14889 , n14888 , n14343 );
and ( n14890 , n14313 , n14324 );
or ( n14891 , n14889 , n14890 );
buf ( n14892 , n14891 );
buf ( n14893 , n14892 );
xor ( n14894 , n14887 , n14893 );
buf ( n14895 , n14894 );
buf ( n14896 , n14895 );
xor ( n14897 , n14858 , n14896 );
not ( n14898 , n14225 );
buf ( n14899 , n14180 );
not ( n14900 , n14899 );
buf ( n14901 , n14900 );
not ( n14902 , n14901 );
or ( n14903 , n14898 , n14902 );
buf ( n14904 , n14225 );
buf ( n14905 , n14901 );
nor ( n14906 , n14904 , n14905 );
buf ( n14907 , n14906 );
or ( n14908 , n14298 , n14907 );
nand ( n14909 , n14903 , n14908 );
buf ( n14910 , n14909 );
xor ( n14911 , n14897 , n14910 );
buf ( n14912 , n14911 );
buf ( n14913 , n14912 );
xor ( n14914 , n14841 , n14913 );
buf ( n14915 , n14299 );
not ( n14916 , n14915 );
buf ( n14917 , n14410 );
not ( n14918 , n14917 );
or ( n14919 , n14916 , n14918 );
buf ( n14920 , n14133 );
nand ( n14921 , n14919 , n14920 );
buf ( n14922 , n14921 );
buf ( n14923 , n14922 );
buf ( n14924 , n14411 );
buf ( n14925 , n14299 );
not ( n14926 , n14925 );
buf ( n14927 , n14926 );
buf ( n14928 , n14927 );
nand ( n14929 , n14924 , n14928 );
buf ( n14930 , n14929 );
buf ( n14931 , n14930 );
nand ( n14932 , n14923 , n14931 );
buf ( n14933 , n14932 );
buf ( n14934 , n14933 );
xor ( n14935 , n14914 , n14934 );
buf ( n14936 , n14935 );
buf ( n14937 , n14936 );
and ( n14938 , n14835 , n14937 );
and ( n14939 , n14828 , n14834 );
or ( n14940 , n14938 , n14939 );
buf ( n14941 , n14940 );
buf ( n14942 , n14941 );
not ( n14943 , n14942 );
buf ( n14944 , n14943 );
buf ( n14945 , n14944 );
not ( n14946 , n14945 );
buf ( n14947 , n14798 );
not ( n14948 , n14947 );
buf ( n14949 , n1931 );
not ( n14950 , n14949 );
or ( n14951 , n14948 , n14950 );
buf ( n14952 , n1940 );
buf ( n14953 , n772 );
buf ( n14954 , n814 );
xor ( n14955 , n14953 , n14954 );
buf ( n14956 , n14955 );
buf ( n14957 , n14956 );
nand ( n14958 , n14952 , n14957 );
buf ( n14959 , n14958 );
buf ( n14960 , n14959 );
nand ( n14961 , n14951 , n14960 );
buf ( n14962 , n14961 );
buf ( n14963 , n14962 );
buf ( n14964 , n14649 );
not ( n14965 , n14964 );
buf ( n14966 , n1480 );
not ( n14967 , n14966 );
or ( n14968 , n14965 , n14967 );
buf ( n14969 , n1496 );
buf ( n14970 , n768 );
buf ( n14971 , n818 );
xor ( n14972 , n14970 , n14971 );
buf ( n14973 , n14972 );
buf ( n14974 , n14973 );
nand ( n14975 , n14969 , n14974 );
buf ( n14976 , n14975 );
buf ( n14977 , n14976 );
nand ( n14978 , n14968 , n14977 );
buf ( n14979 , n14978 );
buf ( n14980 , n14979 );
xor ( n14981 , n14963 , n14980 );
buf ( n14982 , n2671 );
not ( n14983 , n14982 );
buf ( n14984 , n2410 );
not ( n14985 , n14984 );
buf ( n14986 , n14985 );
buf ( n14987 , n14986 );
not ( n14988 , n14987 );
or ( n14989 , n14983 , n14988 );
buf ( n14990 , n820 );
nand ( n14991 , n14989 , n14990 );
buf ( n14992 , n14991 );
buf ( n14993 , n14992 );
xor ( n14994 , n14981 , n14993 );
buf ( n14995 , n14994 );
buf ( n14996 , n14995 );
xor ( n14997 , n14621 , n14638 );
and ( n14998 , n14997 , n14659 );
and ( n14999 , n14621 , n14638 );
or ( n15000 , n14998 , n14999 );
buf ( n15001 , n15000 );
buf ( n15002 , n15001 );
xor ( n15003 , n14996 , n15002 );
not ( n15004 , n14767 );
not ( n15005 , n1737 );
or ( n15006 , n15004 , n15005 );
buf ( n15007 , n1528 );
buf ( n15008 , n782 );
buf ( n15009 , n804 );
xor ( n15010 , n15008 , n15009 );
buf ( n15011 , n15010 );
buf ( n15012 , n15011 );
nand ( n15013 , n15007 , n15012 );
buf ( n15014 , n15013 );
nand ( n15015 , n15006 , n15014 );
not ( n15016 , n14781 );
not ( n15017 , n1403 );
or ( n15018 , n15016 , n15017 );
buf ( n15019 , n1409 );
buf ( n15020 , n780 );
buf ( n15021 , n806 );
xor ( n15022 , n15020 , n15021 );
buf ( n15023 , n15022 );
buf ( n15024 , n15023 );
nand ( n15025 , n15019 , n15024 );
buf ( n15026 , n15025 );
nand ( n15027 , n15018 , n15026 );
xor ( n15028 , n15015 , n15027 );
not ( n15029 , n14594 );
not ( n15030 , n2916 );
or ( n15031 , n15029 , n15030 );
buf ( n15032 , n6446 );
buf ( n15033 , n774 );
buf ( n15034 , n812 );
xor ( n15035 , n15033 , n15034 );
buf ( n15036 , n15035 );
buf ( n15037 , n15036 );
nand ( n15038 , n15032 , n15037 );
buf ( n15039 , n15038 );
nand ( n15040 , n15031 , n15039 );
xor ( n15041 , n15028 , n15040 );
buf ( n15042 , n15041 );
xor ( n15043 , n15003 , n15042 );
buf ( n15044 , n15043 );
buf ( n15045 , n14631 );
not ( n15046 , n15045 );
buf ( n15047 , n11050 );
not ( n15048 , n15047 );
or ( n15049 , n15046 , n15048 );
buf ( n15050 , n5272 );
buf ( n15051 , n776 );
buf ( n15052 , n810 );
xor ( n15053 , n15051 , n15052 );
buf ( n15054 , n15053 );
buf ( n15055 , n15054 );
nand ( n15056 , n15050 , n15055 );
buf ( n15057 , n15056 );
buf ( n15058 , n15057 );
nand ( n15059 , n15049 , n15058 );
buf ( n15060 , n15059 );
buf ( n15061 , n15060 );
buf ( n15062 , n788 );
buf ( n15063 , n800 );
and ( n15064 , n15062 , n15063 );
buf ( n15065 , n15064 );
buf ( n15066 , n15065 );
and ( n15067 , n15061 , n15066 );
not ( n15068 , n15061 );
buf ( n15069 , n788 );
buf ( n15070 , n800 );
nand ( n15071 , n15069 , n15070 );
buf ( n15072 , n15071 );
buf ( n15073 , n15072 );
and ( n15074 , n15068 , n15073 );
nor ( n15075 , n15067 , n15074 );
buf ( n15076 , n15075 );
buf ( n15077 , n15076 );
buf ( n15078 , n14614 );
not ( n15079 , n15078 );
buf ( n15080 , n10674 );
not ( n15081 , n15080 );
or ( n15082 , n15079 , n15081 );
buf ( n15083 , n1309 );
buf ( n15084 , n778 );
buf ( n15085 , n808 );
xor ( n15086 , n15084 , n15085 );
buf ( n15087 , n15086 );
buf ( n15088 , n15087 );
nand ( n15089 , n15083 , n15088 );
buf ( n15090 , n15089 );
buf ( n15091 , n15090 );
nand ( n15092 , n15082 , n15091 );
buf ( n15093 , n15092 );
buf ( n15094 , n15093 );
not ( n15095 , n15094 );
buf ( n15096 , n15095 );
buf ( n15097 , n15096 );
and ( n15098 , n15077 , n15097 );
not ( n15099 , n15077 );
buf ( n15100 , n15093 );
and ( n15101 , n15099 , n15100 );
nor ( n15102 , n15098 , n15101 );
buf ( n15103 , n15102 );
buf ( n15104 , n15103 );
not ( n15105 , n15104 );
xor ( n15106 , n14568 , n14581 );
and ( n15107 , n15106 , n14601 );
and ( n15108 , n14568 , n14581 );
or ( n15109 , n15107 , n15108 );
buf ( n15110 , n15109 );
buf ( n15111 , n15110 );
not ( n15112 , n15111 );
or ( n15113 , n15105 , n15112 );
buf ( n15114 , n15110 );
buf ( n15115 , n15103 );
or ( n15116 , n15114 , n15115 );
nand ( n15117 , n15113 , n15116 );
buf ( n15118 , n15117 );
buf ( n15119 , n15118 );
buf ( n15120 , n14728 );
not ( n15121 , n15120 );
buf ( n15122 , n2526 );
not ( n15123 , n15122 );
or ( n15124 , n15121 , n15123 );
buf ( n15125 , n2535 );
xor ( n15126 , n816 , n770 );
buf ( n15127 , n15126 );
nand ( n15128 , n15125 , n15127 );
buf ( n15129 , n15128 );
buf ( n15130 , n15129 );
nand ( n15131 , n15124 , n15130 );
buf ( n15132 , n15131 );
buf ( n15133 , n14561 );
not ( n15134 , n15133 );
buf ( n15135 , n1551 );
not ( n15136 , n15135 );
or ( n15137 , n15134 , n15136 );
buf ( n15138 , n1560 );
buf ( n15139 , n784 );
buf ( n15140 , n802 );
xor ( n15141 , n15139 , n15140 );
buf ( n15142 , n15141 );
buf ( n15143 , n15142 );
nand ( n15144 , n15138 , n15143 );
buf ( n15145 , n15144 );
buf ( n15146 , n15145 );
nand ( n15147 , n15137 , n15146 );
buf ( n15148 , n15147 );
xor ( n15149 , n15132 , n15148 );
buf ( n15150 , n14576 );
not ( n15151 , n15150 );
buf ( n15152 , n3656 );
not ( n15153 , n15152 );
or ( n15154 , n15151 , n15153 );
buf ( n15155 , n3662 );
buf ( n15156 , n786 );
buf ( n15157 , n800 );
xor ( n15158 , n15156 , n15157 );
buf ( n15159 , n15158 );
buf ( n15160 , n15159 );
nand ( n15161 , n15155 , n15160 );
buf ( n15162 , n15161 );
buf ( n15163 , n15162 );
nand ( n15164 , n15154 , n15163 );
buf ( n15165 , n15164 );
xor ( n15166 , n15149 , n15165 );
buf ( n15167 , n15166 );
not ( n15168 , n15167 );
buf ( n15169 , n15168 );
buf ( n15170 , n15169 );
and ( n15171 , n15119 , n15170 );
not ( n15172 , n15119 );
buf ( n15173 , n15166 );
and ( n15174 , n15172 , n15173 );
nor ( n15175 , n15171 , n15174 );
buf ( n15176 , n15175 );
xor ( n15177 , n15044 , n15176 );
xor ( n15178 , n14604 , n14662 );
and ( n15179 , n15178 , n14669 );
and ( n15180 , n14604 , n14662 );
or ( n15181 , n15179 , n15180 );
buf ( n15182 , n15181 );
buf ( n15183 , n15182 );
not ( n15184 , n15183 );
buf ( n15185 , n15184 );
and ( n15186 , n15177 , n15185 );
not ( n15187 , n15177 );
and ( n15188 , n15187 , n15182 );
nor ( n15189 , n15186 , n15188 );
buf ( n15190 , n15189 );
xor ( n15191 , n14841 , n14913 );
and ( n15192 , n15191 , n14934 );
and ( n15193 , n14841 , n14913 );
or ( n15194 , n15192 , n15193 );
buf ( n15195 , n15194 );
buf ( n15196 , n15195 );
xor ( n15197 , n15190 , n15196 );
xor ( n15198 , n14858 , n14896 );
and ( n15199 , n15198 , n14910 );
and ( n15200 , n14858 , n14896 );
or ( n15201 , n15199 , n15200 );
buf ( n15202 , n15201 );
buf ( n15203 , n15202 );
xor ( n15204 , n14871 , n14886 );
and ( n15205 , n15204 , n14893 );
and ( n15206 , n14871 , n14886 );
or ( n15207 , n15205 , n15206 );
buf ( n15208 , n15207 );
buf ( n15209 , n15208 );
buf ( n15210 , n14655 );
xor ( n15211 , n14718 , n14735 );
and ( n15212 , n15211 , n14749 );
and ( n15213 , n14718 , n14735 );
or ( n15214 , n15212 , n15213 );
buf ( n15215 , n15214 );
buf ( n15216 , n15215 );
xor ( n15217 , n15210 , n15216 );
or ( n15218 , n14771 , n14804 );
nand ( n15219 , n15218 , n14787 );
buf ( n15220 , n15219 );
buf ( n15221 , n14804 );
buf ( n15222 , n14771 );
nand ( n15223 , n15221 , n15222 );
buf ( n15224 , n15223 );
buf ( n15225 , n15224 );
nand ( n15226 , n15220 , n15225 );
buf ( n15227 , n15226 );
buf ( n15228 , n15227 );
xor ( n15229 , n15217 , n15228 );
buf ( n15230 , n15229 );
buf ( n15231 , n15230 );
xor ( n15232 , n15209 , n15231 );
not ( n15233 , n14757 );
not ( n15234 , n14754 );
or ( n15235 , n15233 , n15234 );
nand ( n15236 , n15235 , n14809 );
buf ( n15237 , n15236 );
buf ( n15238 , n14757 );
not ( n15239 , n15238 );
buf ( n15240 , n14751 );
nand ( n15241 , n15239 , n15240 );
buf ( n15242 , n15241 );
buf ( n15243 , n15242 );
nand ( n15244 , n15237 , n15243 );
buf ( n15245 , n15244 );
buf ( n15246 , n15245 );
xor ( n15247 , n15232 , n15246 );
buf ( n15248 , n15247 );
buf ( n15249 , n15248 );
xor ( n15250 , n15203 , n15249 );
not ( n15251 , n14811 );
nor ( n15252 , n15251 , n14671 );
buf ( n15253 , n15252 );
buf ( n15254 , n14698 );
not ( n15255 , n15254 );
buf ( n15256 , n15255 );
buf ( n15257 , n15256 );
or ( n15258 , n15253 , n15257 );
buf ( n15259 , n14671 );
buf ( n15260 , n15251 );
nand ( n15261 , n15259 , n15260 );
buf ( n15262 , n15261 );
buf ( n15263 , n15262 );
nand ( n15264 , n15258 , n15263 );
buf ( n15265 , n15264 );
buf ( n15266 , n15265 );
xor ( n15267 , n15250 , n15266 );
buf ( n15268 , n15267 );
buf ( n15269 , n15268 );
xor ( n15270 , n15197 , n15269 );
buf ( n15271 , n15270 );
buf ( n15272 , n15271 );
not ( n15273 , n15272 );
or ( n15274 , n14946 , n15273 );
buf ( n15275 , n14944 );
buf ( n15276 , n15271 );
or ( n15277 , n15275 , n15276 );
nand ( n15278 , n15274 , n15277 );
buf ( n15279 , n15278 );
buf ( n15280 , n15279 );
not ( n15281 , n15280 );
xor ( n15282 , n14828 , n14834 );
xor ( n15283 , n15282 , n14937 );
buf ( n15284 , n15283 );
buf ( n15285 , n15284 );
xor ( n15286 , n14421 , n14492 );
and ( n15287 , n15286 , n14498 );
and ( n15288 , n14421 , n14492 );
or ( n15289 , n15287 , n15288 );
buf ( n15290 , n15289 );
buf ( n15291 , n15290 );
nand ( n15292 , n15285 , n15291 );
buf ( n15293 , n15292 );
buf ( n15294 , n15293 );
nand ( n15295 , n15281 , n15294 );
buf ( n15296 , n15295 );
buf ( n15297 , n15296 );
not ( n15298 , n15297 );
buf ( n15299 , n15298 );
buf ( n15300 , n15299 );
buf ( n15301 , n14510 );
buf ( n15302 , n14500 );
and ( n15303 , n15301 , n15302 );
buf ( n15304 , n15303 );
buf ( n15305 , n15304 );
buf ( n15306 , n15290 );
buf ( n15307 , n15284 );
and ( n15308 , n15306 , n15307 );
not ( n15309 , n15306 );
buf ( n15310 , n15284 );
not ( n15311 , n15310 );
buf ( n15312 , n15311 );
buf ( n15313 , n15312 );
and ( n15314 , n15309 , n15313 );
nor ( n15315 , n15308 , n15314 );
buf ( n15316 , n15315 );
buf ( n15317 , n15316 );
nor ( n15318 , n15305 , n15317 );
buf ( n15319 , n15318 );
buf ( n15320 , n15319 );
nor ( n15321 , n15300 , n15320 );
buf ( n15322 , n15321 );
buf ( n15323 , n15322 );
nand ( n15324 , n14551 , n15323 );
buf ( n15325 , n15324 );
buf ( n15326 , n15325 );
not ( n15327 , n15326 );
xor ( n15328 , n15190 , n15196 );
and ( n15329 , n15328 , n15269 );
and ( n15330 , n15190 , n15196 );
or ( n15331 , n15329 , n15330 );
buf ( n15332 , n15331 );
buf ( n15333 , n15166 );
buf ( n15334 , n15103 );
not ( n15335 , n15334 );
buf ( n15336 , n15335 );
buf ( n15337 , n15336 );
or ( n15338 , n15333 , n15337 );
buf ( n15339 , n15110 );
nand ( n15340 , n15338 , n15339 );
buf ( n15341 , n15340 );
buf ( n15342 , n15341 );
buf ( n15343 , n15166 );
buf ( n15344 , n15336 );
nand ( n15345 , n15343 , n15344 );
buf ( n15346 , n15345 );
buf ( n15347 , n15346 );
nand ( n15348 , n15342 , n15347 );
buf ( n15349 , n15348 );
buf ( n15350 , n15349 );
xor ( n15351 , n14996 , n15002 );
and ( n15352 , n15351 , n15042 );
and ( n15353 , n14996 , n15002 );
or ( n15354 , n15352 , n15353 );
buf ( n15355 , n15354 );
buf ( n15356 , n15355 );
xor ( n15357 , n15350 , n15356 );
buf ( n15358 , n787 );
buf ( n15359 , n800 );
and ( n15360 , n15358 , n15359 );
buf ( n15361 , n15360 );
buf ( n15362 , n15361 );
buf ( n15363 , n15054 );
not ( n15364 , n15363 );
buf ( n15365 , n11050 );
not ( n15366 , n15365 );
or ( n15367 , n15364 , n15366 );
buf ( n15368 , n3398 );
buf ( n15369 , n775 );
buf ( n15370 , n810 );
xor ( n15371 , n15369 , n15370 );
buf ( n15372 , n15371 );
buf ( n15373 , n15372 );
nand ( n15374 , n15368 , n15373 );
buf ( n15375 , n15374 );
buf ( n15376 , n15375 );
nand ( n15377 , n15367 , n15376 );
buf ( n15378 , n15377 );
buf ( n15379 , n15378 );
xor ( n15380 , n15362 , n15379 );
buf ( n15381 , n15159 );
not ( n15382 , n15381 );
buf ( n15383 , n3656 );
not ( n15384 , n15383 );
or ( n15385 , n15382 , n15384 );
buf ( n15386 , n3662 );
buf ( n15387 , n785 );
buf ( n15388 , n800 );
xor ( n15389 , n15387 , n15388 );
buf ( n15390 , n15389 );
buf ( n15391 , n15390 );
nand ( n15392 , n15386 , n15391 );
buf ( n15393 , n15392 );
buf ( n15394 , n15393 );
nand ( n15395 , n15385 , n15394 );
buf ( n15396 , n15395 );
buf ( n15397 , n15396 );
xor ( n15398 , n15380 , n15397 );
buf ( n15399 , n15398 );
buf ( n15400 , n15142 );
not ( n15401 , n15400 );
buf ( n15402 , n1548 );
not ( n15403 , n15402 );
or ( n15404 , n15401 , n15403 );
buf ( n15405 , n1557 );
buf ( n15406 , n783 );
buf ( n15407 , n802 );
xor ( n15408 , n15406 , n15407 );
buf ( n15409 , n15408 );
buf ( n15410 , n15409 );
nand ( n15411 , n15405 , n15410 );
buf ( n15412 , n15411 );
buf ( n15413 , n15412 );
nand ( n15414 , n15404 , n15413 );
buf ( n15415 , n15414 );
buf ( n15416 , n15415 );
buf ( n15417 , n15011 );
not ( n15418 , n15417 );
buf ( n15419 , n1440 );
not ( n15420 , n15419 );
or ( n15421 , n15418 , n15420 );
buf ( n15422 , n11137 );
buf ( n15423 , n781 );
buf ( n15424 , n804 );
xor ( n15425 , n15423 , n15424 );
buf ( n15426 , n15425 );
buf ( n15427 , n15426 );
nand ( n15428 , n15422 , n15427 );
buf ( n15429 , n15428 );
buf ( n15430 , n15429 );
nand ( n15431 , n15421 , n15430 );
buf ( n15432 , n15431 );
buf ( n15433 , n15432 );
xor ( n15434 , n15416 , n15433 );
buf ( n15435 , n15036 );
not ( n15436 , n15435 );
buf ( n15437 , n2066 );
not ( n15438 , n15437 );
or ( n15439 , n15436 , n15438 );
buf ( n15440 , n14331 );
buf ( n15441 , n773 );
buf ( n15442 , n812 );
xor ( n15443 , n15441 , n15442 );
buf ( n15444 , n15443 );
buf ( n15445 , n15444 );
nand ( n15446 , n15440 , n15445 );
buf ( n15447 , n15446 );
buf ( n15448 , n15447 );
nand ( n15449 , n15439 , n15448 );
buf ( n15450 , n15449 );
buf ( n15451 , n15450 );
xor ( n15452 , n15434 , n15451 );
buf ( n15453 , n15452 );
xor ( n15454 , n15399 , n15453 );
buf ( n15455 , n14956 );
not ( n15456 , n15455 );
buf ( n15457 , n3703 );
not ( n15458 , n15457 );
or ( n15459 , n15456 , n15458 );
buf ( n15460 , n2621 );
buf ( n15461 , n771 );
buf ( n15462 , n814 );
xor ( n15463 , n15461 , n15462 );
buf ( n15464 , n15463 );
buf ( n15465 , n15464 );
nand ( n15466 , n15460 , n15465 );
buf ( n15467 , n15466 );
buf ( n15468 , n15467 );
nand ( n15469 , n15459 , n15468 );
buf ( n15470 , n15469 );
buf ( n15471 , n15470 );
buf ( n15472 , n15087 );
not ( n15473 , n15472 );
buf ( n15474 , n10674 );
not ( n15475 , n15474 );
or ( n15476 , n15473 , n15475 );
buf ( n15477 , n2713 );
buf ( n15478 , n777 );
buf ( n15479 , n808 );
xor ( n15480 , n15478 , n15479 );
buf ( n15481 , n15480 );
buf ( n15482 , n15481 );
nand ( n15483 , n15477 , n15482 );
buf ( n15484 , n15483 );
buf ( n15485 , n15484 );
nand ( n15486 , n15476 , n15485 );
buf ( n15487 , n15486 );
buf ( n15488 , n15487 );
xor ( n15489 , n15471 , n15488 );
buf ( n15490 , n14973 );
not ( n15491 , n15490 );
buf ( n15492 , n2725 );
not ( n15493 , n15492 );
or ( n15494 , n15491 , n15493 );
buf ( n15495 , n818 );
buf ( n15496 , n1496 );
nand ( n15497 , n15495 , n15496 );
buf ( n15498 , n15497 );
buf ( n15499 , n15498 );
nand ( n15500 , n15494 , n15499 );
buf ( n15501 , n15500 );
buf ( n15502 , n15501 );
xor ( n15503 , n15489 , n15502 );
buf ( n15504 , n15503 );
xor ( n15505 , n15454 , n15504 );
buf ( n15506 , n15505 );
xor ( n15507 , n15357 , n15506 );
buf ( n15508 , n15507 );
buf ( n15509 , n15508 );
xor ( n15510 , n15203 , n15249 );
and ( n15511 , n15510 , n15266 );
and ( n15512 , n15203 , n15249 );
or ( n15513 , n15511 , n15512 );
buf ( n15514 , n15513 );
buf ( n15515 , n15514 );
xor ( n15516 , n15509 , n15515 );
buf ( n15517 , n15023 );
not ( n15518 , n15517 );
buf ( n15519 , n1403 );
not ( n15520 , n15519 );
or ( n15521 , n15518 , n15520 );
buf ( n15522 , n2982 );
xor ( n15523 , n806 , n779 );
buf ( n15524 , n15523 );
nand ( n15525 , n15522 , n15524 );
buf ( n15526 , n15525 );
buf ( n15527 , n15526 );
nand ( n15528 , n15521 , n15527 );
buf ( n15529 , n15528 );
not ( n15530 , n15126 );
not ( n15531 , n2526 );
or ( n15532 , n15530 , n15531 );
buf ( n15533 , n2010 );
buf ( n15534 , n769 );
buf ( n15535 , n816 );
xor ( n15536 , n15534 , n15535 );
buf ( n15537 , n15536 );
buf ( n15538 , n15537 );
nand ( n15539 , n15533 , n15538 );
buf ( n15540 , n15539 );
nand ( n15541 , n15532 , n15540 );
xor ( n15542 , n15529 , n15541 );
buf ( n15543 , n15148 );
not ( n15544 , n15543 );
buf ( n15545 , n15165 );
not ( n15546 , n15545 );
or ( n15547 , n15544 , n15546 );
buf ( n15548 , n15165 );
buf ( n15549 , n15148 );
or ( n15550 , n15548 , n15549 );
buf ( n15551 , n15132 );
nand ( n15552 , n15550 , n15551 );
buf ( n15553 , n15552 );
buf ( n15554 , n15553 );
nand ( n15555 , n15547 , n15554 );
buf ( n15556 , n15555 );
xnor ( n15557 , n15542 , n15556 );
buf ( n15558 , n15557 );
xor ( n15559 , n15210 , n15216 );
and ( n15560 , n15559 , n15228 );
and ( n15561 , n15210 , n15216 );
or ( n15562 , n15560 , n15561 );
buf ( n15563 , n15562 );
buf ( n15564 , n15563 );
xor ( n15565 , n15558 , n15564 );
or ( n15566 , n15015 , n15027 );
nand ( n15567 , n15566 , n15040 );
buf ( n15568 , n15567 );
buf ( n15569 , n15027 );
buf ( n15570 , n15015 );
nand ( n15571 , n15569 , n15570 );
buf ( n15572 , n15571 );
buf ( n15573 , n15572 );
nand ( n15574 , n15568 , n15573 );
buf ( n15575 , n15574 );
buf ( n15576 , n15575 );
buf ( n15577 , n15093 );
buf ( n15578 , n15065 );
or ( n15579 , n15577 , n15578 );
buf ( n15580 , n15060 );
nand ( n15581 , n15579 , n15580 );
buf ( n15582 , n15581 );
buf ( n15583 , n15582 );
buf ( n15584 , n15093 );
buf ( n15585 , n15065 );
nand ( n15586 , n15584 , n15585 );
buf ( n15587 , n15586 );
buf ( n15588 , n15587 );
nand ( n15589 , n15583 , n15588 );
buf ( n15590 , n15589 );
buf ( n15591 , n15590 );
xor ( n15592 , n15576 , n15591 );
xor ( n15593 , n14963 , n14980 );
and ( n15594 , n15593 , n14993 );
and ( n15595 , n14963 , n14980 );
or ( n15596 , n15594 , n15595 );
buf ( n15597 , n15596 );
buf ( n15598 , n15597 );
xor ( n15599 , n15592 , n15598 );
buf ( n15600 , n15599 );
buf ( n15601 , n15600 );
xor ( n15602 , n15565 , n15601 );
buf ( n15603 , n15602 );
buf ( n15604 , n15603 );
xor ( n15605 , n15209 , n15231 );
and ( n15606 , n15605 , n15246 );
and ( n15607 , n15209 , n15231 );
or ( n15608 , n15606 , n15607 );
buf ( n15609 , n15608 );
buf ( n15610 , n15609 );
xor ( n15611 , n15604 , n15610 );
buf ( n15612 , n15044 );
not ( n15613 , n15612 );
buf ( n15614 , n15182 );
not ( n15615 , n15614 );
or ( n15616 , n15613 , n15615 );
buf ( n15617 , n15182 );
buf ( n15618 , n15044 );
or ( n15619 , n15617 , n15618 );
buf ( n15620 , n15176 );
not ( n15621 , n15620 );
buf ( n15622 , n15621 );
buf ( n15623 , n15622 );
nand ( n15624 , n15619 , n15623 );
buf ( n15625 , n15624 );
buf ( n15626 , n15625 );
nand ( n15627 , n15616 , n15626 );
buf ( n15628 , n15627 );
buf ( n15629 , n15628 );
xor ( n15630 , n15611 , n15629 );
buf ( n15631 , n15630 );
buf ( n15632 , n15631 );
xor ( n15633 , n15516 , n15632 );
buf ( n15634 , n15633 );
xor ( n15635 , n15332 , n15634 );
buf ( n15636 , n15635 );
not ( n15637 , n15636 );
buf ( n15638 , n15637 );
not ( n15639 , n15638 );
buf ( n15640 , n15271 );
buf ( n15641 , n14941 );
nand ( n15642 , n15640 , n15641 );
buf ( n15643 , n15642 );
not ( n15644 , n15643 );
or ( n15645 , n15639 , n15644 );
xor ( n15646 , n15509 , n15515 );
and ( n15647 , n15646 , n15632 );
and ( n15648 , n15509 , n15515 );
or ( n15649 , n15647 , n15648 );
buf ( n15650 , n15649 );
buf ( n15651 , n15650 );
not ( n15652 , n15651 );
xor ( n15653 , n15350 , n15356 );
and ( n15654 , n15653 , n15506 );
and ( n15655 , n15350 , n15356 );
or ( n15656 , n15654 , n15655 );
buf ( n15657 , n15656 );
buf ( n15658 , n15657 );
xor ( n15659 , n15604 , n15610 );
and ( n15660 , n15659 , n15629 );
and ( n15661 , n15604 , n15610 );
or ( n15662 , n15660 , n15661 );
buf ( n15663 , n15662 );
buf ( n15664 , n15663 );
xor ( n15665 , n15658 , n15664 );
xor ( n15666 , n15558 , n15564 );
and ( n15667 , n15666 , n15601 );
and ( n15668 , n15558 , n15564 );
or ( n15669 , n15667 , n15668 );
buf ( n15670 , n15669 );
buf ( n15671 , n15670 );
not ( n15672 , n15523 );
not ( n15673 , n14278 );
or ( n15674 , n15672 , n15673 );
buf ( n15675 , n14284 );
buf ( n15676 , n778 );
buf ( n15677 , n806 );
xor ( n15678 , n15676 , n15677 );
buf ( n15679 , n15678 );
buf ( n15680 , n15679 );
nand ( n15681 , n15675 , n15680 );
buf ( n15682 , n15681 );
nand ( n15683 , n15674 , n15682 );
xor ( n15684 , n15541 , n15683 );
not ( n15685 , n15481 );
not ( n15686 , n2709 );
or ( n15687 , n15685 , n15686 );
buf ( n15688 , n2713 );
buf ( n15689 , n776 );
buf ( n15690 , n808 );
xor ( n15691 , n15689 , n15690 );
buf ( n15692 , n15691 );
buf ( n15693 , n15692 );
nand ( n15694 , n15688 , n15693 );
buf ( n15695 , n15694 );
nand ( n15696 , n15687 , n15695 );
xor ( n15697 , n15684 , n15696 );
buf ( n15698 , n15697 );
buf ( n15699 , n15529 );
not ( n15700 , n15699 );
buf ( n15701 , n15541 );
nand ( n15702 , n15700 , n15701 );
buf ( n15703 , n15702 );
buf ( n15704 , n15703 );
not ( n15705 , n15704 );
buf ( n15706 , n15556 );
not ( n15707 , n15706 );
or ( n15708 , n15705 , n15707 );
buf ( n15709 , n15541 );
not ( n15710 , n15709 );
buf ( n15711 , n15529 );
nand ( n15712 , n15710 , n15711 );
buf ( n15713 , n15712 );
buf ( n15714 , n15713 );
nand ( n15715 , n15708 , n15714 );
buf ( n15716 , n15715 );
buf ( n15717 , n15716 );
xor ( n15718 , n15698 , n15717 );
xor ( n15719 , n15576 , n15591 );
and ( n15720 , n15719 , n15598 );
and ( n15721 , n15576 , n15591 );
or ( n15722 , n15720 , n15721 );
buf ( n15723 , n15722 );
buf ( n15724 , n15723 );
xor ( n15725 , n15718 , n15724 );
buf ( n15726 , n15725 );
buf ( n15727 , n15726 );
xor ( n15728 , n15671 , n15727 );
not ( n15729 , n15504 );
not ( n15730 , n15453 );
or ( n15731 , n15729 , n15730 );
buf ( n15732 , n15504 );
buf ( n15733 , n15453 );
or ( n15734 , n15732 , n15733 );
buf ( n15735 , n15399 );
nand ( n15736 , n15734 , n15735 );
buf ( n15737 , n15736 );
nand ( n15738 , n15731 , n15737 );
buf ( n15739 , n15738 );
xor ( n15740 , n15362 , n15379 );
and ( n15741 , n15740 , n15397 );
and ( n15742 , n15362 , n15379 );
or ( n15743 , n15741 , n15742 );
buf ( n15744 , n15743 );
buf ( n15745 , n15744 );
xor ( n15746 , n15416 , n15433 );
and ( n15747 , n15746 , n15451 );
and ( n15748 , n15416 , n15433 );
or ( n15749 , n15747 , n15748 );
buf ( n15750 , n15749 );
buf ( n15751 , n15750 );
xor ( n15752 , n15745 , n15751 );
xor ( n15753 , n15471 , n15488 );
and ( n15754 , n15753 , n15502 );
and ( n15755 , n15471 , n15488 );
or ( n15756 , n15754 , n15755 );
buf ( n15757 , n15756 );
buf ( n15758 , n15757 );
xor ( n15759 , n15752 , n15758 );
buf ( n15760 , n15759 );
buf ( n15761 , n15760 );
xor ( n15762 , n15739 , n15761 );
buf ( n15763 , n786 );
buf ( n15764 , n800 );
and ( n15765 , n15763 , n15764 );
buf ( n15766 , n15765 );
buf ( n15767 , n15766 );
buf ( n15768 , n15390 );
not ( n15769 , n15768 );
buf ( n15770 , n3656 );
not ( n15771 , n15770 );
or ( n15772 , n15769 , n15771 );
buf ( n15773 , n3662 );
buf ( n15774 , n784 );
buf ( n15775 , n800 );
xor ( n15776 , n15774 , n15775 );
buf ( n15777 , n15776 );
buf ( n15778 , n15777 );
nand ( n15779 , n15773 , n15778 );
buf ( n15780 , n15779 );
buf ( n15781 , n15780 );
nand ( n15782 , n15772 , n15781 );
buf ( n15783 , n15782 );
buf ( n15784 , n15783 );
xor ( n15785 , n15767 , n15784 );
buf ( n15786 , n15464 );
not ( n15787 , n15786 );
buf ( n15788 , n2612 );
buf ( n15789 , n15788 );
buf ( n15790 , n15789 );
buf ( n15791 , n15790 );
not ( n15792 , n15791 );
or ( n15793 , n15787 , n15792 );
buf ( n15794 , n1940 );
buf ( n15795 , n770 );
buf ( n15796 , n814 );
xor ( n15797 , n15795 , n15796 );
buf ( n15798 , n15797 );
buf ( n15799 , n15798 );
nand ( n15800 , n15794 , n15799 );
buf ( n15801 , n15800 );
buf ( n15802 , n15801 );
nand ( n15803 , n15793 , n15802 );
buf ( n15804 , n15803 );
buf ( n15805 , n15804 );
xor ( n15806 , n15785 , n15805 );
buf ( n15807 , n15806 );
buf ( n15808 , n15807 );
not ( n15809 , n15444 );
not ( n15810 , n2916 );
or ( n15811 , n15809 , n15810 );
buf ( n15812 , n3379 );
buf ( n15813 , n772 );
buf ( n15814 , n812 );
xor ( n15815 , n15813 , n15814 );
buf ( n15816 , n15815 );
buf ( n15817 , n15816 );
nand ( n15818 , n15812 , n15817 );
buf ( n15819 , n15818 );
nand ( n15820 , n15811 , n15819 );
buf ( n15821 , n1496 );
not ( n15822 , n15821 );
buf ( n15823 , n15822 );
buf ( n15824 , n15823 );
not ( n15825 , n15824 );
buf ( n15826 , n1483 );
not ( n15827 , n15826 );
or ( n15828 , n15825 , n15827 );
buf ( n15829 , n818 );
nand ( n15830 , n15828 , n15829 );
buf ( n15831 , n15830 );
xor ( n15832 , n15820 , n15831 );
buf ( n15833 , n15537 );
not ( n15834 , n15833 );
buf ( n15835 , n3719 );
not ( n15836 , n15835 );
or ( n15837 , n15834 , n15836 );
buf ( n15838 , n2010 );
buf ( n15839 , n768 );
buf ( n15840 , n816 );
xor ( n15841 , n15839 , n15840 );
buf ( n15842 , n15841 );
buf ( n15843 , n15842 );
nand ( n15844 , n15838 , n15843 );
buf ( n15845 , n15844 );
buf ( n15846 , n15845 );
nand ( n15847 , n15837 , n15846 );
buf ( n15848 , n15847 );
xor ( n15849 , n15832 , n15848 );
buf ( n15850 , n15849 );
xor ( n15851 , n15808 , n15850 );
buf ( n15852 , n15409 );
not ( n15853 , n15852 );
buf ( n15854 , n1551 );
not ( n15855 , n15854 );
or ( n15856 , n15853 , n15855 );
buf ( n15857 , n1560 );
buf ( n15858 , n782 );
buf ( n15859 , n802 );
xor ( n15860 , n15858 , n15859 );
buf ( n15861 , n15860 );
buf ( n15862 , n15861 );
nand ( n15863 , n15857 , n15862 );
buf ( n15864 , n15863 );
buf ( n15865 , n15864 );
nand ( n15866 , n15856 , n15865 );
buf ( n15867 , n15866 );
buf ( n15868 , n15867 );
buf ( n15869 , n15426 );
not ( n15870 , n15869 );
buf ( n15871 , n1440 );
buf ( n15872 , n15871 );
buf ( n15873 , n15872 );
buf ( n15874 , n15873 );
not ( n15875 , n15874 );
or ( n15876 , n15870 , n15875 );
buf ( n15877 , n11137 );
buf ( n15878 , n780 );
buf ( n15879 , n804 );
xor ( n15880 , n15878 , n15879 );
buf ( n15881 , n15880 );
buf ( n15882 , n15881 );
nand ( n15883 , n15877 , n15882 );
buf ( n15884 , n15883 );
buf ( n15885 , n15884 );
nand ( n15886 , n15876 , n15885 );
buf ( n15887 , n15886 );
buf ( n15888 , n15887 );
xor ( n15889 , n15868 , n15888 );
buf ( n15890 , n15372 );
not ( n15891 , n15890 );
buf ( n15892 , n12889 );
not ( n15893 , n15892 );
or ( n15894 , n15891 , n15893 );
buf ( n15895 , n5272 );
buf ( n15896 , n774 );
buf ( n15897 , n810 );
xor ( n15898 , n15896 , n15897 );
buf ( n15899 , n15898 );
buf ( n15900 , n15899 );
nand ( n15901 , n15895 , n15900 );
buf ( n15902 , n15901 );
buf ( n15903 , n15902 );
nand ( n15904 , n15894 , n15903 );
buf ( n15905 , n15904 );
buf ( n15906 , n15905 );
xor ( n15907 , n15889 , n15906 );
buf ( n15908 , n15907 );
buf ( n15909 , n15908 );
xor ( n15910 , n15851 , n15909 );
buf ( n15911 , n15910 );
buf ( n15912 , n15911 );
xor ( n15913 , n15762 , n15912 );
buf ( n15914 , n15913 );
buf ( n15915 , n15914 );
xor ( n15916 , n15728 , n15915 );
buf ( n15917 , n15916 );
buf ( n15918 , n15917 );
xor ( n15919 , n15665 , n15918 );
buf ( n15920 , n15919 );
buf ( n15921 , n15920 );
not ( n15922 , n15921 );
buf ( n15923 , n15922 );
buf ( n15924 , n15923 );
not ( n15925 , n15924 );
or ( n15926 , n15652 , n15925 );
buf ( n15927 , n15920 );
buf ( n15928 , n15650 );
not ( n15929 , n15928 );
buf ( n15930 , n15929 );
buf ( n15931 , n15930 );
nand ( n15932 , n15927 , n15931 );
buf ( n15933 , n15932 );
buf ( n15934 , n15933 );
nand ( n15935 , n15926 , n15934 );
buf ( n15936 , n15935 );
not ( n15937 , n15936 );
buf ( n15938 , n15332 );
buf ( n15939 , n15634 );
and ( n15940 , n15938 , n15939 );
buf ( n15941 , n15940 );
not ( n15942 , n15941 );
nand ( n15943 , n15937 , n15942 );
nand ( n15944 , n15645 , n15943 );
not ( n15945 , n15944 );
buf ( n15946 , n15945 );
buf ( n15947 , n15920 );
buf ( n15948 , n15947 );
buf ( n15949 , n15948 );
and ( n15950 , n15949 , n15650 );
buf ( n15951 , n15950 );
xor ( n15952 , n15658 , n15664 );
and ( n15953 , n15952 , n15918 );
and ( n15954 , n15658 , n15664 );
or ( n15955 , n15953 , n15954 );
buf ( n15956 , n15955 );
xor ( n15957 , n15767 , n15784 );
and ( n15958 , n15957 , n15805 );
and ( n15959 , n15767 , n15784 );
or ( n15960 , n15958 , n15959 );
buf ( n15961 , n15960 );
buf ( n15962 , n15961 );
buf ( n15963 , n15861 );
not ( n15964 , n15963 );
buf ( n15965 , n1551 );
not ( n15966 , n15965 );
or ( n15967 , n15964 , n15966 );
buf ( n15968 , n1560 );
buf ( n15969 , n781 );
buf ( n15970 , n802 );
xor ( n15971 , n15969 , n15970 );
buf ( n15972 , n15971 );
buf ( n15973 , n15972 );
nand ( n15974 , n15968 , n15973 );
buf ( n15975 , n15974 );
buf ( n15976 , n15975 );
nand ( n15977 , n15967 , n15976 );
buf ( n15978 , n15977 );
buf ( n15979 , n15978 );
buf ( n15980 , n15777 );
not ( n15981 , n15980 );
buf ( n15982 , n10509 );
not ( n15983 , n15982 );
or ( n15984 , n15981 , n15983 );
buf ( n15985 , n3662 );
buf ( n15986 , n783 );
buf ( n15987 , n800 );
xor ( n15988 , n15986 , n15987 );
buf ( n15989 , n15988 );
buf ( n15990 , n15989 );
nand ( n15991 , n15985 , n15990 );
buf ( n15992 , n15991 );
buf ( n15993 , n15992 );
nand ( n15994 , n15984 , n15993 );
buf ( n15995 , n15994 );
buf ( n15996 , n15995 );
xor ( n15997 , n15979 , n15996 );
buf ( n15998 , n12889 );
not ( n15999 , n15998 );
buf ( n16000 , n15999 );
buf ( n16001 , n16000 );
buf ( n16002 , n15899 );
not ( n16003 , n16002 );
buf ( n16004 , n16003 );
buf ( n16005 , n16004 );
or ( n16006 , n16001 , n16005 );
buf ( n16007 , n5272 );
not ( n16008 , n16007 );
buf ( n16009 , n16008 );
buf ( n16010 , n16009 );
buf ( n16011 , n773 );
buf ( n16012 , n810 );
xor ( n16013 , n16011 , n16012 );
buf ( n16014 , n16013 );
buf ( n16015 , n16014 );
not ( n16016 , n16015 );
buf ( n16017 , n16016 );
buf ( n16018 , n16017 );
or ( n16019 , n16010 , n16018 );
nand ( n16020 , n16006 , n16019 );
buf ( n16021 , n16020 );
buf ( n16022 , n16021 );
xor ( n16023 , n15997 , n16022 );
buf ( n16024 , n16023 );
buf ( n16025 , n16024 );
xor ( n16026 , n15962 , n16025 );
buf ( n16027 , n785 );
buf ( n16028 , n800 );
and ( n16029 , n16027 , n16028 );
buf ( n16030 , n16029 );
buf ( n16031 , n16030 );
buf ( n16032 , n15692 );
not ( n16033 , n16032 );
buf ( n16034 , n2709 );
not ( n16035 , n16034 );
or ( n16036 , n16033 , n16035 );
buf ( n16037 , n2713 );
buf ( n16038 , n775 );
buf ( n16039 , n808 );
xor ( n16040 , n16038 , n16039 );
buf ( n16041 , n16040 );
buf ( n16042 , n16041 );
nand ( n16043 , n16037 , n16042 );
buf ( n16044 , n16043 );
buf ( n16045 , n16044 );
nand ( n16046 , n16036 , n16045 );
buf ( n16047 , n16046 );
buf ( n16048 , n16047 );
xor ( n16049 , n16031 , n16048 );
buf ( n16050 , n15798 );
not ( n16051 , n16050 );
buf ( n16052 , n15790 );
not ( n16053 , n16052 );
or ( n16054 , n16051 , n16053 );
buf ( n16055 , n1940 );
buf ( n16056 , n769 );
buf ( n16057 , n814 );
xor ( n16058 , n16056 , n16057 );
buf ( n16059 , n16058 );
buf ( n16060 , n16059 );
nand ( n16061 , n16055 , n16060 );
buf ( n16062 , n16061 );
buf ( n16063 , n16062 );
nand ( n16064 , n16054 , n16063 );
buf ( n16065 , n16064 );
buf ( n16066 , n16065 );
xor ( n16067 , n16049 , n16066 );
buf ( n16068 , n16067 );
buf ( n16069 , n16068 );
xor ( n16070 , n16026 , n16069 );
buf ( n16071 , n16070 );
buf ( n16072 , n15842 );
not ( n16073 , n16072 );
buf ( n16074 , n7628 );
not ( n16075 , n16074 );
or ( n16076 , n16073 , n16075 );
buf ( n16077 , n2010 );
buf ( n16078 , n816 );
nand ( n16079 , n16077 , n16078 );
buf ( n16080 , n16079 );
buf ( n16081 , n16080 );
nand ( n16082 , n16076 , n16081 );
buf ( n16083 , n16082 );
buf ( n16084 , n15831 );
not ( n16085 , n16084 );
buf ( n16086 , n15848 );
not ( n16087 , n16086 );
or ( n16088 , n16085 , n16087 );
buf ( n16089 , n15848 );
buf ( n16090 , n15831 );
or ( n16091 , n16089 , n16090 );
buf ( n16092 , n15820 );
nand ( n16093 , n16091 , n16092 );
buf ( n16094 , n16093 );
buf ( n16095 , n16094 );
nand ( n16096 , n16088 , n16095 );
buf ( n16097 , n16096 );
xor ( n16098 , n16083 , n16097 );
xor ( n16099 , n15868 , n15888 );
and ( n16100 , n16099 , n15906 );
and ( n16101 , n15868 , n15888 );
or ( n16102 , n16100 , n16101 );
buf ( n16103 , n16102 );
xor ( n16104 , n16098 , n16103 );
buf ( n16105 , n16104 );
not ( n16106 , n16105 );
xor ( n16107 , n15808 , n15850 );
and ( n16108 , n16107 , n15909 );
and ( n16109 , n15808 , n15850 );
or ( n16110 , n16108 , n16109 );
buf ( n16111 , n16110 );
buf ( n16112 , n16111 );
not ( n16113 , n16112 );
or ( n16114 , n16106 , n16113 );
buf ( n16115 , n16111 );
buf ( n16116 , n16104 );
or ( n16117 , n16115 , n16116 );
nand ( n16118 , n16114 , n16117 );
buf ( n16119 , n16118 );
xor ( n16120 , n16071 , n16119 );
buf ( n16121 , n16120 );
xor ( n16122 , n15541 , n15683 );
and ( n16123 , n16122 , n15696 );
and ( n16124 , n15541 , n15683 );
or ( n16125 , n16123 , n16124 );
buf ( n16126 , n16125 );
buf ( n16127 , n15881 );
not ( n16128 , n16127 );
buf ( n16129 , n15873 );
not ( n16130 , n16129 );
or ( n16131 , n16128 , n16130 );
buf ( n16132 , n11137 );
buf ( n16133 , n779 );
buf ( n16134 , n804 );
xor ( n16135 , n16133 , n16134 );
buf ( n16136 , n16135 );
buf ( n16137 , n16136 );
nand ( n16138 , n16132 , n16137 );
buf ( n16139 , n16138 );
buf ( n16140 , n16139 );
nand ( n16141 , n16131 , n16140 );
buf ( n16142 , n16141 );
buf ( n16143 , n16142 );
buf ( n16144 , n15816 );
not ( n16145 , n16144 );
buf ( n16146 , n2066 );
not ( n16147 , n16146 );
or ( n16148 , n16145 , n16147 );
buf ( n16149 , n14331 );
buf ( n16150 , n771 );
buf ( n16151 , n812 );
xor ( n16152 , n16150 , n16151 );
buf ( n16153 , n16152 );
buf ( n16154 , n16153 );
nand ( n16155 , n16149 , n16154 );
buf ( n16156 , n16155 );
buf ( n16157 , n16156 );
nand ( n16158 , n16148 , n16157 );
buf ( n16159 , n16158 );
buf ( n16160 , n16159 );
xor ( n16161 , n16143 , n16160 );
buf ( n16162 , n15679 );
not ( n16163 , n16162 );
buf ( n16164 , n14278 );
not ( n16165 , n16164 );
or ( n16166 , n16163 , n16165 );
buf ( n16167 , n14284 );
buf ( n16168 , n777 );
buf ( n16169 , n806 );
xor ( n16170 , n16168 , n16169 );
buf ( n16171 , n16170 );
buf ( n16172 , n16171 );
nand ( n16173 , n16167 , n16172 );
buf ( n16174 , n16173 );
buf ( n16175 , n16174 );
nand ( n16176 , n16166 , n16175 );
buf ( n16177 , n16176 );
buf ( n16178 , n16177 );
xor ( n16179 , n16161 , n16178 );
buf ( n16180 , n16179 );
buf ( n16181 , n16180 );
xor ( n16182 , n16126 , n16181 );
xor ( n16183 , n15745 , n15751 );
and ( n16184 , n16183 , n15758 );
and ( n16185 , n15745 , n15751 );
or ( n16186 , n16184 , n16185 );
buf ( n16187 , n16186 );
buf ( n16188 , n16187 );
xor ( n16189 , n16182 , n16188 );
buf ( n16190 , n16189 );
buf ( n16191 , n16190 );
xor ( n16192 , n15698 , n15717 );
and ( n16193 , n16192 , n15724 );
and ( n16194 , n15698 , n15717 );
or ( n16195 , n16193 , n16194 );
buf ( n16196 , n16195 );
buf ( n16197 , n16196 );
xor ( n16198 , n16191 , n16197 );
xor ( n16199 , n15739 , n15761 );
and ( n16200 , n16199 , n15912 );
and ( n16201 , n15739 , n15761 );
or ( n16202 , n16200 , n16201 );
buf ( n16203 , n16202 );
buf ( n16204 , n16203 );
xor ( n16205 , n16198 , n16204 );
buf ( n16206 , n16205 );
buf ( n16207 , n16206 );
xor ( n16208 , n16121 , n16207 );
xor ( n16209 , n15671 , n15727 );
and ( n16210 , n16209 , n15915 );
and ( n16211 , n15671 , n15727 );
or ( n16212 , n16210 , n16211 );
buf ( n16213 , n16212 );
buf ( n16214 , n16213 );
xor ( n16215 , n16208 , n16214 );
buf ( n16216 , n16215 );
xor ( n16217 , n15956 , n16216 );
buf ( n16218 , n16217 );
nor ( n16219 , n15951 , n16218 );
buf ( n16220 , n16219 );
buf ( n16221 , n16220 );
not ( n16222 , n16221 );
buf ( n16223 , n16222 );
buf ( n16224 , n16223 );
and ( n16225 , n15946 , n16224 );
buf ( n16226 , n16225 );
buf ( n16227 , n16226 );
nand ( n16228 , n15327 , n16227 );
buf ( n16229 , n16228 );
buf ( n16230 , n16229 );
nor ( n16231 , n13772 , n16230 );
buf ( n16232 , n16231 );
buf ( n16233 , n16232 );
not ( n16234 , n16233 );
buf ( n16235 , n10417 );
not ( n16236 , n16235 );
or ( n16237 , n16234 , n16236 );
buf ( n16238 , n16229 );
not ( n16239 , n16238 );
buf ( n16240 , n16239 );
buf ( n16241 , n16240 );
not ( n16242 , n16241 );
buf ( n16243 , n13243 );
buf ( n16244 , n13248 );
nand ( n16245 , n16243 , n16244 );
buf ( n16246 , n16245 );
not ( n16247 , n16246 );
not ( n16248 , n13674 );
and ( n16249 , n16247 , n16248 );
buf ( n16250 , n13671 );
buf ( n16251 , n16250 );
buf ( n16252 , n16251 );
and ( n16253 , n16252 , n13253 );
nor ( n16254 , n16249 , n16253 );
buf ( n16255 , n16254 );
buf ( n16256 , n16255 );
buf ( n16257 , n16256 );
nand ( n16258 , n12807 , n12805 );
not ( n16259 , n16258 );
buf ( n16260 , n16259 );
not ( n16261 , n16260 );
buf ( n16262 , n12575 );
not ( n16263 , n16262 );
buf ( n16264 , n16263 );
buf ( n16265 , n16264 );
buf ( n16266 , n12707 );
not ( n16267 , n16266 );
buf ( n16268 , n16267 );
buf ( n16269 , n16268 );
nand ( n16270 , n16265 , n16269 );
buf ( n16271 , n16270 );
buf ( n16272 , n16271 );
not ( n16273 , n16272 );
or ( n16274 , n16261 , n16273 );
buf ( n16275 , n12575 );
buf ( n16276 , n12707 );
nand ( n16277 , n16275 , n16276 );
buf ( n16278 , n16277 );
buf ( n16279 , n16278 );
nand ( n16280 , n16274 , n16279 );
buf ( n16281 , n16280 );
buf ( n16282 , n16281 );
buf ( n16283 , n13677 );
nand ( n16284 , n16282 , n16283 );
buf ( n16285 , n16284 );
nand ( n16286 , n16257 , n16285 );
not ( n16287 , n16286 );
buf ( n16288 , n13680 );
not ( n16289 , n16288 );
buf ( n16290 , n16289 );
nor ( n16291 , n13752 , n13754 );
or ( n16292 , n4349 , n16291 );
nand ( n16293 , n13754 , n13752 );
nand ( n16294 , n16292 , n16293 );
not ( n16295 , n16294 );
nor ( n16296 , n13732 , n13723 );
not ( n16297 , n16296 );
or ( n16298 , n16295 , n16297 );
not ( n16299 , n13732 );
nand ( n16300 , n13711 , n13722 );
not ( n16301 , n16300 );
and ( n16302 , n16299 , n16301 );
buf ( n16303 , n13729 );
buf ( n16304 , n13727 );
nand ( n16305 , n16303 , n16304 );
buf ( n16306 , n16305 );
buf ( n16307 , n16306 );
not ( n16308 , n16307 );
buf ( n16309 , n16308 );
nor ( n16310 , n16302 , n16309 );
nand ( n16311 , n16298 , n16310 );
nand ( n16312 , n16290 , n16311 );
nand ( n16313 , n16287 , n16312 );
buf ( n16314 , n16313 );
not ( n16315 , n16314 );
or ( n16316 , n16242 , n16315 );
buf ( n16317 , n14523 );
not ( n16318 , n16317 );
buf ( n16319 , n16318 );
buf ( n16320 , n16319 );
buf ( n16321 , n14127 );
not ( n16322 , n16321 );
buf ( n16323 , n16322 );
buf ( n16324 , n16323 );
nand ( n16325 , n16320 , n16324 );
buf ( n16326 , n16325 );
not ( n16327 , n16326 );
nand ( n16328 , n14541 , n14546 );
not ( n16329 , n16328 );
not ( n16330 , n16329 );
or ( n16331 , n16327 , n16330 );
nand ( n16332 , n14523 , n14127 );
nand ( n16333 , n16331 , n16332 );
buf ( n16334 , n16333 );
buf ( n16335 , n15299 );
buf ( n16336 , n15319 );
nor ( n16337 , n16335 , n16336 );
buf ( n16338 , n16337 );
buf ( n16339 , n16338 );
nand ( n16340 , n16334 , n16339 );
buf ( n16341 , n16340 );
buf ( n16342 , n16341 );
buf ( n16343 , n15316 );
not ( n16344 , n16343 );
buf ( n16345 , n16344 );
buf ( n16346 , n16345 );
buf ( n16347 , n15304 );
not ( n16348 , n16347 );
buf ( n16349 , n16348 );
buf ( n16350 , n16349 );
nor ( n16351 , n16346 , n16350 );
buf ( n16352 , n16351 );
buf ( n16353 , n16352 );
not ( n16354 , n16353 );
buf ( n16355 , n15296 );
not ( n16356 , n16355 );
or ( n16357 , n16354 , n16356 );
not ( n16358 , n15293 );
nand ( n16359 , n16358 , n15279 );
buf ( n16360 , n16359 );
nand ( n16361 , n16357 , n16360 );
buf ( n16362 , n16361 );
buf ( n16363 , n16362 );
not ( n16364 , n16363 );
buf ( n16365 , n16364 );
buf ( n16366 , n16365 );
nand ( n16367 , n16342 , n16366 );
buf ( n16368 , n16367 );
and ( n16369 , n16226 , n16368 );
buf ( n16370 , n16223 );
not ( n16371 , n16370 );
buf ( n16372 , n15643 );
buf ( n16373 , n15638 );
nor ( n16374 , n16372 , n16373 );
buf ( n16375 , n16374 );
buf ( n16376 , n16375 );
not ( n16377 , n16376 );
buf ( n16378 , n15937 );
buf ( n16379 , n15942 );
nand ( n16380 , n16378 , n16379 );
buf ( n16381 , n16380 );
buf ( n16382 , n16381 );
not ( n16383 , n16382 );
or ( n16384 , n16377 , n16383 );
buf ( n16385 , n15936 );
buf ( n16386 , n15941 );
nand ( n16387 , n16385 , n16386 );
buf ( n16388 , n16387 );
buf ( n16389 , n16388 );
nand ( n16390 , n16384 , n16389 );
buf ( n16391 , n16390 );
buf ( n16392 , n16391 );
buf ( n16393 , n16392 );
buf ( n16394 , n16393 );
buf ( n16395 , n16394 );
not ( n16396 , n16395 );
or ( n16397 , n16371 , n16396 );
buf ( n16398 , n15950 );
buf ( n16399 , n16217 );
nand ( n16400 , n16398 , n16399 );
buf ( n16401 , n16400 );
buf ( n16402 , n16401 );
nand ( n16403 , n16397 , n16402 );
buf ( n16404 , n16403 );
nor ( n16405 , n16369 , n16404 );
buf ( n16406 , n16405 );
nand ( n16407 , n16316 , n16406 );
buf ( n16408 , n16407 );
buf ( n16409 , n16408 );
not ( n16410 , n16409 );
buf ( n16411 , n16410 );
buf ( n16412 , n16411 );
nand ( n16413 , n16237 , n16412 );
buf ( n16414 , n16413 );
buf ( n16415 , n16414 );
buf ( n16416 , n16216 );
buf ( n16417 , n15956 );
and ( n16418 , n16416 , n16417 );
buf ( n16419 , n16418 );
buf ( n16420 , n16419 );
not ( n16421 , n16103 );
buf ( n16422 , n16083 );
not ( n16423 , n16422 );
buf ( n16424 , n16423 );
not ( n16425 , n16424 );
or ( n16426 , n16421 , n16425 );
buf ( n16427 , n16103 );
buf ( n16428 , n16424 );
nor ( n16429 , n16427 , n16428 );
buf ( n16430 , n16429 );
buf ( n16431 , n16097 );
not ( n16432 , n16431 );
buf ( n16433 , n16432 );
or ( n16434 , n16430 , n16433 );
nand ( n16435 , n16426 , n16434 );
buf ( n16436 , n16435 );
xor ( n16437 , n15962 , n16025 );
and ( n16438 , n16437 , n16069 );
and ( n16439 , n15962 , n16025 );
or ( n16440 , n16438 , n16439 );
buf ( n16441 , n16440 );
buf ( n16442 , n16441 );
xor ( n16443 , n16436 , n16442 );
xor ( n16444 , n16031 , n16048 );
and ( n16445 , n16444 , n16066 );
and ( n16446 , n16031 , n16048 );
or ( n16447 , n16445 , n16446 );
buf ( n16448 , n16447 );
buf ( n16449 , n16448 );
xor ( n16450 , n16143 , n16160 );
and ( n16451 , n16450 , n16178 );
and ( n16452 , n16143 , n16160 );
or ( n16453 , n16451 , n16452 );
buf ( n16454 , n16453 );
buf ( n16455 , n16454 );
xor ( n16456 , n16449 , n16455 );
buf ( n16457 , n784 );
buf ( n16458 , n800 );
and ( n16459 , n16457 , n16458 );
buf ( n16460 , n16459 );
buf ( n16461 , n16460 );
buf ( n16462 , n16171 );
not ( n16463 , n16462 );
buf ( n16464 , n14278 );
not ( n16465 , n16464 );
or ( n16466 , n16463 , n16465 );
buf ( n16467 , n14284 );
buf ( n16468 , n776 );
buf ( n16469 , n806 );
xor ( n16470 , n16468 , n16469 );
buf ( n16471 , n16470 );
buf ( n16472 , n16471 );
nand ( n16473 , n16467 , n16472 );
buf ( n16474 , n16473 );
buf ( n16475 , n16474 );
nand ( n16476 , n16466 , n16475 );
buf ( n16477 , n16476 );
buf ( n16478 , n16477 );
xor ( n16479 , n16461 , n16478 );
buf ( n16480 , n16153 );
not ( n16481 , n16480 );
buf ( n16482 , n2066 );
not ( n16483 , n16482 );
or ( n16484 , n16481 , n16483 );
not ( n16485 , n14588 );
buf ( n16486 , n16485 );
buf ( n16487 , n770 );
buf ( n16488 , n812 );
xor ( n16489 , n16487 , n16488 );
buf ( n16490 , n16489 );
buf ( n16491 , n16490 );
nand ( n16492 , n16486 , n16491 );
buf ( n16493 , n16492 );
buf ( n16494 , n16493 );
nand ( n16495 , n16484 , n16494 );
buf ( n16496 , n16495 );
buf ( n16497 , n16496 );
xor ( n16498 , n16479 , n16497 );
buf ( n16499 , n16498 );
buf ( n16500 , n16499 );
xor ( n16501 , n16456 , n16500 );
buf ( n16502 , n16501 );
buf ( n16503 , n16502 );
xor ( n16504 , n16443 , n16503 );
buf ( n16505 , n16504 );
buf ( n16506 , n16505 );
buf ( n16507 , n16041 );
not ( n16508 , n16507 );
buf ( n16509 , n2709 );
not ( n16510 , n16509 );
or ( n16511 , n16508 , n16510 );
buf ( n16512 , n2713 );
buf ( n16513 , n774 );
buf ( n16514 , n808 );
xor ( n16515 , n16513 , n16514 );
buf ( n16516 , n16515 );
buf ( n16517 , n16516 );
nand ( n16518 , n16512 , n16517 );
buf ( n16519 , n16518 );
buf ( n16520 , n16519 );
nand ( n16521 , n16511 , n16520 );
buf ( n16522 , n16521 );
buf ( n16523 , n16522 );
buf ( n16524 , n15972 );
not ( n16525 , n16524 );
buf ( n16526 , n3109 );
not ( n16527 , n16526 );
or ( n16528 , n16525 , n16527 );
buf ( n16529 , n1560 );
buf ( n16530 , n780 );
buf ( n16531 , n802 );
xor ( n16532 , n16530 , n16531 );
buf ( n16533 , n16532 );
buf ( n16534 , n16533 );
nand ( n16535 , n16529 , n16534 );
buf ( n16536 , n16535 );
buf ( n16537 , n16536 );
nand ( n16538 , n16528 , n16537 );
buf ( n16539 , n16538 );
buf ( n16540 , n16539 );
xor ( n16541 , n16523 , n16540 );
buf ( n16542 , n15989 );
not ( n16543 , n16542 );
buf ( n16544 , n10509 );
not ( n16545 , n16544 );
or ( n16546 , n16543 , n16545 );
buf ( n16547 , n3662 );
buf ( n16548 , n782 );
buf ( n16549 , n800 );
xor ( n16550 , n16548 , n16549 );
buf ( n16551 , n16550 );
buf ( n16552 , n16551 );
nand ( n16553 , n16547 , n16552 );
buf ( n16554 , n16553 );
buf ( n16555 , n16554 );
nand ( n16556 , n16546 , n16555 );
buf ( n16557 , n16556 );
buf ( n16558 , n16557 );
xor ( n16559 , n16541 , n16558 );
buf ( n16560 , n16559 );
buf ( n16561 , n16560 );
buf ( n16562 , n16059 );
not ( n16563 , n16562 );
buf ( n16564 , n15790 );
not ( n16565 , n16564 );
or ( n16566 , n16563 , n16565 );
buf ( n16567 , n1940 );
buf ( n16568 , n768 );
buf ( n16569 , n814 );
xor ( n16570 , n16568 , n16569 );
buf ( n16571 , n16570 );
buf ( n16572 , n16571 );
nand ( n16573 , n16567 , n16572 );
buf ( n16574 , n16573 );
buf ( n16575 , n16574 );
nand ( n16576 , n16566 , n16575 );
buf ( n16577 , n16576 );
buf ( n16578 , n16577 );
buf ( n16579 , n2532 );
buf ( n16580 , n7628 );
or ( n16581 , n16579 , n16580 );
buf ( n16582 , n816 );
nand ( n16583 , n16581 , n16582 );
buf ( n16584 , n16583 );
buf ( n16585 , n16584 );
xor ( n16586 , n16578 , n16585 );
buf ( n16587 , n16014 );
not ( n16588 , n16587 );
buf ( n16589 , n12889 );
not ( n16590 , n16589 );
or ( n16591 , n16588 , n16590 );
buf ( n16592 , n16009 );
not ( n16593 , n16592 );
buf ( n16594 , n16593 );
buf ( n16595 , n16594 );
buf ( n16596 , n772 );
buf ( n16597 , n810 );
xor ( n16598 , n16596 , n16597 );
buf ( n16599 , n16598 );
buf ( n16600 , n16599 );
nand ( n16601 , n16595 , n16600 );
buf ( n16602 , n16601 );
buf ( n16603 , n16602 );
nand ( n16604 , n16591 , n16603 );
buf ( n16605 , n16604 );
buf ( n16606 , n16605 );
xor ( n16607 , n16586 , n16606 );
buf ( n16608 , n16607 );
buf ( n16609 , n16608 );
xor ( n16610 , n16561 , n16609 );
buf ( n16611 , n16083 );
buf ( n16612 , n16136 );
not ( n16613 , n16612 );
buf ( n16614 , n15873 );
not ( n16615 , n16614 );
or ( n16616 , n16613 , n16615 );
buf ( n16617 , n11137 );
buf ( n16618 , n778 );
buf ( n16619 , n804 );
xor ( n16620 , n16618 , n16619 );
buf ( n16621 , n16620 );
buf ( n16622 , n16621 );
nand ( n16623 , n16617 , n16622 );
buf ( n16624 , n16623 );
buf ( n16625 , n16624 );
nand ( n16626 , n16616 , n16625 );
buf ( n16627 , n16626 );
buf ( n16628 , n16627 );
xor ( n16629 , n16611 , n16628 );
xor ( n16630 , n15979 , n15996 );
and ( n16631 , n16630 , n16022 );
and ( n16632 , n15979 , n15996 );
or ( n16633 , n16631 , n16632 );
buf ( n16634 , n16633 );
buf ( n16635 , n16634 );
xor ( n16636 , n16629 , n16635 );
buf ( n16637 , n16636 );
buf ( n16638 , n16637 );
xor ( n16639 , n16610 , n16638 );
buf ( n16640 , n16639 );
buf ( n16641 , n16640 );
xor ( n16642 , n16126 , n16181 );
and ( n16643 , n16642 , n16188 );
and ( n16644 , n16126 , n16181 );
or ( n16645 , n16643 , n16644 );
buf ( n16646 , n16645 );
buf ( n16647 , n16646 );
xor ( n16648 , n16641 , n16647 );
buf ( n16649 , n16111 );
buf ( n16650 , n16104 );
not ( n16651 , n16650 );
buf ( n16652 , n16651 );
buf ( n16653 , n16652 );
or ( n16654 , n16649 , n16653 );
buf ( n16655 , n16071 );
nand ( n16656 , n16654 , n16655 );
buf ( n16657 , n16656 );
buf ( n16658 , n16657 );
buf ( n16659 , n16111 );
buf ( n16660 , n16652 );
nand ( n16661 , n16659 , n16660 );
buf ( n16662 , n16661 );
buf ( n16663 , n16662 );
nand ( n16664 , n16658 , n16663 );
buf ( n16665 , n16664 );
buf ( n16666 , n16665 );
xor ( n16667 , n16648 , n16666 );
buf ( n16668 , n16667 );
buf ( n16669 , n16668 );
xor ( n16670 , n16506 , n16669 );
xor ( n16671 , n16191 , n16197 );
and ( n16672 , n16671 , n16204 );
and ( n16673 , n16191 , n16197 );
or ( n16674 , n16672 , n16673 );
buf ( n16675 , n16674 );
buf ( n16676 , n16675 );
xor ( n16677 , n16670 , n16676 );
buf ( n16678 , n16677 );
buf ( n16679 , n16678 );
xor ( n16680 , n16121 , n16207 );
and ( n16681 , n16680 , n16214 );
and ( n16682 , n16121 , n16207 );
or ( n16683 , n16681 , n16682 );
buf ( n16684 , n16683 );
buf ( n16685 , n16684 );
xor ( n16686 , n16679 , n16685 );
buf ( n16687 , n16686 );
buf ( n16688 , n16687 );
nand ( n16689 , n16420 , n16688 );
buf ( n16690 , n16689 );
buf ( n16691 , n16690 );
not ( n16692 , n16691 );
buf ( n16693 , n16419 );
buf ( n16694 , n16687 );
nor ( n16695 , n16693 , n16694 );
buf ( n16696 , n16695 );
buf ( n16697 , n16696 );
nor ( n16698 , n16692 , n16697 );
buf ( n16699 , n16698 );
buf ( n16700 , n16699 );
and ( n16701 , n16415 , n16700 );
not ( n16702 , n16415 );
buf ( n16703 , n16699 );
not ( n16704 , n16703 );
buf ( n16705 , n16704 );
buf ( n16706 , n16705 );
and ( n16707 , n16702 , n16706 );
nor ( n16708 , n16701 , n16707 );
buf ( n16709 , n16708 );
buf ( n16710 , n16709 );
buf ( n16711 , n13768 );
not ( n16712 , n16711 );
buf ( n16713 , n16712 );
buf ( n16714 , n16713 );
buf ( n16715 , n15325 );
not ( n16716 , n16715 );
not ( n16717 , n15635 );
nand ( n16718 , n16717 , n15643 );
buf ( n16719 , n16718 );
nand ( n16720 , n16716 , n16719 );
buf ( n16721 , n16720 );
buf ( n16722 , n16721 );
nor ( n16723 , n16714 , n16722 );
buf ( n16724 , n16723 );
buf ( n16725 , n16724 );
not ( n16726 , n16725 );
buf ( n16727 , n10427 );
not ( n16728 , n16727 );
or ( n16729 , n16726 , n16728 );
buf ( n16730 , n16721 );
not ( n16731 , n16730 );
buf ( n16732 , n16731 );
buf ( n16733 , n16732 );
not ( n16734 , n16733 );
not ( n16735 , n16286 );
nand ( n16736 , n16735 , n16312 );
buf ( n16737 , n16736 );
not ( n16738 , n16737 );
or ( n16739 , n16734 , n16738 );
buf ( n16740 , n16718 );
not ( n16741 , n16740 );
buf ( n16742 , n16368 );
not ( n16743 , n16742 );
or ( n16744 , n16741 , n16743 );
not ( n16745 , n16375 );
buf ( n16746 , n16745 );
nand ( n16747 , n16744 , n16746 );
buf ( n16748 , n16747 );
buf ( n16749 , n16748 );
not ( n16750 , n16749 );
buf ( n16751 , n16750 );
buf ( n16752 , n16751 );
nand ( n16753 , n16739 , n16752 );
buf ( n16754 , n16753 );
buf ( n16755 , n16754 );
not ( n16756 , n16755 );
buf ( n16757 , n16756 );
buf ( n16758 , n16757 );
nand ( n16759 , n16729 , n16758 );
buf ( n16760 , n16759 );
buf ( n16761 , n16760 );
buf ( n16762 , n16381 );
buf ( n16763 , n16762 );
buf ( n16764 , n16388 );
and ( n16765 , n16763 , n16764 );
buf ( n16766 , n16765 );
buf ( n16767 , n16766 );
and ( n16768 , n16761 , n16767 );
not ( n16769 , n16761 );
buf ( n16770 , n16766 );
not ( n16771 , n16770 );
buf ( n16772 , n16771 );
buf ( n16773 , n16772 );
and ( n16774 , n16769 , n16773 );
nor ( n16775 , n16768 , n16774 );
buf ( n16776 , n16775 );
buf ( n16777 , n16776 );
buf ( n16778 , n16220 );
buf ( n16779 , n16696 );
nor ( n16780 , n16778 , n16779 );
buf ( n16781 , n16780 );
nand ( n16782 , n16781 , n15945 );
not ( n16783 , n16782 );
nand ( n16784 , n15322 , n14550 , n16783 );
not ( n16785 , n16784 );
not ( n16786 , n16341 );
not ( n16787 , n16782 );
and ( n16788 , n16786 , n16787 );
buf ( n16789 , n16362 );
not ( n16790 , n16789 );
buf ( n16791 , n16783 );
not ( n16792 , n16791 );
or ( n16793 , n16790 , n16792 );
not ( n16794 , n16781 );
not ( n16795 , n16391 );
or ( n16796 , n16794 , n16795 );
not ( n16797 , n16401 );
not ( n16798 , n16696 );
and ( n16799 , n16797 , n16798 );
buf ( n16800 , n16690 );
not ( n16801 , n16800 );
buf ( n16802 , n16801 );
nor ( n16803 , n16799 , n16802 );
nand ( n16804 , n16796 , n16803 );
buf ( n16805 , n16804 );
not ( n16806 , n16805 );
buf ( n16807 , n16806 );
buf ( n16808 , n16807 );
nand ( n16809 , n16793 , n16808 );
buf ( n16810 , n16809 );
nor ( n16811 , n16788 , n16810 );
not ( n16812 , n16811 );
or ( n16813 , n16785 , n16812 );
buf ( n16814 , n16285 );
buf ( n16815 , n16807 );
nand ( n16816 , n16814 , n16815 );
buf ( n16817 , n16816 );
not ( n16818 , n16817 );
buf ( n16819 , n16341 );
not ( n16820 , n16819 );
buf ( n16821 , n16254 );
buf ( n16822 , n16365 );
nand ( n16823 , n16821 , n16822 );
buf ( n16824 , n16823 );
buf ( n16825 , n16824 );
nor ( n16826 , n16820 , n16825 );
buf ( n16827 , n16826 );
nand ( n16828 , n16290 , n16311 );
nand ( n16829 , n16818 , n16827 , n16828 );
nand ( n16830 , n16813 , n16829 );
buf ( n16831 , n16830 );
not ( n16832 , n16831 );
buf ( n16833 , n16832 );
buf ( n16834 , n16833 );
buf ( n16835 , n775 );
buf ( n16836 , n804 );
xor ( n16837 , n16835 , n16836 );
buf ( n16838 , n16837 );
buf ( n16839 , n16838 );
not ( n16840 , n16839 );
buf ( n16841 , n15873 );
not ( n16842 , n16841 );
or ( n16843 , n16840 , n16842 );
buf ( n16844 , n11137 );
buf ( n16845 , n774 );
buf ( n16846 , n804 );
xor ( n16847 , n16845 , n16846 );
buf ( n16848 , n16847 );
buf ( n16849 , n16848 );
nand ( n16850 , n16844 , n16849 );
buf ( n16851 , n16850 );
buf ( n16852 , n16851 );
nand ( n16853 , n16843 , n16852 );
buf ( n16854 , n16853 );
buf ( n16855 , n16854 );
buf ( n16856 , n800 );
buf ( n16857 , n780 );
and ( n16858 , n16856 , n16857 );
buf ( n16859 , n16858 );
buf ( n16860 , n16859 );
xor ( n16861 , n16855 , n16860 );
buf ( n16862 , n16861 );
buf ( n16863 , n16862 );
buf ( n16864 , n771 );
buf ( n16865 , n808 );
xor ( n16866 , n16864 , n16865 );
buf ( n16867 , n16866 );
buf ( n16868 , n16867 );
not ( n16869 , n16868 );
buf ( n16870 , n2709 );
not ( n16871 , n16870 );
or ( n16872 , n16869 , n16871 );
buf ( n16873 , n2713 );
xor ( n16874 , n808 , n770 );
buf ( n16875 , n16874 );
nand ( n16876 , n16873 , n16875 );
buf ( n16877 , n16876 );
buf ( n16878 , n16877 );
nand ( n16879 , n16872 , n16878 );
buf ( n16880 , n16879 );
buf ( n16881 , n16880 );
xor ( n16882 , n16863 , n16881 );
buf ( n16883 , n16882 );
buf ( n16884 , n16883 );
buf ( n16885 , n768 );
buf ( n16886 , n812 );
xor ( n16887 , n16885 , n16886 );
buf ( n16888 , n16887 );
buf ( n16889 , n16888 );
not ( n16890 , n16889 );
buf ( n16891 , n2066 );
not ( n16892 , n16891 );
or ( n16893 , n16890 , n16892 );
buf ( n16894 , n14331 );
buf ( n16895 , n812 );
nand ( n16896 , n16894 , n16895 );
buf ( n16897 , n16896 );
buf ( n16898 , n16897 );
nand ( n16899 , n16893 , n16898 );
buf ( n16900 , n16899 );
buf ( n16901 , n16900 );
not ( n16902 , n16901 );
buf ( n16903 , n16902 );
buf ( n16904 , n16903 );
xor ( n16905 , n16856 , n16857 );
buf ( n16906 , n16905 );
buf ( n16907 , n16906 );
not ( n16908 , n16907 );
buf ( n16909 , n10509 );
not ( n16910 , n16909 );
or ( n16911 , n16908 , n16910 );
buf ( n16912 , n3662 );
buf ( n16913 , n800 );
buf ( n16914 , n779 );
xor ( n16915 , n16913 , n16914 );
buf ( n16916 , n16915 );
buf ( n16917 , n16916 );
nand ( n16918 , n16912 , n16917 );
buf ( n16919 , n16918 );
buf ( n16920 , n16919 );
nand ( n16921 , n16911 , n16920 );
buf ( n16922 , n16921 );
buf ( n16923 , n16922 );
xor ( n16924 , n16904 , n16923 );
buf ( n16925 , n15790 );
not ( n16926 , n16925 );
buf ( n16927 , n16926 );
buf ( n16928 , n16927 );
buf ( n16929 , n1940 );
not ( n16930 , n16929 );
buf ( n16931 , n16930 );
buf ( n16932 , n16931 );
and ( n16933 , n16928 , n16932 );
buf ( n16934 , n814 );
not ( n16935 , n16934 );
buf ( n16936 , n16935 );
buf ( n16937 , n16936 );
nor ( n16938 , n16933 , n16937 );
buf ( n16939 , n16938 );
buf ( n16940 , n16939 );
not ( n16941 , n16940 );
buf ( n16942 , n2709 );
buf ( n16943 , n773 );
buf ( n16944 , n808 );
xor ( n16945 , n16943 , n16944 );
buf ( n16946 , n16945 );
buf ( n16947 , n16946 );
and ( n16948 , n16942 , n16947 );
buf ( n16949 , n2713 );
xor ( n16950 , n808 , n772 );
buf ( n16951 , n16950 );
and ( n16952 , n16949 , n16951 );
nor ( n16953 , n16948 , n16952 );
buf ( n16954 , n16953 );
buf ( n16955 , n16954 );
not ( n16956 , n16955 );
or ( n16957 , n16941 , n16956 );
buf ( n16958 , n769 );
buf ( n16959 , n812 );
xor ( n16960 , n16958 , n16959 );
buf ( n16961 , n16960 );
buf ( n16962 , n16961 );
not ( n16963 , n16962 );
buf ( n16964 , n2066 );
not ( n16965 , n16964 );
or ( n16966 , n16963 , n16965 );
buf ( n16967 , n16485 );
buf ( n16968 , n16888 );
nand ( n16969 , n16967 , n16968 );
buf ( n16970 , n16969 );
buf ( n16971 , n16970 );
nand ( n16972 , n16966 , n16971 );
buf ( n16973 , n16972 );
buf ( n16974 , n16973 );
nand ( n16975 , n16957 , n16974 );
buf ( n16976 , n16975 );
buf ( n16977 , n16976 );
buf ( n16978 , n16939 );
not ( n16979 , n16978 );
buf ( n16980 , n16954 );
not ( n16981 , n16980 );
buf ( n16982 , n16981 );
buf ( n16983 , n16982 );
nand ( n16984 , n16979 , n16983 );
buf ( n16985 , n16984 );
buf ( n16986 , n16985 );
nand ( n16987 , n16977 , n16986 );
buf ( n16988 , n16987 );
buf ( n16989 , n16988 );
and ( n16990 , n16924 , n16989 );
and ( n16991 , n16904 , n16923 );
or ( n16992 , n16990 , n16991 );
buf ( n16993 , n16992 );
buf ( n16994 , n16993 );
xor ( n16995 , n16884 , n16994 );
buf ( n16996 , n777 );
buf ( n16997 , n802 );
xor ( n16998 , n16996 , n16997 );
buf ( n16999 , n16998 );
buf ( n17000 , n16999 );
not ( n17001 , n17000 );
buf ( n17002 , n3109 );
not ( n17003 , n17002 );
or ( n17004 , n17001 , n17003 );
buf ( n17005 , n1560 );
xor ( n17006 , n802 , n776 );
buf ( n17007 , n17006 );
nand ( n17008 , n17005 , n17007 );
buf ( n17009 , n17008 );
buf ( n17010 , n17009 );
nand ( n17011 , n17004 , n17010 );
buf ( n17012 , n17011 );
buf ( n17013 , n16916 );
not ( n17014 , n17013 );
buf ( n17015 , n10509 );
not ( n17016 , n17015 );
or ( n17017 , n17014 , n17016 );
buf ( n17018 , n3662 );
buf ( n17019 , n800 );
buf ( n17020 , n778 );
xor ( n17021 , n17019 , n17020 );
buf ( n17022 , n17021 );
buf ( n17023 , n17022 );
nand ( n17024 , n17018 , n17023 );
buf ( n17025 , n17024 );
buf ( n17026 , n17025 );
nand ( n17027 , n17017 , n17026 );
buf ( n17028 , n17027 );
xor ( n17029 , n17012 , n17028 );
buf ( n17030 , n17029 );
buf ( n17031 , n16900 );
and ( n17032 , n17030 , n17031 );
not ( n17033 , n17030 );
buf ( n17034 , n16903 );
and ( n17035 , n17033 , n17034 );
nor ( n17036 , n17032 , n17035 );
buf ( n17037 , n17036 );
buf ( n17038 , n17037 );
xor ( n17039 , n16995 , n17038 );
buf ( n17040 , n17039 );
buf ( n17041 , n17040 );
buf ( n17042 , n16950 );
not ( n17043 , n17042 );
buf ( n17044 , n2709 );
not ( n17045 , n17044 );
or ( n17046 , n17043 , n17045 );
buf ( n17047 , n2713 );
buf ( n17048 , n16867 );
nand ( n17049 , n17047 , n17048 );
buf ( n17050 , n17049 );
buf ( n17051 , n17050 );
nand ( n17052 , n17046 , n17051 );
buf ( n17053 , n17052 );
buf ( n17054 , n776 );
buf ( n17055 , n804 );
xor ( n17056 , n17054 , n17055 );
buf ( n17057 , n17056 );
buf ( n17058 , n17057 );
not ( n17059 , n17058 );
buf ( n17060 , n15873 );
not ( n17061 , n17060 );
or ( n17062 , n17059 , n17061 );
buf ( n17063 , n11137 );
buf ( n17064 , n16838 );
nand ( n17065 , n17063 , n17064 );
buf ( n17066 , n17065 );
buf ( n17067 , n17066 );
nand ( n17068 , n17062 , n17067 );
buf ( n17069 , n17068 );
buf ( n17070 , n17069 );
xor ( n17071 , n17053 , n17070 );
buf ( n17072 , n778 );
buf ( n17073 , n802 );
xor ( n17074 , n17072 , n17073 );
buf ( n17075 , n17074 );
buf ( n17076 , n17075 );
not ( n17077 , n17076 );
buf ( n17078 , n3109 );
not ( n17079 , n17078 );
or ( n17080 , n17077 , n17079 );
buf ( n17081 , n1560 );
buf ( n17082 , n16999 );
nand ( n17083 , n17081 , n17082 );
buf ( n17084 , n17083 );
buf ( n17085 , n17084 );
nand ( n17086 , n17080 , n17085 );
buf ( n17087 , n17086 );
not ( n17088 , n17087 );
xor ( n17089 , n17071 , n17088 );
not ( n17090 , n17089 );
not ( n17091 , n17090 );
buf ( n17092 , n777 );
buf ( n17093 , n804 );
xor ( n17094 , n17092 , n17093 );
buf ( n17095 , n17094 );
buf ( n17096 , n17095 );
not ( n17097 , n17096 );
buf ( n17098 , n15873 );
not ( n17099 , n17098 );
or ( n17100 , n17097 , n17099 );
buf ( n17101 , n11137 );
buf ( n17102 , n17057 );
nand ( n17103 , n17101 , n17102 );
buf ( n17104 , n17103 );
buf ( n17105 , n17104 );
nand ( n17106 , n17100 , n17105 );
buf ( n17107 , n17106 );
buf ( n17108 , n17107 );
buf ( n17109 , n779 );
buf ( n17110 , n802 );
xor ( n17111 , n17109 , n17110 );
buf ( n17112 , n17111 );
buf ( n17113 , n17112 );
not ( n17114 , n17113 );
buf ( n17115 , n3109 );
not ( n17116 , n17115 );
or ( n17117 , n17114 , n17116 );
buf ( n17118 , n1560 );
buf ( n17119 , n17075 );
nand ( n17120 , n17118 , n17119 );
buf ( n17121 , n17120 );
buf ( n17122 , n17121 );
nand ( n17123 , n17117 , n17122 );
buf ( n17124 , n17123 );
buf ( n17125 , n17124 );
xor ( n17126 , n17108 , n17125 );
xor ( n17127 , n810 , n771 );
buf ( n17128 , n17127 );
not ( n17129 , n17128 );
buf ( n17130 , n12889 );
not ( n17131 , n17130 );
or ( n17132 , n17129 , n17131 );
buf ( n17133 , n16594 );
buf ( n17134 , n770 );
buf ( n17135 , n810 );
xor ( n17136 , n17134 , n17135 );
buf ( n17137 , n17136 );
buf ( n17138 , n17137 );
nand ( n17139 , n17133 , n17138 );
buf ( n17140 , n17139 );
buf ( n17141 , n17140 );
nand ( n17142 , n17132 , n17141 );
buf ( n17143 , n17142 );
buf ( n17144 , n17143 );
and ( n17145 , n17126 , n17144 );
and ( n17146 , n17108 , n17125 );
or ( n17147 , n17145 , n17146 );
buf ( n17148 , n17147 );
buf ( n17149 , n17148 );
not ( n17150 , n17149 );
buf ( n17151 , n782 );
buf ( n17152 , n800 );
and ( n17153 , n17151 , n17152 );
buf ( n17154 , n17153 );
buf ( n17155 , n17154 );
buf ( n17156 , n781 );
buf ( n17157 , n800 );
xor ( n17158 , n17156 , n17157 );
buf ( n17159 , n17158 );
buf ( n17160 , n17159 );
not ( n17161 , n17160 );
buf ( n17162 , n10509 );
not ( n17163 , n17162 );
or ( n17164 , n17161 , n17163 );
buf ( n17165 , n3662 );
buf ( n17166 , n16906 );
nand ( n17167 , n17165 , n17166 );
buf ( n17168 , n17167 );
buf ( n17169 , n17168 );
nand ( n17170 , n17164 , n17169 );
buf ( n17171 , n17170 );
buf ( n17172 , n17171 );
xor ( n17173 , n17155 , n17172 );
xor ( n17174 , n806 , n775 );
buf ( n17175 , n17174 );
not ( n17176 , n17175 );
buf ( n17177 , n14278 );
not ( n17178 , n17177 );
or ( n17179 , n17176 , n17178 );
buf ( n17180 , n14284 );
buf ( n17181 , n774 );
buf ( n17182 , n806 );
xor ( n17183 , n17181 , n17182 );
buf ( n17184 , n17183 );
buf ( n17185 , n17184 );
nand ( n17186 , n17180 , n17185 );
buf ( n17187 , n17186 );
buf ( n17188 , n17187 );
nand ( n17189 , n17179 , n17188 );
buf ( n17190 , n17189 );
buf ( n17191 , n17190 );
and ( n17192 , n17173 , n17191 );
and ( n17193 , n17155 , n17172 );
or ( n17194 , n17192 , n17193 );
buf ( n17195 , n17194 );
buf ( n17196 , n17195 );
not ( n17197 , n17196 );
nand ( n17198 , n17150 , n17197 );
not ( n17199 , n17198 );
or ( n17200 , n17091 , n17199 );
nand ( n17201 , n17196 , n17149 );
nand ( n17202 , n17200 , n17201 );
buf ( n17203 , n17202 );
not ( n17204 , n17053 );
not ( n17205 , n17204 );
not ( n17206 , n17088 );
or ( n17207 , n17205 , n17206 );
nand ( n17208 , n17207 , n17070 );
or ( n17209 , n17088 , n17204 );
nand ( n17210 , n17208 , n17209 );
buf ( n17211 , n781 );
buf ( n17212 , n800 );
and ( n17213 , n17211 , n17212 );
buf ( n17214 , n17213 );
buf ( n17215 , n17214 );
buf ( n17216 , n17184 );
not ( n17217 , n17216 );
buf ( n17218 , n1403 );
not ( n17219 , n17218 );
or ( n17220 , n17217 , n17219 );
buf ( n17221 , n14284 );
buf ( n17222 , n773 );
buf ( n17223 , n806 );
xor ( n17224 , n17222 , n17223 );
buf ( n17225 , n17224 );
buf ( n17226 , n17225 );
nand ( n17227 , n17221 , n17226 );
buf ( n17228 , n17227 );
buf ( n17229 , n17228 );
nand ( n17230 , n17220 , n17229 );
buf ( n17231 , n17230 );
buf ( n17232 , n17231 );
xor ( n17233 , n17215 , n17232 );
buf ( n17234 , n17137 );
not ( n17235 , n17234 );
buf ( n17236 , n12889 );
not ( n17237 , n17236 );
or ( n17238 , n17235 , n17237 );
buf ( n17239 , n16594 );
buf ( n17240 , n769 );
buf ( n17241 , n810 );
xor ( n17242 , n17240 , n17241 );
buf ( n17243 , n17242 );
buf ( n17244 , n17243 );
nand ( n17245 , n17239 , n17244 );
buf ( n17246 , n17245 );
buf ( n17247 , n17246 );
nand ( n17248 , n17238 , n17247 );
buf ( n17249 , n17248 );
buf ( n17250 , n17249 );
and ( n17251 , n17233 , n17250 );
and ( n17252 , n17215 , n17232 );
or ( n17253 , n17251 , n17252 );
buf ( n17254 , n17253 );
buf ( n17255 , n17254 );
xor ( n17256 , n17210 , n17255 );
not ( n17257 , n1713 );
not ( n17258 , n14588 );
or ( n17259 , n17257 , n17258 );
nand ( n17260 , n17259 , n812 );
buf ( n17261 , n17260 );
buf ( n17262 , n17243 );
not ( n17263 , n17262 );
buf ( n17264 , n12889 );
not ( n17265 , n17264 );
or ( n17266 , n17263 , n17265 );
buf ( n17267 , n16594 );
buf ( n17268 , n768 );
buf ( n17269 , n810 );
xor ( n17270 , n17268 , n17269 );
buf ( n17271 , n17270 );
buf ( n17272 , n17271 );
nand ( n17273 , n17267 , n17272 );
buf ( n17274 , n17273 );
buf ( n17275 , n17274 );
nand ( n17276 , n17266 , n17275 );
buf ( n17277 , n17276 );
buf ( n17278 , n17277 );
xor ( n17279 , n17261 , n17278 );
buf ( n17280 , n17225 );
not ( n17281 , n17280 );
buf ( n17282 , n14278 );
not ( n17283 , n17282 );
or ( n17284 , n17281 , n17283 );
buf ( n17285 , n14284 );
xor ( n17286 , n806 , n772 );
buf ( n17287 , n17286 );
nand ( n17288 , n17285 , n17287 );
buf ( n17289 , n17288 );
buf ( n17290 , n17289 );
nand ( n17291 , n17284 , n17290 );
buf ( n17292 , n17291 );
buf ( n17293 , n17292 );
xor ( n17294 , n17279 , n17293 );
buf ( n17295 , n17294 );
xor ( n17296 , n17256 , n17295 );
buf ( n17297 , n17296 );
xor ( n17298 , n17203 , n17297 );
xor ( n17299 , n17215 , n17232 );
xor ( n17300 , n17299 , n17250 );
buf ( n17301 , n17300 );
buf ( n17302 , n17301 );
xor ( n17303 , n16904 , n16923 );
xor ( n17304 , n17303 , n16989 );
buf ( n17305 , n17304 );
buf ( n17306 , n17305 );
xor ( n17307 , n17302 , n17306 );
buf ( n17308 , n16571 );
not ( n17309 , n17308 );
buf ( n17310 , n15790 );
not ( n17311 , n17310 );
or ( n17312 , n17309 , n17311 );
buf ( n17313 , n16931 );
not ( n17314 , n17313 );
buf ( n17315 , n814 );
nand ( n17316 , n17314 , n17315 );
buf ( n17317 , n17316 );
buf ( n17318 , n17317 );
nand ( n17319 , n17312 , n17318 );
buf ( n17320 , n17319 );
buf ( n17321 , n17320 );
buf ( n17322 , n16471 );
not ( n17323 , n17322 );
buf ( n17324 , n14278 );
not ( n17325 , n17324 );
or ( n17326 , n17323 , n17325 );
buf ( n17327 , n14284 );
buf ( n17328 , n17174 );
nand ( n17329 , n17327 , n17328 );
buf ( n17330 , n17329 );
buf ( n17331 , n17330 );
nand ( n17332 , n17326 , n17331 );
buf ( n17333 , n17332 );
buf ( n17334 , n17333 );
not ( n17335 , n17334 );
not ( n17336 , n16594 );
not ( n17337 , n17127 );
or ( n17338 , n17336 , n17337 );
nand ( n17339 , n16599 , n12889 );
nand ( n17340 , n17338 , n17339 );
buf ( n17341 , n17340 );
not ( n17342 , n17341 );
or ( n17343 , n17335 , n17342 );
buf ( n17344 , n17340 );
buf ( n17345 , n17333 );
or ( n17346 , n17344 , n17345 );
buf ( n17347 , n16490 );
not ( n17348 , n17347 );
buf ( n17349 , n2916 );
not ( n17350 , n17349 );
or ( n17351 , n17348 , n17350 );
buf ( n17352 , n14589 );
buf ( n17353 , n16961 );
nand ( n17354 , n17352 , n17353 );
buf ( n17355 , n17354 );
buf ( n17356 , n17355 );
nand ( n17357 , n17351 , n17356 );
buf ( n17358 , n17357 );
buf ( n17359 , n17358 );
nand ( n17360 , n17346 , n17359 );
buf ( n17361 , n17360 );
buf ( n17362 , n17361 );
nand ( n17363 , n17343 , n17362 );
buf ( n17364 , n17363 );
buf ( n17365 , n17364 );
xor ( n17366 , n17321 , n17365 );
buf ( n17367 , n783 );
buf ( n17368 , n800 );
and ( n17369 , n17367 , n17368 );
buf ( n17370 , n17369 );
buf ( n17371 , n17370 );
buf ( n17372 , n16516 );
not ( n17373 , n17372 );
buf ( n17374 , n2709 );
not ( n17375 , n17374 );
or ( n17376 , n17373 , n17375 );
buf ( n17377 , n2713 );
buf ( n17378 , n16946 );
nand ( n17379 , n17377 , n17378 );
buf ( n17380 , n17379 );
buf ( n17381 , n17380 );
nand ( n17382 , n17376 , n17381 );
buf ( n17383 , n17382 );
buf ( n17384 , n17383 );
xor ( n17385 , n17371 , n17384 );
buf ( n17386 , n16551 );
not ( n17387 , n17386 );
buf ( n17388 , n10509 );
not ( n17389 , n17388 );
or ( n17390 , n17387 , n17389 );
buf ( n17391 , n3662 );
buf ( n17392 , n17159 );
nand ( n17393 , n17391 , n17392 );
buf ( n17394 , n17393 );
buf ( n17395 , n17394 );
nand ( n17396 , n17390 , n17395 );
buf ( n17397 , n17396 );
buf ( n17398 , n17397 );
and ( n17399 , n17385 , n17398 );
and ( n17400 , n17371 , n17384 );
or ( n17401 , n17399 , n17400 );
buf ( n17402 , n17401 );
buf ( n17403 , n17402 );
and ( n17404 , n17366 , n17403 );
and ( n17405 , n17321 , n17365 );
or ( n17406 , n17404 , n17405 );
buf ( n17407 , n17406 );
buf ( n17408 , n17407 );
and ( n17409 , n17307 , n17408 );
and ( n17410 , n17302 , n17306 );
or ( n17411 , n17409 , n17410 );
buf ( n17412 , n17411 );
buf ( n17413 , n17412 );
xor ( n17414 , n17298 , n17413 );
buf ( n17415 , n17414 );
buf ( n17416 , n17415 );
xor ( n17417 , n17041 , n17416 );
xor ( n17418 , n17155 , n17172 );
xor ( n17419 , n17418 , n17191 );
buf ( n17420 , n17419 );
buf ( n17421 , n17420 );
xor ( n17422 , n17108 , n17125 );
xor ( n17423 , n17422 , n17144 );
buf ( n17424 , n17423 );
buf ( n17425 , n17424 );
xor ( n17426 , n17421 , n17425 );
xor ( n17427 , n16939 , n16973 );
buf ( n17428 , n17427 );
buf ( n17429 , n16954 );
and ( n17430 , n17428 , n17429 );
not ( n17431 , n17428 );
buf ( n17432 , n16982 );
and ( n17433 , n17431 , n17432 );
nor ( n17434 , n17430 , n17433 );
buf ( n17435 , n17434 );
buf ( n17436 , n17435 );
and ( n17437 , n17426 , n17436 );
and ( n17438 , n17421 , n17425 );
or ( n17439 , n17437 , n17438 );
buf ( n17440 , n17439 );
buf ( n17441 , n17440 );
and ( n17442 , n17149 , n17197 , n17089 );
not ( n17443 , n17442 );
nand ( n17444 , n17196 , n17149 , n17090 );
nand ( n17445 , n17197 , n17150 , n17090 );
not ( n17446 , n17149 );
nand ( n17447 , n17446 , n17196 , n17089 );
nand ( n17448 , n17443 , n17444 , n17445 , n17447 );
buf ( n17449 , n17448 );
xor ( n17450 , n17441 , n17449 );
xor ( n17451 , n17302 , n17306 );
xor ( n17452 , n17451 , n17408 );
buf ( n17453 , n17452 );
buf ( n17454 , n17453 );
and ( n17455 , n17450 , n17454 );
and ( n17456 , n17441 , n17449 );
or ( n17457 , n17455 , n17456 );
buf ( n17458 , n17457 );
buf ( n17459 , n17458 );
xor ( n17460 , n17417 , n17459 );
buf ( n17461 , n17460 );
buf ( n17462 , n17461 );
buf ( n17463 , n16621 );
not ( n17464 , n17463 );
buf ( n17465 , n15873 );
not ( n17466 , n17465 );
or ( n17467 , n17464 , n17466 );
buf ( n17468 , n11137 );
buf ( n17469 , n17095 );
nand ( n17470 , n17468 , n17469 );
buf ( n17471 , n17470 );
buf ( n17472 , n17471 );
nand ( n17473 , n17467 , n17472 );
buf ( n17474 , n17473 );
buf ( n17475 , n17474 );
buf ( n17476 , n16533 );
not ( n17477 , n17476 );
buf ( n17478 , n3109 );
not ( n17479 , n17478 );
or ( n17480 , n17477 , n17479 );
buf ( n17481 , n1560 );
buf ( n17482 , n17112 );
nand ( n17483 , n17481 , n17482 );
buf ( n17484 , n17483 );
buf ( n17485 , n17484 );
nand ( n17486 , n17480 , n17485 );
buf ( n17487 , n17486 );
buf ( n17488 , n17487 );
xor ( n17489 , n17475 , n17488 );
buf ( n17490 , n17320 );
not ( n17491 , n17490 );
buf ( n17492 , n17491 );
buf ( n17493 , n17492 );
and ( n17494 , n17489 , n17493 );
and ( n17495 , n17475 , n17488 );
or ( n17496 , n17494 , n17495 );
buf ( n17497 , n17496 );
buf ( n17498 , n17497 );
xor ( n17499 , n17321 , n17365 );
xor ( n17500 , n17499 , n17403 );
buf ( n17501 , n17500 );
buf ( n17502 , n17501 );
xor ( n17503 , n17498 , n17502 );
xor ( n17504 , n16461 , n16478 );
and ( n17505 , n17504 , n16497 );
and ( n17506 , n16461 , n16478 );
or ( n17507 , n17505 , n17506 );
buf ( n17508 , n17507 );
buf ( n17509 , n17508 );
xor ( n17510 , n16523 , n16540 );
and ( n17511 , n17510 , n16558 );
and ( n17512 , n16523 , n16540 );
or ( n17513 , n17511 , n17512 );
buf ( n17514 , n17513 );
buf ( n17515 , n17514 );
xor ( n17516 , n17509 , n17515 );
xor ( n17517 , n16578 , n16585 );
and ( n17518 , n17517 , n16606 );
and ( n17519 , n16578 , n16585 );
or ( n17520 , n17518 , n17519 );
buf ( n17521 , n17520 );
buf ( n17522 , n17521 );
and ( n17523 , n17516 , n17522 );
and ( n17524 , n17509 , n17515 );
or ( n17525 , n17523 , n17524 );
buf ( n17526 , n17525 );
buf ( n17527 , n17526 );
and ( n17528 , n17503 , n17527 );
and ( n17529 , n17498 , n17502 );
or ( n17530 , n17528 , n17529 );
buf ( n17531 , n17530 );
buf ( n17532 , n17531 );
xor ( n17533 , n17441 , n17449 );
xor ( n17534 , n17533 , n17454 );
buf ( n17535 , n17534 );
buf ( n17536 , n17535 );
xor ( n17537 , n17532 , n17536 );
xor ( n17538 , n17371 , n17384 );
xor ( n17539 , n17538 , n17398 );
buf ( n17540 , n17539 );
buf ( n17541 , n17540 );
xor ( n17542 , n17340 , n17333 );
xor ( n17543 , n17542 , n17358 );
buf ( n17544 , n17543 );
xor ( n17545 , n17541 , n17544 );
xor ( n17546 , n17475 , n17488 );
xor ( n17547 , n17546 , n17493 );
buf ( n17548 , n17547 );
buf ( n17549 , n17548 );
and ( n17550 , n17545 , n17549 );
and ( n17551 , n17541 , n17544 );
or ( n17552 , n17550 , n17551 );
buf ( n17553 , n17552 );
buf ( n17554 , n17553 );
xor ( n17555 , n17421 , n17425 );
xor ( n17556 , n17555 , n17436 );
buf ( n17557 , n17556 );
buf ( n17558 , n17557 );
xor ( n17559 , n17554 , n17558 );
xor ( n17560 , n16611 , n16628 );
and ( n17561 , n17560 , n16635 );
and ( n17562 , n16611 , n16628 );
or ( n17563 , n17561 , n17562 );
buf ( n17564 , n17563 );
buf ( n17565 , n17564 );
xor ( n17566 , n16449 , n16455 );
and ( n17567 , n17566 , n16500 );
and ( n17568 , n16449 , n16455 );
or ( n17569 , n17567 , n17568 );
buf ( n17570 , n17569 );
buf ( n17571 , n17570 );
xor ( n17572 , n17565 , n17571 );
xor ( n17573 , n17509 , n17515 );
xor ( n17574 , n17573 , n17522 );
buf ( n17575 , n17574 );
buf ( n17576 , n17575 );
and ( n17577 , n17572 , n17576 );
and ( n17578 , n17565 , n17571 );
or ( n17579 , n17577 , n17578 );
buf ( n17580 , n17579 );
buf ( n17581 , n17580 );
and ( n17582 , n17559 , n17581 );
and ( n17583 , n17554 , n17558 );
or ( n17584 , n17582 , n17583 );
buf ( n17585 , n17584 );
buf ( n17586 , n17585 );
and ( n17587 , n17537 , n17586 );
and ( n17588 , n17532 , n17536 );
or ( n17589 , n17587 , n17588 );
buf ( n17590 , n17589 );
buf ( n17591 , n17590 );
xor ( n17592 , n17462 , n17591 );
buf ( n17593 , n17592 );
buf ( n17594 , n17593 );
not ( n17595 , n17594 );
buf ( n17596 , n17595 );
buf ( n17597 , n17596 );
xor ( n17598 , n17532 , n17536 );
xor ( n17599 , n17598 , n17586 );
buf ( n17600 , n17599 );
buf ( n17601 , n17600 );
xor ( n17602 , n17498 , n17502 );
xor ( n17603 , n17602 , n17527 );
buf ( n17604 , n17603 );
buf ( n17605 , n17604 );
xor ( n17606 , n16561 , n16609 );
and ( n17607 , n17606 , n16638 );
and ( n17608 , n16561 , n16609 );
or ( n17609 , n17607 , n17608 );
buf ( n17610 , n17609 );
buf ( n17611 , n17610 );
xor ( n17612 , n17541 , n17544 );
xor ( n17613 , n17612 , n17549 );
buf ( n17614 , n17613 );
buf ( n17615 , n17614 );
xor ( n17616 , n17611 , n17615 );
xor ( n17617 , n16436 , n16442 );
and ( n17618 , n17617 , n16503 );
and ( n17619 , n16436 , n16442 );
or ( n17620 , n17618 , n17619 );
buf ( n17621 , n17620 );
buf ( n17622 , n17621 );
and ( n17623 , n17616 , n17622 );
and ( n17624 , n17611 , n17615 );
or ( n17625 , n17623 , n17624 );
buf ( n17626 , n17625 );
buf ( n17627 , n17626 );
xor ( n17628 , n17605 , n17627 );
xor ( n17629 , n17554 , n17558 );
xor ( n17630 , n17629 , n17581 );
buf ( n17631 , n17630 );
buf ( n17632 , n17631 );
and ( n17633 , n17628 , n17632 );
and ( n17634 , n17605 , n17627 );
or ( n17635 , n17633 , n17634 );
buf ( n17636 , n17635 );
buf ( n17637 , n17636 );
and ( n17638 , n17601 , n17637 );
buf ( n17639 , n17638 );
buf ( n17640 , n17639 );
not ( n17641 , n17640 );
buf ( n17642 , n17641 );
buf ( n17643 , n17642 );
nand ( n17644 , n17597 , n17643 );
buf ( n17645 , n17644 );
buf ( n17646 , n17645 );
xor ( n17647 , n17605 , n17627 );
xor ( n17648 , n17647 , n17632 );
buf ( n17649 , n17648 );
buf ( n17650 , n17649 );
xor ( n17651 , n17565 , n17571 );
xor ( n17652 , n17651 , n17576 );
buf ( n17653 , n17652 );
buf ( n17654 , n17653 );
xor ( n17655 , n17611 , n17615 );
xor ( n17656 , n17655 , n17622 );
buf ( n17657 , n17656 );
buf ( n17658 , n17657 );
xor ( n17659 , n17654 , n17658 );
xor ( n17660 , n16641 , n16647 );
and ( n17661 , n17660 , n16666 );
and ( n17662 , n16641 , n16647 );
or ( n17663 , n17661 , n17662 );
buf ( n17664 , n17663 );
buf ( n17665 , n17664 );
and ( n17666 , n17659 , n17665 );
and ( n17667 , n17654 , n17658 );
or ( n17668 , n17666 , n17667 );
buf ( n17669 , n17668 );
buf ( n17670 , n17669 );
and ( n17671 , n17650 , n17670 );
buf ( n17672 , n17671 );
buf ( n17673 , n17672 );
not ( n17674 , n17673 );
xor ( n17675 , n17601 , n17637 );
buf ( n17676 , n17675 );
buf ( n17677 , n17676 );
not ( n17678 , n17677 );
buf ( n17679 , n17678 );
buf ( n17680 , n17679 );
nand ( n17681 , n17674 , n17680 );
buf ( n17682 , n17681 );
buf ( n17683 , n17682 );
and ( n17684 , n17646 , n17683 );
buf ( n17685 , n17684 );
buf ( n17686 , n17685 );
xor ( n17687 , n16506 , n16669 );
and ( n17688 , n17687 , n16676 );
and ( n17689 , n16506 , n16669 );
or ( n17690 , n17688 , n17689 );
buf ( n17691 , n17690 );
xor ( n17692 , n17654 , n17658 );
xor ( n17693 , n17692 , n17665 );
buf ( n17694 , n17693 );
xor ( n17695 , n17691 , n17694 );
buf ( n17696 , n17695 );
and ( n17697 , n16679 , n16685 );
buf ( n17698 , n17697 );
buf ( n17699 , n17698 );
nor ( n17700 , n17696 , n17699 );
buf ( n17701 , n17700 );
buf ( n17702 , n17701 );
buf ( n17703 , n17694 );
buf ( n17704 , n17691 );
and ( n17705 , n17703 , n17704 );
buf ( n17706 , n17705 );
buf ( n17707 , n17706 );
buf ( n17708 , n17669 );
not ( n17709 , n17708 );
buf ( n17710 , n17649 );
not ( n17711 , n17710 );
buf ( n17712 , n17711 );
buf ( n17713 , n17712 );
not ( n17714 , n17713 );
or ( n17715 , n17709 , n17714 );
buf ( n17716 , n17669 );
not ( n17717 , n17716 );
buf ( n17718 , n17649 );
nand ( n17719 , n17717 , n17718 );
buf ( n17720 , n17719 );
buf ( n17721 , n17720 );
nand ( n17722 , n17715 , n17721 );
buf ( n17723 , n17722 );
buf ( n17724 , n17723 );
nor ( n17725 , n17707 , n17724 );
buf ( n17726 , n17725 );
buf ( n17727 , n17726 );
nor ( n17728 , n17702 , n17727 );
buf ( n17729 , n17728 );
buf ( n17730 , n17729 );
nand ( n17731 , n17686 , n17730 );
buf ( n17732 , n17731 );
buf ( n17733 , n17732 );
buf ( n17734 , n17733 );
buf ( n17735 , n17734 );
buf ( n17736 , n17735 );
not ( n17737 , n17736 );
buf ( n17738 , n17737 );
buf ( n17739 , n17738 );
and ( n17740 , n17462 , n17591 );
buf ( n17741 , n17740 );
buf ( n17742 , n17741 );
not ( n17743 , n17742 );
xor ( n17744 , n17041 , n17416 );
and ( n17745 , n17744 , n17459 );
and ( n17746 , n17041 , n17416 );
or ( n17747 , n17745 , n17746 );
buf ( n17748 , n17747 );
buf ( n17749 , n17748 );
xor ( n17750 , n16884 , n16994 );
and ( n17751 , n17750 , n17038 );
and ( n17752 , n16884 , n16994 );
or ( n17753 , n17751 , n17752 );
buf ( n17754 , n17753 );
buf ( n17755 , n17754 );
xor ( n17756 , n17203 , n17297 );
and ( n17757 , n17756 , n17413 );
and ( n17758 , n17203 , n17297 );
or ( n17759 , n17757 , n17758 );
buf ( n17760 , n17759 );
buf ( n17761 , n17760 );
xor ( n17762 , n17755 , n17761 );
buf ( n17763 , n17271 );
not ( n17764 , n17763 );
buf ( n17765 , n11050 );
not ( n17766 , n17765 );
or ( n17767 , n17764 , n17766 );
buf ( n17768 , n16594 );
buf ( n17769 , n810 );
nand ( n17770 , n17768 , n17769 );
buf ( n17771 , n17770 );
buf ( n17772 , n17771 );
nand ( n17773 , n17767 , n17772 );
buf ( n17774 , n17773 );
buf ( n17775 , n17774 );
not ( n17776 , n17775 );
buf ( n17777 , n17776 );
buf ( n17778 , n17777 );
buf ( n17779 , n16880 );
buf ( n17780 , n16859 );
or ( n17781 , n17779 , n17780 );
buf ( n17782 , n16854 );
nand ( n17783 , n17781 , n17782 );
buf ( n17784 , n17783 );
buf ( n17785 , n17784 );
buf ( n17786 , n16859 );
buf ( n17787 , n16880 );
nand ( n17788 , n17786 , n17787 );
buf ( n17789 , n17788 );
buf ( n17790 , n17789 );
nand ( n17791 , n17785 , n17790 );
buf ( n17792 , n17791 );
buf ( n17793 , n17792 );
xor ( n17794 , n17778 , n17793 );
xor ( n17795 , n17261 , n17278 );
and ( n17796 , n17795 , n17293 );
and ( n17797 , n17261 , n17278 );
or ( n17798 , n17796 , n17797 );
buf ( n17799 , n17798 );
buf ( n17800 , n17799 );
xor ( n17801 , n17794 , n17800 );
buf ( n17802 , n17801 );
buf ( n17803 , n17802 );
not ( n17804 , n17295 );
or ( n17805 , n17210 , n17255 );
not ( n17806 , n17805 );
or ( n17807 , n17804 , n17806 );
nand ( n17808 , n17255 , n17210 );
nand ( n17809 , n17807 , n17808 );
buf ( n17810 , n17809 );
xor ( n17811 , n17803 , n17810 );
buf ( n17812 , n17012 );
buf ( n17813 , n17028 );
or ( n17814 , n17812 , n17813 );
buf ( n17815 , n16900 );
nand ( n17816 , n17814 , n17815 );
buf ( n17817 , n17816 );
buf ( n17818 , n17817 );
buf ( n17819 , n17028 );
buf ( n17820 , n17012 );
nand ( n17821 , n17819 , n17820 );
buf ( n17822 , n17821 );
buf ( n17823 , n17822 );
nand ( n17824 , n17818 , n17823 );
buf ( n17825 , n17824 );
buf ( n17826 , n17825 );
buf ( n17827 , n16848 );
not ( n17828 , n17827 );
buf ( n17829 , n15873 );
not ( n17830 , n17829 );
or ( n17831 , n17828 , n17830 );
buf ( n17832 , n11137 );
buf ( n17833 , n773 );
buf ( n17834 , n804 );
xor ( n17835 , n17833 , n17834 );
buf ( n17836 , n17835 );
buf ( n17837 , n17836 );
nand ( n17838 , n17832 , n17837 );
buf ( n17839 , n17838 );
buf ( n17840 , n17839 );
nand ( n17841 , n17831 , n17840 );
buf ( n17842 , n17841 );
buf ( n17843 , n17842 );
buf ( n17844 , n17006 );
not ( n17845 , n17844 );
buf ( n17846 , n3109 );
not ( n17847 , n17846 );
or ( n17848 , n17845 , n17847 );
buf ( n17849 , n1560 );
xor ( n17850 , n802 , n775 );
buf ( n17851 , n17850 );
nand ( n17852 , n17849 , n17851 );
buf ( n17853 , n17852 );
buf ( n17854 , n17853 );
nand ( n17855 , n17848 , n17854 );
buf ( n17856 , n17855 );
buf ( n17857 , n17856 );
xor ( n17858 , n17843 , n17857 );
buf ( n17859 , n16874 );
not ( n17860 , n17859 );
buf ( n17861 , n2709 );
not ( n17862 , n17861 );
or ( n17863 , n17860 , n17862 );
buf ( n17864 , n2713 );
buf ( n17865 , n769 );
buf ( n17866 , n808 );
xor ( n17867 , n17865 , n17866 );
buf ( n17868 , n17867 );
buf ( n17869 , n17868 );
nand ( n17870 , n17864 , n17869 );
buf ( n17871 , n17870 );
buf ( n17872 , n17871 );
nand ( n17873 , n17863 , n17872 );
buf ( n17874 , n17873 );
buf ( n17875 , n17874 );
xor ( n17876 , n17858 , n17875 );
buf ( n17877 , n17876 );
buf ( n17878 , n17877 );
xor ( n17879 , n17826 , n17878 );
and ( n17880 , n16913 , n16914 );
buf ( n17881 , n17880 );
buf ( n17882 , n17286 );
not ( n17883 , n17882 );
buf ( n17884 , n14278 );
not ( n17885 , n17884 );
or ( n17886 , n17883 , n17885 );
buf ( n17887 , n14284 );
xor ( n17888 , n806 , n771 );
buf ( n17889 , n17888 );
nand ( n17890 , n17887 , n17889 );
buf ( n17891 , n17890 );
buf ( n17892 , n17891 );
nand ( n17893 , n17886 , n17892 );
buf ( n17894 , n17893 );
xor ( n17895 , n17881 , n17894 );
buf ( n17896 , n17022 );
not ( n17897 , n17896 );
buf ( n17898 , n10509 );
not ( n17899 , n17898 );
or ( n17900 , n17897 , n17899 );
buf ( n17901 , n3662 );
buf ( n17902 , n800 );
buf ( n17903 , n777 );
xor ( n17904 , n17902 , n17903 );
buf ( n17905 , n17904 );
buf ( n17906 , n17905 );
nand ( n17907 , n17901 , n17906 );
buf ( n17908 , n17907 );
buf ( n17909 , n17908 );
nand ( n17910 , n17900 , n17909 );
buf ( n17911 , n17910 );
xor ( n17912 , n17895 , n17911 );
buf ( n17913 , n17912 );
xor ( n17914 , n17879 , n17913 );
buf ( n17915 , n17914 );
buf ( n17916 , n17915 );
xor ( n17917 , n17811 , n17916 );
buf ( n17918 , n17917 );
buf ( n17919 , n17918 );
xor ( n17920 , n17762 , n17919 );
buf ( n17921 , n17920 );
buf ( n17922 , n17921 );
xor ( n17923 , n17749 , n17922 );
buf ( n17924 , n17923 );
buf ( n17925 , n17924 );
not ( n17926 , n17925 );
buf ( n17927 , n17926 );
buf ( n17928 , n17927 );
nand ( n17929 , n17743 , n17928 );
buf ( n17930 , n17929 );
buf ( n17931 , n17930 );
and ( n17932 , n17749 , n17922 );
buf ( n17933 , n17932 );
nand ( n17934 , n17881 , n17894 );
nand ( n17935 , n17881 , n17911 );
nand ( n17936 , n17894 , n17911 );
nand ( n17937 , n17934 , n17935 , n17936 );
buf ( n17938 , n17937 );
buf ( n17939 , n17868 );
not ( n17940 , n17939 );
buf ( n17941 , n2709 );
not ( n17942 , n17941 );
or ( n17943 , n17940 , n17942 );
buf ( n17944 , n2713 );
buf ( n17945 , n768 );
buf ( n17946 , n808 );
xor ( n17947 , n17945 , n17946 );
buf ( n17948 , n17947 );
buf ( n17949 , n17948 );
nand ( n17950 , n17944 , n17949 );
buf ( n17951 , n17950 );
buf ( n17952 , n17951 );
nand ( n17953 , n17943 , n17952 );
buf ( n17954 , n17953 );
buf ( n17955 , n17954 );
buf ( n17956 , n16009 );
not ( n17957 , n17956 );
buf ( n17958 , n16000 );
not ( n17959 , n17958 );
or ( n17960 , n17957 , n17959 );
buf ( n17961 , n810 );
nand ( n17962 , n17960 , n17961 );
buf ( n17963 , n17962 );
buf ( n17964 , n17963 );
xor ( n17965 , n17955 , n17964 );
buf ( n17966 , n17836 );
not ( n17967 , n17966 );
buf ( n17968 , n15873 );
not ( n17969 , n17968 );
or ( n17970 , n17967 , n17969 );
buf ( n17971 , n11137 );
buf ( n17972 , n772 );
buf ( n17973 , n804 );
xor ( n17974 , n17972 , n17973 );
buf ( n17975 , n17974 );
buf ( n17976 , n17975 );
nand ( n17977 , n17971 , n17976 );
buf ( n17978 , n17977 );
buf ( n17979 , n17978 );
nand ( n17980 , n17970 , n17979 );
buf ( n17981 , n17980 );
buf ( n17982 , n17981 );
xor ( n17983 , n17965 , n17982 );
buf ( n17984 , n17983 );
buf ( n17985 , n17984 );
xor ( n17986 , n17938 , n17985 );
buf ( n17987 , n17905 );
not ( n17988 , n17987 );
buf ( n17989 , n10509 );
not ( n17990 , n17989 );
or ( n17991 , n17988 , n17990 );
buf ( n17992 , n3662 );
buf ( n17993 , n800 );
buf ( n17994 , n776 );
xor ( n17995 , n17993 , n17994 );
buf ( n17996 , n17995 );
buf ( n17997 , n17996 );
nand ( n17998 , n17992 , n17997 );
buf ( n17999 , n17998 );
buf ( n18000 , n17999 );
nand ( n18001 , n17991 , n18000 );
buf ( n18002 , n18001 );
buf ( n18003 , n18002 );
buf ( n18004 , n17850 );
not ( n18005 , n18004 );
buf ( n18006 , n3109 );
not ( n18007 , n18006 );
or ( n18008 , n18005 , n18007 );
buf ( n18009 , n1560 );
buf ( n18010 , n802 );
buf ( n18011 , n774 );
xor ( n18012 , n18010 , n18011 );
buf ( n18013 , n18012 );
buf ( n18014 , n18013 );
nand ( n18015 , n18009 , n18014 );
buf ( n18016 , n18015 );
buf ( n18017 , n18016 );
nand ( n18018 , n18008 , n18017 );
buf ( n18019 , n18018 );
buf ( n18020 , n18019 );
xor ( n18021 , n18003 , n18020 );
buf ( n18022 , n17888 );
not ( n18023 , n18022 );
buf ( n18024 , n14278 );
not ( n18025 , n18024 );
or ( n18026 , n18023 , n18025 );
buf ( n18027 , n14284 );
buf ( n18028 , n770 );
buf ( n18029 , n806 );
xor ( n18030 , n18028 , n18029 );
buf ( n18031 , n18030 );
buf ( n18032 , n18031 );
nand ( n18033 , n18027 , n18032 );
buf ( n18034 , n18033 );
buf ( n18035 , n18034 );
nand ( n18036 , n18026 , n18035 );
buf ( n18037 , n18036 );
buf ( n18038 , n18037 );
xor ( n18039 , n18021 , n18038 );
buf ( n18040 , n18039 );
buf ( n18041 , n18040 );
xor ( n18042 , n17986 , n18041 );
buf ( n18043 , n18042 );
buf ( n18044 , n18043 );
and ( n18045 , n17019 , n17020 );
buf ( n18046 , n18045 );
buf ( n18047 , n18046 );
buf ( n18048 , n17774 );
xor ( n18049 , n18047 , n18048 );
xor ( n18050 , n17843 , n17857 );
and ( n18051 , n18050 , n17875 );
and ( n18052 , n17843 , n17857 );
or ( n18053 , n18051 , n18052 );
buf ( n18054 , n18053 );
buf ( n18055 , n18054 );
xor ( n18056 , n18049 , n18055 );
buf ( n18057 , n18056 );
buf ( n18058 , n18057 );
xor ( n18059 , n17778 , n17793 );
and ( n18060 , n18059 , n17800 );
and ( n18061 , n17778 , n17793 );
or ( n18062 , n18060 , n18061 );
buf ( n18063 , n18062 );
buf ( n18064 , n18063 );
xor ( n18065 , n18058 , n18064 );
xor ( n18066 , n17826 , n17878 );
and ( n18067 , n18066 , n17913 );
and ( n18068 , n17826 , n17878 );
or ( n18069 , n18067 , n18068 );
buf ( n18070 , n18069 );
buf ( n18071 , n18070 );
xor ( n18072 , n18065 , n18071 );
buf ( n18073 , n18072 );
buf ( n18074 , n18073 );
xor ( n18075 , n18044 , n18074 );
xor ( n18076 , n17803 , n17810 );
and ( n18077 , n18076 , n17916 );
and ( n18078 , n17803 , n17810 );
or ( n18079 , n18077 , n18078 );
buf ( n18080 , n18079 );
buf ( n18081 , n18080 );
xor ( n18082 , n18075 , n18081 );
buf ( n18083 , n18082 );
buf ( n18084 , n18083 );
xor ( n18085 , n17755 , n17761 );
and ( n18086 , n18085 , n17919 );
and ( n18087 , n17755 , n17761 );
or ( n18088 , n18086 , n18087 );
buf ( n18089 , n18088 );
buf ( n18090 , n18089 );
xor ( n18091 , n18084 , n18090 );
buf ( n18092 , n18091 );
or ( n18093 , n17933 , n18092 );
buf ( n18094 , n18093 );
and ( n18095 , n17931 , n18094 );
buf ( n18096 , n18095 );
buf ( n18097 , n18096 );
nand ( n18098 , n17739 , n18097 );
buf ( n18099 , n18098 );
buf ( n18100 , n18099 );
not ( n18101 , n18100 );
buf ( n18102 , n18101 );
buf ( n18103 , n18102 );
nand ( n18104 , n16834 , n18103 );
buf ( n18105 , n18104 );
buf ( n18106 , n10417 );
nand ( n18107 , n14550 , n15322 );
buf ( n18108 , n18107 );
not ( n18109 , n18108 );
buf ( n18110 , n13733 );
buf ( n18111 , n13677 );
and ( n18112 , n18110 , n18111 );
buf ( n18113 , n18112 );
buf ( n18114 , n18113 );
buf ( n18115 , n16781 );
buf ( n18116 , n15945 );
buf ( n18117 , n16271 );
buf ( n18118 , n18117 );
buf ( n18119 , n18118 );
buf ( n18120 , n18119 );
and ( n18121 , n18115 , n18116 , n18120 );
buf ( n18122 , n18121 );
buf ( n18123 , n18122 );
buf ( n18124 , n13759 );
buf ( n18125 , n12808 );
nor ( n18126 , n18124 , n18125 );
buf ( n18127 , n18126 );
buf ( n18128 , n18127 );
nand ( n18129 , n18109 , n18114 , n18123 , n18128 );
buf ( n18130 , n18129 );
buf ( n18131 , n18130 );
not ( n18132 , n18131 );
buf ( n18133 , n18132 );
buf ( n18134 , n18133 );
not ( n18135 , n18134 );
buf ( n18136 , n18135 );
buf ( n18137 , n18136 );
buf ( n18138 , n18099 );
nor ( n18139 , n18137 , n18138 );
buf ( n18140 , n18139 );
buf ( n18141 , n18140 );
nand ( n18142 , n18106 , n18141 );
buf ( n18143 , n18142 );
buf ( n18144 , n18096 );
not ( n18145 , n18144 );
buf ( n18146 , n17685 );
not ( n18147 , n18146 );
buf ( n18148 , n17695 );
buf ( n18149 , n17698 );
nand ( n18150 , n18148 , n18149 );
buf ( n18151 , n18150 );
not ( n18152 , n18151 );
not ( n18153 , n18152 );
not ( n18154 , n17726 );
not ( n18155 , n18154 );
or ( n18156 , n18153 , n18155 );
nand ( n18157 , n17706 , n17723 );
nand ( n18158 , n18156 , n18157 );
buf ( n18159 , n18158 );
not ( n18160 , n18159 );
or ( n18161 , n18147 , n18160 );
buf ( n18162 , n17645 );
buf ( n18163 , n17672 );
buf ( n18164 , n17676 );
nand ( n18165 , n18163 , n18164 );
buf ( n18166 , n18165 );
buf ( n18167 , n18166 );
not ( n18168 , n18167 );
buf ( n18169 , n18168 );
buf ( n18170 , n18169 );
and ( n18171 , n18162 , n18170 );
buf ( n18172 , n17596 );
buf ( n18173 , n17642 );
nor ( n18174 , n18172 , n18173 );
buf ( n18175 , n18174 );
buf ( n18176 , n18175 );
nor ( n18177 , n18171 , n18176 );
buf ( n18178 , n18177 );
buf ( n18179 , n18178 );
nand ( n18180 , n18161 , n18179 );
buf ( n18181 , n18180 );
buf ( n18182 , n18181 );
buf ( n18183 , n18182 );
buf ( n18184 , n18183 );
buf ( n18185 , n18184 );
not ( n18186 , n18185 );
or ( n18187 , n18145 , n18186 );
buf ( n18188 , n18093 );
not ( n18189 , n18188 );
buf ( n18190 , n17741 );
buf ( n18191 , n18190 );
buf ( n18192 , n18191 );
buf ( n18193 , n18192 );
buf ( n18194 , n17924 );
nand ( n18195 , n18193 , n18194 );
buf ( n18196 , n18195 );
buf ( n18197 , n18196 );
not ( n18198 , n18197 );
buf ( n18199 , n18198 );
buf ( n18200 , n18199 );
not ( n18201 , n18200 );
or ( n18202 , n18189 , n18201 );
buf ( n18203 , n17933 );
buf ( n18204 , n18092 );
nand ( n18205 , n18203 , n18204 );
buf ( n18206 , n18205 );
buf ( n18207 , n18206 );
nand ( n18208 , n18202 , n18207 );
buf ( n18209 , n18208 );
buf ( n18210 , n18209 );
not ( n18211 , n18210 );
buf ( n18212 , n18211 );
buf ( n18213 , n18212 );
nand ( n18214 , n18187 , n18213 );
buf ( n18215 , n18214 );
buf ( n18216 , n18215 );
not ( n18217 , n18216 );
buf ( n18218 , n18217 );
nand ( n18219 , n18105 , n18143 , n18218 );
and ( n18220 , n18084 , n18090 );
buf ( n18221 , n18220 );
buf ( n18222 , n18221 );
xor ( n18223 , n17955 , n17964 );
and ( n18224 , n18223 , n17982 );
and ( n18225 , n17955 , n17964 );
or ( n18226 , n18224 , n18225 );
buf ( n18227 , n18226 );
buf ( n18228 , n18227 );
xor ( n18229 , n18003 , n18020 );
and ( n18230 , n18229 , n18038 );
and ( n18231 , n18003 , n18020 );
or ( n18232 , n18230 , n18231 );
buf ( n18233 , n18232 );
buf ( n18234 , n18233 );
xor ( n18235 , n18228 , n18234 );
buf ( n18236 , n17996 );
not ( n18237 , n18236 );
buf ( n18238 , n10509 );
not ( n18239 , n18238 );
or ( n18240 , n18237 , n18239 );
buf ( n18241 , n3662 );
buf ( n18242 , n775 );
buf ( n18243 , n800 );
xor ( n18244 , n18242 , n18243 );
buf ( n18245 , n18244 );
buf ( n18246 , n18245 );
nand ( n18247 , n18241 , n18246 );
buf ( n18248 , n18247 );
buf ( n18249 , n18248 );
nand ( n18250 , n18240 , n18249 );
buf ( n18251 , n18250 );
buf ( n18252 , n17948 );
not ( n18253 , n18252 );
buf ( n18254 , n2709 );
not ( n18255 , n18254 );
or ( n18256 , n18253 , n18255 );
buf ( n18257 , n2713 );
buf ( n18258 , n808 );
nand ( n18259 , n18257 , n18258 );
buf ( n18260 , n18259 );
buf ( n18261 , n18260 );
nand ( n18262 , n18256 , n18261 );
buf ( n18263 , n18262 );
xor ( n18264 , n18251 , n18263 );
buf ( n18265 , n18013 );
not ( n18266 , n18265 );
buf ( n18267 , n3109 );
not ( n18268 , n18267 );
or ( n18269 , n18266 , n18268 );
buf ( n18270 , n1560 );
buf ( n18271 , n802 );
buf ( n18272 , n773 );
xor ( n18273 , n18271 , n18272 );
buf ( n18274 , n18273 );
buf ( n18275 , n18274 );
nand ( n18276 , n18270 , n18275 );
buf ( n18277 , n18276 );
buf ( n18278 , n18277 );
nand ( n18279 , n18269 , n18278 );
buf ( n18280 , n18279 );
xor ( n18281 , n18264 , n18280 );
buf ( n18282 , n18281 );
xor ( n18283 , n18235 , n18282 );
buf ( n18284 , n18283 );
buf ( n18285 , n18284 );
and ( n18286 , n17902 , n17903 );
buf ( n18287 , n18286 );
buf ( n18288 , n18287 );
buf ( n18289 , n17975 );
not ( n18290 , n18289 );
buf ( n18291 , n15873 );
not ( n18292 , n18291 );
or ( n18293 , n18290 , n18292 );
buf ( n18294 , n11137 );
buf ( n18295 , n771 );
buf ( n18296 , n804 );
xor ( n18297 , n18295 , n18296 );
buf ( n18298 , n18297 );
buf ( n18299 , n18298 );
nand ( n18300 , n18294 , n18299 );
buf ( n18301 , n18300 );
buf ( n18302 , n18301 );
nand ( n18303 , n18293 , n18302 );
buf ( n18304 , n18303 );
buf ( n18305 , n18304 );
xor ( n18306 , n18288 , n18305 );
buf ( n18307 , n18031 );
not ( n18308 , n18307 );
buf ( n18309 , n14278 );
not ( n18310 , n18309 );
or ( n18311 , n18308 , n18310 );
buf ( n18312 , n14284 );
xor ( n18313 , n806 , n769 );
buf ( n18314 , n18313 );
nand ( n18315 , n18312 , n18314 );
buf ( n18316 , n18315 );
buf ( n18317 , n18316 );
nand ( n18318 , n18311 , n18317 );
buf ( n18319 , n18318 );
buf ( n18320 , n18319 );
not ( n18321 , n18320 );
buf ( n18322 , n18321 );
buf ( n18323 , n18322 );
xor ( n18324 , n18306 , n18323 );
buf ( n18325 , n18324 );
buf ( n18326 , n18325 );
xor ( n18327 , n18047 , n18048 );
and ( n18328 , n18327 , n18055 );
and ( n18329 , n18047 , n18048 );
or ( n18330 , n18328 , n18329 );
buf ( n18331 , n18330 );
buf ( n18332 , n18331 );
xor ( n18333 , n18326 , n18332 );
xor ( n18334 , n17938 , n17985 );
and ( n18335 , n18334 , n18041 );
and ( n18336 , n17938 , n17985 );
or ( n18337 , n18335 , n18336 );
buf ( n18338 , n18337 );
buf ( n18339 , n18338 );
xor ( n18340 , n18333 , n18339 );
buf ( n18341 , n18340 );
buf ( n18342 , n18341 );
xor ( n18343 , n18285 , n18342 );
xor ( n18344 , n18058 , n18064 );
and ( n18345 , n18344 , n18071 );
and ( n18346 , n18058 , n18064 );
or ( n18347 , n18345 , n18346 );
buf ( n18348 , n18347 );
buf ( n18349 , n18348 );
xor ( n18350 , n18343 , n18349 );
buf ( n18351 , n18350 );
buf ( n18352 , n18351 );
xor ( n18353 , n18044 , n18074 );
and ( n18354 , n18353 , n18081 );
and ( n18355 , n18044 , n18074 );
or ( n18356 , n18354 , n18355 );
buf ( n18357 , n18356 );
buf ( n18358 , n18357 );
xor ( n18359 , n18352 , n18358 );
buf ( n18360 , n18359 );
buf ( n18361 , n18360 );
nor ( n18362 , n18222 , n18361 );
buf ( n18363 , n18362 );
buf ( n18364 , n18363 );
not ( n18365 , n18364 );
buf ( n18366 , n18365 );
buf ( n18367 , n18221 );
buf ( n18368 , n18360 );
nand ( n18369 , n18367 , n18368 );
buf ( n18370 , n18369 );
nand ( n18371 , n18366 , n18370 );
not ( n18372 , n18371 );
and ( n18373 , n18219 , n18372 );
not ( n18374 , n18219 );
and ( n18375 , n18374 , n18371 );
nor ( n18376 , n18373 , n18375 );
buf ( n18377 , n18376 );
buf ( n18378 , n13771 );
buf ( n18379 , n15325 );
nor ( n18380 , n18378 , n18379 );
buf ( n18381 , n18380 );
buf ( n18382 , n18381 );
not ( n18383 , n18382 );
buf ( n18384 , n10417 );
not ( n18385 , n18384 );
or ( n18386 , n18383 , n18385 );
buf ( n18387 , n15325 );
not ( n18388 , n18387 );
buf ( n18389 , n18388 );
buf ( n18390 , n18389 );
not ( n18391 , n18390 );
buf ( n18392 , n16313 );
not ( n18393 , n18392 );
or ( n18394 , n18391 , n18393 );
buf ( n18395 , n16368 );
not ( n18396 , n18395 );
buf ( n18397 , n18396 );
buf ( n18398 , n18397 );
nand ( n18399 , n18394 , n18398 );
buf ( n18400 , n18399 );
buf ( n18401 , n18400 );
not ( n18402 , n18401 );
buf ( n18403 , n18402 );
buf ( n18404 , n18403 );
nand ( n18405 , n18386 , n18404 );
buf ( n18406 , n18405 );
buf ( n18407 , n18406 );
buf ( n18408 , n16718 );
buf ( n18409 , n16745 );
nand ( n18410 , n18408 , n18409 );
buf ( n18411 , n18410 );
buf ( n18412 , n18411 );
not ( n18413 , n18412 );
buf ( n18414 , n18413 );
buf ( n18415 , n18414 );
and ( n18416 , n18407 , n18415 );
not ( n18417 , n18407 );
buf ( n18418 , n18411 );
and ( n18419 , n18417 , n18418 );
nor ( n18420 , n18416 , n18419 );
buf ( n18421 , n18420 );
buf ( n18422 , n18421 );
buf ( n18423 , n10359 );
not ( n18424 , n18423 );
nor ( n18425 , n7956 , n7727 );
nor ( n18426 , n8891 , n18425 );
buf ( n18427 , n18426 );
not ( n18428 , n18427 );
or ( n18429 , n18424 , n18428 );
not ( n18430 , n18425 );
not ( n18431 , n18430 );
not ( n18432 , n8798 );
or ( n18433 , n18431 , n18432 );
nand ( n18434 , n7956 , n7727 );
nand ( n18435 , n18433 , n18434 );
buf ( n18436 , n18435 );
not ( n18437 , n18436 );
buf ( n18438 , n18437 );
buf ( n18439 , n18438 );
nand ( n18440 , n18429 , n18439 );
buf ( n18441 , n18440 );
buf ( n18442 , n18441 );
buf ( n18443 , n8820 );
buf ( n18444 , n8825 );
and ( n18445 , n18443 , n18444 );
buf ( n18446 , n18445 );
buf ( n18447 , n18446 );
and ( n18448 , n18442 , n18447 );
not ( n18449 , n18442 );
buf ( n18450 , n18446 );
not ( n18451 , n18450 );
buf ( n18452 , n18451 );
buf ( n18453 , n18452 );
and ( n18454 , n18449 , n18453 );
nor ( n18455 , n18448 , n18454 );
buf ( n18456 , n18455 );
buf ( n18457 , n18456 );
buf ( n18458 , n4347 );
not ( n18459 , n18458 );
buf ( n18460 , n10417 );
not ( n18461 , n18460 );
or ( n18462 , n18459 , n18461 );
buf ( n18463 , n4352 );
nand ( n18464 , n18462 , n18463 );
buf ( n18465 , n18464 );
buf ( n18466 , n18465 );
nand ( n18467 , n13756 , n16293 );
buf ( n18468 , n18467 );
not ( n18469 , n18468 );
buf ( n18470 , n18469 );
buf ( n18471 , n18470 );
and ( n18472 , n18466 , n18471 );
not ( n18473 , n18466 );
buf ( n18474 , n18467 );
and ( n18475 , n18473 , n18474 );
nor ( n18476 , n18472 , n18475 );
buf ( n18477 , n18476 );
buf ( n18478 , n18477 );
buf ( n18479 , n13762 );
buf ( n18480 , n18479 );
buf ( n18481 , n18480 );
buf ( n18482 , n18481 );
not ( n18483 , n18482 );
buf ( n18484 , n18483 );
buf ( n18485 , n18484 );
buf ( n18486 , n12809 );
buf ( n18487 , n18486 );
buf ( n18488 , n18487 );
buf ( n18489 , n18488 );
buf ( n18490 , n13251 );
not ( n18491 , n18490 );
buf ( n18492 , n18491 );
buf ( n18493 , n18492 );
nand ( n18494 , n18489 , n18493 );
buf ( n18495 , n18494 );
buf ( n18496 , n18495 );
nor ( n18497 , n18485 , n18496 );
buf ( n18498 , n18497 );
buf ( n18499 , n18498 );
not ( n18500 , n18499 );
buf ( n18501 , n10427 );
not ( n18502 , n18501 );
or ( n18503 , n18500 , n18502 );
buf ( n18504 , n16311 );
buf ( n18505 , n18504 );
not ( n18506 , n18505 );
buf ( n18507 , n18495 );
not ( n18508 , n18507 );
buf ( n18509 , n18508 );
buf ( n18510 , n18509 );
not ( n18511 , n18510 );
or ( n18512 , n18506 , n18511 );
buf ( n18513 , n18492 );
not ( n18514 , n18513 );
buf ( n18515 , n16281 );
buf ( n18516 , n18515 );
buf ( n18517 , n18516 );
buf ( n18518 , n18517 );
not ( n18519 , n18518 );
or ( n18520 , n18514 , n18519 );
buf ( n18521 , n16246 );
nand ( n18522 , n18520 , n18521 );
buf ( n18523 , n18522 );
buf ( n18524 , n18523 );
not ( n18525 , n18524 );
buf ( n18526 , n18525 );
buf ( n18527 , n18526 );
nand ( n18528 , n18512 , n18527 );
buf ( n18529 , n18528 );
not ( n18530 , n18529 );
buf ( n18531 , n18530 );
nand ( n18532 , n18503 , n18531 );
buf ( n18533 , n18532 );
buf ( n18534 , n13674 );
and ( n18535 , n16252 , n13253 );
buf ( n18536 , n18535 );
or ( n18537 , n18534 , n18536 );
buf ( n18538 , n18537 );
xnor ( n18539 , n18533 , n18538 );
buf ( n18540 , n18539 );
not ( n18541 , n10307 );
buf ( n18542 , n9367 );
not ( n18543 , n18542 );
buf ( n18544 , n18543 );
buf ( n18545 , n18544 );
buf ( n18546 , n10319 );
nand ( n18547 , n18545 , n18546 );
buf ( n18548 , n18547 );
not ( n18549 , n18548 );
or ( n18550 , n18541 , n18549 );
not ( n18551 , n18548 );
nand ( n18552 , n18551 , n10256 , n10306 );
nand ( n18553 , n18550 , n18552 );
buf ( n18554 , n18553 );
buf ( n18555 , n17682 );
buf ( n18556 , n18555 );
buf ( n18557 , n18556 );
buf ( n18558 , n18557 );
buf ( n18559 , n18558 );
not ( n18560 , n18559 );
buf ( n18561 , n18158 );
not ( n18562 , n18561 );
or ( n18563 , n18560 , n18562 );
buf ( n18564 , n18166 );
nand ( n18565 , n18563 , n18564 );
buf ( n18566 , n18565 );
not ( n18567 , n18566 );
buf ( n18568 , n10430 );
buf ( n18569 , n18130 );
not ( n18570 , n18569 );
buf ( n18571 , n18570 );
buf ( n18572 , n18571 );
buf ( n18573 , n17729 );
buf ( n18574 , n18558 );
and ( n18575 , n18573 , n18574 );
buf ( n18576 , n18575 );
buf ( n18577 , n18576 );
and ( n18578 , n18572 , n18577 );
buf ( n18579 , n18578 );
buf ( n18580 , n18579 );
nand ( n18581 , n18568 , n18580 );
buf ( n18582 , n18581 );
buf ( n18583 , n16830 );
not ( n18584 , n18583 );
buf ( n18585 , n18584 );
buf ( n18586 , n18585 );
buf ( n18587 , n18576 );
nand ( n18588 , n18586 , n18587 );
buf ( n18589 , n18588 );
nand ( n18590 , n18567 , n18582 , n18589 );
buf ( n18591 , n18590 );
buf ( n18592 , n17645 );
not ( n18593 , n18592 );
buf ( n18594 , n18175 );
nor ( n18595 , n18593 , n18594 );
buf ( n18596 , n18595 );
buf ( n18597 , n18596 );
and ( n18598 , n18591 , n18597 );
not ( n18599 , n18591 );
buf ( n18600 , n18596 );
not ( n18601 , n18600 );
buf ( n18602 , n18601 );
buf ( n18603 , n18602 );
and ( n18604 , n18599 , n18603 );
nor ( n18605 , n18598 , n18604 );
buf ( n18606 , n18605 );
buf ( n18607 , n18606 );
buf ( n18608 , n18488 );
not ( n18609 , n18608 );
buf ( n18610 , n18484 );
nor ( n18611 , n18609 , n18610 );
buf ( n18612 , n18611 );
buf ( n18613 , n18612 );
not ( n18614 , n18613 );
buf ( n18615 , n10427 );
not ( n18616 , n18615 );
or ( n18617 , n18614 , n18616 );
buf ( n18618 , n18488 );
buf ( n18619 , n18504 );
and ( n18620 , n18618 , n18619 );
buf ( n18621 , n18517 );
nor ( n18622 , n18620 , n18621 );
buf ( n18623 , n18622 );
buf ( n18624 , n18623 );
nand ( n18625 , n18617 , n18624 );
buf ( n18626 , n18625 );
buf ( n18627 , n18626 );
buf ( n18628 , n18492 );
buf ( n18629 , n16246 );
nand ( n18630 , n18628 , n18629 );
buf ( n18631 , n18630 );
buf ( n18632 , n18631 );
not ( n18633 , n18632 );
buf ( n18634 , n18633 );
buf ( n18635 , n18634 );
and ( n18636 , n18627 , n18635 );
not ( n18637 , n18627 );
buf ( n18638 , n18631 );
and ( n18639 , n18637 , n18638 );
nor ( n18640 , n18636 , n18639 );
buf ( n18641 , n18640 );
buf ( n18642 , n18641 );
buf ( n18643 , n18481 );
not ( n18644 , n18643 );
buf ( n18645 , n10417 );
not ( n18646 , n18645 );
or ( n18647 , n18644 , n18646 );
buf ( n18648 , n18504 );
not ( n18649 , n18648 );
buf ( n18650 , n18649 );
buf ( n18651 , n18650 );
nand ( n18652 , n18647 , n18651 );
buf ( n18653 , n18652 );
buf ( n18654 , n18653 );
or ( n18655 , n12807 , n12805 );
buf ( n18656 , n18655 );
buf ( n18657 , n16258 );
nand ( n18658 , n18656 , n18657 );
buf ( n18659 , n18658 );
buf ( n18660 , n18659 );
not ( n18661 , n18660 );
buf ( n18662 , n18661 );
buf ( n18663 , n18662 );
and ( n18664 , n18654 , n18663 );
not ( n18665 , n18654 );
buf ( n18666 , n18659 );
and ( n18667 , n18665 , n18666 );
nor ( n18668 , n18664 , n18667 );
buf ( n18669 , n18668 );
buf ( n18670 , n18669 );
buf ( n18671 , n13759 );
buf ( n18672 , n18671 );
buf ( n18673 , n18672 );
buf ( n18674 , n18673 );
buf ( n18675 , n13723 );
buf ( n18676 , n18675 );
buf ( n18677 , n18676 );
buf ( n18678 , n18677 );
nor ( n18679 , n18674 , n18678 );
buf ( n18680 , n18679 );
nand ( n18681 , n18680 , n10417 );
not ( n18682 , n18681 );
buf ( n18683 , n16294 );
not ( n18684 , n18683 );
nor ( n18685 , n18684 , n18677 );
nand ( n18686 , n16299 , n16306 );
buf ( n18687 , n16300 );
buf ( n18688 , n18687 );
buf ( n18689 , n18688 );
buf ( n18690 , n18689 );
not ( n18691 , n18690 );
buf ( n18692 , n18691 );
nor ( n18693 , n18685 , n18686 , n18692 );
not ( n18694 , n18693 );
or ( n18695 , n18682 , n18694 );
nor ( n18696 , n18685 , n18692 );
not ( n18697 , n18696 );
not ( n18698 , n18681 );
or ( n18699 , n18697 , n18698 );
nand ( n18700 , n18699 , n18686 );
nand ( n18701 , n18695 , n18700 );
buf ( n18702 , n18701 );
buf ( n18703 , n17701 );
buf ( n18704 , n16784 );
nor ( n18705 , n18703 , n18704 );
buf ( n18706 , n18705 );
not ( n18707 , n18706 );
not ( n18708 , n16313 );
buf ( n18709 , n8862 );
buf ( n18710 , n6857 );
and ( n18711 , n18709 , n18710 );
buf ( n18712 , n18711 );
buf ( n18713 , n18712 );
buf ( n18714 , n18713 );
buf ( n18715 , n18714 );
buf ( n18716 , n18715 );
not ( n18717 , n18716 );
buf ( n18718 , n8799 );
buf ( n18719 , n8854 );
not ( n18720 , n18719 );
buf ( n18721 , n18720 );
buf ( n18722 , n18721 );
nand ( n18723 , n18718 , n18722 );
buf ( n18724 , n18723 );
buf ( n18725 , n18724 );
not ( n18726 , n18725 );
buf ( n18727 , n10359 );
not ( n18728 , n18727 );
nand ( n18729 , n8895 , n8888 );
buf ( n18730 , n18729 );
nor ( n18731 , n18728 , n18730 );
buf ( n18732 , n18731 );
buf ( n18733 , n18732 );
not ( n18734 , n18733 );
buf ( n18735 , n18734 );
buf ( n18736 , n18735 );
nand ( n18737 , n18726 , n18736 );
buf ( n18738 , n18737 );
buf ( n18739 , n18738 );
not ( n18740 , n18739 );
or ( n18741 , n18717 , n18740 );
buf ( n18742 , n10408 );
buf ( n18743 , n18742 );
buf ( n18744 , n18743 );
buf ( n18745 , n18744 );
not ( n18746 , n6884 );
not ( n18747 , n8862 );
or ( n18748 , n18746 , n18747 );
not ( n18749 , n6353 );
nand ( n18750 , n18748 , n18749 );
buf ( n18751 , n18750 );
buf ( n18752 , n18751 );
buf ( n18753 , n18752 );
buf ( n18754 , n18753 );
nor ( n18755 , n18745 , n18754 );
buf ( n18756 , n18755 );
buf ( n18757 , n18756 );
nand ( n18758 , n18741 , n18757 );
buf ( n18759 , n18758 );
buf ( n18760 , n18759 );
buf ( n18761 , n5887 );
not ( n18762 , n18761 );
buf ( n18763 , n18744 );
nor ( n18764 , n18762 , n18763 );
buf ( n18765 , n18764 );
buf ( n18766 , n18765 );
buf ( n18767 , n13765 );
nor ( n18768 , n18766 , n18767 );
buf ( n18769 , n18768 );
buf ( n18770 , n18769 );
nand ( n18771 , n18760 , n18770 );
buf ( n18772 , n18771 );
nand ( n18773 , n18708 , n18772 );
not ( n18774 , n18773 );
or ( n18775 , n18707 , n18774 );
buf ( n18776 , n16783 );
not ( n18777 , n18776 );
buf ( n18778 , n16368 );
not ( n18779 , n18778 );
or ( n18780 , n18777 , n18779 );
buf ( n18781 , n16807 );
nand ( n18782 , n18780 , n18781 );
buf ( n18783 , n18782 );
buf ( n18784 , n18783 );
buf ( n18785 , n17701 );
not ( n18786 , n18785 );
buf ( n18787 , n18786 );
buf ( n18788 , n18787 );
nand ( n18789 , n18784 , n18788 );
buf ( n18790 , n18789 );
buf ( n18791 , n18790 );
buf ( n18792 , n18151 );
and ( n18793 , n18791 , n18792 );
buf ( n18794 , n18793 );
nand ( n18795 , n18775 , n18794 );
and ( n18796 , n18157 , n18154 );
and ( n18797 , n18795 , n18796 );
not ( n18798 , n18795 );
not ( n18799 , n18796 );
and ( n18800 , n18798 , n18799 );
nor ( n18801 , n18797 , n18800 );
buf ( n18802 , n18801 );
not ( n18803 , n8884 );
not ( n18804 , n10307 );
not ( n18805 , n9371 );
or ( n18806 , n18804 , n18805 );
nand ( n18807 , n18806 , n10356 );
not ( n18808 , n18807 );
or ( n18809 , n18803 , n18808 );
buf ( n18810 , n8772 );
buf ( n18811 , n18810 );
buf ( n18812 , n18811 );
not ( n18813 , n18812 );
nand ( n18814 , n18809 , n18813 );
buf ( n18815 , n18814 );
buf ( n18816 , n8788 );
not ( n18817 , n18816 );
buf ( n18818 , n8875 );
buf ( n18819 , n18818 );
buf ( n18820 , n18819 );
buf ( n18821 , n18820 );
nand ( n18822 , n18817 , n18821 );
buf ( n18823 , n18822 );
buf ( n18824 , n18823 );
not ( n18825 , n18824 );
buf ( n18826 , n18825 );
buf ( n18827 , n18826 );
and ( n18828 , n18815 , n18827 );
not ( n18829 , n18815 );
buf ( n18830 , n18823 );
and ( n18831 , n18829 , n18830 );
nor ( n18832 , n18828 , n18831 );
buf ( n18833 , n18832 );
buf ( n18834 , n18833 );
buf ( n18835 , n832 );
buf ( n18836 , n880 );
xor ( n18837 , n18835 , n18836 );
buf ( n18838 , n18837 );
buf ( n18839 , n18838 );
not ( n18840 , n18839 );
not ( n18841 , n880 );
not ( n18842 , n881 );
or ( n18843 , n18841 , n18842 );
not ( n18844 , n880 );
not ( n18845 , n881 );
nand ( n18846 , n18844 , n18845 );
nand ( n18847 , n18843 , n18846 );
xor ( n18848 , n881 , n882 );
nor ( n18849 , n18847 , n18848 );
buf ( n18850 , n18849 );
buf ( n18851 , n18850 );
not ( n18852 , n18851 );
or ( n18853 , n18840 , n18852 );
not ( n18854 , n882 );
not ( n18855 , n881 );
not ( n18856 , n18855 );
or ( n18857 , n18854 , n18856 );
not ( n18858 , n882 );
nand ( n18859 , n18858 , n881 );
nand ( n18860 , n18857 , n18859 );
buf ( n18861 , n18860 );
buf ( n18862 , n880 );
nand ( n18863 , n18861 , n18862 );
buf ( n18864 , n18863 );
buf ( n18865 , n18864 );
nand ( n18866 , n18853 , n18865 );
buf ( n18867 , n18866 );
buf ( n18868 , n18867 );
buf ( n18869 , n843 );
buf ( n18870 , n868 );
xor ( n18871 , n18869 , n18870 );
buf ( n18872 , n18871 );
buf ( n18873 , n18872 );
not ( n18874 , n18873 );
xor ( n18875 , n869 , n870 );
not ( n18876 , n18875 );
buf ( n18877 , n18876 );
buf ( n18878 , n868 );
buf ( n18879 , n869 );
xor ( n18880 , n18878 , n18879 );
buf ( n18881 , n18880 );
buf ( n18882 , n18881 );
and ( n18883 , n18877 , n18882 );
buf ( n18884 , n18883 );
buf ( n18885 , n18884 );
buf ( n18886 , n18885 );
buf ( n18887 , n18886 );
buf ( n18888 , n18887 );
not ( n18889 , n18888 );
or ( n18890 , n18874 , n18889 );
not ( n18891 , n18875 );
not ( n18892 , n18891 );
buf ( n18893 , n18892 );
not ( n18894 , n18893 );
buf ( n18895 , n18894 );
buf ( n18896 , n18895 );
not ( n18897 , n18896 );
buf ( n18898 , n18897 );
buf ( n18899 , n18898 );
buf ( n18900 , n842 );
buf ( n18901 , n868 );
xor ( n18902 , n18900 , n18901 );
buf ( n18903 , n18902 );
buf ( n18904 , n18903 );
nand ( n18905 , n18899 , n18904 );
buf ( n18906 , n18905 );
buf ( n18907 , n18906 );
nand ( n18908 , n18890 , n18907 );
buf ( n18909 , n18908 );
buf ( n18910 , n18909 );
xor ( n18911 , n18868 , n18910 );
buf ( n18912 , n846 );
buf ( n18913 , n866 );
xor ( n18914 , n18912 , n18913 );
buf ( n18915 , n18914 );
buf ( n18916 , n18915 );
not ( n18917 , n18916 );
and ( n18918 , n867 , n866 );
not ( n18919 , n867 );
not ( n18920 , n866 );
and ( n18921 , n18919 , n18920 );
nor ( n18922 , n18918 , n18921 );
not ( n18923 , n18922 );
buf ( n18924 , n867 );
buf ( n18925 , n868 );
xor ( n18926 , n18924 , n18925 );
buf ( n18927 , n18926 );
nor ( n18928 , n18923 , n18927 );
buf ( n18929 , n18928 );
buf ( n18930 , n18929 );
buf ( n18931 , n18930 );
buf ( n18932 , n18931 );
not ( n18933 , n18932 );
or ( n18934 , n18917 , n18933 );
buf ( n18935 , n867 );
buf ( n18936 , n868 );
xor ( n18937 , n18935 , n18936 );
buf ( n18938 , n18937 );
buf ( n18939 , n18938 );
not ( n18940 , n18939 );
buf ( n18941 , n18940 );
buf ( n18942 , n18941 );
not ( n18943 , n18942 );
buf ( n18944 , n18943 );
buf ( n18945 , n18944 );
buf ( n18946 , n845 );
buf ( n18947 , n866 );
xor ( n18948 , n18946 , n18947 );
buf ( n18949 , n18948 );
buf ( n18950 , n18949 );
nand ( n18951 , n18945 , n18950 );
buf ( n18952 , n18951 );
buf ( n18953 , n18952 );
nand ( n18954 , n18934 , n18953 );
buf ( n18955 , n18954 );
buf ( n18956 , n18955 );
buf ( n18957 , n838 );
buf ( n18958 , n874 );
xor ( n18959 , n18957 , n18958 );
buf ( n18960 , n18959 );
buf ( n18961 , n18960 );
not ( n18962 , n18961 );
buf ( n18963 , n875 );
not ( n18964 , n18963 );
buf ( n18965 , n876 );
nand ( n18966 , n18964 , n18965 );
buf ( n18967 , n18966 );
buf ( n18968 , n876 );
not ( n18969 , n18968 );
buf ( n18970 , n875 );
nand ( n18971 , n18969 , n18970 );
buf ( n18972 , n18971 );
xor ( n18973 , n874 , n875 );
and ( n18974 , n18967 , n18972 , n18973 );
buf ( n18975 , n18974 );
buf ( n18976 , n18975 );
buf ( n18977 , n18976 );
buf ( n18978 , n18977 );
not ( n18979 , n18978 );
or ( n18980 , n18962 , n18979 );
xor ( n18981 , n876 , n875 );
buf ( n18982 , n18981 );
not ( n18983 , n18982 );
buf ( n18984 , n18983 );
buf ( n18985 , n18984 );
not ( n18986 , n18985 );
buf ( n18987 , n18986 );
buf ( n18988 , n18987 );
buf ( n18989 , n837 );
buf ( n18990 , n874 );
xor ( n18991 , n18989 , n18990 );
buf ( n18992 , n18991 );
buf ( n18993 , n18992 );
nand ( n18994 , n18988 , n18993 );
buf ( n18995 , n18994 );
buf ( n18996 , n18995 );
nand ( n18997 , n18980 , n18996 );
buf ( n18998 , n18997 );
buf ( n18999 , n18998 );
xor ( n19000 , n18956 , n18999 );
not ( n19001 , n865 );
not ( n19002 , n864 );
not ( n19003 , n19002 );
or ( n19004 , n19001 , n19003 );
nand ( n19005 , n19004 , n866 );
not ( n19006 , n864 );
not ( n19007 , n865 );
not ( n19008 , n19007 );
or ( n19009 , n19006 , n19008 );
not ( n19010 , n866 );
nand ( n19011 , n19009 , n19010 );
nand ( n19012 , n19005 , n19011 );
not ( n19013 , n19012 );
buf ( n19014 , n19013 );
not ( n19015 , n19014 );
buf ( n19016 , n19015 );
buf ( n19017 , n19016 );
buf ( n19018 , n848 );
buf ( n19019 , n864 );
xnor ( n19020 , n19018 , n19019 );
buf ( n19021 , n19020 );
buf ( n19022 , n19021 );
or ( n19023 , n19017 , n19022 );
buf ( n19024 , n865 );
buf ( n19025 , n866 );
xor ( n19026 , n19024 , n19025 );
buf ( n19027 , n19026 );
buf ( n19028 , n19027 );
buf ( n19029 , n19028 );
buf ( n19030 , n19029 );
buf ( n19031 , n19030 );
not ( n19032 , n19031 );
buf ( n19033 , n19032 );
buf ( n19034 , n19033 );
buf ( n19035 , n847 );
buf ( n19036 , n864 );
xor ( n19037 , n19035 , n19036 );
buf ( n19038 , n19037 );
buf ( n19039 , n19038 );
not ( n19040 , n19039 );
buf ( n19041 , n19040 );
buf ( n19042 , n19041 );
or ( n19043 , n19034 , n19042 );
nand ( n19044 , n19023 , n19043 );
buf ( n19045 , n19044 );
buf ( n19046 , n19045 );
and ( n19047 , n19000 , n19046 );
and ( n19048 , n18956 , n18999 );
or ( n19049 , n19047 , n19048 );
buf ( n19050 , n19049 );
buf ( n19051 , n19050 );
and ( n19052 , n18911 , n19051 );
and ( n19053 , n18868 , n18910 );
or ( n19054 , n19052 , n19053 );
buf ( n19055 , n19054 );
buf ( n19056 , n19055 );
buf ( n19057 , n848 );
buf ( n19058 , n864 );
and ( n19059 , n19057 , n19058 );
buf ( n19060 , n19059 );
not ( n19061 , n19060 );
buf ( n19062 , n835 );
buf ( n19063 , n876 );
xor ( n19064 , n19062 , n19063 );
buf ( n19065 , n19064 );
buf ( n19066 , n19065 );
not ( n19067 , n19066 );
not ( n19068 , n876 );
not ( n19069 , n19068 );
nand ( n19070 , n877 , n878 );
not ( n19071 , n19070 );
or ( n19072 , n19069 , n19071 );
or ( n19073 , n877 , n878 );
nand ( n19074 , n19073 , n876 );
nand ( n19075 , n19072 , n19074 );
not ( n19076 , n19075 );
buf ( n19077 , n19076 );
buf ( n19078 , n19077 );
not ( n19079 , n19078 );
or ( n19080 , n19067 , n19079 );
xor ( n19081 , n877 , n878 );
buf ( n19082 , n19081 );
buf ( n19083 , n19082 );
buf ( n19084 , n19083 );
buf ( n19085 , n19084 );
buf ( n19086 , n19085 );
buf ( n19087 , n834 );
buf ( n19088 , n876 );
xor ( n19089 , n19087 , n19088 );
buf ( n19090 , n19089 );
buf ( n19091 , n19090 );
nand ( n19092 , n19086 , n19091 );
buf ( n19093 , n19092 );
buf ( n19094 , n19093 );
nand ( n19095 , n19080 , n19094 );
buf ( n19096 , n19095 );
not ( n19097 , n19096 );
xor ( n19098 , n19061 , n19097 );
buf ( n19099 , n841 );
buf ( n19100 , n870 );
xor ( n19101 , n19099 , n19100 );
buf ( n19102 , n19101 );
buf ( n19103 , n19102 );
not ( n19104 , n19103 );
not ( n19105 , n871 );
not ( n19106 , n872 );
not ( n19107 , n19106 );
or ( n19108 , n19105 , n19107 );
buf ( n19109 , n871 );
not ( n19110 , n19109 );
buf ( n19111 , n872 );
nand ( n19112 , n19110 , n19111 );
buf ( n19113 , n19112 );
nand ( n19114 , n19108 , n19113 );
buf ( n19115 , n19114 );
xnor ( n19116 , n870 , n871 );
buf ( n19117 , n19116 );
nor ( n19118 , n19115 , n19117 );
buf ( n19119 , n19118 );
buf ( n19120 , n19119 );
buf ( n19121 , n19120 );
buf ( n19122 , n19121 );
buf ( n19123 , n19122 );
buf ( n19124 , n19123 );
buf ( n19125 , n19124 );
buf ( n19126 , n19125 );
not ( n19127 , n19126 );
or ( n19128 , n19104 , n19127 );
buf ( n19129 , n19114 );
buf ( n19130 , n19129 );
buf ( n19131 , n19130 );
buf ( n19132 , n19131 );
buf ( n19133 , n19132 );
buf ( n19134 , n19133 );
buf ( n19135 , n19134 );
buf ( n19136 , n840 );
buf ( n19137 , n870 );
xor ( n19138 , n19136 , n19137 );
buf ( n19139 , n19138 );
buf ( n19140 , n19139 );
nand ( n19141 , n19135 , n19140 );
buf ( n19142 , n19141 );
buf ( n19143 , n19142 );
nand ( n19144 , n19128 , n19143 );
buf ( n19145 , n19144 );
xor ( n19146 , n19098 , n19145 );
buf ( n19147 , n836 );
buf ( n19148 , n876 );
xor ( n19149 , n19147 , n19148 );
buf ( n19150 , n19149 );
buf ( n19151 , n19150 );
not ( n19152 , n19151 );
buf ( n19153 , n19076 );
buf ( n19154 , n19153 );
not ( n19155 , n19154 );
or ( n19156 , n19152 , n19155 );
buf ( n19157 , n19085 );
buf ( n19158 , n19065 );
nand ( n19159 , n19157 , n19158 );
buf ( n19160 , n19159 );
buf ( n19161 , n19160 );
nand ( n19162 , n19156 , n19161 );
buf ( n19163 , n19162 );
not ( n19164 , n19163 );
buf ( n19165 , n844 );
buf ( n19166 , n868 );
xor ( n19167 , n19165 , n19166 );
buf ( n19168 , n19167 );
buf ( n19169 , n19168 );
not ( n19170 , n19169 );
buf ( n19171 , n18887 );
not ( n19172 , n19171 );
or ( n19173 , n19170 , n19172 );
buf ( n19174 , n18892 );
buf ( n19175 , n19174 );
buf ( n19176 , n18872 );
nand ( n19177 , n19175 , n19176 );
buf ( n19178 , n19177 );
buf ( n19179 , n19178 );
nand ( n19180 , n19173 , n19179 );
buf ( n19181 , n19180 );
buf ( n19182 , n19181 );
not ( n19183 , n19182 );
buf ( n19184 , n19183 );
nand ( n19185 , n19164 , n19184 );
not ( n19186 , n19185 );
buf ( n19187 , n842 );
buf ( n19188 , n870 );
xor ( n19189 , n19187 , n19188 );
buf ( n19190 , n19189 );
buf ( n19191 , n19190 );
not ( n19192 , n19191 );
buf ( n19193 , n19125 );
not ( n19194 , n19193 );
or ( n19195 , n19192 , n19194 );
buf ( n19196 , n19134 );
buf ( n19197 , n19102 );
nand ( n19198 , n19196 , n19197 );
buf ( n19199 , n19198 );
buf ( n19200 , n19199 );
nand ( n19201 , n19195 , n19200 );
buf ( n19202 , n19201 );
not ( n19203 , n19202 );
or ( n19204 , n19186 , n19203 );
buf ( n19205 , n19163 );
buf ( n19206 , n19181 );
nand ( n19207 , n19205 , n19206 );
buf ( n19208 , n19207 );
nand ( n19209 , n19204 , n19208 );
or ( n19210 , n19146 , n19209 );
buf ( n19211 , n849 );
buf ( n19212 , n864 );
and ( n19213 , n19211 , n19212 );
buf ( n19214 , n19213 );
buf ( n19215 , n840 );
buf ( n19216 , n872 );
xor ( n19217 , n19215 , n19216 );
buf ( n19218 , n19217 );
buf ( n19219 , n19218 );
not ( n19220 , n19219 );
xor ( n19221 , n873 , n874 );
buf ( n19222 , n19221 );
not ( n19223 , n19222 );
buf ( n19224 , n19223 );
buf ( n19225 , n872 );
buf ( n19226 , n873 );
xor ( n19227 , n19225 , n19226 );
buf ( n19228 , n19227 );
nand ( n19229 , n19224 , n19228 );
not ( n19230 , n19229 );
buf ( n19231 , n19230 );
not ( n19232 , n19231 );
or ( n19233 , n19220 , n19232 );
buf ( n19234 , n19221 );
buf ( n19235 , n19234 );
buf ( n19236 , n19235 );
buf ( n19237 , n839 );
buf ( n19238 , n872 );
xor ( n19239 , n19237 , n19238 );
buf ( n19240 , n19239 );
buf ( n19241 , n19240 );
nand ( n19242 , n19236 , n19241 );
buf ( n19243 , n19242 );
buf ( n19244 , n19243 );
nand ( n19245 , n19233 , n19244 );
buf ( n19246 , n19245 );
xor ( n19247 , n19214 , n19246 );
buf ( n19248 , n834 );
buf ( n19249 , n878 );
xor ( n19250 , n19248 , n19249 );
buf ( n19251 , n19250 );
buf ( n19252 , n19251 );
not ( n19253 , n19252 );
xnor ( n19254 , n879 , n878 );
xor ( n19255 , n879 , n880 );
nor ( n19256 , n19254 , n19255 );
buf ( n19257 , n19256 );
buf ( n19258 , n19257 );
buf ( n19259 , n19258 );
buf ( n19260 , n19259 );
not ( n19261 , n19260 );
or ( n19262 , n19253 , n19261 );
buf ( n19263 , n19255 );
buf ( n19264 , n19263 );
buf ( n19265 , n19264 );
buf ( n19266 , n19265 );
buf ( n19267 , n833 );
buf ( n19268 , n878 );
xor ( n19269 , n19267 , n19268 );
buf ( n19270 , n19269 );
buf ( n19271 , n19270 );
nand ( n19272 , n19266 , n19271 );
buf ( n19273 , n19272 );
buf ( n19274 , n19273 );
nand ( n19275 , n19262 , n19274 );
buf ( n19276 , n19275 );
and ( n19277 , n19247 , n19276 );
and ( n19278 , n19214 , n19246 );
or ( n19279 , n19277 , n19278 );
nand ( n19280 , n19210 , n19279 );
nand ( n19281 , n19209 , n19146 );
nand ( n19282 , n19280 , n19281 );
buf ( n19283 , n19282 );
xor ( n19284 , n19056 , n19283 );
buf ( n19285 , n19060 );
not ( n19286 , n19285 );
buf ( n19287 , n19096 );
not ( n19288 , n19287 );
or ( n19289 , n19286 , n19288 );
buf ( n19290 , n19096 );
buf ( n19291 , n19060 );
or ( n19292 , n19290 , n19291 );
buf ( n19293 , n19145 );
nand ( n19294 , n19292 , n19293 );
buf ( n19295 , n19294 );
buf ( n19296 , n19295 );
nand ( n19297 , n19289 , n19296 );
buf ( n19298 , n19297 );
buf ( n19299 , n19298 );
buf ( n19300 , n18949 );
not ( n19301 , n19300 );
buf ( n19302 , n18931 );
not ( n19303 , n19302 );
or ( n19304 , n19301 , n19303 );
buf ( n19305 , n18944 );
buf ( n19306 , n844 );
buf ( n19307 , n866 );
xor ( n19308 , n19306 , n19307 );
buf ( n19309 , n19308 );
buf ( n19310 , n19309 );
nand ( n19311 , n19305 , n19310 );
buf ( n19312 , n19311 );
buf ( n19313 , n19312 );
nand ( n19314 , n19304 , n19313 );
buf ( n19315 , n19314 );
buf ( n19316 , n19315 );
not ( n19317 , n19235 );
buf ( n19318 , n838 );
buf ( n19319 , n872 );
xor ( n19320 , n19318 , n19319 );
buf ( n19321 , n19320 );
not ( n19322 , n19321 );
or ( n19323 , n19317 , n19322 );
nand ( n19324 , n19240 , n19230 );
nand ( n19325 , n19323 , n19324 );
buf ( n19326 , n19325 );
xor ( n19327 , n19316 , n19326 );
buf ( n19328 , n19038 );
not ( n19329 , n19328 );
buf ( n19330 , n19013 );
buf ( n19331 , n19330 );
not ( n19332 , n19331 );
or ( n19333 , n19329 , n19332 );
buf ( n19334 , n19030 );
xor ( n19335 , n864 , n846 );
buf ( n19336 , n19335 );
nand ( n19337 , n19334 , n19336 );
buf ( n19338 , n19337 );
buf ( n19339 , n19338 );
nand ( n19340 , n19333 , n19339 );
buf ( n19341 , n19340 );
buf ( n19342 , n19341 );
and ( n19343 , n19327 , n19342 );
and ( n19344 , n19316 , n19326 );
or ( n19345 , n19343 , n19344 );
buf ( n19346 , n19345 );
buf ( n19347 , n19346 );
xor ( n19348 , n19299 , n19347 );
buf ( n19349 , n19270 );
not ( n19350 , n19349 );
buf ( n19351 , n19259 );
not ( n19352 , n19351 );
or ( n19353 , n19350 , n19352 );
buf ( n19354 , n19265 );
buf ( n19355 , n832 );
buf ( n19356 , n878 );
xor ( n19357 , n19355 , n19356 );
buf ( n19358 , n19357 );
buf ( n19359 , n19358 );
nand ( n19360 , n19354 , n19359 );
buf ( n19361 , n19360 );
buf ( n19362 , n19361 );
nand ( n19363 , n19353 , n19362 );
buf ( n19364 , n19363 );
buf ( n19365 , n19364 );
buf ( n19366 , n18860 );
buf ( n19367 , n18850 );
or ( n19368 , n19366 , n19367 );
buf ( n19369 , n880 );
nand ( n19370 , n19368 , n19369 );
buf ( n19371 , n19370 );
buf ( n19372 , n19371 );
xor ( n19373 , n19365 , n19372 );
buf ( n19374 , n18992 );
not ( n19375 , n19374 );
buf ( n19376 , n18977 );
not ( n19377 , n19376 );
or ( n19378 , n19375 , n19377 );
buf ( n19379 , n18987 );
buf ( n19380 , n836 );
buf ( n19381 , n874 );
xor ( n19382 , n19380 , n19381 );
buf ( n19383 , n19382 );
buf ( n19384 , n19383 );
nand ( n19385 , n19379 , n19384 );
buf ( n19386 , n19385 );
buf ( n19387 , n19386 );
nand ( n19388 , n19378 , n19387 );
buf ( n19389 , n19388 );
buf ( n19390 , n19389 );
and ( n19391 , n19373 , n19390 );
and ( n19392 , n19365 , n19372 );
or ( n19393 , n19391 , n19392 );
buf ( n19394 , n19393 );
buf ( n19395 , n19394 );
xor ( n19396 , n19348 , n19395 );
buf ( n19397 , n19396 );
buf ( n19398 , n19397 );
xor ( n19399 , n19284 , n19398 );
buf ( n19400 , n19399 );
buf ( n19401 , n19400 );
buf ( n19402 , n847 );
buf ( n19403 , n864 );
and ( n19404 , n19402 , n19403 );
buf ( n19405 , n19404 );
buf ( n19406 , n19405 );
buf ( n19407 , n19335 );
not ( n19408 , n19407 );
buf ( n19409 , n19013 );
not ( n19410 , n19409 );
or ( n19411 , n19408 , n19410 );
buf ( n19412 , n19030 );
xor ( n19413 , n864 , n845 );
buf ( n19414 , n19413 );
nand ( n19415 , n19412 , n19414 );
buf ( n19416 , n19415 );
buf ( n19417 , n19416 );
nand ( n19418 , n19411 , n19417 );
buf ( n19419 , n19418 );
buf ( n19420 , n19419 );
xor ( n19421 , n19406 , n19420 );
buf ( n19422 , n19321 );
not ( n19423 , n19422 );
buf ( n19424 , n19230 );
not ( n19425 , n19424 );
or ( n19426 , n19423 , n19425 );
buf ( n19427 , n19235 );
xor ( n19428 , n872 , n837 );
buf ( n19429 , n19428 );
nand ( n19430 , n19427 , n19429 );
buf ( n19431 , n19430 );
buf ( n19432 , n19431 );
nand ( n19433 , n19426 , n19432 );
buf ( n19434 , n19433 );
buf ( n19435 , n19434 );
xor ( n19436 , n19421 , n19435 );
buf ( n19437 , n19436 );
buf ( n19438 , n19437 );
buf ( n19439 , n19309 );
not ( n19440 , n19439 );
buf ( n19441 , n18931 );
not ( n19442 , n19441 );
or ( n19443 , n19440 , n19442 );
buf ( n19444 , n18944 );
buf ( n19445 , n843 );
buf ( n19446 , n866 );
xor ( n19447 , n19445 , n19446 );
buf ( n19448 , n19447 );
buf ( n19449 , n19448 );
nand ( n19450 , n19444 , n19449 );
buf ( n19451 , n19450 );
buf ( n19452 , n19451 );
nand ( n19453 , n19443 , n19452 );
buf ( n19454 , n19453 );
buf ( n19455 , n19454 );
buf ( n19456 , n18903 );
not ( n19457 , n19456 );
buf ( n19458 , n18887 );
not ( n19459 , n19458 );
or ( n19460 , n19457 , n19459 );
buf ( n19461 , n18892 );
buf ( n19462 , n19461 );
buf ( n19463 , n841 );
buf ( n19464 , n868 );
xor ( n19465 , n19463 , n19464 );
buf ( n19466 , n19465 );
buf ( n19467 , n19466 );
nand ( n19468 , n19462 , n19467 );
buf ( n19469 , n19468 );
buf ( n19470 , n19469 );
nand ( n19471 , n19460 , n19470 );
buf ( n19472 , n19471 );
buf ( n19473 , n19472 );
xor ( n19474 , n19455 , n19473 );
buf ( n19475 , n19358 );
not ( n19476 , n19475 );
buf ( n19477 , n19259 );
buf ( n19478 , n19477 );
buf ( n19479 , n19478 );
buf ( n19480 , n19479 );
not ( n19481 , n19480 );
or ( n19482 , n19476 , n19481 );
buf ( n19483 , n19265 );
buf ( n19484 , n878 );
nand ( n19485 , n19483 , n19484 );
buf ( n19486 , n19485 );
buf ( n19487 , n19486 );
nand ( n19488 , n19482 , n19487 );
buf ( n19489 , n19488 );
buf ( n19490 , n19489 );
not ( n19491 , n19490 );
buf ( n19492 , n19491 );
buf ( n19493 , n19492 );
xor ( n19494 , n19474 , n19493 );
buf ( n19495 , n19494 );
buf ( n19496 , n19495 );
xor ( n19497 , n19438 , n19496 );
buf ( n19498 , n19139 );
not ( n19499 , n19498 );
buf ( n19500 , n19125 );
not ( n19501 , n19500 );
or ( n19502 , n19499 , n19501 );
buf ( n19503 , n19134 );
xor ( n19504 , n870 , n839 );
buf ( n19505 , n19504 );
nand ( n19506 , n19503 , n19505 );
buf ( n19507 , n19506 );
buf ( n19508 , n19507 );
nand ( n19509 , n19502 , n19508 );
buf ( n19510 , n19509 );
buf ( n19511 , n19510 );
buf ( n19512 , n19383 );
not ( n19513 , n19512 );
buf ( n19514 , n18977 );
not ( n19515 , n19514 );
or ( n19516 , n19513 , n19515 );
buf ( n19517 , n18987 );
xor ( n19518 , n874 , n835 );
buf ( n19519 , n19518 );
nand ( n19520 , n19517 , n19519 );
buf ( n19521 , n19520 );
buf ( n19522 , n19521 );
nand ( n19523 , n19516 , n19522 );
buf ( n19524 , n19523 );
buf ( n19525 , n19524 );
xor ( n19526 , n19511 , n19525 );
buf ( n19527 , n19090 );
not ( n19528 , n19527 );
buf ( n19529 , n19153 );
not ( n19530 , n19529 );
or ( n19531 , n19528 , n19530 );
buf ( n19532 , n19085 );
xor ( n19533 , n876 , n833 );
buf ( n19534 , n19533 );
nand ( n19535 , n19532 , n19534 );
buf ( n19536 , n19535 );
buf ( n19537 , n19536 );
nand ( n19538 , n19531 , n19537 );
buf ( n19539 , n19538 );
buf ( n19540 , n19539 );
xor ( n19541 , n19526 , n19540 );
buf ( n19542 , n19541 );
buf ( n19543 , n19542 );
xor ( n19544 , n19497 , n19543 );
buf ( n19545 , n19544 );
buf ( n19546 , n19545 );
xor ( n19547 , n19316 , n19326 );
xor ( n19548 , n19547 , n19342 );
buf ( n19549 , n19548 );
buf ( n19550 , n19549 );
xor ( n19551 , n19365 , n19372 );
xor ( n19552 , n19551 , n19390 );
buf ( n19553 , n19552 );
buf ( n19554 , n19553 );
xor ( n19555 , n19550 , n19554 );
xor ( n19556 , n18868 , n18910 );
xor ( n19557 , n19556 , n19051 );
buf ( n19558 , n19557 );
buf ( n19559 , n19558 );
and ( n19560 , n19555 , n19559 );
and ( n19561 , n19550 , n19554 );
or ( n19562 , n19560 , n19561 );
buf ( n19563 , n19562 );
buf ( n19564 , n19563 );
xor ( n19565 , n19546 , n19564 );
buf ( n19566 , n18867 );
not ( n19567 , n19566 );
xor ( n19568 , n883 , n884 );
not ( n19569 , n19568 );
buf ( n19570 , n19569 );
not ( n19571 , n19570 );
and ( n19572 , n883 , n882 );
not ( n19573 , n883 );
not ( n19574 , n882 );
and ( n19575 , n19573 , n19574 );
nor ( n19576 , n19572 , n19575 );
not ( n19577 , n19576 );
xor ( n19578 , n883 , n884 );
nor ( n19579 , n19577 , n19578 );
buf ( n19580 , n19579 );
buf ( n19581 , n19580 );
not ( n19582 , n19581 );
buf ( n19583 , n19582 );
buf ( n19584 , n19583 );
not ( n19585 , n19584 );
or ( n19586 , n19571 , n19585 );
buf ( n19587 , n882 );
nand ( n19588 , n19586 , n19587 );
buf ( n19589 , n19588 );
buf ( n19590 , n19589 );
buf ( n19591 , n837 );
buf ( n19592 , n876 );
xor ( n19593 , n19591 , n19592 );
buf ( n19594 , n19593 );
buf ( n19595 , n19594 );
not ( n19596 , n19595 );
buf ( n19597 , n19077 );
not ( n19598 , n19597 );
or ( n19599 , n19596 , n19598 );
buf ( n19600 , n19085 );
buf ( n19601 , n19150 );
nand ( n19602 , n19600 , n19601 );
buf ( n19603 , n19602 );
buf ( n19604 , n19603 );
nand ( n19605 , n19599 , n19604 );
buf ( n19606 , n19605 );
buf ( n19607 , n19606 );
xor ( n19608 , n19590 , n19607 );
xor ( n19609 , n880 , n833 );
buf ( n19610 , n19609 );
not ( n19611 , n19610 );
buf ( n19612 , n18850 );
buf ( n19613 , n19612 );
buf ( n19614 , n19613 );
buf ( n19615 , n19614 );
not ( n19616 , n19615 );
or ( n19617 , n19611 , n19616 );
buf ( n19618 , n18860 );
buf ( n19619 , n18838 );
nand ( n19620 , n19618 , n19619 );
buf ( n19621 , n19620 );
buf ( n19622 , n19621 );
nand ( n19623 , n19617 , n19622 );
buf ( n19624 , n19623 );
buf ( n19625 , n19624 );
and ( n19626 , n19608 , n19625 );
and ( n19627 , n19590 , n19607 );
or ( n19628 , n19626 , n19627 );
buf ( n19629 , n19628 );
buf ( n19630 , n19629 );
not ( n19631 , n19630 );
buf ( n19632 , n19631 );
buf ( n19633 , n19632 );
not ( n19634 , n19633 );
or ( n19635 , n19567 , n19634 );
xor ( n19636 , n868 , n845 );
buf ( n19637 , n19636 );
not ( n19638 , n19637 );
buf ( n19639 , n18887 );
not ( n19640 , n19639 );
or ( n19641 , n19638 , n19640 );
buf ( n19642 , n18892 );
buf ( n19643 , n19168 );
nand ( n19644 , n19642 , n19643 );
buf ( n19645 , n19644 );
buf ( n19646 , n19645 );
nand ( n19647 , n19641 , n19646 );
buf ( n19648 , n19647 );
buf ( n19649 , n19648 );
not ( n19650 , n19649 );
buf ( n19651 , n847 );
buf ( n19652 , n866 );
xor ( n19653 , n19651 , n19652 );
buf ( n19654 , n19653 );
buf ( n19655 , n19654 );
not ( n19656 , n19655 );
buf ( n19657 , n18931 );
not ( n19658 , n19657 );
or ( n19659 , n19656 , n19658 );
buf ( n19660 , n18944 );
buf ( n19661 , n18915 );
nand ( n19662 , n19660 , n19661 );
buf ( n19663 , n19662 );
buf ( n19664 , n19663 );
nand ( n19665 , n19659 , n19664 );
buf ( n19666 , n19665 );
buf ( n19667 , n19666 );
not ( n19668 , n19667 );
or ( n19669 , n19650 , n19668 );
buf ( n19670 , n19648 );
not ( n19671 , n19670 );
buf ( n19672 , n19671 );
buf ( n19673 , n19672 );
not ( n19674 , n19673 );
buf ( n19675 , n19666 );
not ( n19676 , n19675 );
buf ( n19677 , n19676 );
buf ( n19678 , n19677 );
not ( n19679 , n19678 );
or ( n19680 , n19674 , n19679 );
buf ( n19681 , n839 );
buf ( n19682 , n874 );
xor ( n19683 , n19681 , n19682 );
buf ( n19684 , n19683 );
buf ( n19685 , n19684 );
not ( n19686 , n19685 );
buf ( n19687 , n18977 );
not ( n19688 , n19687 );
or ( n19689 , n19686 , n19688 );
buf ( n19690 , n18987 );
buf ( n19691 , n18960 );
nand ( n19692 , n19690 , n19691 );
buf ( n19693 , n19692 );
buf ( n19694 , n19693 );
nand ( n19695 , n19689 , n19694 );
buf ( n19696 , n19695 );
buf ( n19697 , n19696 );
nand ( n19698 , n19680 , n19697 );
buf ( n19699 , n19698 );
buf ( n19700 , n19699 );
nand ( n19701 , n19669 , n19700 );
buf ( n19702 , n19701 );
buf ( n19703 , n19702 );
nand ( n19704 , n19635 , n19703 );
buf ( n19705 , n19704 );
buf ( n19706 , n19705 );
buf ( n19707 , n18867 );
not ( n19708 , n19707 );
buf ( n19709 , n19629 );
nand ( n19710 , n19708 , n19709 );
buf ( n19711 , n19710 );
buf ( n19712 , n19711 );
nand ( n19713 , n19706 , n19712 );
buf ( n19714 , n19713 );
buf ( n19715 , n19714 );
xor ( n19716 , n19214 , n19246 );
xor ( n19717 , n19716 , n19276 );
not ( n19718 , n19717 );
not ( n19719 , n19718 );
xor ( n19720 , n18956 , n18999 );
xor ( n19721 , n19720 , n19046 );
buf ( n19722 , n19721 );
not ( n19723 , n19722 );
not ( n19724 , n19723 );
or ( n19725 , n19719 , n19724 );
and ( n19726 , n850 , n864 );
buf ( n19727 , n849 );
buf ( n19728 , n864 );
xor ( n19729 , n19727 , n19728 );
buf ( n19730 , n19729 );
not ( n19731 , n19730 );
not ( n19732 , n19013 );
or ( n19733 , n19731 , n19732 );
buf ( n19734 , n19021 );
not ( n19735 , n19734 );
buf ( n19736 , n19030 );
nand ( n19737 , n19735 , n19736 );
buf ( n19738 , n19737 );
nand ( n19739 , n19733 , n19738 );
xor ( n19740 , n19726 , n19739 );
not ( n19741 , n19479 );
buf ( n19742 , n835 );
buf ( n19743 , n878 );
xor ( n19744 , n19742 , n19743 );
buf ( n19745 , n19744 );
not ( n19746 , n19745 );
or ( n19747 , n19741 , n19746 );
buf ( n19748 , n19265 );
buf ( n19749 , n19251 );
nand ( n19750 , n19748 , n19749 );
buf ( n19751 , n19750 );
nand ( n19752 , n19747 , n19751 );
and ( n19753 , n19740 , n19752 );
and ( n19754 , n19726 , n19739 );
or ( n19755 , n19753 , n19754 );
nand ( n19756 , n19725 , n19755 );
not ( n19757 , n19723 );
nand ( n19758 , n19757 , n19717 );
nand ( n19759 , n19756 , n19758 );
buf ( n19760 , n19759 );
xor ( n19761 , n19715 , n19760 );
nand ( n19762 , n19209 , n19146 , n19279 );
not ( n19763 , n19209 );
xor ( n19764 , n19061 , n19097 );
xnor ( n19765 , n19764 , n19145 );
nand ( n19766 , n19763 , n19765 , n19279 );
nor ( n19767 , n19765 , n19279 );
nand ( n19768 , n19767 , n19763 );
not ( n19769 , n19279 );
nand ( n19770 , n19769 , n19209 , n19765 );
nand ( n19771 , n19762 , n19766 , n19768 , n19770 );
buf ( n19772 , n19771 );
and ( n19773 , n19761 , n19772 );
and ( n19774 , n19715 , n19760 );
or ( n19775 , n19773 , n19774 );
buf ( n19776 , n19775 );
buf ( n19777 , n19776 );
xor ( n19778 , n19565 , n19777 );
buf ( n19779 , n19778 );
buf ( n19780 , n19779 );
xor ( n19781 , n19401 , n19780 );
xor ( n19782 , n19550 , n19554 );
xor ( n19783 , n19782 , n19559 );
buf ( n19784 , n19783 );
buf ( n19785 , n19784 );
buf ( n19786 , n19614 );
buf ( n19787 , n834 );
buf ( n19788 , n880 );
xor ( n19789 , n19787 , n19788 );
buf ( n19790 , n19789 );
buf ( n19791 , n19790 );
and ( n19792 , n19786 , n19791 );
buf ( n19793 , n18860 );
buf ( n19794 , n19609 );
and ( n19795 , n19793 , n19794 );
nor ( n19796 , n19792 , n19795 );
buf ( n19797 , n19796 );
buf ( n19798 , n19797 );
not ( n19799 , n19798 );
buf ( n19800 , n19799 );
buf ( n19801 , n19800 );
xor ( n19802 , n870 , n843 );
buf ( n19803 , n19802 );
not ( n19804 , n19803 );
buf ( n19805 , n19125 );
not ( n19806 , n19805 );
or ( n19807 , n19804 , n19806 );
buf ( n19808 , n19134 );
buf ( n19809 , n19190 );
nand ( n19810 , n19808 , n19809 );
buf ( n19811 , n19810 );
buf ( n19812 , n19811 );
nand ( n19813 , n19807 , n19812 );
buf ( n19814 , n19813 );
buf ( n19815 , n19814 );
xor ( n19816 , n19801 , n19815 );
buf ( n19817 , n841 );
buf ( n19818 , n872 );
xor ( n19819 , n19817 , n19818 );
buf ( n19820 , n19819 );
buf ( n19821 , n19820 );
not ( n19822 , n19821 );
buf ( n19823 , n19230 );
not ( n19824 , n19823 );
or ( n19825 , n19822 , n19824 );
buf ( n19826 , n19235 );
buf ( n19827 , n19218 );
nand ( n19828 , n19826 , n19827 );
buf ( n19829 , n19828 );
buf ( n19830 , n19829 );
nand ( n19831 , n19825 , n19830 );
buf ( n19832 , n19831 );
buf ( n19833 , n19832 );
and ( n19834 , n19816 , n19833 );
and ( n19835 , n19801 , n19815 );
or ( n19836 , n19834 , n19835 );
buf ( n19837 , n19836 );
buf ( n19838 , n19837 );
xor ( n19839 , n19184 , n19163 );
xnor ( n19840 , n19839 , n19202 );
buf ( n19841 , n19840 );
xor ( n19842 , n19838 , n19841 );
buf ( n19843 , n848 );
buf ( n19844 , n866 );
xor ( n19845 , n19843 , n19844 );
buf ( n19846 , n19845 );
buf ( n19847 , n19846 );
not ( n19848 , n19847 );
buf ( n19849 , n18931 );
not ( n19850 , n19849 );
or ( n19851 , n19848 , n19850 );
buf ( n19852 , n18944 );
buf ( n19853 , n19654 );
nand ( n19854 , n19852 , n19853 );
buf ( n19855 , n19854 );
buf ( n19856 , n19855 );
nand ( n19857 , n19851 , n19856 );
buf ( n19858 , n19857 );
buf ( n19859 , n19858 );
xor ( n19860 , n868 , n846 );
buf ( n19861 , n19860 );
not ( n19862 , n19861 );
buf ( n19863 , n18887 );
not ( n19864 , n19863 );
or ( n19865 , n19862 , n19864 );
buf ( n19866 , n19461 );
buf ( n19867 , n19636 );
nand ( n19868 , n19866 , n19867 );
buf ( n19869 , n19868 );
buf ( n19870 , n19869 );
nand ( n19871 , n19865 , n19870 );
buf ( n19872 , n19871 );
buf ( n19873 , n19872 );
xor ( n19874 , n19859 , n19873 );
xor ( n19875 , n876 , n838 );
buf ( n19876 , n19875 );
not ( n19877 , n19876 );
buf ( n19878 , n19153 );
not ( n19879 , n19878 );
or ( n19880 , n19877 , n19879 );
buf ( n19881 , n19085 );
buf ( n19882 , n19594 );
nand ( n19883 , n19881 , n19882 );
buf ( n19884 , n19883 );
buf ( n19885 , n19884 );
nand ( n19886 , n19880 , n19885 );
buf ( n19887 , n19886 );
buf ( n19888 , n19887 );
and ( n19889 , n19874 , n19888 );
and ( n19890 , n19859 , n19873 );
or ( n19891 , n19889 , n19890 );
buf ( n19892 , n19891 );
buf ( n19893 , n19892 );
buf ( n19894 , n832 );
buf ( n19895 , n882 );
xor ( n19896 , n19894 , n19895 );
buf ( n19897 , n19896 );
buf ( n19898 , n19897 );
not ( n19899 , n19898 );
buf ( n19900 , n19580 );
not ( n19901 , n19900 );
or ( n19902 , n19899 , n19901 );
not ( n19903 , n883 );
not ( n19904 , n884 );
not ( n19905 , n19904 );
or ( n19906 , n19903 , n19905 );
not ( n19907 , n883 );
nand ( n19908 , n19907 , n884 );
nand ( n19909 , n19906 , n19908 );
buf ( n19910 , n19909 );
buf ( n19911 , n19910 );
buf ( n19912 , n882 );
nand ( n19913 , n19911 , n19912 );
buf ( n19914 , n19913 );
buf ( n19915 , n19914 );
nand ( n19916 , n19902 , n19915 );
buf ( n19917 , n19916 );
buf ( n19918 , n19917 );
buf ( n19919 , n842 );
buf ( n19920 , n872 );
xor ( n19921 , n19919 , n19920 );
buf ( n19922 , n19921 );
buf ( n19923 , n19922 );
not ( n19924 , n19923 );
buf ( n19925 , n19230 );
not ( n19926 , n19925 );
or ( n19927 , n19924 , n19926 );
buf ( n19928 , n19235 );
buf ( n19929 , n19820 );
nand ( n19930 , n19928 , n19929 );
buf ( n19931 , n19930 );
buf ( n19932 , n19931 );
nand ( n19933 , n19927 , n19932 );
buf ( n19934 , n19933 );
buf ( n19935 , n19934 );
xor ( n19936 , n19918 , n19935 );
buf ( n19937 , n836 );
buf ( n19938 , n878 );
xor ( n19939 , n19937 , n19938 );
buf ( n19940 , n19939 );
buf ( n19941 , n19940 );
not ( n19942 , n19941 );
buf ( n19943 , n19479 );
not ( n19944 , n19943 );
or ( n19945 , n19942 , n19944 );
buf ( n19946 , n19265 );
buf ( n19947 , n19745 );
nand ( n19948 , n19946 , n19947 );
buf ( n19949 , n19948 );
buf ( n19950 , n19949 );
nand ( n19951 , n19945 , n19950 );
buf ( n19952 , n19951 );
buf ( n19953 , n19952 );
and ( n19954 , n19936 , n19953 );
and ( n19955 , n19918 , n19935 );
or ( n19956 , n19954 , n19955 );
buf ( n19957 , n19956 );
buf ( n19958 , n19957 );
xor ( n19959 , n19893 , n19958 );
buf ( n19960 , n851 );
buf ( n19961 , n864 );
and ( n19962 , n19960 , n19961 );
buf ( n19963 , n19962 );
buf ( n19964 , n19963 );
buf ( n19965 , n850 );
buf ( n19966 , n864 );
xor ( n19967 , n19965 , n19966 );
buf ( n19968 , n19967 );
buf ( n19969 , n19968 );
not ( n19970 , n19969 );
buf ( n19971 , n19013 );
not ( n19972 , n19971 );
or ( n19973 , n19970 , n19972 );
buf ( n19974 , n19030 );
buf ( n19975 , n19730 );
nand ( n19976 , n19974 , n19975 );
buf ( n19977 , n19976 );
buf ( n19978 , n19977 );
nand ( n19979 , n19973 , n19978 );
buf ( n19980 , n19979 );
buf ( n19981 , n19980 );
xor ( n19982 , n19964 , n19981 );
buf ( n19983 , n840 );
buf ( n19984 , n874 );
xor ( n19985 , n19983 , n19984 );
buf ( n19986 , n19985 );
buf ( n19987 , n19986 );
not ( n19988 , n19987 );
buf ( n19989 , n18977 );
not ( n19990 , n19989 );
or ( n19991 , n19988 , n19990 );
buf ( n19992 , n18987 );
buf ( n19993 , n19684 );
nand ( n19994 , n19992 , n19993 );
buf ( n19995 , n19994 );
buf ( n19996 , n19995 );
nand ( n19997 , n19991 , n19996 );
buf ( n19998 , n19997 );
buf ( n19999 , n19998 );
and ( n20000 , n19982 , n19999 );
and ( n20001 , n19964 , n19981 );
or ( n20002 , n20000 , n20001 );
buf ( n20003 , n20002 );
buf ( n20004 , n20003 );
and ( n20005 , n19959 , n20004 );
and ( n20006 , n19893 , n19958 );
or ( n20007 , n20005 , n20006 );
buf ( n20008 , n20007 );
buf ( n20009 , n20008 );
and ( n20010 , n19842 , n20009 );
and ( n20011 , n19838 , n19841 );
or ( n20012 , n20010 , n20011 );
buf ( n20013 , n20012 );
buf ( n20014 , n20013 );
xor ( n20015 , n19785 , n20014 );
xor ( n20016 , n19726 , n19739 );
xor ( n20017 , n20016 , n19752 );
xor ( n20018 , n19590 , n19607 );
xor ( n20019 , n20018 , n19625 );
buf ( n20020 , n20019 );
xor ( n20021 , n20017 , n20020 );
buf ( n20022 , n19696 );
not ( n20023 , n20022 );
buf ( n20024 , n19672 );
not ( n20025 , n20024 );
buf ( n20026 , n19666 );
not ( n20027 , n20026 );
and ( n20028 , n20025 , n20027 );
buf ( n20029 , n19666 );
buf ( n20030 , n19672 );
and ( n20031 , n20029 , n20030 );
nor ( n20032 , n20028 , n20031 );
buf ( n20033 , n20032 );
buf ( n20034 , n20033 );
not ( n20035 , n20034 );
or ( n20036 , n20023 , n20035 );
buf ( n20037 , n20033 );
buf ( n20038 , n19696 );
or ( n20039 , n20037 , n20038 );
nand ( n20040 , n20036 , n20039 );
buf ( n20041 , n20040 );
and ( n20042 , n20021 , n20041 );
and ( n20043 , n20017 , n20020 );
or ( n20044 , n20042 , n20043 );
buf ( n20045 , n20044 );
and ( n20046 , n19755 , n19717 );
not ( n20047 , n19755 );
and ( n20048 , n20047 , n19718 );
nor ( n20049 , n20046 , n20048 );
and ( n20050 , n20049 , n19757 );
not ( n20051 , n20049 );
and ( n20052 , n20051 , n19723 );
nor ( n20053 , n20050 , n20052 );
buf ( n20054 , n20053 );
or ( n20055 , n20045 , n20054 );
buf ( n20056 , n19702 );
not ( n20057 , n20056 );
buf ( n20058 , n18867 );
not ( n20059 , n20058 );
and ( n20060 , n20057 , n20059 );
buf ( n20061 , n19702 );
buf ( n20062 , n18867 );
and ( n20063 , n20061 , n20062 );
nor ( n20064 , n20060 , n20063 );
buf ( n20065 , n20064 );
buf ( n20066 , n20065 );
buf ( n20067 , n19629 );
and ( n20068 , n20066 , n20067 );
not ( n20069 , n20066 );
buf ( n20070 , n19632 );
and ( n20071 , n20069 , n20070 );
nor ( n20072 , n20068 , n20071 );
buf ( n20073 , n20072 );
buf ( n20074 , n20073 );
not ( n20075 , n20074 );
buf ( n20076 , n20075 );
buf ( n20077 , n20076 );
nand ( n20078 , n20055 , n20077 );
buf ( n20079 , n20078 );
buf ( n20080 , n20079 );
buf ( n20081 , n20053 );
buf ( n20082 , n20044 );
nand ( n20083 , n20081 , n20082 );
buf ( n20084 , n20083 );
buf ( n20085 , n20084 );
nand ( n20086 , n20080 , n20085 );
buf ( n20087 , n20086 );
buf ( n20088 , n20087 );
and ( n20089 , n20015 , n20088 );
and ( n20090 , n19785 , n20014 );
or ( n20091 , n20089 , n20090 );
buf ( n20092 , n20091 );
buf ( n20093 , n20092 );
xor ( n20094 , n19781 , n20093 );
buf ( n20095 , n20094 );
buf ( n20096 , n20095 );
buf ( n20097 , n894 );
buf ( n20098 , n859 );
buf ( n20099 , n866 );
xor ( n20100 , n20098 , n20099 );
buf ( n20101 , n20100 );
buf ( n20102 , n20101 );
not ( n20103 , n20102 );
buf ( n20104 , n18931 );
not ( n20105 , n20104 );
or ( n20106 , n20103 , n20105 );
buf ( n20107 , n18944 );
buf ( n20108 , n858 );
buf ( n20109 , n866 );
xor ( n20110 , n20108 , n20109 );
buf ( n20111 , n20110 );
buf ( n20112 , n20111 );
nand ( n20113 , n20107 , n20112 );
buf ( n20114 , n20113 );
buf ( n20115 , n20114 );
nand ( n20116 , n20106 , n20115 );
buf ( n20117 , n20116 );
buf ( n20118 , n20117 );
xor ( n20119 , n20097 , n20118 );
buf ( n20120 , n863 );
buf ( n20121 , n864 );
and ( n20122 , n20120 , n20121 );
buf ( n20123 , n20122 );
buf ( n20124 , n20123 );
and ( n20125 , n832 , n894 );
not ( n20126 , n832 );
not ( n20127 , n894 );
and ( n20128 , n20126 , n20127 );
nor ( n20129 , n20125 , n20128 );
not ( n20130 , n20129 );
not ( n20131 , n894 );
nor ( n20132 , n20131 , n895 );
not ( n20133 , n20132 );
or ( n20134 , n20130 , n20133 );
nand ( n20135 , n894 , n895 );
nand ( n20136 , n20134 , n20135 );
buf ( n20137 , n20136 );
xor ( n20138 , n20124 , n20137 );
buf ( n20139 , n834 );
buf ( n20140 , n892 );
xor ( n20141 , n20139 , n20140 );
buf ( n20142 , n20141 );
buf ( n20143 , n20142 );
not ( n20144 , n20143 );
and ( n20145 , n893 , n20127 );
not ( n20146 , n893 );
and ( n20147 , n20146 , n894 );
nor ( n20148 , n20145 , n20147 );
not ( n20149 , n892 );
not ( n20150 , n893 );
not ( n20151 , n20150 );
or ( n20152 , n20149 , n20151 );
not ( n20153 , n892 );
nand ( n20154 , n20153 , n893 );
nand ( n20155 , n20152 , n20154 );
nand ( n20156 , n20148 , n20155 );
buf ( n20157 , n20156 );
not ( n20158 , n20157 );
buf ( n20159 , n20158 );
buf ( n20160 , n20159 );
not ( n20161 , n20160 );
or ( n20162 , n20144 , n20161 );
xor ( n20163 , n893 , n894 );
not ( n20164 , n20163 );
buf ( n20165 , n20164 );
not ( n20166 , n20165 );
buf ( n20167 , n20166 );
buf ( n20168 , n20167 );
xor ( n20169 , n892 , n833 );
buf ( n20170 , n20169 );
nand ( n20171 , n20168 , n20170 );
buf ( n20172 , n20171 );
buf ( n20173 , n20172 );
nand ( n20174 , n20162 , n20173 );
buf ( n20175 , n20174 );
buf ( n20176 , n20175 );
and ( n20177 , n20138 , n20176 );
and ( n20178 , n20124 , n20137 );
or ( n20179 , n20177 , n20178 );
buf ( n20180 , n20179 );
buf ( n20181 , n20180 );
and ( n20182 , n20119 , n20181 );
and ( n20183 , n20097 , n20118 );
or ( n20184 , n20182 , n20183 );
buf ( n20185 , n20184 );
buf ( n20186 , n20185 );
not ( n20187 , n20186 );
xor ( n20188 , n882 , n844 );
not ( n20189 , n20188 );
buf ( n20190 , n882 );
buf ( n20191 , n883 );
xnor ( n20192 , n20190 , n20191 );
buf ( n20193 , n20192 );
buf ( n20194 , n20193 );
buf ( n20195 , n19568 );
nor ( n20196 , n20194 , n20195 );
buf ( n20197 , n20196 );
not ( n20198 , n20197 );
or ( n20199 , n20189 , n20198 );
buf ( n20200 , n19568 );
xor ( n20201 , n882 , n843 );
buf ( n20202 , n20201 );
nand ( n20203 , n20200 , n20202 );
buf ( n20204 , n20203 );
nand ( n20205 , n20199 , n20204 );
not ( n20206 , n20205 );
xor ( n20207 , n872 , n854 );
not ( n20208 , n20207 );
xnor ( n20209 , n873 , n874 );
nand ( n20210 , n20209 , n19228 );
not ( n20211 , n20210 );
not ( n20212 , n20211 );
or ( n20213 , n20208 , n20212 );
buf ( n20214 , n19234 );
xor ( n20215 , n872 , n853 );
buf ( n20216 , n20215 );
nand ( n20217 , n20214 , n20216 );
buf ( n20218 , n20217 );
nand ( n20219 , n20213 , n20218 );
not ( n20220 , n20219 );
or ( n20221 , n20206 , n20220 );
or ( n20222 , n20219 , n20205 );
and ( n20223 , n871 , n872 );
not ( n20224 , n871 );
and ( n20225 , n20224 , n19106 );
nor ( n20226 , n20223 , n20225 );
not ( n20227 , n20226 );
buf ( n20228 , n855 );
buf ( n20229 , n870 );
xor ( n20230 , n20228 , n20229 );
buf ( n20231 , n20230 );
not ( n20232 , n20231 );
or ( n20233 , n20227 , n20232 );
not ( n20234 , n20226 );
not ( n20235 , n19116 );
xor ( n20236 , n856 , n870 );
nand ( n20237 , n20234 , n20235 , n20236 );
nand ( n20238 , n20233 , n20237 );
nand ( n20239 , n20222 , n20238 );
nand ( n20240 , n20221 , n20239 );
xor ( n20241 , n876 , n850 );
not ( n20242 , n20241 );
not ( n20243 , n19075 );
not ( n20244 , n20243 );
or ( n20245 , n20242 , n20244 );
buf ( n20246 , n19081 );
buf ( n20247 , n20246 );
xor ( n20248 , n876 , n849 );
buf ( n20249 , n20248 );
nand ( n20250 , n20247 , n20249 );
buf ( n20251 , n20250 );
nand ( n20252 , n20245 , n20251 );
buf ( n20253 , n20252 );
not ( n20254 , n20253 );
xor ( n20255 , n887 , n888 );
not ( n20256 , n20255 );
xor ( n20257 , n886 , n839 );
not ( n20258 , n20257 );
or ( n20259 , n20256 , n20258 );
xor ( n20260 , n887 , n888 );
not ( n20261 , n20260 );
xor ( n20262 , n887 , n886 );
and ( n20263 , n840 , n886 );
not ( n20264 , n840 );
not ( n20265 , n886 );
and ( n20266 , n20264 , n20265 );
nor ( n20267 , n20263 , n20266 );
nand ( n20268 , n20261 , n20262 , n20267 );
nand ( n20269 , n20259 , n20268 );
buf ( n20270 , n20269 );
not ( n20271 , n20270 );
or ( n20272 , n20254 , n20271 );
buf ( n20273 , n20269 );
buf ( n20274 , n20252 );
or ( n20275 , n20273 , n20274 );
buf ( n20276 , n847 );
buf ( n20277 , n878 );
xor ( n20278 , n20276 , n20277 );
buf ( n20279 , n20278 );
not ( n20280 , n20279 );
not ( n20281 , n19265 );
or ( n20282 , n20280 , n20281 );
buf ( n20283 , n848 );
buf ( n20284 , n878 );
xor ( n20285 , n20283 , n20284 );
buf ( n20286 , n20285 );
nand ( n20287 , n20286 , n19256 );
nand ( n20288 , n20282 , n20287 );
buf ( n20289 , n20288 );
nand ( n20290 , n20275 , n20289 );
buf ( n20291 , n20290 );
buf ( n20292 , n20291 );
nand ( n20293 , n20272 , n20292 );
buf ( n20294 , n20293 );
xor ( n20295 , n20240 , n20294 );
buf ( n20296 , n862 );
buf ( n20297 , n864 );
xor ( n20298 , n20296 , n20297 );
buf ( n20299 , n20298 );
buf ( n20300 , n20299 );
not ( n20301 , n20300 );
not ( n20302 , n19012 );
buf ( n20303 , n20302 );
not ( n20304 , n20303 );
or ( n20305 , n20301 , n20304 );
xor ( n20306 , n861 , n864 );
nand ( n20307 , n19027 , n20306 );
buf ( n20308 , n20307 );
nand ( n20309 , n20305 , n20308 );
buf ( n20310 , n20309 );
buf ( n20311 , n20310 );
not ( n20312 , n20311 );
buf ( n20313 , n20312 );
buf ( n20314 , n20313 );
not ( n20315 , n20314 );
buf ( n20316 , n846 );
buf ( n20317 , n880 );
xor ( n20318 , n20316 , n20317 );
buf ( n20319 , n20318 );
buf ( n20320 , n20319 );
not ( n20321 , n20320 );
buf ( n20322 , n18850 );
not ( n20323 , n20322 );
or ( n20324 , n20321 , n20323 );
xor ( n20325 , n881 , n882 );
buf ( n20326 , n20325 );
buf ( n20327 , n845 );
buf ( n20328 , n880 );
xor ( n20329 , n20327 , n20328 );
buf ( n20330 , n20329 );
buf ( n20331 , n20330 );
nand ( n20332 , n20326 , n20331 );
buf ( n20333 , n20332 );
buf ( n20334 , n20333 );
nand ( n20335 , n20324 , n20334 );
buf ( n20336 , n20335 );
buf ( n20337 , n20336 );
not ( n20338 , n20337 );
buf ( n20339 , n20338 );
buf ( n20340 , n20339 );
not ( n20341 , n20340 );
or ( n20342 , n20315 , n20341 );
buf ( n20343 , n838 );
buf ( n20344 , n888 );
xor ( n20345 , n20343 , n20344 );
buf ( n20346 , n20345 );
buf ( n20347 , n20346 );
not ( n20348 , n20347 );
not ( n20349 , n888 );
not ( n20350 , n20349 );
nand ( n20351 , n889 , n890 );
not ( n20352 , n20351 );
not ( n20353 , n20352 );
or ( n20354 , n20350 , n20353 );
nor ( n20355 , n889 , n890 );
nand ( n20356 , n888 , n20355 );
nand ( n20357 , n20354 , n20356 );
buf ( n20358 , n20357 );
buf ( n20359 , n20358 );
not ( n20360 , n20359 );
or ( n20361 , n20348 , n20360 );
xor ( n20362 , n889 , n890 );
buf ( n20363 , n20362 );
buf ( n20364 , n20363 );
xor ( n20365 , n888 , n837 );
buf ( n20366 , n20365 );
nand ( n20367 , n20364 , n20366 );
buf ( n20368 , n20367 );
buf ( n20369 , n20368 );
nand ( n20370 , n20361 , n20369 );
buf ( n20371 , n20370 );
buf ( n20372 , n20371 );
nand ( n20373 , n20342 , n20372 );
buf ( n20374 , n20373 );
buf ( n20375 , n20374 );
buf ( n20376 , n20310 );
buf ( n20377 , n20336 );
nand ( n20378 , n20376 , n20377 );
buf ( n20379 , n20378 );
buf ( n20380 , n20379 );
nand ( n20381 , n20375 , n20380 );
buf ( n20382 , n20381 );
and ( n20383 , n20295 , n20382 );
and ( n20384 , n20240 , n20294 );
or ( n20385 , n20383 , n20384 );
not ( n20386 , n20385 );
not ( n20387 , n20386 );
buf ( n20388 , n20387 );
not ( n20389 , n20388 );
or ( n20390 , n20187 , n20389 );
buf ( n20391 , n20185 );
not ( n20392 , n20391 );
buf ( n20393 , n20392 );
buf ( n20394 , n20393 );
not ( n20395 , n20394 );
buf ( n20396 , n20386 );
not ( n20397 , n20396 );
or ( n20398 , n20395 , n20397 );
xor ( n20399 , n890 , n835 );
buf ( n20400 , n20399 );
not ( n20401 , n20400 );
xnor ( n20402 , n891 , n890 );
xor ( n20403 , n891 , n892 );
nor ( n20404 , n20402 , n20403 );
buf ( n20405 , n20404 );
not ( n20406 , n20405 );
or ( n20407 , n20401 , n20406 );
xor ( n20408 , n890 , n834 );
buf ( n20409 , n20408 );
buf ( n20410 , n20403 );
nand ( n20411 , n20409 , n20410 );
buf ( n20412 , n20411 );
buf ( n20413 , n20412 );
nand ( n20414 , n20407 , n20413 );
buf ( n20415 , n20414 );
buf ( n20416 , n20415 );
xor ( n20417 , n884 , n841 );
buf ( n20418 , n20417 );
not ( n20419 , n20418 );
buf ( n20420 , n885 );
buf ( n20421 , n886 );
xor ( n20422 , n20420 , n20421 );
buf ( n20423 , n20422 );
and ( n20424 , n885 , n884 );
not ( n20425 , n885 );
not ( n20426 , n884 );
and ( n20427 , n20425 , n20426 );
nor ( n20428 , n20424 , n20427 );
not ( n20429 , n20428 );
nor ( n20430 , n20423 , n20429 );
buf ( n20431 , n20430 );
not ( n20432 , n20431 );
or ( n20433 , n20419 , n20432 );
buf ( n20434 , n20423 );
xor ( n20435 , n884 , n840 );
buf ( n20436 , n20435 );
nand ( n20437 , n20434 , n20436 );
buf ( n20438 , n20437 );
buf ( n20439 , n20438 );
nand ( n20440 , n20433 , n20439 );
buf ( n20441 , n20440 );
buf ( n20442 , n20441 );
or ( n20443 , n20416 , n20442 );
buf ( n20444 , n20215 );
not ( n20445 , n20444 );
buf ( n20446 , n20211 );
not ( n20447 , n20446 );
or ( n20448 , n20445 , n20447 );
buf ( n20449 , n19234 );
buf ( n20450 , n852 );
buf ( n20451 , n872 );
xor ( n20452 , n20450 , n20451 );
buf ( n20453 , n20452 );
buf ( n20454 , n20453 );
nand ( n20455 , n20449 , n20454 );
buf ( n20456 , n20455 );
buf ( n20457 , n20456 );
nand ( n20458 , n20448 , n20457 );
buf ( n20459 , n20458 );
buf ( n20460 , n20459 );
nand ( n20461 , n20443 , n20460 );
buf ( n20462 , n20461 );
buf ( n20463 , n20462 );
buf ( n20464 , n20415 );
buf ( n20465 , n20441 );
nand ( n20466 , n20464 , n20465 );
buf ( n20467 , n20466 );
buf ( n20468 , n20467 );
nand ( n20469 , n20463 , n20468 );
buf ( n20470 , n20469 );
buf ( n20471 , n20470 );
buf ( n20472 , n20169 );
not ( n20473 , n20472 );
buf ( n20474 , n20159 );
not ( n20475 , n20474 );
or ( n20476 , n20473 , n20475 );
buf ( n20477 , n20167 );
xor ( n20478 , n892 , n832 );
buf ( n20479 , n20478 );
nand ( n20480 , n20477 , n20479 );
buf ( n20481 , n20480 );
buf ( n20482 , n20481 );
nand ( n20483 , n20476 , n20482 );
buf ( n20484 , n20483 );
buf ( n20485 , n20365 );
not ( n20486 , n20485 );
buf ( n20487 , n20358 );
not ( n20488 , n20487 );
or ( n20489 , n20486 , n20488 );
buf ( n20490 , n20363 );
buf ( n20491 , n836 );
buf ( n20492 , n888 );
xor ( n20493 , n20491 , n20492 );
buf ( n20494 , n20493 );
buf ( n20495 , n20494 );
nand ( n20496 , n20490 , n20495 );
buf ( n20497 , n20496 );
buf ( n20498 , n20497 );
nand ( n20499 , n20489 , n20498 );
buf ( n20500 , n20499 );
xor ( n20501 , n20484 , n20500 );
buf ( n20502 , n20279 );
not ( n20503 , n20502 );
buf ( n20504 , n19259 );
not ( n20505 , n20504 );
or ( n20506 , n20503 , n20505 );
xnor ( n20507 , n878 , n846 );
not ( n20508 , n20507 );
nand ( n20509 , n20508 , n19265 );
buf ( n20510 , n20509 );
nand ( n20511 , n20506 , n20510 );
buf ( n20512 , n20511 );
and ( n20513 , n20501 , n20512 );
and ( n20514 , n20484 , n20500 );
or ( n20515 , n20513 , n20514 );
buf ( n20516 , n20515 );
xor ( n20517 , n20471 , n20516 );
buf ( n20518 , n20257 );
not ( n20519 , n20518 );
nand ( n20520 , n20261 , n20262 );
not ( n20521 , n20520 );
buf ( n20522 , n20521 );
not ( n20523 , n20522 );
or ( n20524 , n20519 , n20523 );
buf ( n20525 , n20255 );
buf ( n20526 , n20525 );
buf ( n20527 , n838 );
buf ( n20528 , n886 );
xor ( n20529 , n20527 , n20528 );
buf ( n20530 , n20529 );
buf ( n20531 , n20530 );
nand ( n20532 , n20526 , n20531 );
buf ( n20533 , n20532 );
buf ( n20534 , n20533 );
nand ( n20535 , n20524 , n20534 );
buf ( n20536 , n20535 );
not ( n20537 , n20536 );
buf ( n20538 , n851 );
buf ( n20539 , n874 );
xor ( n20540 , n20538 , n20539 );
buf ( n20541 , n20540 );
buf ( n20542 , n20541 );
not ( n20543 , n20542 );
buf ( n20544 , n876 );
not ( n20545 , n20544 );
buf ( n20546 , n875 );
nand ( n20547 , n20545 , n20546 );
buf ( n20548 , n20547 );
and ( n20549 , n20548 , n18967 , n18973 );
buf ( n20550 , n20549 );
not ( n20551 , n20550 );
or ( n20552 , n20543 , n20551 );
buf ( n20553 , n18984 );
not ( n20554 , n20553 );
buf ( n20555 , n20554 );
buf ( n20556 , n20555 );
xor ( n20557 , n874 , n850 );
buf ( n20558 , n20557 );
nand ( n20559 , n20556 , n20558 );
buf ( n20560 , n20559 );
buf ( n20561 , n20560 );
nand ( n20562 , n20552 , n20561 );
buf ( n20563 , n20562 );
not ( n20564 , n20563 );
buf ( n20565 , n20248 );
not ( n20566 , n20565 );
buf ( n20567 , n19153 );
not ( n20568 , n20567 );
or ( n20569 , n20566 , n20568 );
buf ( n20570 , n19082 );
xor ( n20571 , n876 , n848 );
buf ( n20572 , n20571 );
nand ( n20573 , n20570 , n20572 );
buf ( n20574 , n20573 );
buf ( n20575 , n20574 );
nand ( n20576 , n20569 , n20575 );
buf ( n20577 , n20576 );
not ( n20578 , n20577 );
nand ( n20579 , n20564 , n20578 );
not ( n20580 , n20579 );
or ( n20581 , n20537 , n20580 );
nand ( n20582 , n20577 , n20563 );
nand ( n20583 , n20581 , n20582 );
buf ( n20584 , n20583 );
xor ( n20585 , n20517 , n20584 );
buf ( n20586 , n20585 );
buf ( n20587 , n20586 );
nand ( n20588 , n20398 , n20587 );
buf ( n20589 , n20588 );
buf ( n20590 , n20589 );
nand ( n20591 , n20390 , n20590 );
buf ( n20592 , n20591 );
buf ( n20593 , n20592 );
buf ( n20594 , n894 );
not ( n20595 , n20594 );
buf ( n20596 , n20595 );
buf ( n20597 , n20596 );
not ( n20598 , n20478 );
not ( n20599 , n20156 );
not ( n20600 , n20599 );
or ( n20601 , n20598 , n20600 );
buf ( n20602 , n20167 );
buf ( n20603 , n20602 );
buf ( n20604 , n892 );
nand ( n20605 , n20603 , n20604 );
buf ( n20606 , n20605 );
nand ( n20607 , n20601 , n20606 );
not ( n20608 , n20607 );
buf ( n20609 , n20608 );
xor ( n20610 , n20597 , n20609 );
buf ( n20611 , n862 );
buf ( n20612 , n864 );
nand ( n20613 , n20611 , n20612 );
buf ( n20614 , n20613 );
buf ( n20615 , n20614 );
not ( n20616 , n20615 );
buf ( n20617 , n20616 );
buf ( n20618 , n20617 );
not ( n20619 , n20618 );
buf ( n20620 , n20306 );
not ( n20621 , n20620 );
buf ( n20622 , n19013 );
not ( n20623 , n20622 );
or ( n20624 , n20621 , n20623 );
buf ( n20625 , n19027 );
xor ( n20626 , n864 , n860 );
buf ( n20627 , n20626 );
nand ( n20628 , n20625 , n20627 );
buf ( n20629 , n20628 );
buf ( n20630 , n20629 );
nand ( n20631 , n20624 , n20630 );
buf ( n20632 , n20631 );
buf ( n20633 , n20632 );
not ( n20634 , n20633 );
or ( n20635 , n20619 , n20634 );
buf ( n20636 , n20330 );
not ( n20637 , n20636 );
nand ( n20638 , n18855 , n882 );
nand ( n20639 , n18844 , n18845 );
nand ( n20640 , n880 , n881 );
nand ( n20641 , n20638 , n20639 , n18859 , n20640 );
not ( n20642 , n20641 );
buf ( n20643 , n20642 );
not ( n20644 , n20643 );
or ( n20645 , n20637 , n20644 );
not ( n20646 , n18859 );
not ( n20647 , n20638 );
or ( n20648 , n20646 , n20647 );
xor ( n20649 , n880 , n844 );
nand ( n20650 , n20648 , n20649 );
buf ( n20651 , n20650 );
nand ( n20652 , n20645 , n20651 );
buf ( n20653 , n20652 );
buf ( n20654 , n20653 );
buf ( n20655 , n19013 );
buf ( n20656 , n20306 );
nand ( n20657 , n20655 , n20656 );
buf ( n20658 , n20657 );
buf ( n20659 , n20658 );
buf ( n20660 , n20629 );
buf ( n20661 , n20614 );
nand ( n20662 , n20659 , n20660 , n20661 );
buf ( n20663 , n20662 );
buf ( n20664 , n20663 );
nand ( n20665 , n20654 , n20664 );
buf ( n20666 , n20665 );
buf ( n20667 , n20666 );
nand ( n20668 , n20635 , n20667 );
buf ( n20669 , n20668 );
buf ( n20670 , n20669 );
xor ( n20671 , n20610 , n20670 );
buf ( n20672 , n20671 );
buf ( n20673 , n20672 );
buf ( n20674 , n20673 );
not ( n20675 , n20674 );
buf ( n20676 , n20614 );
buf ( n20677 , n20653 );
xor ( n20678 , n20676 , n20677 );
buf ( n20679 , n20632 );
xor ( n20680 , n20678 , n20679 );
buf ( n20681 , n20680 );
buf ( n20682 , n20681 );
not ( n20683 , n20682 );
buf ( n20684 , n20683 );
not ( n20685 , n20684 );
buf ( n20686 , n842 );
buf ( n20687 , n884 );
xor ( n20688 , n20686 , n20687 );
buf ( n20689 , n20688 );
buf ( n20690 , n20689 );
not ( n20691 , n20690 );
xnor ( n20692 , n885 , n884 );
nor ( n20693 , n20692 , n20423 );
buf ( n20694 , n20693 );
buf ( n20695 , n20694 );
not ( n20696 , n20695 );
or ( n20697 , n20691 , n20696 );
buf ( n20698 , n20423 );
buf ( n20699 , n20698 );
buf ( n20700 , n20699 );
buf ( n20701 , n20700 );
buf ( n20702 , n20417 );
nand ( n20703 , n20701 , n20702 );
buf ( n20704 , n20703 );
buf ( n20705 , n20704 );
nand ( n20706 , n20697 , n20705 );
buf ( n20707 , n20706 );
not ( n20708 , n20707 );
buf ( n20709 , n836 );
buf ( n20710 , n890 );
xor ( n20711 , n20709 , n20710 );
buf ( n20712 , n20711 );
buf ( n20713 , n20712 );
not ( n20714 , n20713 );
buf ( n20715 , n20404 );
not ( n20716 , n20715 );
or ( n20717 , n20714 , n20716 );
buf ( n20718 , n20399 );
buf ( n20719 , n20403 );
nand ( n20720 , n20718 , n20719 );
buf ( n20721 , n20720 );
buf ( n20722 , n20721 );
nand ( n20723 , n20717 , n20722 );
buf ( n20724 , n20723 );
buf ( n20725 , n20724 );
not ( n20726 , n20725 );
buf ( n20727 , n20726 );
nand ( n20728 , n20708 , n20727 );
not ( n20729 , n20728 );
buf ( n20730 , n852 );
buf ( n20731 , n874 );
xor ( n20732 , n20730 , n20731 );
buf ( n20733 , n20732 );
buf ( n20734 , n20733 );
not ( n20735 , n20734 );
and ( n20736 , n18973 , n18967 , n20548 );
buf ( n20737 , n20736 );
not ( n20738 , n20737 );
or ( n20739 , n20735 , n20738 );
buf ( n20740 , n18981 );
buf ( n20741 , n20541 );
nand ( n20742 , n20740 , n20741 );
buf ( n20743 , n20742 );
buf ( n20744 , n20743 );
nand ( n20745 , n20739 , n20744 );
buf ( n20746 , n20745 );
not ( n20747 , n20746 );
or ( n20748 , n20729 , n20747 );
buf ( n20749 , n20724 );
buf ( n20750 , n20707 );
nand ( n20751 , n20749 , n20750 );
buf ( n20752 , n20751 );
nand ( n20753 , n20748 , n20752 );
not ( n20754 , n20753 );
or ( n20755 , n20685 , n20754 );
not ( n20756 , n20681 );
buf ( n20757 , n20753 );
not ( n20758 , n20757 );
buf ( n20759 , n20758 );
not ( n20760 , n20759 );
or ( n20761 , n20756 , n20760 );
not ( n20762 , n20201 );
not ( n20763 , n19576 );
nor ( n20764 , n20763 , n19909 );
not ( n20765 , n20764 );
or ( n20766 , n20762 , n20765 );
not ( n20767 , n19569 );
buf ( n20768 , n20767 );
buf ( n20769 , n842 );
buf ( n20770 , n882 );
xor ( n20771 , n20769 , n20770 );
buf ( n20772 , n20771 );
buf ( n20773 , n20772 );
nand ( n20774 , n20768 , n20773 );
buf ( n20775 , n20774 );
nand ( n20776 , n20766 , n20775 );
not ( n20777 , n18881 );
nor ( n20778 , n20777 , n18875 );
not ( n20779 , n20778 );
buf ( n20780 , n857 );
buf ( n20781 , n868 );
xor ( n20782 , n20780 , n20781 );
buf ( n20783 , n20782 );
not ( n20784 , n20783 );
or ( n20785 , n20779 , n20784 );
not ( n20786 , n18891 );
buf ( n20787 , n20786 );
buf ( n20788 , n856 );
buf ( n20789 , n868 );
xor ( n20790 , n20788 , n20789 );
buf ( n20791 , n20790 );
buf ( n20792 , n20791 );
nand ( n20793 , n20787 , n20792 );
buf ( n20794 , n20793 );
nand ( n20795 , n20785 , n20794 );
xor ( n20796 , n20776 , n20795 );
buf ( n20797 , n19131 );
buf ( n20798 , n854 );
buf ( n20799 , n870 );
xor ( n20800 , n20798 , n20799 );
buf ( n20801 , n20800 );
buf ( n20802 , n20801 );
nand ( n20803 , n20797 , n20802 );
buf ( n20804 , n20803 );
nor ( n20805 , n20226 , n19116 );
nand ( n20806 , n20231 , n20805 );
nand ( n20807 , n20804 , n20806 );
xor ( n20808 , n20796 , n20807 );
nand ( n20809 , n20761 , n20808 );
nand ( n20810 , n20755 , n20809 );
buf ( n20811 , n20810 );
not ( n20812 , n20811 );
or ( n20813 , n20675 , n20812 );
or ( n20814 , n20810 , n20672 );
xor ( n20815 , n20484 , n20500 );
xor ( n20816 , n20815 , n20512 );
xor ( n20817 , n20441 , n20415 );
and ( n20818 , n20817 , n20459 );
not ( n20819 , n20817 );
not ( n20820 , n20459 );
and ( n20821 , n20819 , n20820 );
nor ( n20822 , n20818 , n20821 );
buf ( n20823 , n20822 );
or ( n20824 , n20816 , n20823 );
xor ( n20825 , n20563 , n20578 );
xnor ( n20826 , n20825 , n20536 );
nand ( n20827 , n20824 , n20826 );
nand ( n20828 , n20816 , n20823 );
nand ( n20829 , n20827 , n20828 );
nand ( n20830 , n20814 , n20829 );
buf ( n20831 , n20830 );
nand ( n20832 , n20813 , n20831 );
buf ( n20833 , n20832 );
buf ( n20834 , n20833 );
xor ( n20835 , n20593 , n20834 );
buf ( n20836 , n20835 );
buf ( n20837 , n20836 );
buf ( n20838 , n861 );
buf ( n20839 , n864 );
and ( n20840 , n20838 , n20839 );
buf ( n20841 , n20840 );
buf ( n20842 , n20530 );
not ( n20843 , n20842 );
and ( n20844 , n20261 , n20262 );
buf ( n20845 , n20844 );
not ( n20846 , n20845 );
or ( n20847 , n20843 , n20846 );
buf ( n20848 , n20255 );
buf ( n20849 , n837 );
buf ( n20850 , n886 );
xor ( n20851 , n20849 , n20850 );
buf ( n20852 , n20851 );
buf ( n20853 , n20852 );
nand ( n20854 , n20848 , n20853 );
buf ( n20855 , n20854 );
buf ( n20856 , n20855 );
nand ( n20857 , n20847 , n20856 );
buf ( n20858 , n20857 );
xor ( n20859 , n20841 , n20858 );
buf ( n20860 , n20408 );
not ( n20861 , n20860 );
buf ( n20862 , n20404 );
not ( n20863 , n20862 );
or ( n20864 , n20861 , n20863 );
buf ( n20865 , n833 );
buf ( n20866 , n890 );
xor ( n20867 , n20865 , n20866 );
buf ( n20868 , n20867 );
buf ( n20869 , n20403 );
nand ( n20870 , n20868 , n20869 );
buf ( n20871 , n20870 );
nand ( n20872 , n20864 , n20871 );
buf ( n20873 , n20872 );
xor ( n20874 , n20859 , n20873 );
buf ( n20875 , n20874 );
not ( n20876 , n20875 );
not ( n20877 , n20494 );
not ( n20878 , n20357 );
or ( n20879 , n20877 , n20878 );
buf ( n20880 , n20363 );
buf ( n20881 , n835 );
buf ( n20882 , n888 );
xor ( n20883 , n20881 , n20882 );
buf ( n20884 , n20883 );
buf ( n20885 , n20884 );
nand ( n20886 , n20880 , n20885 );
buf ( n20887 , n20886 );
nand ( n20888 , n20879 , n20887 );
not ( n20889 , n20888 );
buf ( n20890 , n20557 );
not ( n20891 , n20890 );
buf ( n20892 , n20736 );
not ( n20893 , n20892 );
or ( n20894 , n20891 , n20893 );
xor ( n20895 , n874 , n849 );
nand ( n20896 , n18981 , n20895 );
buf ( n20897 , n20896 );
nand ( n20898 , n20894 , n20897 );
buf ( n20899 , n20898 );
not ( n20900 , n20899 );
buf ( n20901 , n20453 );
not ( n20902 , n20901 );
buf ( n20903 , n19224 );
buf ( n20904 , n19228 );
and ( n20905 , n20903 , n20904 );
buf ( n20906 , n20905 );
buf ( n20907 , n20906 );
not ( n20908 , n20907 );
or ( n20909 , n20902 , n20908 );
buf ( n20910 , n19234 );
buf ( n20911 , n851 );
buf ( n20912 , n872 );
xor ( n20913 , n20911 , n20912 );
buf ( n20914 , n20913 );
buf ( n20915 , n20914 );
nand ( n20916 , n20910 , n20915 );
buf ( n20917 , n20916 );
buf ( n20918 , n20917 );
nand ( n20919 , n20909 , n20918 );
buf ( n20920 , n20919 );
nand ( n20921 , n20900 , n20920 );
buf ( n20922 , n20453 );
not ( n20923 , n20922 );
buf ( n20924 , n20906 );
not ( n20925 , n20924 );
or ( n20926 , n20923 , n20925 );
buf ( n20927 , n20917 );
nand ( n20928 , n20926 , n20927 );
buf ( n20929 , n20928 );
buf ( n20930 , n20929 );
not ( n20931 , n20930 );
buf ( n20932 , n20931 );
buf ( n20933 , n20932 );
buf ( n20934 , n20899 );
nand ( n20935 , n20933 , n20934 );
buf ( n20936 , n20935 );
nand ( n20937 , n20921 , n20936 );
not ( n20938 , n20937 );
or ( n20939 , n20889 , n20938 );
buf ( n20940 , n20888 );
not ( n20941 , n20940 );
buf ( n20942 , n20941 );
nand ( n20943 , n20921 , n20936 , n20942 );
nand ( n20944 , n20939 , n20943 );
buf ( n20945 , n20944 );
not ( n20946 , n20945 );
buf ( n20947 , n20946 );
buf ( n20948 , n20947 );
not ( n20949 , n20948 );
or ( n20950 , n20876 , n20949 );
buf ( n20951 , n20944 );
not ( n20952 , n20951 );
not ( n20953 , n20874 );
buf ( n20954 , n20953 );
not ( n20955 , n20954 );
or ( n20956 , n20952 , n20955 );
not ( n20957 , n20778 );
not ( n20958 , n20791 );
or ( n20959 , n20957 , n20958 );
buf ( n20960 , n18875 );
xor ( n20961 , n855 , n868 );
nand ( n20962 , n20960 , n20961 );
nand ( n20963 , n20959 , n20962 );
not ( n20964 , n20805 );
not ( n20965 , n20801 );
or ( n20966 , n20964 , n20965 );
buf ( n20967 , n19131 );
buf ( n20968 , n853 );
buf ( n20969 , n870 );
xor ( n20970 , n20968 , n20969 );
buf ( n20971 , n20970 );
buf ( n20972 , n20971 );
nand ( n20973 , n20967 , n20972 );
buf ( n20974 , n20973 );
nand ( n20975 , n20966 , n20974 );
xor ( n20976 , n20963 , n20975 );
not ( n20977 , n20772 );
not ( n20978 , n20197 );
or ( n20979 , n20977 , n20978 );
buf ( n20980 , n19568 );
buf ( n20981 , n841 );
buf ( n20982 , n882 );
xor ( n20983 , n20981 , n20982 );
buf ( n20984 , n20983 );
buf ( n20985 , n20984 );
nand ( n20986 , n20980 , n20985 );
buf ( n20987 , n20986 );
nand ( n20988 , n20979 , n20987 );
xor ( n20989 , n20976 , n20988 );
buf ( n20990 , n20989 );
nand ( n20991 , n20956 , n20990 );
buf ( n20992 , n20991 );
buf ( n20993 , n20992 );
nand ( n20994 , n20950 , n20993 );
buf ( n20995 , n20994 );
not ( n20996 , n20995 );
or ( n20997 , n20776 , n20795 );
nand ( n20998 , n20997 , n20807 );
buf ( n20999 , n20776 );
buf ( n21000 , n20795 );
nand ( n21001 , n20999 , n21000 );
buf ( n21002 , n21001 );
nand ( n21003 , n20998 , n21002 );
not ( n21004 , n21003 );
and ( n21005 , n879 , n878 );
not ( n21006 , n879 );
not ( n21007 , n878 );
and ( n21008 , n21006 , n21007 );
nor ( n21009 , n21005 , n21008 );
not ( n21010 , n21009 );
not ( n21011 , n21010 );
not ( n21012 , n19255 );
nand ( n21013 , n21011 , n21012 );
not ( n21014 , n21013 );
not ( n21015 , n20507 );
and ( n21016 , n21014 , n21015 );
xor ( n21017 , n878 , n845 );
not ( n21018 , n21017 );
nor ( n21019 , n21018 , n21012 );
nor ( n21020 , n21016 , n21019 );
not ( n21021 , n21020 );
not ( n21022 , n21021 );
buf ( n21023 , n20571 );
not ( n21024 , n21023 );
buf ( n21025 , n20243 );
not ( n21026 , n21025 );
or ( n21027 , n21024 , n21026 );
buf ( n21028 , n20246 );
xor ( n21029 , n876 , n847 );
buf ( n21030 , n21029 );
nand ( n21031 , n21028 , n21030 );
buf ( n21032 , n21031 );
buf ( n21033 , n21032 );
nand ( n21034 , n21027 , n21033 );
buf ( n21035 , n21034 );
not ( n21036 , n21035 );
not ( n21037 , n21036 );
or ( n21038 , n21022 , n21037 );
nand ( n21039 , n21020 , n21035 );
nand ( n21040 , n21038 , n21039 );
not ( n21041 , n20435 );
not ( n21042 , n20430 );
or ( n21043 , n21041 , n21042 );
buf ( n21044 , n20423 );
xor ( n21045 , n884 , n839 );
buf ( n21046 , n21045 );
nand ( n21047 , n21044 , n21046 );
buf ( n21048 , n21047 );
nand ( n21049 , n21043 , n21048 );
not ( n21050 , n21049 );
and ( n21051 , n21040 , n21050 );
not ( n21052 , n21040 );
and ( n21053 , n21052 , n21049 );
nor ( n21054 , n21051 , n21053 );
not ( n21055 , n21054 );
not ( n21056 , n21055 );
or ( n21057 , n21004 , n21056 );
buf ( n21058 , n21003 );
not ( n21059 , n21058 );
buf ( n21060 , n21059 );
not ( n21061 , n21060 );
not ( n21062 , n21054 );
or ( n21063 , n21061 , n21062 );
buf ( n21064 , n20111 );
not ( n21065 , n21064 );
buf ( n21066 , n18928 );
not ( n21067 , n21066 );
or ( n21068 , n21065 , n21067 );
buf ( n21069 , n18938 );
buf ( n21070 , n857 );
buf ( n21071 , n866 );
xor ( n21072 , n21070 , n21071 );
buf ( n21073 , n21072 );
buf ( n21074 , n21073 );
nand ( n21075 , n21069 , n21074 );
buf ( n21076 , n21075 );
buf ( n21077 , n21076 );
nand ( n21078 , n21068 , n21077 );
buf ( n21079 , n21078 );
buf ( n21080 , n21079 );
not ( n21081 , n21080 );
and ( n21082 , n20642 , n20649 );
nand ( n21083 , n18859 , n20638 );
xor ( n21084 , n880 , n843 );
and ( n21085 , n21083 , n21084 );
nor ( n21086 , n21082 , n21085 );
buf ( n21087 , n21086 );
not ( n21088 , n21087 );
or ( n21089 , n21081 , n21088 );
buf ( n21090 , n21086 );
buf ( n21091 , n21079 );
or ( n21092 , n21090 , n21091 );
nand ( n21093 , n21089 , n21092 );
buf ( n21094 , n21093 );
buf ( n21095 , n21094 );
buf ( n21096 , n20626 );
not ( n21097 , n21096 );
buf ( n21098 , n19013 );
not ( n21099 , n21098 );
or ( n21100 , n21097 , n21099 );
buf ( n21101 , n19027 );
buf ( n21102 , n859 );
buf ( n21103 , n864 );
xor ( n21104 , n21102 , n21103 );
buf ( n21105 , n21104 );
buf ( n21106 , n21105 );
nand ( n21107 , n21101 , n21106 );
buf ( n21108 , n21107 );
buf ( n21109 , n21108 );
nand ( n21110 , n21100 , n21109 );
buf ( n21111 , n21110 );
buf ( n21112 , n21111 );
not ( n21113 , n21112 );
buf ( n21114 , n21113 );
buf ( n21115 , n21114 );
and ( n21116 , n21095 , n21115 );
not ( n21117 , n21095 );
buf ( n21118 , n21111 );
and ( n21119 , n21117 , n21118 );
nor ( n21120 , n21116 , n21119 );
buf ( n21121 , n21120 );
buf ( n21122 , n21121 );
not ( n21123 , n21122 );
buf ( n21124 , n21123 );
nand ( n21125 , n21063 , n21124 );
nand ( n21126 , n21057 , n21125 );
not ( n21127 , n21126 );
not ( n21128 , n21127 );
and ( n21129 , n20996 , n21128 );
and ( n21130 , n21127 , n20995 );
nor ( n21131 , n21129 , n21130 );
buf ( n21132 , n20932 );
not ( n21133 , n21132 );
buf ( n21134 , n20942 );
not ( n21135 , n21134 );
or ( n21136 , n21133 , n21135 );
buf ( n21137 , n20899 );
nand ( n21138 , n21136 , n21137 );
buf ( n21139 , n21138 );
buf ( n21140 , n21139 );
buf ( n21141 , n20888 );
buf ( n21142 , n20929 );
nand ( n21143 , n21141 , n21142 );
buf ( n21144 , n21143 );
buf ( n21145 , n21144 );
nand ( n21146 , n21140 , n21145 );
buf ( n21147 , n21146 );
not ( n21148 , n21049 );
not ( n21149 , n21035 );
or ( n21150 , n21148 , n21149 );
or ( n21151 , n21049 , n21035 );
nand ( n21152 , n21151 , n21021 );
nand ( n21153 , n21150 , n21152 );
and ( n21154 , n21147 , n21153 );
not ( n21155 , n21147 );
buf ( n21156 , n21153 );
not ( n21157 , n21156 );
buf ( n21158 , n21157 );
and ( n21159 , n21155 , n21158 );
nor ( n21160 , n21154 , n21159 );
or ( n21161 , n20963 , n20988 );
nand ( n21162 , n21161 , n20975 );
nand ( n21163 , n20963 , n20988 );
nand ( n21164 , n21162 , n21163 );
not ( n21165 , n21164 );
and ( n21166 , n21160 , n21165 );
not ( n21167 , n21160 );
and ( n21168 , n21167 , n21164 );
nor ( n21169 , n21166 , n21168 );
buf ( n21170 , n21169 );
and ( n21171 , n21131 , n21170 );
not ( n21172 , n21131 );
buf ( n21173 , n21169 );
not ( n21174 , n21173 );
buf ( n21175 , n21174 );
and ( n21176 , n21172 , n21175 );
nor ( n21177 , n21171 , n21176 );
buf ( n21178 , n21177 );
and ( n21179 , n20837 , n21178 );
not ( n21180 , n20837 );
buf ( n21181 , n21177 );
not ( n21182 , n21181 );
buf ( n21183 , n21182 );
buf ( n21184 , n21183 );
and ( n21185 , n21180 , n21184 );
nor ( n21186 , n21179 , n21185 );
buf ( n21187 , n21186 );
buf ( n21188 , n21187 );
not ( n21189 , n21188 );
buf ( n21190 , n21189 );
buf ( n21191 , n21190 );
not ( n21192 , n21191 );
xor ( n21193 , n20822 , n20816 );
xor ( n21194 , n21193 , n20826 );
not ( n21195 , n21194 );
buf ( n21196 , n20759 );
not ( n21197 , n21196 );
buf ( n21198 , n20684 );
not ( n21199 , n21198 );
or ( n21200 , n21197 , n21199 );
buf ( n21201 , n20681 );
buf ( n21202 , n20753 );
nand ( n21203 , n21201 , n21202 );
buf ( n21204 , n21203 );
buf ( n21205 , n21204 );
nand ( n21206 , n21200 , n21205 );
buf ( n21207 , n21206 );
buf ( n21208 , n21207 );
buf ( n21209 , n20808 );
not ( n21210 , n21209 );
buf ( n21211 , n21210 );
buf ( n21212 , n21211 );
and ( n21213 , n21208 , n21212 );
not ( n21214 , n21208 );
buf ( n21215 , n20808 );
and ( n21216 , n21214 , n21215 );
nor ( n21217 , n21213 , n21216 );
buf ( n21218 , n21217 );
buf ( n21219 , n21218 );
not ( n21220 , n21219 );
buf ( n21221 , n21220 );
not ( n21222 , n21221 );
or ( n21223 , n21195 , n21222 );
nor ( n21224 , n21194 , n21221 );
and ( n21225 , n20371 , n20310 );
not ( n21226 , n20371 );
and ( n21227 , n21226 , n20313 );
nor ( n21228 , n21225 , n21227 );
buf ( n21229 , n21228 );
buf ( n21230 , n20339 );
and ( n21231 , n21229 , n21230 );
not ( n21232 , n21229 );
buf ( n21233 , n20336 );
and ( n21234 , n21232 , n21233 );
or ( n21235 , n21231 , n21234 );
buf ( n21236 , n21235 );
buf ( n21237 , n21236 );
buf ( n21238 , n860 );
buf ( n21239 , n866 );
xor ( n21240 , n21238 , n21239 );
buf ( n21241 , n21240 );
buf ( n21242 , n21241 );
not ( n21243 , n21242 );
buf ( n21244 , n18931 );
not ( n21245 , n21244 );
or ( n21246 , n21243 , n21245 );
buf ( n21247 , n18938 );
buf ( n21248 , n21247 );
buf ( n21249 , n21248 );
buf ( n21250 , n21249 );
buf ( n21251 , n20101 );
nand ( n21252 , n21250 , n21251 );
buf ( n21253 , n21252 );
buf ( n21254 , n21253 );
nand ( n21255 , n21246 , n21254 );
buf ( n21256 , n21255 );
buf ( n21257 , n21256 );
buf ( n21258 , n858 );
buf ( n21259 , n868 );
xor ( n21260 , n21258 , n21259 );
buf ( n21261 , n21260 );
buf ( n21262 , n21261 );
not ( n21263 , n21262 );
buf ( n21264 , n18887 );
not ( n21265 , n21264 );
or ( n21266 , n21263 , n21265 );
buf ( n21267 , n19461 );
buf ( n21268 , n20783 );
nand ( n21269 , n21267 , n21268 );
buf ( n21270 , n21269 );
buf ( n21271 , n21270 );
nand ( n21272 , n21266 , n21271 );
buf ( n21273 , n21272 );
buf ( n21274 , n21273 );
xor ( n21275 , n21257 , n21274 );
buf ( n21276 , n863 );
buf ( n21277 , n865 );
or ( n21278 , n21276 , n21277 );
buf ( n21279 , n866 );
nand ( n21280 , n21278 , n21279 );
buf ( n21281 , n21280 );
buf ( n21282 , n21281 );
buf ( n21283 , n863 );
buf ( n21284 , n865 );
nand ( n21285 , n21283 , n21284 );
buf ( n21286 , n21285 );
buf ( n21287 , n21286 );
buf ( n21288 , n864 );
and ( n21289 , n21282 , n21287 , n21288 );
buf ( n21290 , n21289 );
buf ( n21291 , n21290 );
xor ( n21292 , n894 , n833 );
buf ( n21293 , n21292 );
not ( n21294 , n21293 );
not ( n21295 , n895 );
nand ( n21296 , n21295 , n894 );
not ( n21297 , n21296 );
buf ( n21298 , n21297 );
not ( n21299 , n21298 );
or ( n21300 , n21294 , n21299 );
buf ( n21301 , n20129 );
buf ( n21302 , n895 );
nand ( n21303 , n21301 , n21302 );
buf ( n21304 , n21303 );
buf ( n21305 , n21304 );
nand ( n21306 , n21300 , n21305 );
buf ( n21307 , n21306 );
buf ( n21308 , n21307 );
and ( n21309 , n21291 , n21308 );
buf ( n21310 , n21309 );
buf ( n21311 , n21310 );
xor ( n21312 , n21275 , n21311 );
buf ( n21313 , n21312 );
buf ( n21314 , n21313 );
xor ( n21315 , n21237 , n21314 );
buf ( n21316 , n860 );
buf ( n21317 , n868 );
xor ( n21318 , n21316 , n21317 );
buf ( n21319 , n21318 );
buf ( n21320 , n21319 );
not ( n21321 , n21320 );
buf ( n21322 , n20778 );
not ( n21323 , n21322 );
or ( n21324 , n21321 , n21323 );
buf ( n21325 , n20786 );
buf ( n21326 , n859 );
buf ( n21327 , n868 );
xor ( n21328 , n21326 , n21327 );
buf ( n21329 , n21328 );
buf ( n21330 , n21329 );
nand ( n21331 , n21325 , n21330 );
buf ( n21332 , n21331 );
buf ( n21333 , n21332 );
nand ( n21334 , n21324 , n21333 );
buf ( n21335 , n21334 );
buf ( n21336 , n21335 );
not ( n21337 , n21336 );
buf ( n21338 , n21337 );
buf ( n21339 , n21338 );
not ( n21340 , n21339 );
buf ( n21341 , n846 );
buf ( n21342 , n882 );
xor ( n21343 , n21341 , n21342 );
buf ( n21344 , n21343 );
buf ( n21345 , n21344 );
not ( n21346 , n21345 );
buf ( n21347 , n20197 );
not ( n21348 , n21347 );
or ( n21349 , n21346 , n21348 );
buf ( n21350 , n19909 );
buf ( n21351 , n845 );
buf ( n21352 , n882 );
xor ( n21353 , n21351 , n21352 );
buf ( n21354 , n21353 );
buf ( n21355 , n21354 );
nand ( n21356 , n21350 , n21355 );
buf ( n21357 , n21356 );
buf ( n21358 , n21357 );
nand ( n21359 , n21349 , n21358 );
buf ( n21360 , n21359 );
buf ( n21361 , n21360 );
not ( n21362 , n21361 );
buf ( n21363 , n21362 );
buf ( n21364 , n21363 );
not ( n21365 , n21364 );
or ( n21366 , n21340 , n21365 );
xor ( n21367 , n870 , n858 );
buf ( n21368 , n21367 );
not ( n21369 , n21368 );
buf ( n21370 , n19122 );
not ( n21371 , n21370 );
or ( n21372 , n21369 , n21371 );
buf ( n21373 , n19131 );
buf ( n21374 , n857 );
buf ( n21375 , n870 );
xor ( n21376 , n21374 , n21375 );
buf ( n21377 , n21376 );
buf ( n21378 , n21377 );
nand ( n21379 , n21373 , n21378 );
buf ( n21380 , n21379 );
buf ( n21381 , n21380 );
nand ( n21382 , n21372 , n21381 );
buf ( n21383 , n21382 );
buf ( n21384 , n21383 );
nand ( n21385 , n21366 , n21384 );
buf ( n21386 , n21385 );
buf ( n21387 , n21386 );
buf ( n21388 , n21360 );
buf ( n21389 , n21335 );
nand ( n21390 , n21388 , n21389 );
buf ( n21391 , n21390 );
buf ( n21392 , n21391 );
nand ( n21393 , n21387 , n21392 );
buf ( n21394 , n21393 );
buf ( n21395 , n21394 );
buf ( n21396 , n844 );
buf ( n21397 , n884 );
xor ( n21398 , n21396 , n21397 );
buf ( n21399 , n21398 );
not ( n21400 , n21399 );
not ( n21401 , n20430 );
or ( n21402 , n21400 , n21401 );
buf ( n21403 , n20423 );
buf ( n21404 , n843 );
buf ( n21405 , n884 );
xor ( n21406 , n21404 , n21405 );
buf ( n21407 , n21406 );
buf ( n21408 , n21407 );
nand ( n21409 , n21403 , n21408 );
buf ( n21410 , n21409 );
nand ( n21411 , n21402 , n21410 );
buf ( n21412 , n856 );
buf ( n21413 , n872 );
xor ( n21414 , n21412 , n21413 );
buf ( n21415 , n21414 );
not ( n21416 , n21415 );
not ( n21417 , n20211 );
or ( n21418 , n21416 , n21417 );
buf ( n21419 , n19234 );
buf ( n21420 , n855 );
buf ( n21421 , n872 );
xor ( n21422 , n21420 , n21421 );
buf ( n21423 , n21422 );
buf ( n21424 , n21423 );
nand ( n21425 , n21419 , n21424 );
buf ( n21426 , n21425 );
nand ( n21427 , n21418 , n21426 );
xor ( n21428 , n21411 , n21427 );
buf ( n21429 , n838 );
buf ( n21430 , n890 );
xor ( n21431 , n21429 , n21430 );
buf ( n21432 , n21431 );
not ( n21433 , n21432 );
nor ( n21434 , n890 , n891 );
not ( n21435 , n21434 );
nand ( n21436 , n890 , n891 );
nand ( n21437 , n21435 , n21436 );
nor ( n21438 , n20403 , n21437 );
buf ( n21439 , n21438 );
buf ( n21440 , n21439 );
buf ( n21441 , n21440 );
not ( n21442 , n21441 );
or ( n21443 , n21433 , n21442 );
buf ( n21444 , n20869 );
buf ( n21445 , n837 );
buf ( n21446 , n890 );
xor ( n21447 , n21445 , n21446 );
buf ( n21448 , n21447 );
buf ( n21449 , n21448 );
nand ( n21450 , n21444 , n21449 );
buf ( n21451 , n21450 );
nand ( n21452 , n21443 , n21451 );
and ( n21453 , n21428 , n21452 );
and ( n21454 , n21411 , n21427 );
or ( n21455 , n21453 , n21454 );
buf ( n21456 , n21455 );
or ( n21457 , n21395 , n21456 );
buf ( n21458 , n852 );
buf ( n21459 , n876 );
xor ( n21460 , n21458 , n21459 );
buf ( n21461 , n21460 );
buf ( n21462 , n21461 );
not ( n21463 , n21462 );
buf ( n21464 , n20243 );
not ( n21465 , n21464 );
or ( n21466 , n21463 , n21465 );
buf ( n21467 , n19082 );
buf ( n21468 , n851 );
buf ( n21469 , n876 );
xor ( n21470 , n21468 , n21469 );
buf ( n21471 , n21470 );
buf ( n21472 , n21471 );
nand ( n21473 , n21467 , n21472 );
buf ( n21474 , n21473 );
buf ( n21475 , n21474 );
nand ( n21476 , n21466 , n21475 );
buf ( n21477 , n21476 );
not ( n21478 , n21477 );
not ( n21479 , n20255 );
buf ( n21480 , n841 );
buf ( n21481 , n886 );
xor ( n21482 , n21480 , n21481 );
buf ( n21483 , n21482 );
not ( n21484 , n21483 );
or ( n21485 , n21479 , n21484 );
buf ( n21486 , n20261 );
and ( n21487 , n842 , n886 );
not ( n21488 , n842 );
and ( n21489 , n21488 , n20265 );
nor ( n21490 , n21487 , n21489 );
nand ( n21491 , n20262 , n21486 , n21490 );
nand ( n21492 , n21485 , n21491 );
not ( n21493 , n21492 );
or ( n21494 , n21478 , n21493 );
buf ( n21495 , n21477 );
not ( n21496 , n21495 );
buf ( n21497 , n21496 );
not ( n21498 , n21497 );
not ( n21499 , n21492 );
not ( n21500 , n21499 );
or ( n21501 , n21498 , n21500 );
buf ( n21502 , n854 );
buf ( n21503 , n874 );
xor ( n21504 , n21502 , n21503 );
buf ( n21505 , n21504 );
buf ( n21506 , n21505 );
not ( n21507 , n21506 );
buf ( n21508 , n18974 );
not ( n21509 , n21508 );
or ( n21510 , n21507 , n21509 );
buf ( n21511 , n18984 );
not ( n21512 , n21511 );
buf ( n21513 , n21512 );
buf ( n21514 , n21513 );
buf ( n21515 , n853 );
buf ( n21516 , n874 );
xor ( n21517 , n21515 , n21516 );
buf ( n21518 , n21517 );
buf ( n21519 , n21518 );
nand ( n21520 , n21514 , n21519 );
buf ( n21521 , n21520 );
buf ( n21522 , n21521 );
nand ( n21523 , n21510 , n21522 );
buf ( n21524 , n21523 );
nand ( n21525 , n21501 , n21524 );
nand ( n21526 , n21494 , n21525 );
buf ( n21527 , n21526 );
nand ( n21528 , n21457 , n21527 );
buf ( n21529 , n21528 );
buf ( n21530 , n21529 );
buf ( n21531 , n21394 );
buf ( n21532 , n21455 );
nand ( n21533 , n21531 , n21532 );
buf ( n21534 , n21533 );
buf ( n21535 , n21534 );
nand ( n21536 , n21530 , n21535 );
buf ( n21537 , n21536 );
buf ( n21538 , n21537 );
and ( n21539 , n21315 , n21538 );
and ( n21540 , n21237 , n21314 );
or ( n21541 , n21539 , n21540 );
buf ( n21542 , n21541 );
not ( n21543 , n21542 );
or ( n21544 , n21224 , n21543 );
nand ( n21545 , n21223 , n21544 );
buf ( n21546 , n21545 );
buf ( n21547 , n20989 );
not ( n21548 , n21547 );
buf ( n21549 , n21548 );
buf ( n21550 , n21549 );
not ( n21551 , n21550 );
and ( n21552 , n20944 , n20953 );
not ( n21553 , n20944 );
and ( n21554 , n21553 , n20874 );
nor ( n21555 , n21552 , n21554 );
buf ( n21556 , n21555 );
not ( n21557 , n21556 );
or ( n21558 , n21551 , n21557 );
buf ( n21559 , n21555 );
buf ( n21560 , n21549 );
or ( n21561 , n21559 , n21560 );
nand ( n21562 , n21558 , n21561 );
buf ( n21563 , n21562 );
buf ( n21564 , n21563 );
buf ( n21565 , n21003 );
not ( n21566 , n21565 );
buf ( n21567 , n21121 );
not ( n21568 , n21567 );
or ( n21569 , n21566 , n21568 );
buf ( n21570 , n21003 );
buf ( n21571 , n21121 );
or ( n21572 , n21570 , n21571 );
nand ( n21573 , n21569 , n21572 );
buf ( n21574 , n21573 );
and ( n21575 , n21574 , n21054 );
not ( n21576 , n21574 );
and ( n21577 , n21576 , n21055 );
or ( n21578 , n21575 , n21577 );
buf ( n21579 , n21578 );
xor ( n21580 , n21564 , n21579 );
xor ( n21581 , n20097 , n20118 );
xor ( n21582 , n21581 , n20181 );
buf ( n21583 , n21582 );
buf ( n21584 , n21583 );
xor ( n21585 , n20240 , n20294 );
xor ( n21586 , n21585 , n20382 );
buf ( n21587 , n21586 );
xor ( n21588 , n21584 , n21587 );
xor ( n21589 , n20746 , n20727 );
buf ( n21590 , n20707 );
buf ( n21591 , n21590 );
buf ( n21592 , n21591 );
xor ( n21593 , n21589 , n21592 );
buf ( n21594 , n21593 );
not ( n21595 , n21594 );
buf ( n21596 , n21595 );
not ( n21597 , n21596 );
buf ( n21598 , n20238 );
not ( n21599 , n21598 );
not ( n21600 , n21599 );
not ( n21601 , n20205 );
not ( n21602 , n21601 );
not ( n21603 , n20219 );
not ( n21604 , n21603 );
or ( n21605 , n21602 , n21604 );
or ( n21606 , n21601 , n21603 );
nand ( n21607 , n21605 , n21606 );
not ( n21608 , n21607 );
or ( n21609 , n21600 , n21608 );
or ( n21610 , n21599 , n21607 );
nand ( n21611 , n21609 , n21610 );
buf ( n21612 , n21611 );
not ( n21613 , n21612 );
buf ( n21614 , n21613 );
not ( n21615 , n21614 );
or ( n21616 , n21597 , n21615 );
not ( n21617 , n21611 );
not ( n21618 , n21593 );
or ( n21619 , n21617 , n21618 );
xor ( n21620 , n20269 , n20288 );
xor ( n21621 , n21620 , n20252 );
nand ( n21622 , n21619 , n21621 );
nand ( n21623 , n21616 , n21622 );
buf ( n21624 , n21623 );
and ( n21625 , n21588 , n21624 );
and ( n21626 , n21584 , n21587 );
or ( n21627 , n21625 , n21626 );
buf ( n21628 , n21627 );
buf ( n21629 , n21628 );
xor ( n21630 , n21580 , n21629 );
buf ( n21631 , n21630 );
buf ( n21632 , n21631 );
xor ( n21633 , n21546 , n21632 );
xor ( n21634 , n21257 , n21274 );
and ( n21635 , n21634 , n21311 );
and ( n21636 , n21257 , n21274 );
or ( n21637 , n21635 , n21636 );
buf ( n21638 , n21637 );
xor ( n21639 , n20124 , n20137 );
xor ( n21640 , n21639 , n20176 );
buf ( n21641 , n21640 );
buf ( n21642 , n21641 );
buf ( n21643 , n21329 );
not ( n21644 , n21643 );
buf ( n21645 , n20778 );
not ( n21646 , n21645 );
or ( n21647 , n21644 , n21646 );
buf ( n21648 , n20960 );
buf ( n21649 , n21261 );
nand ( n21650 , n21648 , n21649 );
buf ( n21651 , n21650 );
buf ( n21652 , n21651 );
nand ( n21653 , n21647 , n21652 );
buf ( n21654 , n21653 );
buf ( n21655 , n21654 );
not ( n21656 , n21655 );
buf ( n21657 , n21354 );
not ( n21658 , n21657 );
buf ( n21659 , n20197 );
not ( n21660 , n21659 );
or ( n21661 , n21658 , n21660 );
buf ( n21662 , n20188 );
buf ( n21663 , n19568 );
nand ( n21664 , n21662 , n21663 );
buf ( n21665 , n21664 );
buf ( n21666 , n21665 );
nand ( n21667 , n21661 , n21666 );
buf ( n21668 , n21667 );
buf ( n21669 , n21668 );
not ( n21670 , n21669 );
or ( n21671 , n21656 , n21670 );
buf ( n21672 , n21654 );
not ( n21673 , n21672 );
buf ( n21674 , n21673 );
buf ( n21675 , n21674 );
not ( n21676 , n21675 );
not ( n21677 , n21668 );
buf ( n21678 , n21677 );
not ( n21679 , n21678 );
or ( n21680 , n21676 , n21679 );
buf ( n21681 , n861 );
buf ( n21682 , n866 );
xor ( n21683 , n21681 , n21682 );
buf ( n21684 , n21683 );
buf ( n21685 , n21684 );
not ( n21686 , n21685 );
buf ( n21687 , n18931 );
not ( n21688 , n21687 );
or ( n21689 , n21686 , n21688 );
buf ( n21690 , n21249 );
buf ( n21691 , n21241 );
nand ( n21692 , n21690 , n21691 );
buf ( n21693 , n21692 );
buf ( n21694 , n21693 );
nand ( n21695 , n21689 , n21694 );
buf ( n21696 , n21695 );
buf ( n21697 , n21696 );
nand ( n21698 , n21680 , n21697 );
buf ( n21699 , n21698 );
buf ( n21700 , n21699 );
nand ( n21701 , n21671 , n21700 );
buf ( n21702 , n21701 );
buf ( n21703 , n21702 );
xor ( n21704 , n21642 , n21703 );
not ( n21705 , n21423 );
not ( n21706 , n20211 );
or ( n21707 , n21705 , n21706 );
buf ( n21708 , n19234 );
buf ( n21709 , n20207 );
nand ( n21710 , n21708 , n21709 );
buf ( n21711 , n21710 );
nand ( n21712 , n21707 , n21711 );
not ( n21713 , n21407 );
not ( n21714 , n20694 );
or ( n21715 , n21713 , n21714 );
buf ( n21716 , n20700 );
buf ( n21717 , n20689 );
nand ( n21718 , n21716 , n21717 );
buf ( n21719 , n21718 );
nand ( n21720 , n21715 , n21719 );
nor ( n21721 , n21712 , n21720 );
buf ( n21722 , n19114 );
not ( n21723 , n21722 );
buf ( n21724 , n21723 );
buf ( n21725 , n21724 );
not ( n21726 , n21725 );
buf ( n21727 , n21726 );
buf ( n21728 , n21727 );
buf ( n21729 , n20236 );
nand ( n21730 , n21728 , n21729 );
buf ( n21731 , n21730 );
nand ( n21732 , n19122 , n21377 );
and ( n21733 , n21731 , n21732 );
or ( n21734 , n21721 , n21733 );
nand ( n21735 , n21712 , n21720 );
nand ( n21736 , n21734 , n21735 );
buf ( n21737 , n21736 );
and ( n21738 , n21704 , n21737 );
and ( n21739 , n21642 , n21703 );
or ( n21740 , n21738 , n21739 );
buf ( n21741 , n21740 );
xor ( n21742 , n21638 , n21741 );
buf ( n21743 , n839 );
buf ( n21744 , n888 );
xor ( n21745 , n21743 , n21744 );
buf ( n21746 , n21745 );
not ( n21747 , n21746 );
not ( n21748 , n20357 );
or ( n21749 , n21747 , n21748 );
buf ( n21750 , n20363 );
buf ( n21751 , n20346 );
nand ( n21752 , n21750 , n21751 );
buf ( n21753 , n21752 );
nand ( n21754 , n21749 , n21753 );
not ( n21755 , n21754 );
not ( n21756 , n21755 );
buf ( n21757 , n835 );
buf ( n21758 , n892 );
xor ( n21759 , n21757 , n21758 );
buf ( n21760 , n21759 );
not ( n21761 , n21760 );
nand ( n21762 , n20164 , n20155 );
not ( n21763 , n21762 );
not ( n21764 , n21763 );
or ( n21765 , n21761 , n21764 );
buf ( n21766 , n20167 );
buf ( n21767 , n20142 );
nand ( n21768 , n21766 , n21767 );
buf ( n21769 , n21768 );
nand ( n21770 , n21765 , n21769 );
not ( n21771 , n21770 );
not ( n21772 , n21771 );
or ( n21773 , n21756 , n21772 );
buf ( n21774 , n863 );
buf ( n21775 , n864 );
xor ( n21776 , n21774 , n21775 );
buf ( n21777 , n21776 );
buf ( n21778 , n21777 );
not ( n21779 , n21778 );
buf ( n21780 , n19013 );
not ( n21781 , n21780 );
or ( n21782 , n21779 , n21781 );
buf ( n21783 , n19030 );
buf ( n21784 , n20299 );
nand ( n21785 , n21783 , n21784 );
buf ( n21786 , n21785 );
buf ( n21787 , n21786 );
nand ( n21788 , n21782 , n21787 );
buf ( n21789 , n21788 );
nand ( n21790 , n21773 , n21789 );
buf ( n21791 , n21790 );
nand ( n21792 , n21754 , n21770 );
buf ( n21793 , n21792 );
nand ( n21794 , n21791 , n21793 );
buf ( n21795 , n21794 );
buf ( n21796 , n21795 );
buf ( n21797 , n847 );
buf ( n21798 , n880 );
xor ( n21799 , n21797 , n21798 );
buf ( n21800 , n21799 );
buf ( n21801 , n21800 );
not ( n21802 , n21801 );
buf ( n21803 , n20642 );
not ( n21804 , n21803 );
or ( n21805 , n21802 , n21804 );
buf ( n21806 , n20325 );
buf ( n21807 , n20319 );
nand ( n21808 , n21806 , n21807 );
buf ( n21809 , n21808 );
buf ( n21810 , n21809 );
nand ( n21811 , n21805 , n21810 );
buf ( n21812 , n21811 );
buf ( n21813 , n21812 );
not ( n21814 , n21813 );
buf ( n21815 , n21483 );
not ( n21816 , n21815 );
and ( n21817 , n20261 , n20262 );
buf ( n21818 , n21817 );
not ( n21819 , n21818 );
or ( n21820 , n21816 , n21819 );
buf ( n21821 , n20525 );
buf ( n21822 , n20267 );
nand ( n21823 , n21821 , n21822 );
buf ( n21824 , n21823 );
buf ( n21825 , n21824 );
nand ( n21826 , n21820 , n21825 );
buf ( n21827 , n21826 );
buf ( n21828 , n21827 );
not ( n21829 , n21828 );
or ( n21830 , n21814 , n21829 );
buf ( n21831 , n21812 );
buf ( n21832 , n21827 );
or ( n21833 , n21831 , n21832 );
buf ( n21834 , n849 );
buf ( n21835 , n878 );
xor ( n21836 , n21834 , n21835 );
buf ( n21837 , n21836 );
buf ( n21838 , n21837 );
not ( n21839 , n21838 );
buf ( n21840 , n19259 );
not ( n21841 , n21840 );
or ( n21842 , n21839 , n21841 );
buf ( n21843 , n19265 );
buf ( n21844 , n20286 );
nand ( n21845 , n21843 , n21844 );
buf ( n21846 , n21845 );
buf ( n21847 , n21846 );
nand ( n21848 , n21842 , n21847 );
buf ( n21849 , n21848 );
buf ( n21850 , n21849 );
nand ( n21851 , n21833 , n21850 );
buf ( n21852 , n21851 );
buf ( n21853 , n21852 );
nand ( n21854 , n21830 , n21853 );
buf ( n21855 , n21854 );
buf ( n21856 , n21855 );
or ( n21857 , n21796 , n21856 );
buf ( n21858 , n21448 );
not ( n21859 , n21858 );
buf ( n21860 , n21441 );
not ( n21861 , n21860 );
or ( n21862 , n21859 , n21861 );
buf ( n21863 , n20869 );
buf ( n21864 , n20712 );
nand ( n21865 , n21863 , n21864 );
buf ( n21866 , n21865 );
buf ( n21867 , n21866 );
nand ( n21868 , n21862 , n21867 );
buf ( n21869 , n21868 );
buf ( n21870 , n21869 );
not ( n21871 , n21870 );
buf ( n21872 , n21471 );
not ( n21873 , n21872 );
buf ( n21874 , n19153 );
not ( n21875 , n21874 );
or ( n21876 , n21873 , n21875 );
buf ( n21877 , n20246 );
buf ( n21878 , n20241 );
nand ( n21879 , n21877 , n21878 );
buf ( n21880 , n21879 );
buf ( n21881 , n21880 );
nand ( n21882 , n21876 , n21881 );
buf ( n21883 , n21882 );
buf ( n21884 , n21883 );
not ( n21885 , n21884 );
or ( n21886 , n21871 , n21885 );
or ( n21887 , n21869 , n21883 );
buf ( n21888 , n21518 );
not ( n21889 , n21888 );
buf ( n21890 , n20549 );
not ( n21891 , n21890 );
or ( n21892 , n21889 , n21891 );
buf ( n21893 , n20555 );
buf ( n21894 , n20733 );
nand ( n21895 , n21893 , n21894 );
buf ( n21896 , n21895 );
buf ( n21897 , n21896 );
nand ( n21898 , n21892 , n21897 );
buf ( n21899 , n21898 );
nand ( n21900 , n21887 , n21899 );
buf ( n21901 , n21900 );
nand ( n21902 , n21886 , n21901 );
buf ( n21903 , n21902 );
buf ( n21904 , n21903 );
nand ( n21905 , n21857 , n21904 );
buf ( n21906 , n21905 );
buf ( n21907 , n21906 );
buf ( n21908 , n21795 );
buf ( n21909 , n21855 );
nand ( n21910 , n21908 , n21909 );
buf ( n21911 , n21910 );
buf ( n21912 , n21911 );
nand ( n21913 , n21907 , n21912 );
buf ( n21914 , n21913 );
xor ( n21915 , n21742 , n21914 );
buf ( n21916 , n21915 );
xor ( n21917 , n21291 , n21308 );
buf ( n21918 , n21917 );
buf ( n21919 , n21918 );
not ( n21920 , n21292 );
not ( n21921 , n895 );
or ( n21922 , n21920 , n21921 );
buf ( n21923 , n895 );
not ( n21924 , n21923 );
buf ( n21925 , n894 );
nand ( n21926 , n21924 , n21925 );
buf ( n21927 , n21926 );
buf ( n21928 , n834 );
buf ( n21929 , n894 );
xor ( n21930 , n21928 , n21929 );
buf ( n21931 , n21930 );
buf ( n21932 , n21931 );
not ( n21933 , n21932 );
buf ( n21934 , n21933 );
or ( n21935 , n21927 , n21934 );
nand ( n21936 , n21922 , n21935 );
buf ( n21937 , n21936 );
buf ( n21938 , n19027 );
buf ( n21939 , n863 );
and ( n21940 , n21938 , n21939 );
buf ( n21941 , n21940 );
buf ( n21942 , n21941 );
xor ( n21943 , n21937 , n21942 );
buf ( n21944 , n836 );
buf ( n21945 , n892 );
xor ( n21946 , n21944 , n21945 );
buf ( n21947 , n21946 );
buf ( n21948 , n21947 );
not ( n21949 , n21948 );
buf ( n21950 , n20159 );
not ( n21951 , n21950 );
or ( n21952 , n21949 , n21951 );
buf ( n21953 , n20167 );
buf ( n21954 , n21760 );
nand ( n21955 , n21953 , n21954 );
buf ( n21956 , n21955 );
buf ( n21957 , n21956 );
nand ( n21958 , n21952 , n21957 );
buf ( n21959 , n21958 );
buf ( n21960 , n21959 );
and ( n21961 , n21943 , n21960 );
and ( n21962 , n21937 , n21942 );
or ( n21963 , n21961 , n21962 );
buf ( n21964 , n21963 );
buf ( n21965 , n21964 );
xor ( n21966 , n21919 , n21965 );
buf ( n21967 , n840 );
buf ( n21968 , n888 );
xor ( n21969 , n21967 , n21968 );
buf ( n21970 , n21969 );
buf ( n21971 , n21970 );
not ( n21972 , n21971 );
buf ( n21973 , n20358 );
not ( n21974 , n21973 );
or ( n21975 , n21972 , n21974 );
buf ( n21976 , n20362 );
buf ( n21977 , n21976 );
buf ( n21978 , n21746 );
nand ( n21979 , n21977 , n21978 );
buf ( n21980 , n21979 );
buf ( n21981 , n21980 );
nand ( n21982 , n21975 , n21981 );
buf ( n21983 , n21982 );
buf ( n21984 , n21983 );
not ( n21985 , n21984 );
and ( n21986 , n848 , n880 );
not ( n21987 , n848 );
and ( n21988 , n21987 , n18844 );
nor ( n21989 , n21986 , n21988 );
buf ( n21990 , n21989 );
not ( n21991 , n21990 );
buf ( n21992 , n18850 );
not ( n21993 , n21992 );
or ( n21994 , n21991 , n21993 );
buf ( n21995 , n20325 );
buf ( n21996 , n21800 );
nand ( n21997 , n21995 , n21996 );
buf ( n21998 , n21997 );
buf ( n21999 , n21998 );
nand ( n22000 , n21994 , n21999 );
buf ( n22001 , n22000 );
buf ( n22002 , n22001 );
not ( n22003 , n22002 );
or ( n22004 , n21985 , n22003 );
buf ( n22005 , n22001 );
not ( n22006 , n22005 );
buf ( n22007 , n22006 );
buf ( n22008 , n22007 );
not ( n22009 , n22008 );
buf ( n22010 , n21983 );
not ( n22011 , n22010 );
buf ( n22012 , n22011 );
buf ( n22013 , n22012 );
not ( n22014 , n22013 );
or ( n22015 , n22009 , n22014 );
buf ( n22016 , n850 );
buf ( n22017 , n878 );
xor ( n22018 , n22016 , n22017 );
buf ( n22019 , n22018 );
buf ( n22020 , n22019 );
not ( n22021 , n22020 );
buf ( n22022 , n19259 );
not ( n22023 , n22022 );
or ( n22024 , n22021 , n22023 );
buf ( n22025 , n19265 );
buf ( n22026 , n21837 );
nand ( n22027 , n22025 , n22026 );
buf ( n22028 , n22027 );
buf ( n22029 , n22028 );
nand ( n22030 , n22024 , n22029 );
buf ( n22031 , n22030 );
buf ( n22032 , n22031 );
nand ( n22033 , n22015 , n22032 );
buf ( n22034 , n22033 );
buf ( n22035 , n22034 );
nand ( n22036 , n22004 , n22035 );
buf ( n22037 , n22036 );
buf ( n22038 , n22037 );
and ( n22039 , n21966 , n22038 );
and ( n22040 , n21919 , n21965 );
or ( n22041 , n22039 , n22040 );
buf ( n22042 , n22041 );
not ( n22043 , n22042 );
xor ( n22044 , n21642 , n21703 );
xor ( n22045 , n22044 , n21737 );
buf ( n22046 , n22045 );
not ( n22047 , n22046 );
not ( n22048 , n22047 );
not ( n22049 , n22048 );
or ( n22050 , n22043 , n22049 );
not ( n22051 , n22042 );
not ( n22052 , n22051 );
not ( n22053 , n22047 );
or ( n22054 , n22052 , n22053 );
not ( n22055 , n21789 );
and ( n22056 , n21770 , n21754 );
not ( n22057 , n21770 );
and ( n22058 , n22057 , n21755 );
nor ( n22059 , n22056 , n22058 );
not ( n22060 , n22059 );
or ( n22061 , n22055 , n22060 );
or ( n22062 , n21789 , n22059 );
nand ( n22063 , n22061 , n22062 );
buf ( n22064 , n22063 );
not ( n22065 , n22064 );
not ( n22066 , n21668 );
not ( n22067 , n21654 );
or ( n22068 , n22066 , n22067 );
nand ( n22069 , n21674 , n21677 );
nand ( n22070 , n22068 , n22069 );
not ( n22071 , n21696 );
and ( n22072 , n22070 , n22071 );
not ( n22073 , n22070 );
and ( n22074 , n22073 , n21696 );
nor ( n22075 , n22072 , n22074 );
not ( n22076 , n22075 );
buf ( n22077 , n22076 );
not ( n22078 , n22077 );
or ( n22079 , n22065 , n22078 );
xor ( n22080 , n21849 , n21827 );
xor ( n22081 , n22080 , n21812 );
buf ( n22082 , n22081 );
nand ( n22083 , n22079 , n22082 );
buf ( n22084 , n22083 );
buf ( n22085 , n22084 );
buf ( n22086 , n22063 );
not ( n22087 , n22086 );
not ( n22088 , n22076 );
buf ( n22089 , n22088 );
nand ( n22090 , n22087 , n22089 );
buf ( n22091 , n22090 );
buf ( n22092 , n22091 );
nand ( n22093 , n22085 , n22092 );
buf ( n22094 , n22093 );
nand ( n22095 , n22054 , n22094 );
nand ( n22096 , n22050 , n22095 );
buf ( n22097 , n22096 );
or ( n22098 , n21916 , n22097 );
xor ( n22099 , n21584 , n21587 );
xor ( n22100 , n22099 , n21624 );
buf ( n22101 , n22100 );
buf ( n22102 , n22101 );
nand ( n22103 , n22098 , n22102 );
buf ( n22104 , n22103 );
buf ( n22105 , n22104 );
buf ( n22106 , n22096 );
buf ( n22107 , n21915 );
nand ( n22108 , n22106 , n22107 );
buf ( n22109 , n22108 );
buf ( n22110 , n22109 );
nand ( n22111 , n22105 , n22110 );
buf ( n22112 , n22111 );
buf ( n22113 , n22112 );
and ( n22114 , n21633 , n22113 );
and ( n22115 , n21546 , n21632 );
or ( n22116 , n22114 , n22115 );
buf ( n22117 , n22116 );
buf ( n22118 , n22117 );
not ( n22119 , n22118 );
buf ( n22120 , n22119 );
buf ( n22121 , n22120 );
not ( n22122 , n22121 );
or ( n22123 , n21192 , n22122 );
xor ( n22124 , n21564 , n21579 );
and ( n22125 , n22124 , n21629 );
and ( n22126 , n21564 , n21579 );
or ( n22127 , n22125 , n22126 );
buf ( n22128 , n22127 );
buf ( n22129 , n22128 );
buf ( n22130 , n860 );
buf ( n22131 , n864 );
and ( n22132 , n22130 , n22131 );
buf ( n22133 , n22132 );
buf ( n22134 , n22133 );
buf ( n22135 , n21029 );
not ( n22136 , n22135 );
buf ( n22137 , n20243 );
not ( n22138 , n22137 );
or ( n22139 , n22136 , n22138 );
buf ( n22140 , n20246 );
xor ( n22141 , n876 , n846 );
buf ( n22142 , n22141 );
nand ( n22143 , n22140 , n22142 );
buf ( n22144 , n22143 );
buf ( n22145 , n22144 );
nand ( n22146 , n22139 , n22145 );
buf ( n22147 , n22146 );
buf ( n22148 , n22147 );
xor ( n22149 , n22134 , n22148 );
not ( n22150 , n21017 );
not ( n22151 , n21013 );
not ( n22152 , n22151 );
or ( n22153 , n22150 , n22152 );
buf ( n22154 , n19265 );
buf ( n22155 , n844 );
buf ( n22156 , n878 );
xor ( n22157 , n22155 , n22156 );
buf ( n22158 , n22157 );
buf ( n22159 , n22158 );
nand ( n22160 , n22154 , n22159 );
buf ( n22161 , n22160 );
nand ( n22162 , n22153 , n22161 );
buf ( n22163 , n22162 );
xor ( n22164 , n22149 , n22163 );
buf ( n22165 , n22164 );
buf ( n22166 , n22165 );
buf ( n22167 , n20164 );
not ( n22168 , n22167 );
buf ( n22169 , n21762 );
not ( n22170 , n22169 );
or ( n22171 , n22168 , n22170 );
buf ( n22172 , n892 );
nand ( n22173 , n22171 , n22172 );
buf ( n22174 , n22173 );
buf ( n22175 , n22174 );
buf ( n22176 , n20852 );
not ( n22177 , n22176 );
buf ( n22178 , n21817 );
not ( n22179 , n22178 );
or ( n22180 , n22177 , n22179 );
buf ( n22181 , n20255 );
buf ( n22182 , n836 );
buf ( n22183 , n886 );
xor ( n22184 , n22182 , n22183 );
buf ( n22185 , n22184 );
buf ( n22186 , n22185 );
nand ( n22187 , n22181 , n22186 );
buf ( n22188 , n22187 );
buf ( n22189 , n22188 );
nand ( n22190 , n22180 , n22189 );
buf ( n22191 , n22190 );
buf ( n22192 , n22191 );
xor ( n22193 , n22175 , n22192 );
buf ( n22194 , n20868 );
not ( n22195 , n22194 );
buf ( n22196 , n21441 );
not ( n22197 , n22196 );
or ( n22198 , n22195 , n22197 );
buf ( n22199 , n20869 );
buf ( n22200 , n832 );
buf ( n22201 , n890 );
xor ( n22202 , n22200 , n22201 );
buf ( n22203 , n22202 );
buf ( n22204 , n22203 );
nand ( n22205 , n22199 , n22204 );
buf ( n22206 , n22205 );
buf ( n22207 , n22206 );
nand ( n22208 , n22198 , n22207 );
buf ( n22209 , n22208 );
buf ( n22210 , n22209 );
xor ( n22211 , n22193 , n22210 );
buf ( n22212 , n22211 );
buf ( n22213 , n22212 );
xor ( n22214 , n22166 , n22213 );
buf ( n22215 , n21086 );
buf ( n22216 , n22215 );
not ( n22217 , n22216 );
buf ( n22218 , n21114 );
not ( n22219 , n22218 );
or ( n22220 , n22217 , n22219 );
buf ( n22221 , n21079 );
nand ( n22222 , n22220 , n22221 );
buf ( n22223 , n22222 );
buf ( n22224 , n22223 );
not ( n22225 , n22215 );
nand ( n22226 , n22225 , n21111 );
buf ( n22227 , n22226 );
nand ( n22228 , n22224 , n22227 );
buf ( n22229 , n22228 );
buf ( n22230 , n22229 );
xor ( n22231 , n22214 , n22230 );
buf ( n22232 , n22231 );
buf ( n22233 , n22232 );
buf ( n22234 , n21073 );
not ( n22235 , n22234 );
buf ( n22236 , n18923 );
buf ( n22237 , n18927 );
nor ( n22238 , n22236 , n22237 );
buf ( n22239 , n22238 );
buf ( n22240 , n22239 );
not ( n22241 , n22240 );
or ( n22242 , n22235 , n22241 );
buf ( n22243 , n18938 );
buf ( n22244 , n856 );
buf ( n22245 , n866 );
xor ( n22246 , n22244 , n22245 );
buf ( n22247 , n22246 );
buf ( n22248 , n22247 );
nand ( n22249 , n22243 , n22248 );
buf ( n22250 , n22249 );
buf ( n22251 , n22250 );
nand ( n22252 , n22242 , n22251 );
buf ( n22253 , n22252 );
buf ( n22254 , n22253 );
not ( n22255 , n20961 );
not ( n22256 , n18884 );
or ( n22257 , n22255 , n22256 );
buf ( n22258 , n20786 );
xor ( n22259 , n868 , n854 );
buf ( n22260 , n22259 );
nand ( n22261 , n22258 , n22260 );
buf ( n22262 , n22261 );
nand ( n22263 , n22257 , n22262 );
buf ( n22264 , n22263 );
xor ( n22265 , n22254 , n22264 );
buf ( n22266 , n21084 );
not ( n22267 , n22266 );
buf ( n22268 , n18850 );
not ( n22269 , n22268 );
or ( n22270 , n22267 , n22269 );
buf ( n22271 , n21083 );
buf ( n22272 , n22271 );
xor ( n22273 , n880 , n842 );
buf ( n22274 , n22273 );
nand ( n22275 , n22272 , n22274 );
buf ( n22276 , n22275 );
buf ( n22277 , n22276 );
nand ( n22278 , n22270 , n22277 );
buf ( n22279 , n22278 );
buf ( n22280 , n22279 );
xor ( n22281 , n22265 , n22280 );
buf ( n22282 , n22281 );
buf ( n22283 , n22282 );
not ( n22284 , n22283 );
not ( n22285 , n20984 );
not ( n22286 , n20197 );
or ( n22287 , n22285 , n22286 );
buf ( n22288 , n19568 );
buf ( n22289 , n840 );
buf ( n22290 , n882 );
xor ( n22291 , n22289 , n22290 );
buf ( n22292 , n22291 );
buf ( n22293 , n22292 );
nand ( n22294 , n22288 , n22293 );
buf ( n22295 , n22294 );
nand ( n22296 , n22287 , n22295 );
not ( n22297 , n20884 );
not ( n22298 , n20349 );
nand ( n22299 , n889 , n890 );
not ( n22300 , n22299 );
not ( n22301 , n22300 );
or ( n22302 , n22298 , n22301 );
nand ( n22303 , n22302 , n20356 );
not ( n22304 , n22303 );
or ( n22305 , n22297 , n22304 );
buf ( n22306 , n20363 );
buf ( n22307 , n834 );
buf ( n22308 , n888 );
xor ( n22309 , n22307 , n22308 );
buf ( n22310 , n22309 );
buf ( n22311 , n22310 );
nand ( n22312 , n22306 , n22311 );
buf ( n22313 , n22312 );
nand ( n22314 , n22305 , n22313 );
not ( n22315 , n22314 );
xor ( n22316 , n22296 , n22315 );
buf ( n22317 , n20971 );
not ( n22318 , n22317 );
buf ( n22319 , n19122 );
not ( n22320 , n22319 );
or ( n22321 , n22318 , n22320 );
buf ( n22322 , n19131 );
xor ( n22323 , n870 , n852 );
buf ( n22324 , n22323 );
nand ( n22325 , n22322 , n22324 );
buf ( n22326 , n22325 );
buf ( n22327 , n22326 );
nand ( n22328 , n22321 , n22327 );
buf ( n22329 , n22328 );
xor ( n22330 , n22316 , n22329 );
buf ( n22331 , n22330 );
not ( n22332 , n22331 );
and ( n22333 , n22284 , n22332 );
buf ( n22334 , n22282 );
buf ( n22335 , n22330 );
and ( n22336 , n22334 , n22335 );
nor ( n22337 , n22333 , n22336 );
buf ( n22338 , n22337 );
buf ( n22339 , n22338 );
not ( n22340 , n20895 );
not ( n22341 , n20736 );
or ( n22342 , n22340 , n22341 );
buf ( n22343 , n18981 );
buf ( n22344 , n848 );
buf ( n22345 , n874 );
xor ( n22346 , n22344 , n22345 );
buf ( n22347 , n22346 );
buf ( n22348 , n22347 );
nand ( n22349 , n22343 , n22348 );
buf ( n22350 , n22349 );
nand ( n22351 , n22342 , n22350 );
buf ( n22352 , n22351 );
not ( n22353 , n22352 );
buf ( n22354 , n21045 );
not ( n22355 , n22354 );
buf ( n22356 , n20430 );
not ( n22357 , n22356 );
or ( n22358 , n22355 , n22357 );
buf ( n22359 , n20700 );
buf ( n22360 , n838 );
buf ( n22361 , n884 );
xor ( n22362 , n22360 , n22361 );
buf ( n22363 , n22362 );
buf ( n22364 , n22363 );
nand ( n22365 , n22359 , n22364 );
buf ( n22366 , n22365 );
buf ( n22367 , n22366 );
nand ( n22368 , n22358 , n22367 );
buf ( n22369 , n22368 );
buf ( n22370 , n22369 );
not ( n22371 , n22370 );
buf ( n22372 , n22371 );
buf ( n22373 , n22372 );
not ( n22374 , n22373 );
or ( n22375 , n22353 , n22374 );
buf ( n22376 , n22351 );
not ( n22377 , n22376 );
buf ( n22378 , n22369 );
nand ( n22379 , n22377 , n22378 );
buf ( n22380 , n22379 );
buf ( n22381 , n22380 );
nand ( n22382 , n22375 , n22381 );
buf ( n22383 , n22382 );
buf ( n22384 , n22383 );
buf ( n22385 , n20914 );
not ( n22386 , n22385 );
buf ( n22387 , n20211 );
not ( n22388 , n22387 );
or ( n22389 , n22386 , n22388 );
buf ( n22390 , n850 );
buf ( n22391 , n872 );
xor ( n22392 , n22390 , n22391 );
buf ( n22393 , n22392 );
buf ( n22394 , n22393 );
buf ( n22395 , n19234 );
nand ( n22396 , n22394 , n22395 );
buf ( n22397 , n22396 );
buf ( n22398 , n22397 );
nand ( n22399 , n22389 , n22398 );
buf ( n22400 , n22399 );
buf ( n22401 , n22400 );
not ( n22402 , n22401 );
buf ( n22403 , n22402 );
buf ( n22404 , n22403 );
and ( n22405 , n22384 , n22404 );
not ( n22406 , n22384 );
buf ( n22407 , n22400 );
and ( n22408 , n22406 , n22407 );
nor ( n22409 , n22405 , n22408 );
buf ( n22410 , n22409 );
buf ( n22411 , n22410 );
and ( n22412 , n22339 , n22411 );
not ( n22413 , n22339 );
buf ( n22414 , n22410 );
not ( n22415 , n22414 );
buf ( n22416 , n22415 );
buf ( n22417 , n22416 );
and ( n22418 , n22413 , n22417 );
nor ( n22419 , n22412 , n22418 );
buf ( n22420 , n22419 );
buf ( n22421 , n22420 );
xor ( n22422 , n22233 , n22421 );
xor ( n22423 , n20597 , n20609 );
and ( n22424 , n22423 , n20670 );
and ( n22425 , n20597 , n20609 );
or ( n22426 , n22424 , n22425 );
buf ( n22427 , n22426 );
buf ( n22428 , n22427 );
buf ( n22429 , n20607 );
buf ( n22430 , n21105 );
not ( n22431 , n22430 );
buf ( n22432 , n19013 );
not ( n22433 , n22432 );
or ( n22434 , n22431 , n22433 );
buf ( n22435 , n19030 );
buf ( n22436 , n858 );
buf ( n22437 , n864 );
xor ( n22438 , n22436 , n22437 );
buf ( n22439 , n22438 );
buf ( n22440 , n22439 );
nand ( n22441 , n22435 , n22440 );
buf ( n22442 , n22441 );
buf ( n22443 , n22442 );
nand ( n22444 , n22434 , n22443 );
buf ( n22445 , n22444 );
buf ( n22446 , n22445 );
xor ( n22447 , n22429 , n22446 );
xor ( n22448 , n20841 , n20858 );
and ( n22449 , n22448 , n20873 );
and ( n22450 , n20841 , n20858 );
or ( n22451 , n22449 , n22450 );
buf ( n22452 , n22451 );
xor ( n22453 , n22447 , n22452 );
buf ( n22454 , n22453 );
buf ( n22455 , n22454 );
xor ( n22456 , n22428 , n22455 );
xor ( n22457 , n20471 , n20516 );
and ( n22458 , n22457 , n20584 );
and ( n22459 , n20471 , n20516 );
or ( n22460 , n22458 , n22459 );
buf ( n22461 , n22460 );
buf ( n22462 , n22461 );
xor ( n22463 , n22456 , n22462 );
buf ( n22464 , n22463 );
buf ( n22465 , n22464 );
xor ( n22466 , n22422 , n22465 );
buf ( n22467 , n22466 );
buf ( n22468 , n22467 );
xor ( n22469 , n22129 , n22468 );
buf ( n22470 , n20386 );
buf ( n22471 , n20393 );
and ( n22472 , n22470 , n22471 );
not ( n22473 , n22470 );
buf ( n22474 , n20185 );
and ( n22475 , n22473 , n22474 );
nor ( n22476 , n22472 , n22475 );
buf ( n22477 , n22476 );
buf ( n22478 , n22477 );
not ( n22479 , n20586 );
buf ( n22480 , n22479 );
and ( n22481 , n22478 , n22480 );
not ( n22482 , n22478 );
buf ( n22483 , n20586 );
and ( n22484 , n22482 , n22483 );
nor ( n22485 , n22481 , n22484 );
buf ( n22486 , n22485 );
buf ( n22487 , n22486 );
not ( n22488 , n22487 );
buf ( n22489 , n22488 );
not ( n22490 , n22489 );
buf ( n22491 , n20672 );
buf ( n22492 , n20810 );
xor ( n22493 , n22491 , n22492 );
buf ( n22494 , n20829 );
xnor ( n22495 , n22493 , n22494 );
buf ( n22496 , n22495 );
buf ( n22497 , n22496 );
not ( n22498 , n22497 );
buf ( n22499 , n22498 );
not ( n22500 , n22499 );
or ( n22501 , n22490 , n22500 );
not ( n22502 , n22486 );
not ( n22503 , n22496 );
or ( n22504 , n22502 , n22503 );
xor ( n22505 , n21638 , n21741 );
and ( n22506 , n22505 , n21914 );
and ( n22507 , n21638 , n21741 );
or ( n22508 , n22506 , n22507 );
nand ( n22509 , n22504 , n22508 );
nand ( n22510 , n22501 , n22509 );
buf ( n22511 , n22510 );
xor ( n22512 , n22469 , n22511 );
buf ( n22513 , n22512 );
buf ( n22514 , n22513 );
nand ( n22515 , n22123 , n22514 );
buf ( n22516 , n22515 );
buf ( n22517 , n22516 );
buf ( n22518 , n21190 );
not ( n22519 , n22518 );
buf ( n22520 , n22117 );
nand ( n22521 , n22519 , n22520 );
buf ( n22522 , n22521 );
buf ( n22523 , n22522 );
nand ( n22524 , n22517 , n22523 );
buf ( n22525 , n22524 );
buf ( n22526 , n22525 );
buf ( n22527 , n22496 );
buf ( n22528 , n22527 );
buf ( n22529 , n22528 );
buf ( n22530 , n22529 );
buf ( n22531 , n22486 );
not ( n22532 , n22531 );
buf ( n22533 , n22508 );
not ( n22534 , n22533 );
and ( n22535 , n22532 , n22534 );
buf ( n22536 , n22486 );
buf ( n22537 , n22508 );
and ( n22538 , n22536 , n22537 );
nor ( n22539 , n22535 , n22538 );
buf ( n22540 , n22539 );
buf ( n22541 , n22540 );
xor ( n22542 , n22530 , n22541 );
buf ( n22543 , n22542 );
buf ( n22544 , n22543 );
xor ( n22545 , n21546 , n21632 );
xor ( n22546 , n22545 , n22113 );
buf ( n22547 , n22546 );
buf ( n22548 , n22547 );
xor ( n22549 , n22544 , n22548 );
xor ( n22550 , n21899 , n21883 );
not ( n22551 , n21869 );
xor ( n22552 , n22550 , n22551 );
buf ( n22553 , n22552 );
not ( n22554 , n22553 );
buf ( n22555 , n22554 );
not ( n22556 , n22555 );
not ( n22557 , n21720 );
not ( n22558 , n21712 );
or ( n22559 , n22557 , n22558 );
or ( n22560 , n21712 , n21720 );
nand ( n22561 , n22559 , n22560 );
not ( n22562 , n21733 );
and ( n22563 , n22561 , n22562 );
not ( n22564 , n22561 );
and ( n22565 , n22564 , n21733 );
nor ( n22566 , n22563 , n22565 );
not ( n22567 , n22566 );
not ( n22568 , n22567 );
or ( n22569 , n22556 , n22568 );
not ( n22570 , n22566 );
not ( n22571 , n22552 );
or ( n22572 , n22570 , n22571 );
xor ( n22573 , n870 , n859 );
buf ( n22574 , n22573 );
not ( n22575 , n22574 );
buf ( n22576 , n20805 );
not ( n22577 , n22576 );
or ( n22578 , n22575 , n22577 );
buf ( n22579 , n19114 );
buf ( n22580 , n21367 );
nand ( n22581 , n22579 , n22580 );
buf ( n22582 , n22581 );
buf ( n22583 , n22582 );
nand ( n22584 , n22578 , n22583 );
buf ( n22585 , n22584 );
not ( n22586 , n22585 );
buf ( n22587 , n847 );
buf ( n22588 , n882 );
xor ( n22589 , n22587 , n22588 );
buf ( n22590 , n22589 );
buf ( n22591 , n22590 );
not ( n22592 , n22591 );
buf ( n22593 , n19580 );
not ( n22594 , n22593 );
or ( n22595 , n22592 , n22594 );
buf ( n22596 , n19909 );
buf ( n22597 , n21344 );
nand ( n22598 , n22596 , n22597 );
buf ( n22599 , n22598 );
buf ( n22600 , n22599 );
nand ( n22601 , n22595 , n22600 );
buf ( n22602 , n22601 );
not ( n22603 , n22602 );
or ( n22604 , n22586 , n22603 );
buf ( n22605 , n22602 );
buf ( n22606 , n22585 );
or ( n22607 , n22605 , n22606 );
buf ( n22608 , n857 );
buf ( n22609 , n872 );
xor ( n22610 , n22608 , n22609 );
buf ( n22611 , n22610 );
buf ( n22612 , n22611 );
not ( n22613 , n22612 );
buf ( n22614 , n20211 );
not ( n22615 , n22614 );
or ( n22616 , n22613 , n22615 );
buf ( n22617 , n19234 );
buf ( n22618 , n21415 );
nand ( n22619 , n22617 , n22618 );
buf ( n22620 , n22619 );
buf ( n22621 , n22620 );
nand ( n22622 , n22616 , n22621 );
buf ( n22623 , n22622 );
buf ( n22624 , n22623 );
nand ( n22625 , n22607 , n22624 );
buf ( n22626 , n22625 );
nand ( n22627 , n22604 , n22626 );
buf ( n22628 , n851 );
buf ( n22629 , n878 );
xor ( n22630 , n22628 , n22629 );
buf ( n22631 , n22630 );
buf ( n22632 , n22631 );
not ( n22633 , n22632 );
buf ( n22634 , n19259 );
not ( n22635 , n22634 );
or ( n22636 , n22633 , n22635 );
buf ( n22637 , n19265 );
buf ( n22638 , n22019 );
nand ( n22639 , n22637 , n22638 );
buf ( n22640 , n22639 );
buf ( n22641 , n22640 );
nand ( n22642 , n22636 , n22641 );
buf ( n22643 , n22642 );
not ( n22644 , n22643 );
buf ( n22645 , n843 );
buf ( n22646 , n886 );
xor ( n22647 , n22645 , n22646 );
buf ( n22648 , n22647 );
nand ( n22649 , n22648 , n20521 );
nand ( n22650 , n20255 , n21490 );
buf ( n22651 , n21461 );
buf ( n22652 , n20246 );
nand ( n22653 , n22651 , n22652 );
buf ( n22654 , n22653 );
buf ( n22655 , n853 );
buf ( n22656 , n876 );
xor ( n22657 , n22655 , n22656 );
buf ( n22658 , n22657 );
nand ( n22659 , n19153 , n22658 );
nand ( n22660 , n22649 , n22650 , n22654 , n22659 );
not ( n22661 , n22660 );
or ( n22662 , n22644 , n22661 );
and ( n22663 , n22659 , n22654 );
not ( n22664 , n22663 );
nand ( n22665 , n22649 , n22650 );
nand ( n22666 , n22664 , n22665 );
nand ( n22667 , n22662 , n22666 );
nor ( n22668 , n22627 , n22667 );
buf ( n22669 , n845 );
buf ( n22670 , n884 );
xor ( n22671 , n22669 , n22670 );
buf ( n22672 , n22671 );
buf ( n22673 , n22672 );
not ( n22674 , n22673 );
buf ( n22675 , n20694 );
not ( n22676 , n22675 );
or ( n22677 , n22674 , n22676 );
buf ( n22678 , n20700 );
buf ( n22679 , n21399 );
nand ( n22680 , n22678 , n22679 );
buf ( n22681 , n22680 );
buf ( n22682 , n22681 );
nand ( n22683 , n22677 , n22682 );
buf ( n22684 , n22683 );
not ( n22685 , n22684 );
buf ( n22686 , n839 );
buf ( n22687 , n890 );
xor ( n22688 , n22686 , n22687 );
buf ( n22689 , n22688 );
buf ( n22690 , n22689 );
not ( n22691 , n22690 );
buf ( n22692 , n21441 );
not ( n22693 , n22692 );
or ( n22694 , n22691 , n22693 );
buf ( n22695 , n20869 );
buf ( n22696 , n21432 );
nand ( n22697 , n22695 , n22696 );
buf ( n22698 , n22697 );
buf ( n22699 , n22698 );
nand ( n22700 , n22694 , n22699 );
buf ( n22701 , n22700 );
not ( n22702 , n22701 );
or ( n22703 , n22685 , n22702 );
buf ( n22704 , n22701 );
buf ( n22705 , n22684 );
or ( n22706 , n22704 , n22705 );
buf ( n22707 , n855 );
buf ( n22708 , n874 );
xor ( n22709 , n22707 , n22708 );
buf ( n22710 , n22709 );
buf ( n22711 , n22710 );
not ( n22712 , n22711 );
buf ( n22713 , n20549 );
not ( n22714 , n22713 );
or ( n22715 , n22712 , n22714 );
buf ( n22716 , n20555 );
buf ( n22717 , n21505 );
nand ( n22718 , n22716 , n22717 );
buf ( n22719 , n22718 );
buf ( n22720 , n22719 );
nand ( n22721 , n22715 , n22720 );
buf ( n22722 , n22721 );
buf ( n22723 , n22722 );
nand ( n22724 , n22706 , n22723 );
buf ( n22725 , n22724 );
nand ( n22726 , n22703 , n22725 );
not ( n22727 , n22726 );
or ( n22728 , n22668 , n22727 );
nand ( n22729 , n22627 , n22667 );
nand ( n22730 , n22728 , n22729 );
nand ( n22731 , n22572 , n22730 );
nand ( n22732 , n22569 , n22731 );
buf ( n22733 , n22732 );
xor ( n22734 , n21903 , n21855 );
xor ( n22735 , n22734 , n21795 );
buf ( n22736 , n22735 );
xor ( n22737 , n22733 , n22736 );
xor ( n22738 , n21614 , n21596 );
xor ( n22739 , n22738 , n21621 );
buf ( n22740 , n22739 );
and ( n22741 , n22737 , n22740 );
and ( n22742 , n22733 , n22736 );
or ( n22743 , n22741 , n22742 );
buf ( n22744 , n22743 );
buf ( n22745 , n22744 );
xor ( n22746 , n21218 , n21194 );
xnor ( n22747 , n22746 , n21542 );
buf ( n22748 , n22747 );
xor ( n22749 , n22745 , n22748 );
xor ( n22750 , n21237 , n21314 );
xor ( n22751 , n22750 , n21538 );
buf ( n22752 , n22751 );
buf ( n22753 , n22752 );
buf ( n22754 , n863 );
buf ( n22755 , n867 );
or ( n22756 , n22754 , n22755 );
buf ( n22757 , n868 );
nand ( n22758 , n22756 , n22757 );
buf ( n22759 , n22758 );
buf ( n22760 , n22759 );
buf ( n22761 , n863 );
buf ( n22762 , n867 );
nand ( n22763 , n22761 , n22762 );
buf ( n22764 , n22763 );
buf ( n22765 , n22764 );
buf ( n22766 , n866 );
and ( n22767 , n22760 , n22765 , n22766 );
buf ( n22768 , n22767 );
buf ( n22769 , n22768 );
buf ( n22770 , n835 );
buf ( n22771 , n894 );
xor ( n22772 , n22770 , n22771 );
buf ( n22773 , n22772 );
buf ( n22774 , n22773 );
not ( n22775 , n22774 );
not ( n22776 , n21296 );
buf ( n22777 , n22776 );
not ( n22778 , n22777 );
or ( n22779 , n22775 , n22778 );
buf ( n22780 , n21931 );
buf ( n22781 , n895 );
nand ( n22782 , n22780 , n22781 );
buf ( n22783 , n22782 );
buf ( n22784 , n22783 );
nand ( n22785 , n22779 , n22784 );
buf ( n22786 , n22785 );
buf ( n22787 , n22786 );
and ( n22788 , n22769 , n22787 );
buf ( n22789 , n22788 );
buf ( n22790 , n22789 );
buf ( n22791 , n862 );
buf ( n22792 , n866 );
xor ( n22793 , n22791 , n22792 );
buf ( n22794 , n22793 );
buf ( n22795 , n22794 );
not ( n22796 , n22795 );
buf ( n22797 , n18931 );
not ( n22798 , n22797 );
or ( n22799 , n22796 , n22798 );
buf ( n22800 , n18944 );
buf ( n22801 , n21684 );
nand ( n22802 , n22800 , n22801 );
buf ( n22803 , n22802 );
buf ( n22804 , n22803 );
nand ( n22805 , n22799 , n22804 );
buf ( n22806 , n22805 );
buf ( n22807 , n22806 );
xor ( n22808 , n22790 , n22807 );
buf ( n22809 , n837 );
buf ( n22810 , n892 );
xor ( n22811 , n22809 , n22810 );
buf ( n22812 , n22811 );
not ( n22813 , n22812 );
not ( n22814 , n20599 );
or ( n22815 , n22813 , n22814 );
buf ( n22816 , n20167 );
buf ( n22817 , n22816 );
buf ( n22818 , n22817 );
buf ( n22819 , n22818 );
buf ( n22820 , n21947 );
nand ( n22821 , n22819 , n22820 );
buf ( n22822 , n22821 );
nand ( n22823 , n22815 , n22822 );
not ( n22824 , n22823 );
not ( n22825 , n21083 );
not ( n22826 , n21989 );
or ( n22827 , n22825 , n22826 );
not ( n22828 , n18848 );
xor ( n22829 , n880 , n849 );
and ( n22830 , n881 , n880 );
not ( n22831 , n881 );
and ( n22832 , n22831 , n18844 );
nor ( n22833 , n22830 , n22832 );
nand ( n22834 , n22828 , n22829 , n22833 );
nand ( n22835 , n22827 , n22834 );
not ( n22836 , n22835 );
or ( n22837 , n22824 , n22836 );
nor ( n22838 , n22823 , n22835 );
buf ( n22839 , n20363 );
buf ( n22840 , n21970 );
nand ( n22841 , n22839 , n22840 );
buf ( n22842 , n22841 );
buf ( n22843 , n841 );
buf ( n22844 , n888 );
xor ( n22845 , n22843 , n22844 );
buf ( n22846 , n22845 );
nand ( n22847 , n22846 , n22303 );
and ( n22848 , n22842 , n22847 );
or ( n22849 , n22838 , n22848 );
nand ( n22850 , n22837 , n22849 );
buf ( n22851 , n22850 );
and ( n22852 , n22808 , n22851 );
and ( n22853 , n22790 , n22807 );
or ( n22854 , n22852 , n22853 );
buf ( n22855 , n22854 );
buf ( n22856 , n22855 );
xor ( n22857 , n21919 , n21965 );
xor ( n22858 , n22857 , n22038 );
buf ( n22859 , n22858 );
buf ( n22860 , n22859 );
xor ( n22861 , n22856 , n22860 );
buf ( n22862 , n21526 );
buf ( n22863 , n21394 );
xor ( n22864 , n22862 , n22863 );
buf ( n22865 , n22864 );
buf ( n22866 , n22865 );
buf ( n22867 , n21455 );
xor ( n22868 , n22866 , n22867 );
buf ( n22869 , n22868 );
buf ( n22870 , n22869 );
and ( n22871 , n22861 , n22870 );
and ( n22872 , n22856 , n22860 );
or ( n22873 , n22871 , n22872 );
buf ( n22874 , n22873 );
buf ( n22875 , n22874 );
xor ( n22876 , n22753 , n22875 );
xor ( n22877 , n21411 , n21427 );
xor ( n22878 , n22877 , n21452 );
xor ( n22879 , n21937 , n21942 );
xor ( n22880 , n22879 , n21960 );
buf ( n22881 , n22880 );
or ( n22882 , n22878 , n22881 );
xor ( n22883 , n21360 , n21338 );
xnor ( n22884 , n22883 , n21383 );
nand ( n22885 , n22882 , n22884 );
buf ( n22886 , n22885 );
buf ( n22887 , n22878 );
buf ( n22888 , n22881 );
nand ( n22889 , n22887 , n22888 );
buf ( n22890 , n22889 );
buf ( n22891 , n22890 );
nand ( n22892 , n22886 , n22891 );
buf ( n22893 , n22892 );
buf ( n22894 , n22893 );
buf ( n22895 , n21524 );
not ( n22896 , n22895 );
buf ( n22897 , n22896 );
not ( n22898 , n21497 );
not ( n22899 , n21499 );
or ( n22900 , n22898 , n22899 );
or ( n22901 , n21497 , n21499 );
nand ( n22902 , n22900 , n22901 );
or ( n22903 , n22897 , n22902 );
nand ( n22904 , n22902 , n22897 );
nand ( n22905 , n22903 , n22904 );
not ( n22906 , n22905 );
buf ( n22907 , n861 );
buf ( n22908 , n868 );
xor ( n22909 , n22907 , n22908 );
buf ( n22910 , n22909 );
buf ( n22911 , n22910 );
not ( n22912 , n22911 );
buf ( n22913 , n18887 );
not ( n22914 , n22913 );
or ( n22915 , n22912 , n22914 );
buf ( n22916 , n20786 );
buf ( n22917 , n22916 );
buf ( n22918 , n21319 );
nand ( n22919 , n22917 , n22918 );
buf ( n22920 , n22919 );
buf ( n22921 , n22920 );
nand ( n22922 , n22915 , n22921 );
buf ( n22923 , n22922 );
buf ( n22924 , n22923 );
not ( n22925 , n22924 );
xor ( n22926 , n22769 , n22787 );
buf ( n22927 , n22926 );
buf ( n22928 , n22927 );
not ( n22929 , n22928 );
or ( n22930 , n22925 , n22929 );
buf ( n22931 , n22910 );
not ( n22932 , n22931 );
buf ( n22933 , n18887 );
not ( n22934 , n22933 );
or ( n22935 , n22932 , n22934 );
buf ( n22936 , n22920 );
nand ( n22937 , n22935 , n22936 );
buf ( n22938 , n22937 );
buf ( n22939 , n22938 );
buf ( n22940 , n22927 );
or ( n22941 , n22939 , n22940 );
buf ( n22942 , n863 );
buf ( n22943 , n866 );
xor ( n22944 , n22942 , n22943 );
buf ( n22945 , n22944 );
not ( n22946 , n22945 );
not ( n22947 , n18931 );
or ( n22948 , n22946 , n22947 );
buf ( n22949 , n18944 );
buf ( n22950 , n22794 );
nand ( n22951 , n22949 , n22950 );
buf ( n22952 , n22951 );
nand ( n22953 , n22948 , n22952 );
buf ( n22954 , n22953 );
nand ( n22955 , n22941 , n22954 );
buf ( n22956 , n22955 );
buf ( n22957 , n22956 );
nand ( n22958 , n22930 , n22957 );
buf ( n22959 , n22958 );
not ( n22960 , n22959 );
not ( n22961 , n22960 );
or ( n22962 , n22906 , n22961 );
buf ( n22963 , n21983 );
not ( n22964 , n22963 );
buf ( n22965 , n22007 );
not ( n22966 , n22965 );
or ( n22967 , n22964 , n22966 );
buf ( n22968 , n22007 );
buf ( n22969 , n21983 );
or ( n22970 , n22968 , n22969 );
nand ( n22971 , n22967 , n22970 );
buf ( n22972 , n22971 );
xor ( n22973 , n22031 , n22972 );
nand ( n22974 , n22962 , n22973 );
buf ( n22975 , n22974 );
not ( n22976 , n22905 );
nand ( n22977 , n22959 , n22976 );
buf ( n22978 , n22977 );
nand ( n22979 , n22975 , n22978 );
buf ( n22980 , n22979 );
buf ( n22981 , n22980 );
xor ( n22982 , n22894 , n22981 );
buf ( n22983 , n22081 );
buf ( n22984 , n22075 );
not ( n22985 , n22984 );
buf ( n22986 , n22063 );
not ( n22987 , n22986 );
or ( n22988 , n22985 , n22987 );
buf ( n22989 , n22075 );
buf ( n22990 , n22063 );
or ( n22991 , n22989 , n22990 );
nand ( n22992 , n22988 , n22991 );
buf ( n22993 , n22992 );
buf ( n22994 , n22993 );
xor ( n22995 , n22983 , n22994 );
buf ( n22996 , n22995 );
buf ( n22997 , n22996 );
and ( n22998 , n22982 , n22997 );
and ( n22999 , n22894 , n22981 );
or ( n23000 , n22998 , n22999 );
buf ( n23001 , n23000 );
buf ( n23002 , n23001 );
and ( n23003 , n22876 , n23002 );
and ( n23004 , n22753 , n22875 );
or ( n23005 , n23003 , n23004 );
buf ( n23006 , n23005 );
buf ( n23007 , n23006 );
and ( n23008 , n22749 , n23007 );
and ( n23009 , n22745 , n22748 );
or ( n23010 , n23008 , n23009 );
buf ( n23011 , n23010 );
buf ( n23012 , n23011 );
xor ( n23013 , n22549 , n23012 );
buf ( n23014 , n23013 );
buf ( n23015 , n23014 );
buf ( n23016 , n862 );
buf ( n23017 , n886 );
xor ( n23018 , n23016 , n23017 );
buf ( n23019 , n23018 );
buf ( n23020 , n23019 );
not ( n23021 , n23020 );
buf ( n23022 , n21817 );
not ( n23023 , n23022 );
buf ( n23024 , n23023 );
buf ( n23025 , n23024 );
not ( n23026 , n23025 );
buf ( n23027 , n23026 );
buf ( n23028 , n23027 );
not ( n23029 , n23028 );
or ( n23030 , n23021 , n23029 );
buf ( n23031 , n20525 );
buf ( n23032 , n861 );
buf ( n23033 , n886 );
xor ( n23034 , n23032 , n23033 );
buf ( n23035 , n23034 );
buf ( n23036 , n23035 );
nand ( n23037 , n23031 , n23036 );
buf ( n23038 , n23037 );
buf ( n23039 , n23038 );
nand ( n23040 , n23030 , n23039 );
buf ( n23041 , n23040 );
buf ( n23042 , n854 );
buf ( n23043 , n894 );
xor ( n23044 , n23042 , n23043 );
buf ( n23045 , n23044 );
buf ( n23046 , n23045 );
not ( n23047 , n23046 );
buf ( n23048 , n22776 );
not ( n23049 , n23048 );
or ( n23050 , n23047 , n23049 );
buf ( n23051 , n853 );
buf ( n23052 , n894 );
xor ( n23053 , n23051 , n23052 );
buf ( n23054 , n23053 );
buf ( n23055 , n23054 );
buf ( n23056 , n895 );
nand ( n23057 , n23055 , n23056 );
buf ( n23058 , n23057 );
buf ( n23059 , n23058 );
nand ( n23060 , n23050 , n23059 );
buf ( n23061 , n23060 );
xor ( n23062 , n23041 , n23061 );
buf ( n23063 , n858 );
buf ( n23064 , n890 );
xor ( n23065 , n23063 , n23064 );
buf ( n23066 , n23065 );
buf ( n23067 , n23066 );
not ( n23068 , n23067 );
buf ( n23069 , n21441 );
not ( n23070 , n23069 );
or ( n23071 , n23068 , n23070 );
buf ( n23072 , n20869 );
buf ( n23073 , n857 );
buf ( n23074 , n890 );
xor ( n23075 , n23073 , n23074 );
buf ( n23076 , n23075 );
buf ( n23077 , n23076 );
nand ( n23078 , n23072 , n23077 );
buf ( n23079 , n23078 );
buf ( n23080 , n23079 );
nand ( n23081 , n23071 , n23080 );
buf ( n23082 , n23081 );
xor ( n23083 , n23062 , n23082 );
buf ( n23084 , n23083 );
buf ( n23085 , n859 );
buf ( n23086 , n890 );
xor ( n23087 , n23085 , n23086 );
buf ( n23088 , n23087 );
buf ( n23089 , n23088 );
not ( n23090 , n23089 );
buf ( n23091 , n21441 );
not ( n23092 , n23091 );
or ( n23093 , n23090 , n23092 );
buf ( n23094 , n20869 );
buf ( n23095 , n23094 );
buf ( n23096 , n23066 );
nand ( n23097 , n23095 , n23096 );
buf ( n23098 , n23097 );
buf ( n23099 , n23098 );
nand ( n23100 , n23093 , n23099 );
buf ( n23101 , n23100 );
buf ( n23102 , n23101 );
buf ( n23103 , n20525 );
buf ( n23104 , n863 );
nand ( n23105 , n23103 , n23104 );
buf ( n23106 , n23105 );
buf ( n23107 , n23106 );
not ( n23108 , n23107 );
buf ( n23109 , n23108 );
buf ( n23110 , n23109 );
not ( n23111 , n23110 );
not ( n23112 , n21927 );
buf ( n23113 , n856 );
buf ( n23114 , n894 );
xor ( n23115 , n23113 , n23114 );
buf ( n23116 , n23115 );
buf ( n23117 , n23116 );
not ( n23118 , n23117 );
buf ( n23119 , n23118 );
not ( n23120 , n23119 );
and ( n23121 , n23112 , n23120 );
xor ( n23122 , n894 , n855 );
and ( n23123 , n23122 , n895 );
nor ( n23124 , n23121 , n23123 );
buf ( n23125 , n23124 );
not ( n23126 , n23125 );
buf ( n23127 , n23126 );
buf ( n23128 , n23127 );
not ( n23129 , n23128 );
or ( n23130 , n23111 , n23129 );
buf ( n23131 , n23106 );
not ( n23132 , n23131 );
buf ( n23133 , n23124 );
not ( n23134 , n23133 );
or ( n23135 , n23132 , n23134 );
buf ( n23136 , n862 );
buf ( n23137 , n888 );
xor ( n23138 , n23136 , n23137 );
buf ( n23139 , n23138 );
buf ( n23140 , n23139 );
not ( n23141 , n23140 );
buf ( n23142 , n22303 );
buf ( n23143 , n23142 );
buf ( n23144 , n23143 );
buf ( n23145 , n23144 );
not ( n23146 , n23145 );
or ( n23147 , n23141 , n23146 );
buf ( n23148 , n20363 );
buf ( n23149 , n861 );
buf ( n23150 , n888 );
xor ( n23151 , n23149 , n23150 );
buf ( n23152 , n23151 );
buf ( n23153 , n23152 );
nand ( n23154 , n23148 , n23153 );
buf ( n23155 , n23154 );
buf ( n23156 , n23155 );
nand ( n23157 , n23147 , n23156 );
buf ( n23158 , n23157 );
buf ( n23159 , n23158 );
nand ( n23160 , n23135 , n23159 );
buf ( n23161 , n23160 );
buf ( n23162 , n23161 );
nand ( n23163 , n23130 , n23162 );
buf ( n23164 , n23163 );
buf ( n23165 , n23164 );
xor ( n23166 , n23102 , n23165 );
buf ( n23167 , n857 );
buf ( n23168 , n892 );
xor ( n23169 , n23167 , n23168 );
buf ( n23170 , n23169 );
buf ( n23171 , n23170 );
not ( n23172 , n23171 );
buf ( n23173 , n20159 );
buf ( n23174 , n23173 );
buf ( n23175 , n23174 );
buf ( n23176 , n23175 );
not ( n23177 , n23176 );
or ( n23178 , n23172 , n23177 );
buf ( n23179 , n20164 );
not ( n23180 , n23179 );
buf ( n23181 , n23180 );
buf ( n23182 , n23181 );
buf ( n23183 , n856 );
buf ( n23184 , n892 );
xor ( n23185 , n23183 , n23184 );
buf ( n23186 , n23185 );
buf ( n23187 , n23186 );
nand ( n23188 , n23182 , n23187 );
buf ( n23189 , n23188 );
buf ( n23190 , n23189 );
nand ( n23191 , n23178 , n23190 );
buf ( n23192 , n23191 );
buf ( n23193 , n23192 );
not ( n23194 , n23193 );
buf ( n23195 , n863 );
buf ( n23196 , n887 );
or ( n23197 , n23195 , n23196 );
buf ( n23198 , n888 );
nand ( n23199 , n23197 , n23198 );
buf ( n23200 , n23199 );
buf ( n23201 , n23200 );
buf ( n23202 , n863 );
buf ( n23203 , n887 );
nand ( n23204 , n23202 , n23203 );
buf ( n23205 , n23204 );
buf ( n23206 , n23205 );
buf ( n23207 , n886 );
nand ( n23208 , n23201 , n23206 , n23207 );
buf ( n23209 , n23208 );
buf ( n23210 , n23209 );
not ( n23211 , n23210 );
or ( n23212 , n23194 , n23211 );
buf ( n23213 , n23209 );
buf ( n23214 , n23192 );
or ( n23215 , n23213 , n23214 );
nand ( n23216 , n23212 , n23215 );
buf ( n23217 , n23216 );
buf ( n23218 , n23217 );
and ( n23219 , n23166 , n23218 );
and ( n23220 , n23102 , n23165 );
or ( n23221 , n23219 , n23220 );
buf ( n23222 , n23221 );
buf ( n23223 , n23222 );
xor ( n23224 , n23084 , n23223 );
buf ( n23225 , n23192 );
not ( n23226 , n23225 );
buf ( n23227 , n23209 );
nor ( n23228 , n23226 , n23227 );
buf ( n23229 , n23228 );
buf ( n23230 , n23229 );
buf ( n23231 , n20700 );
buf ( n23232 , n23231 );
buf ( n23233 , n23232 );
buf ( n23234 , n23233 );
not ( n23235 , n23234 );
buf ( n23236 , n863 );
not ( n23237 , n23236 );
buf ( n23238 , n23237 );
buf ( n23239 , n23238 );
nor ( n23240 , n23235 , n23239 );
buf ( n23241 , n23240 );
buf ( n23242 , n23241 );
buf ( n23243 , n860 );
buf ( n23244 , n888 );
xor ( n23245 , n23243 , n23244 );
buf ( n23246 , n23245 );
buf ( n23247 , n23246 );
not ( n23248 , n23247 );
buf ( n23249 , n23144 );
not ( n23250 , n23249 );
or ( n23251 , n23248 , n23250 );
buf ( n23252 , n20363 );
buf ( n23253 , n859 );
buf ( n23254 , n888 );
xor ( n23255 , n23253 , n23254 );
buf ( n23256 , n23255 );
buf ( n23257 , n23256 );
nand ( n23258 , n23252 , n23257 );
buf ( n23259 , n23258 );
buf ( n23260 , n23259 );
nand ( n23261 , n23251 , n23260 );
buf ( n23262 , n23261 );
buf ( n23263 , n23262 );
xor ( n23264 , n23242 , n23263 );
buf ( n23265 , n23186 );
not ( n23266 , n23265 );
buf ( n23267 , n23175 );
not ( n23268 , n23267 );
or ( n23269 , n23266 , n23268 );
buf ( n23270 , n23181 );
buf ( n23271 , n855 );
buf ( n23272 , n892 );
xor ( n23273 , n23271 , n23272 );
buf ( n23274 , n23273 );
buf ( n23275 , n23274 );
nand ( n23276 , n23270 , n23275 );
buf ( n23277 , n23276 );
buf ( n23278 , n23277 );
nand ( n23279 , n23269 , n23278 );
buf ( n23280 , n23279 );
buf ( n23281 , n23280 );
xor ( n23282 , n23264 , n23281 );
buf ( n23283 , n23282 );
buf ( n23284 , n23283 );
xor ( n23285 , n23230 , n23284 );
buf ( n23286 , n23122 );
not ( n23287 , n23286 );
buf ( n23288 , n20132 );
buf ( n23289 , n23288 );
not ( n23290 , n23289 );
or ( n23291 , n23287 , n23290 );
buf ( n23292 , n23045 );
buf ( n23293 , n895 );
nand ( n23294 , n23292 , n23293 );
buf ( n23295 , n23294 );
buf ( n23296 , n23295 );
nand ( n23297 , n23291 , n23296 );
buf ( n23298 , n23297 );
buf ( n23299 , n23298 );
buf ( n23300 , n23152 );
not ( n23301 , n23300 );
buf ( n23302 , n23144 );
not ( n23303 , n23302 );
or ( n23304 , n23301 , n23303 );
buf ( n23305 , n20363 );
buf ( n23306 , n23246 );
nand ( n23307 , n23305 , n23306 );
buf ( n23308 , n23307 );
buf ( n23309 , n23308 );
nand ( n23310 , n23304 , n23309 );
buf ( n23311 , n23310 );
buf ( n23312 , n23311 );
xor ( n23313 , n23299 , n23312 );
xor ( n23314 , n886 , n863 );
buf ( n23315 , n23314 );
not ( n23316 , n23315 );
buf ( n23317 , n23027 );
not ( n23318 , n23317 );
or ( n23319 , n23316 , n23318 );
buf ( n23320 , n20260 );
buf ( n23321 , n23320 );
buf ( n23322 , n23019 );
nand ( n23323 , n23321 , n23322 );
buf ( n23324 , n23323 );
buf ( n23325 , n23324 );
nand ( n23326 , n23319 , n23325 );
buf ( n23327 , n23326 );
buf ( n23328 , n23327 );
and ( n23329 , n23313 , n23328 );
and ( n23330 , n23299 , n23312 );
or ( n23331 , n23329 , n23330 );
buf ( n23332 , n23331 );
buf ( n23333 , n23332 );
xor ( n23334 , n23285 , n23333 );
buf ( n23335 , n23334 );
buf ( n23336 , n23335 );
xor ( n23337 , n23224 , n23336 );
buf ( n23338 , n23337 );
buf ( n23339 , n23338 );
buf ( n23340 , n859 );
buf ( n23341 , n864 );
and ( n23342 , n23340 , n23341 );
buf ( n23343 , n23342 );
buf ( n23344 , n23343 );
buf ( n23345 , n22439 );
not ( n23346 , n23345 );
buf ( n23347 , n20302 );
not ( n23348 , n23347 );
or ( n23349 , n23346 , n23348 );
buf ( n23350 , n19030 );
buf ( n23351 , n857 );
buf ( n23352 , n864 );
xor ( n23353 , n23351 , n23352 );
buf ( n23354 , n23353 );
buf ( n23355 , n23354 );
nand ( n23356 , n23350 , n23355 );
buf ( n23357 , n23356 );
buf ( n23358 , n23357 );
nand ( n23359 , n23349 , n23358 );
buf ( n23360 , n23359 );
buf ( n23361 , n23360 );
xor ( n23362 , n23344 , n23361 );
buf ( n23363 , n22203 );
not ( n23364 , n23363 );
buf ( n23365 , n20404 );
not ( n23366 , n23365 );
or ( n23367 , n23364 , n23366 );
buf ( n23368 , n20869 );
buf ( n23369 , n890 );
nand ( n23370 , n23368 , n23369 );
buf ( n23371 , n23370 );
buf ( n23372 , n23371 );
nand ( n23373 , n23367 , n23372 );
buf ( n23374 , n23373 );
buf ( n23375 , n23374 );
not ( n23376 , n23375 );
buf ( n23377 , n23376 );
buf ( n23378 , n23377 );
xor ( n23379 , n23362 , n23378 );
buf ( n23380 , n23379 );
buf ( n23381 , n23380 );
xor ( n23382 , n22429 , n22446 );
and ( n23383 , n23382 , n22452 );
and ( n23384 , n22429 , n22446 );
or ( n23385 , n23383 , n23384 );
buf ( n23386 , n23385 );
buf ( n23387 , n23386 );
xor ( n23388 , n23381 , n23387 );
not ( n23389 , n21153 );
not ( n23390 , n21164 );
or ( n23391 , n23389 , n23390 );
not ( n23392 , n21158 );
not ( n23393 , n21165 );
or ( n23394 , n23392 , n23393 );
nand ( n23395 , n23394 , n21147 );
nand ( n23396 , n23391 , n23395 );
buf ( n23397 , n23396 );
and ( n23398 , n23388 , n23397 );
and ( n23399 , n23381 , n23387 );
or ( n23400 , n23398 , n23399 );
buf ( n23401 , n23400 );
xor ( n23402 , n22254 , n22264 );
and ( n23403 , n23402 , n22280 );
and ( n23404 , n22254 , n22264 );
or ( n23405 , n23403 , n23404 );
buf ( n23406 , n23405 );
not ( n23407 , n22296 );
not ( n23408 , n22314 );
or ( n23409 , n23407 , n23408 );
not ( n23410 , n22296 );
not ( n23411 , n23410 );
not ( n23412 , n22315 );
or ( n23413 , n23411 , n23412 );
nand ( n23414 , n23413 , n22329 );
nand ( n23415 , n23409 , n23414 );
or ( n23416 , n23406 , n23415 );
buf ( n23417 , n22363 );
not ( n23418 , n23417 );
buf ( n23419 , n20694 );
not ( n23420 , n23419 );
or ( n23421 , n23418 , n23420 );
buf ( n23422 , n23233 );
buf ( n23423 , n837 );
buf ( n23424 , n884 );
xor ( n23425 , n23423 , n23424 );
buf ( n23426 , n23425 );
buf ( n23427 , n23426 );
nand ( n23428 , n23422 , n23427 );
buf ( n23429 , n23428 );
buf ( n23430 , n23429 );
nand ( n23431 , n23421 , n23430 );
buf ( n23432 , n23431 );
buf ( n23433 , n23432 );
buf ( n23434 , n22310 );
not ( n23435 , n23434 );
buf ( n23436 , n20358 );
not ( n23437 , n23436 );
or ( n23438 , n23435 , n23437 );
buf ( n23439 , n833 );
buf ( n23440 , n888 );
xor ( n23441 , n23439 , n23440 );
buf ( n23442 , n23441 );
buf ( n23443 , n23442 );
buf ( n23444 , n20363 );
nand ( n23445 , n23443 , n23444 );
buf ( n23446 , n23445 );
buf ( n23447 , n23446 );
nand ( n23448 , n23438 , n23447 );
buf ( n23449 , n23448 );
buf ( n23450 , n23449 );
buf ( n23451 , n22141 );
not ( n23452 , n23451 );
buf ( n23453 , n20243 );
not ( n23454 , n23453 );
or ( n23455 , n23452 , n23454 );
and ( n23456 , n845 , n876 );
not ( n23457 , n845 );
and ( n23458 , n23457 , n19068 );
nor ( n23459 , n23456 , n23458 );
nand ( n23460 , n20246 , n23459 );
buf ( n23461 , n23460 );
nand ( n23462 , n23455 , n23461 );
buf ( n23463 , n23462 );
buf ( n23464 , n23463 );
and ( n23465 , n23450 , n23464 );
not ( n23466 , n23450 );
buf ( n23467 , n23463 );
not ( n23468 , n23467 );
buf ( n23469 , n23468 );
buf ( n23470 , n23469 );
and ( n23471 , n23466 , n23470 );
nor ( n23472 , n23465 , n23471 );
buf ( n23473 , n23472 );
buf ( n23474 , n23473 );
xor ( n23475 , n23433 , n23474 );
buf ( n23476 , n23475 );
nand ( n23477 , n23416 , n23476 );
buf ( n23478 , n23406 );
buf ( n23479 , n23415 );
nand ( n23480 , n23478 , n23479 );
buf ( n23481 , n23480 );
nand ( n23482 , n23477 , n23481 );
buf ( n23483 , n23374 );
buf ( n23484 , n23463 );
not ( n23485 , n23484 );
buf ( n23486 , n23449 );
not ( n23487 , n23486 );
or ( n23488 , n23485 , n23487 );
buf ( n23489 , n23449 );
buf ( n23490 , n23463 );
or ( n23491 , n23489 , n23490 );
buf ( n23492 , n23432 );
nand ( n23493 , n23491 , n23492 );
buf ( n23494 , n23493 );
buf ( n23495 , n23494 );
nand ( n23496 , n23488 , n23495 );
buf ( n23497 , n23496 );
buf ( n23498 , n23497 );
xor ( n23499 , n23483 , n23498 );
not ( n23500 , n20767 );
xor ( n23501 , n882 , n839 );
not ( n23502 , n23501 );
or ( n23503 , n23500 , n23502 );
nand ( n23504 , n22292 , n19569 , n19576 );
nand ( n23505 , n23503 , n23504 );
buf ( n23506 , n23505 );
not ( n23507 , n22347 );
not ( n23508 , n20736 );
or ( n23509 , n23507 , n23508 );
buf ( n23510 , n20555 );
buf ( n23511 , n847 );
buf ( n23512 , n874 );
xor ( n23513 , n23511 , n23512 );
buf ( n23514 , n23513 );
buf ( n23515 , n23514 );
nand ( n23516 , n23510 , n23515 );
buf ( n23517 , n23516 );
nand ( n23518 , n23509 , n23517 );
buf ( n23519 , n23518 );
xor ( n23520 , n23506 , n23519 );
buf ( n23521 , n22393 );
not ( n23522 , n23521 );
buf ( n23523 , n19230 );
not ( n23524 , n23523 );
or ( n23525 , n23522 , n23524 );
buf ( n23526 , n19235 );
buf ( n23527 , n849 );
buf ( n23528 , n872 );
xor ( n23529 , n23527 , n23528 );
buf ( n23530 , n23529 );
buf ( n23531 , n23530 );
nand ( n23532 , n23526 , n23531 );
buf ( n23533 , n23532 );
buf ( n23534 , n23533 );
nand ( n23535 , n23525 , n23534 );
buf ( n23536 , n23535 );
buf ( n23537 , n23536 );
and ( n23538 , n23520 , n23537 );
and ( n23539 , n23506 , n23519 );
or ( n23540 , n23538 , n23539 );
buf ( n23541 , n23540 );
buf ( n23542 , n23541 );
xor ( n23543 , n23499 , n23542 );
buf ( n23544 , n23543 );
xor ( n23545 , n23482 , n23544 );
not ( n23546 , n22247 );
not ( n23547 , n22239 );
or ( n23548 , n23546 , n23547 );
buf ( n23549 , n18938 );
xor ( n23550 , n866 , n855 );
buf ( n23551 , n23550 );
nand ( n23552 , n23549 , n23551 );
buf ( n23553 , n23552 );
nand ( n23554 , n23548 , n23553 );
not ( n23555 , n22259 );
not ( n23556 , n18884 );
or ( n23557 , n23555 , n23556 );
buf ( n23558 , n20786 );
xor ( n23559 , n868 , n853 );
buf ( n23560 , n23559 );
nand ( n23561 , n23558 , n23560 );
buf ( n23562 , n23561 );
nand ( n23563 , n23557 , n23562 );
xor ( n23564 , n23554 , n23563 );
not ( n23565 , n22158 );
buf ( n23566 , n21010 );
buf ( n23567 , n19255 );
nor ( n23568 , n23566 , n23567 );
buf ( n23569 , n23568 );
not ( n23570 , n23569 );
or ( n23571 , n23565 , n23570 );
buf ( n23572 , n843 );
buf ( n23573 , n878 );
xor ( n23574 , n23572 , n23573 );
buf ( n23575 , n23574 );
nand ( n23576 , n23575 , n19265 );
nand ( n23577 , n23571 , n23576 );
and ( n23578 , n23564 , n23577 );
and ( n23579 , n23554 , n23563 );
or ( n23580 , n23578 , n23579 );
not ( n23581 , n23580 );
buf ( n23582 , n22273 );
not ( n23583 , n23582 );
buf ( n23584 , n20642 );
not ( n23585 , n23584 );
or ( n23586 , n23583 , n23585 );
xor ( n23587 , n880 , n841 );
nand ( n23588 , n21083 , n23587 );
buf ( n23589 , n23588 );
nand ( n23590 , n23586 , n23589 );
buf ( n23591 , n23590 );
buf ( n23592 , n23591 );
buf ( n23593 , n22323 );
not ( n23594 , n23593 );
buf ( n23595 , n19119 );
not ( n23596 , n23595 );
or ( n23597 , n23594 , n23596 );
xor ( n23598 , n870 , n851 );
nand ( n23599 , n23598 , n20226 );
buf ( n23600 , n23599 );
nand ( n23601 , n23597 , n23600 );
buf ( n23602 , n23601 );
buf ( n23603 , n23602 );
xor ( n23604 , n23592 , n23603 );
buf ( n23605 , n22185 );
not ( n23606 , n23605 );
buf ( n23607 , n20521 );
not ( n23608 , n23607 );
or ( n23609 , n23606 , n23608 );
buf ( n23610 , n20525 );
xor ( n23611 , n886 , n835 );
buf ( n23612 , n23611 );
nand ( n23613 , n23610 , n23612 );
buf ( n23614 , n23613 );
buf ( n23615 , n23614 );
nand ( n23616 , n23609 , n23615 );
buf ( n23617 , n23616 );
buf ( n23618 , n23617 );
and ( n23619 , n23604 , n23618 );
and ( n23620 , n23592 , n23603 );
or ( n23621 , n23619 , n23620 );
buf ( n23622 , n23621 );
not ( n23623 , n23622 );
not ( n23624 , n23623 );
or ( n23625 , n23581 , n23624 );
not ( n23626 , n23580 );
nand ( n23627 , n23622 , n23626 );
nand ( n23628 , n23625 , n23627 );
buf ( n23629 , n23514 );
not ( n23630 , n23629 );
buf ( n23631 , n20549 );
not ( n23632 , n23631 );
or ( n23633 , n23630 , n23632 );
buf ( n23634 , n20555 );
buf ( n23635 , n846 );
buf ( n23636 , n874 );
xor ( n23637 , n23635 , n23636 );
buf ( n23638 , n23637 );
buf ( n23639 , n23638 );
nand ( n23640 , n23634 , n23639 );
buf ( n23641 , n23640 );
buf ( n23642 , n23641 );
nand ( n23643 , n23633 , n23642 );
buf ( n23644 , n23643 );
buf ( n23645 , n23501 );
not ( n23646 , n23645 );
buf ( n23647 , n19580 );
not ( n23648 , n23647 );
or ( n23649 , n23646 , n23648 );
buf ( n23650 , n19909 );
buf ( n23651 , n838 );
buf ( n23652 , n882 );
xor ( n23653 , n23651 , n23652 );
buf ( n23654 , n23653 );
buf ( n23655 , n23654 );
nand ( n23656 , n23650 , n23655 );
buf ( n23657 , n23656 );
buf ( n23658 , n23657 );
nand ( n23659 , n23649 , n23658 );
buf ( n23660 , n23659 );
not ( n23661 , n23660 );
and ( n23662 , n23644 , n23661 );
not ( n23663 , n23644 );
and ( n23664 , n23663 , n23660 );
nor ( n23665 , n23662 , n23664 );
buf ( n23666 , n19082 );
buf ( n23667 , n844 );
buf ( n23668 , n876 );
xor ( n23669 , n23667 , n23668 );
buf ( n23670 , n23669 );
buf ( n23671 , n23670 );
nand ( n23672 , n23666 , n23671 );
buf ( n23673 , n23672 );
nand ( n23674 , n23459 , n19077 );
nand ( n23675 , n23673 , n23674 );
not ( n23676 , n23675 );
xor ( n23677 , n23665 , n23676 );
and ( n23678 , n23628 , n23677 );
not ( n23679 , n23628 );
not ( n23680 , n23677 );
and ( n23681 , n23679 , n23680 );
nor ( n23682 , n23678 , n23681 );
xor ( n23683 , n23545 , n23682 );
xor ( n23684 , n23401 , n23683 );
xor ( n23685 , n22134 , n22148 );
and ( n23686 , n23685 , n22163 );
and ( n23687 , n22134 , n22148 );
or ( n23688 , n23686 , n23687 );
buf ( n23689 , n23688 );
buf ( n23690 , n23689 );
xor ( n23691 , n22175 , n22192 );
and ( n23692 , n23691 , n22210 );
and ( n23693 , n22175 , n22192 );
or ( n23694 , n23692 , n23693 );
buf ( n23695 , n23694 );
buf ( n23696 , n23695 );
xor ( n23697 , n23690 , n23696 );
buf ( n23698 , n22372 );
not ( n23699 , n23698 );
buf ( n23700 , n22403 );
not ( n23701 , n23700 );
or ( n23702 , n23699 , n23701 );
buf ( n23703 , n22351 );
nand ( n23704 , n23702 , n23703 );
buf ( n23705 , n23704 );
buf ( n23706 , n23705 );
buf ( n23707 , n22400 );
buf ( n23708 , n22369 );
nand ( n23709 , n23707 , n23708 );
buf ( n23710 , n23709 );
buf ( n23711 , n23710 );
nand ( n23712 , n23706 , n23711 );
buf ( n23713 , n23712 );
buf ( n23714 , n23713 );
xor ( n23715 , n23697 , n23714 );
buf ( n23716 , n23715 );
buf ( n23717 , n23716 );
xor ( n23718 , n22166 , n22213 );
and ( n23719 , n23718 , n22230 );
and ( n23720 , n22166 , n22213 );
or ( n23721 , n23719 , n23720 );
buf ( n23722 , n23721 );
buf ( n23723 , n23722 );
xor ( n23724 , n23717 , n23723 );
xor ( n23725 , n23415 , n23406 );
buf ( n23726 , n23725 );
buf ( n23727 , n23476 );
and ( n23728 , n23726 , n23727 );
not ( n23729 , n23726 );
buf ( n23730 , n23476 );
not ( n23731 , n23730 );
buf ( n23732 , n23731 );
buf ( n23733 , n23732 );
and ( n23734 , n23729 , n23733 );
nor ( n23735 , n23728 , n23734 );
buf ( n23736 , n23735 );
buf ( n23737 , n23736 );
and ( n23738 , n23724 , n23737 );
and ( n23739 , n23717 , n23723 );
or ( n23740 , n23738 , n23739 );
buf ( n23741 , n23740 );
xor ( n23742 , n23684 , n23741 );
not ( n23743 , n23742 );
not ( n23744 , n23743 );
buf ( n23745 , n22410 );
not ( n23746 , n23745 );
buf ( n23747 , n22330 );
not ( n23748 , n23747 );
or ( n23749 , n23746 , n23748 );
buf ( n23750 , n22282 );
nand ( n23751 , n23749 , n23750 );
buf ( n23752 , n23751 );
buf ( n23753 , n23752 );
buf ( n23754 , n22330 );
not ( n23755 , n23754 );
buf ( n23756 , n22416 );
nand ( n23757 , n23755 , n23756 );
buf ( n23758 , n23757 );
buf ( n23759 , n23758 );
nand ( n23760 , n23753 , n23759 );
buf ( n23761 , n23760 );
buf ( n23762 , n23761 );
xor ( n23763 , n23554 , n23563 );
xor ( n23764 , n23763 , n23577 );
buf ( n23765 , n23764 );
xor ( n23766 , n23506 , n23519 );
xor ( n23767 , n23766 , n23537 );
buf ( n23768 , n23767 );
buf ( n23769 , n23768 );
xor ( n23770 , n23765 , n23769 );
xor ( n23771 , n23592 , n23603 );
xor ( n23772 , n23771 , n23618 );
buf ( n23773 , n23772 );
buf ( n23774 , n23773 );
xor ( n23775 , n23770 , n23774 );
buf ( n23776 , n23775 );
buf ( n23777 , n23776 );
xor ( n23778 , n23762 , n23777 );
xor ( n23779 , n22428 , n22455 );
and ( n23780 , n23779 , n22462 );
and ( n23781 , n22428 , n22455 );
or ( n23782 , n23780 , n23781 );
buf ( n23783 , n23782 );
buf ( n23784 , n23783 );
and ( n23785 , n23778 , n23784 );
and ( n23786 , n23762 , n23777 );
or ( n23787 , n23785 , n23786 );
buf ( n23788 , n23787 );
xor ( n23789 , n23765 , n23769 );
and ( n23790 , n23789 , n23774 );
and ( n23791 , n23765 , n23769 );
or ( n23792 , n23790 , n23791 );
buf ( n23793 , n23792 );
buf ( n23794 , n23793 );
buf ( n23795 , n858 );
buf ( n23796 , n864 );
and ( n23797 , n23795 , n23796 );
buf ( n23798 , n23797 );
buf ( n23799 , n23798 );
buf ( n23800 , n23354 );
not ( n23801 , n23800 );
buf ( n23802 , n20302 );
not ( n23803 , n23802 );
or ( n23804 , n23801 , n23803 );
buf ( n23805 , n19027 );
buf ( n23806 , n856 );
buf ( n23807 , n864 );
xor ( n23808 , n23806 , n23807 );
buf ( n23809 , n23808 );
buf ( n23810 , n23809 );
nand ( n23811 , n23805 , n23810 );
buf ( n23812 , n23811 );
buf ( n23813 , n23812 );
nand ( n23814 , n23804 , n23813 );
buf ( n23815 , n23814 );
buf ( n23816 , n23815 );
xor ( n23817 , n23799 , n23816 );
buf ( n23818 , n23575 );
not ( n23819 , n23818 );
buf ( n23820 , n19259 );
not ( n23821 , n23820 );
or ( n23822 , n23819 , n23821 );
buf ( n23823 , n19265 );
buf ( n23824 , n842 );
buf ( n23825 , n878 );
xor ( n23826 , n23824 , n23825 );
buf ( n23827 , n23826 );
buf ( n23828 , n23827 );
nand ( n23829 , n23823 , n23828 );
buf ( n23830 , n23829 );
buf ( n23831 , n23830 );
nand ( n23832 , n23822 , n23831 );
buf ( n23833 , n23832 );
buf ( n23834 , n23833 );
xor ( n23835 , n23817 , n23834 );
buf ( n23836 , n23835 );
buf ( n23837 , n20404 );
not ( n23838 , n23837 );
buf ( n23839 , n23838 );
not ( n23840 , n20869 );
nand ( n23841 , n23839 , n23840 );
nand ( n23842 , n23841 , n890 );
nand ( n23843 , n22303 , n23442 );
buf ( n23844 , n20363 );
buf ( n23845 , n832 );
buf ( n23846 , n888 );
xor ( n23847 , n23845 , n23846 );
buf ( n23848 , n23847 );
buf ( n23849 , n23848 );
nand ( n23850 , n23844 , n23849 );
buf ( n23851 , n23850 );
nand ( n23852 , n23843 , n23851 );
not ( n23853 , n23852 );
and ( n23854 , n23842 , n23853 );
not ( n23855 , n23842 );
and ( n23856 , n23855 , n23852 );
nor ( n23857 , n23854 , n23856 );
not ( n23858 , n23426 );
not ( n23859 , n20694 );
or ( n23860 , n23858 , n23859 );
buf ( n23861 , n20700 );
buf ( n23862 , n836 );
buf ( n23863 , n884 );
xor ( n23864 , n23862 , n23863 );
buf ( n23865 , n23864 );
buf ( n23866 , n23865 );
nand ( n23867 , n23861 , n23866 );
buf ( n23868 , n23867 );
nand ( n23869 , n23860 , n23868 );
xnor ( n23870 , n23857 , n23869 );
xor ( n23871 , n23836 , n23870 );
buf ( n23872 , n23550 );
not ( n23873 , n23872 );
buf ( n23874 , n18931 );
not ( n23875 , n23874 );
or ( n23876 , n23873 , n23875 );
buf ( n23877 , n21249 );
buf ( n23878 , n854 );
buf ( n23879 , n866 );
xor ( n23880 , n23878 , n23879 );
buf ( n23881 , n23880 );
buf ( n23882 , n23881 );
nand ( n23883 , n23877 , n23882 );
buf ( n23884 , n23883 );
buf ( n23885 , n23884 );
nand ( n23886 , n23876 , n23885 );
buf ( n23887 , n23886 );
buf ( n23888 , n23559 );
not ( n23889 , n23888 );
buf ( n23890 , n18876 );
buf ( n23891 , n18881 );
and ( n23892 , n23890 , n23891 );
buf ( n23893 , n23892 );
buf ( n23894 , n23893 );
not ( n23895 , n23894 );
or ( n23896 , n23889 , n23895 );
buf ( n23897 , n18892 );
buf ( n23898 , n852 );
buf ( n23899 , n868 );
xor ( n23900 , n23898 , n23899 );
buf ( n23901 , n23900 );
buf ( n23902 , n23901 );
nand ( n23903 , n23897 , n23902 );
buf ( n23904 , n23903 );
buf ( n23905 , n23904 );
nand ( n23906 , n23896 , n23905 );
buf ( n23907 , n23906 );
xor ( n23908 , n23887 , n23907 );
buf ( n23909 , n23908 );
buf ( n23910 , n23587 );
not ( n23911 , n23910 );
buf ( n23912 , n19614 );
not ( n23913 , n23912 );
or ( n23914 , n23911 , n23913 );
buf ( n23915 , n20325 );
buf ( n23916 , n23915 );
buf ( n23917 , n23916 );
buf ( n23918 , n23917 );
buf ( n23919 , n840 );
buf ( n23920 , n880 );
xor ( n23921 , n23919 , n23920 );
buf ( n23922 , n23921 );
buf ( n23923 , n23922 );
nand ( n23924 , n23918 , n23923 );
buf ( n23925 , n23924 );
buf ( n23926 , n23925 );
nand ( n23927 , n23914 , n23926 );
buf ( n23928 , n23927 );
buf ( n23929 , n23928 );
xor ( n23930 , n23909 , n23929 );
buf ( n23931 , n23930 );
xor ( n23932 , n23871 , n23931 );
buf ( n23933 , n23932 );
xor ( n23934 , n23794 , n23933 );
xor ( n23935 , n23344 , n23361 );
and ( n23936 , n23935 , n23378 );
and ( n23937 , n23344 , n23361 );
or ( n23938 , n23936 , n23937 );
buf ( n23939 , n23938 );
buf ( n23940 , n23939 );
buf ( n23941 , n23598 );
not ( n23942 , n23941 );
buf ( n23943 , n19122 );
not ( n23944 , n23943 );
or ( n23945 , n23942 , n23944 );
buf ( n23946 , n19131 );
buf ( n23947 , n850 );
buf ( n23948 , n870 );
xor ( n23949 , n23947 , n23948 );
buf ( n23950 , n23949 );
buf ( n23951 , n23950 );
nand ( n23952 , n23946 , n23951 );
buf ( n23953 , n23952 );
buf ( n23954 , n23953 );
nand ( n23955 , n23945 , n23954 );
buf ( n23956 , n23955 );
buf ( n23957 , n23530 );
not ( n23958 , n23957 );
buf ( n23959 , n20211 );
not ( n23960 , n23959 );
or ( n23961 , n23958 , n23960 );
buf ( n23962 , n19234 );
buf ( n23963 , n848 );
buf ( n23964 , n872 );
xor ( n23965 , n23963 , n23964 );
buf ( n23966 , n23965 );
buf ( n23967 , n23966 );
nand ( n23968 , n23962 , n23967 );
buf ( n23969 , n23968 );
buf ( n23970 , n23969 );
nand ( n23971 , n23961 , n23970 );
buf ( n23972 , n23971 );
xor ( n23973 , n23956 , n23972 );
buf ( n23974 , n23611 );
not ( n23975 , n23974 );
buf ( n23976 , n20521 );
not ( n23977 , n23976 );
or ( n23978 , n23975 , n23977 );
buf ( n23979 , n20525 );
buf ( n23980 , n834 );
buf ( n23981 , n886 );
xor ( n23982 , n23980 , n23981 );
buf ( n23983 , n23982 );
buf ( n23984 , n23983 );
nand ( n23985 , n23979 , n23984 );
buf ( n23986 , n23985 );
buf ( n23987 , n23986 );
nand ( n23988 , n23978 , n23987 );
buf ( n23989 , n23988 );
xor ( n23990 , n23973 , n23989 );
buf ( n23991 , n23990 );
xor ( n23992 , n23940 , n23991 );
xor ( n23993 , n23690 , n23696 );
and ( n23994 , n23993 , n23714 );
and ( n23995 , n23690 , n23696 );
or ( n23996 , n23994 , n23995 );
buf ( n23997 , n23996 );
buf ( n23998 , n23997 );
xor ( n23999 , n23992 , n23998 );
buf ( n24000 , n23999 );
buf ( n24001 , n24000 );
xor ( n24002 , n23934 , n24001 );
buf ( n24003 , n24002 );
xor ( n24004 , n23788 , n24003 );
xor ( n24005 , n23381 , n23387 );
xor ( n24006 , n24005 , n23397 );
buf ( n24007 , n24006 );
buf ( n24008 , n24007 );
not ( n24009 , n21175 );
not ( n24010 , n21126 );
or ( n24011 , n24009 , n24010 );
not ( n24012 , n21127 );
not ( n24013 , n21169 );
or ( n24014 , n24012 , n24013 );
nand ( n24015 , n24014 , n20995 );
nand ( n24016 , n24011 , n24015 );
buf ( n24017 , n24016 );
xor ( n24018 , n24008 , n24017 );
xor ( n24019 , n23717 , n23723 );
xor ( n24020 , n24019 , n23737 );
buf ( n24021 , n24020 );
buf ( n24022 , n24021 );
and ( n24023 , n24018 , n24022 );
and ( n24024 , n24008 , n24017 );
or ( n24025 , n24023 , n24024 );
buf ( n24026 , n24025 );
xor ( n24027 , n24004 , n24026 );
not ( n24028 , n24027 );
not ( n24029 , n24028 );
or ( n24030 , n23744 , n24029 );
xor ( n24031 , n23762 , n23777 );
xor ( n24032 , n24031 , n23784 );
buf ( n24033 , n24032 );
not ( n24034 , n24033 );
xor ( n24035 , n22233 , n22421 );
and ( n24036 , n24035 , n22465 );
and ( n24037 , n22233 , n22421 );
or ( n24038 , n24036 , n24037 );
buf ( n24039 , n24038 );
not ( n24040 , n24039 );
or ( n24041 , n24034 , n24040 );
not ( n24042 , n24039 );
not ( n24043 , n24042 );
not ( n24044 , n24033 );
not ( n24045 , n24044 );
or ( n24046 , n24043 , n24045 );
buf ( n24047 , n20833 );
buf ( n24048 , n20592 );
or ( n24049 , n24047 , n24048 );
buf ( n24050 , n21177 );
nand ( n24051 , n24049 , n24050 );
buf ( n24052 , n24051 );
buf ( n24053 , n24052 );
buf ( n24054 , n20833 );
buf ( n24055 , n20185 );
not ( n24056 , n24055 );
buf ( n24057 , n20387 );
not ( n24058 , n24057 );
or ( n24059 , n24056 , n24058 );
buf ( n24060 , n20589 );
nand ( n24061 , n24059 , n24060 );
buf ( n24062 , n24061 );
buf ( n24063 , n24062 );
nand ( n24064 , n24054 , n24063 );
buf ( n24065 , n24064 );
buf ( n24066 , n24065 );
nand ( n24067 , n24053 , n24066 );
buf ( n24068 , n24067 );
nand ( n24069 , n24046 , n24068 );
nand ( n24070 , n24041 , n24069 );
buf ( n24071 , n24070 );
nand ( n24072 , n24030 , n24071 );
nand ( n24073 , n24027 , n23742 );
nand ( n24074 , n24072 , n24073 );
buf ( n24075 , n24074 );
buf ( n24076 , n22730 );
not ( n24077 , n24076 );
not ( n24078 , n22567 );
not ( n24079 , n22555 );
or ( n24080 , n24078 , n24079 );
or ( n24081 , n22555 , n22567 );
nand ( n24082 , n24080 , n24081 );
buf ( n24083 , n24082 );
not ( n24084 , n24083 );
or ( n24085 , n24077 , n24084 );
buf ( n24086 , n24082 );
buf ( n24087 , n22730 );
or ( n24088 , n24086 , n24087 );
nand ( n24089 , n24085 , n24088 );
buf ( n24090 , n24089 );
buf ( n24091 , n24090 );
xor ( n24092 , n22790 , n22807 );
xor ( n24093 , n24092 , n22851 );
buf ( n24094 , n24093 );
buf ( n24095 , n24094 );
buf ( n24096 , n842 );
buf ( n24097 , n888 );
xor ( n24098 , n24096 , n24097 );
buf ( n24099 , n24098 );
buf ( n24100 , n24099 );
not ( n24101 , n24100 );
buf ( n24102 , n23144 );
not ( n24103 , n24102 );
or ( n24104 , n24101 , n24103 );
buf ( n24105 , n20363 );
buf ( n24106 , n22846 );
nand ( n24107 , n24105 , n24106 );
buf ( n24108 , n24107 );
buf ( n24109 , n24108 );
nand ( n24110 , n24104 , n24109 );
buf ( n24111 , n24110 );
not ( n24112 , n24111 );
buf ( n24113 , n21249 );
buf ( n24114 , n863 );
and ( n24115 , n24113 , n24114 );
buf ( n24116 , n24115 );
not ( n24117 , n24116 );
or ( n24118 , n24112 , n24117 );
buf ( n24119 , n24111 );
buf ( n24120 , n24116 );
nor ( n24121 , n24119 , n24120 );
buf ( n24122 , n24121 );
buf ( n24123 , n838 );
buf ( n24124 , n892 );
xor ( n24125 , n24123 , n24124 );
buf ( n24126 , n24125 );
buf ( n24127 , n24126 );
not ( n24128 , n24127 );
buf ( n24129 , n23175 );
not ( n24130 , n24129 );
or ( n24131 , n24128 , n24130 );
buf ( n24132 , n23181 );
buf ( n24133 , n22812 );
nand ( n24134 , n24132 , n24133 );
buf ( n24135 , n24134 );
buf ( n24136 , n24135 );
nand ( n24137 , n24131 , n24136 );
buf ( n24138 , n24137 );
buf ( n24139 , n24138 );
not ( n24140 , n24139 );
buf ( n24141 , n24140 );
or ( n24142 , n24122 , n24141 );
nand ( n24143 , n24118 , n24142 );
not ( n24144 , n24143 );
buf ( n24145 , n24144 );
not ( n24146 , n24145 );
buf ( n24147 , n850 );
buf ( n24148 , n880 );
xor ( n24149 , n24147 , n24148 );
buf ( n24150 , n24149 );
buf ( n24151 , n24150 );
not ( n24152 , n24151 );
buf ( n24153 , n18850 );
not ( n24154 , n24153 );
or ( n24155 , n24152 , n24154 );
nand ( n24156 , n22271 , n22829 );
buf ( n24157 , n24156 );
nand ( n24158 , n24155 , n24157 );
buf ( n24159 , n24158 );
buf ( n24160 , n24159 );
buf ( n24161 , n852 );
buf ( n24162 , n878 );
xor ( n24163 , n24161 , n24162 );
buf ( n24164 , n24163 );
buf ( n24165 , n24164 );
not ( n24166 , n24165 );
buf ( n24167 , n19259 );
not ( n24168 , n24167 );
or ( n24169 , n24166 , n24168 );
buf ( n24170 , n19265 );
buf ( n24171 , n22631 );
nand ( n24172 , n24170 , n24171 );
buf ( n24173 , n24172 );
buf ( n24174 , n24173 );
nand ( n24175 , n24169 , n24174 );
buf ( n24176 , n24175 );
buf ( n24177 , n24176 );
xor ( n24178 , n24160 , n24177 );
buf ( n24179 , n844 );
buf ( n24180 , n886 );
xor ( n24181 , n24179 , n24180 );
buf ( n24182 , n24181 );
buf ( n24183 , n24182 );
not ( n24184 , n24183 );
buf ( n24185 , n20521 );
not ( n24186 , n24185 );
or ( n24187 , n24184 , n24186 );
buf ( n24188 , n20525 );
buf ( n24189 , n22648 );
nand ( n24190 , n24188 , n24189 );
buf ( n24191 , n24190 );
buf ( n24192 , n24191 );
nand ( n24193 , n24187 , n24192 );
buf ( n24194 , n24193 );
buf ( n24195 , n24194 );
and ( n24196 , n24178 , n24195 );
and ( n24197 , n24160 , n24177 );
or ( n24198 , n24196 , n24197 );
buf ( n24199 , n24198 );
buf ( n24200 , n24199 );
not ( n24201 , n24200 );
buf ( n24202 , n24201 );
buf ( n24203 , n24202 );
not ( n24204 , n24203 );
or ( n24205 , n24146 , n24204 );
buf ( n24206 , n836 );
buf ( n24207 , n894 );
xor ( n24208 , n24206 , n24207 );
buf ( n24209 , n24208 );
buf ( n24210 , n24209 );
not ( n24211 , n24210 );
buf ( n24212 , n22776 );
not ( n24213 , n24212 );
or ( n24214 , n24211 , n24213 );
buf ( n24215 , n22773 );
buf ( n24216 , n895 );
nand ( n24217 , n24215 , n24216 );
buf ( n24218 , n24217 );
buf ( n24219 , n24218 );
nand ( n24220 , n24214 , n24219 );
buf ( n24221 , n24220 );
not ( n24222 , n24221 );
buf ( n24223 , n854 );
buf ( n24224 , n876 );
xor ( n24225 , n24223 , n24224 );
buf ( n24226 , n24225 );
not ( n24227 , n24226 );
not ( n24228 , n19153 );
or ( n24229 , n24227 , n24228 );
buf ( n24230 , n20246 );
buf ( n24231 , n22658 );
nand ( n24232 , n24230 , n24231 );
buf ( n24233 , n24232 );
nand ( n24234 , n24229 , n24233 );
not ( n24235 , n24234 );
or ( n24236 , n24222 , n24235 );
buf ( n24237 , n24234 );
buf ( n24238 , n24221 );
nor ( n24239 , n24237 , n24238 );
buf ( n24240 , n24239 );
buf ( n24241 , n20549 );
buf ( n24242 , n856 );
buf ( n24243 , n874 );
xor ( n24244 , n24242 , n24243 );
buf ( n24245 , n24244 );
buf ( n24246 , n24245 );
and ( n24247 , n24241 , n24246 );
buf ( n24248 , n20555 );
buf ( n24249 , n22710 );
and ( n24250 , n24248 , n24249 );
nor ( n24251 , n24247 , n24250 );
buf ( n24252 , n24251 );
or ( n24253 , n24240 , n24252 );
nand ( n24254 , n24236 , n24253 );
buf ( n24255 , n24254 );
buf ( n24256 , n24255 );
nand ( n24257 , n24205 , n24256 );
buf ( n24258 , n24257 );
buf ( n24259 , n24258 );
buf ( n24260 , n24199 );
buf ( n24261 , n24143 );
nand ( n24262 , n24260 , n24261 );
buf ( n24263 , n24262 );
buf ( n24264 , n24263 );
nand ( n24265 , n24259 , n24264 );
buf ( n24266 , n24265 );
buf ( n24267 , n24266 );
xor ( n24268 , n24095 , n24267 );
not ( n24269 , n22585 );
not ( n24270 , n22623 );
not ( n24271 , n24270 );
or ( n24272 , n24269 , n24271 );
not ( n24273 , n22585 );
nand ( n24274 , n24273 , n22623 );
nand ( n24275 , n24272 , n24274 );
and ( n24276 , n24275 , n22602 );
not ( n24277 , n24275 );
not ( n24278 , n22602 );
and ( n24279 , n24277 , n24278 );
nor ( n24280 , n24276 , n24279 );
not ( n24281 , n22664 );
not ( n24282 , n22665 );
not ( n24283 , n24282 );
or ( n24284 , n24281 , n24283 );
nand ( n24285 , n22665 , n22663 );
nand ( n24286 , n24284 , n24285 );
buf ( n24287 , n24286 );
buf ( n24288 , n22643 );
xor ( n24289 , n24287 , n24288 );
buf ( n24290 , n24289 );
xor ( n24291 , n24280 , n24290 );
buf ( n24292 , n22701 );
buf ( n24293 , n22722 );
xor ( n24294 , n24292 , n24293 );
buf ( n24295 , n24294 );
buf ( n24296 , n24295 );
buf ( n24297 , n22684 );
xor ( n24298 , n24296 , n24297 );
buf ( n24299 , n24298 );
and ( n24300 , n24291 , n24299 );
and ( n24301 , n24280 , n24290 );
or ( n24302 , n24300 , n24301 );
buf ( n24303 , n24302 );
and ( n24304 , n24268 , n24303 );
and ( n24305 , n24095 , n24267 );
or ( n24306 , n24304 , n24305 );
buf ( n24307 , n24306 );
buf ( n24308 , n24307 );
xor ( n24309 , n24091 , n24308 );
not ( n24310 , n22667 );
not ( n24311 , n22726 );
and ( n24312 , n24310 , n24311 );
and ( n24313 , n22667 , n22726 );
nor ( n24314 , n24312 , n24313 );
and ( n24315 , n24314 , n22627 );
not ( n24316 , n24314 );
buf ( n24317 , n22627 );
not ( n24318 , n24317 );
buf ( n24319 , n24318 );
and ( n24320 , n24316 , n24319 );
nor ( n24321 , n24315 , n24320 );
buf ( n24322 , n24321 );
buf ( n24323 , n848 );
buf ( n24324 , n882 );
xor ( n24325 , n24323 , n24324 );
buf ( n24326 , n24325 );
not ( n24327 , n24326 );
not ( n24328 , n19580 );
or ( n24329 , n24327 , n24328 );
buf ( n24330 , n20767 );
buf ( n24331 , n22590 );
nand ( n24332 , n24330 , n24331 );
buf ( n24333 , n24332 );
nand ( n24334 , n24329 , n24333 );
not ( n24335 , n24334 );
buf ( n24336 , n862 );
buf ( n24337 , n868 );
xor ( n24338 , n24336 , n24337 );
buf ( n24339 , n24338 );
buf ( n24340 , n24339 );
not ( n24341 , n24340 );
buf ( n24342 , n23893 );
not ( n24343 , n24342 );
or ( n24344 , n24341 , n24343 );
buf ( n24345 , n18892 );
buf ( n24346 , n22910 );
nand ( n24347 , n24345 , n24346 );
buf ( n24348 , n24347 );
buf ( n24349 , n24348 );
nand ( n24350 , n24344 , n24349 );
buf ( n24351 , n24350 );
not ( n24352 , n24351 );
or ( n24353 , n24335 , n24352 );
or ( n24354 , n24351 , n24334 );
buf ( n24355 , n840 );
buf ( n24356 , n890 );
xor ( n24357 , n24355 , n24356 );
buf ( n24358 , n24357 );
buf ( n24359 , n24358 );
not ( n24360 , n24359 );
buf ( n24361 , n21441 );
not ( n24362 , n24361 );
or ( n24363 , n24360 , n24362 );
buf ( n24364 , n20869 );
buf ( n24365 , n22689 );
nand ( n24366 , n24364 , n24365 );
buf ( n24367 , n24366 );
buf ( n24368 , n24367 );
nand ( n24369 , n24363 , n24368 );
buf ( n24370 , n24369 );
nand ( n24371 , n24354 , n24370 );
nand ( n24372 , n24353 , n24371 );
buf ( n24373 , n858 );
buf ( n24374 , n872 );
xor ( n24375 , n24373 , n24374 );
buf ( n24376 , n24375 );
buf ( n24377 , n24376 );
not ( n24378 , n24377 );
buf ( n24379 , n20211 );
not ( n24380 , n24379 );
or ( n24381 , n24378 , n24380 );
buf ( n24382 , n22611 );
buf ( n24383 , n19234 );
nand ( n24384 , n24382 , n24383 );
buf ( n24385 , n24384 );
buf ( n24386 , n24385 );
nand ( n24387 , n24381 , n24386 );
buf ( n24388 , n24387 );
buf ( n24389 , n24388 );
not ( n24390 , n24389 );
buf ( n24391 , n846 );
buf ( n24392 , n884 );
xor ( n24393 , n24391 , n24392 );
buf ( n24394 , n24393 );
buf ( n24395 , n24394 );
not ( n24396 , n24395 );
buf ( n24397 , n20694 );
not ( n24398 , n24397 );
or ( n24399 , n24396 , n24398 );
buf ( n24400 , n20700 );
buf ( n24401 , n22672 );
nand ( n24402 , n24400 , n24401 );
buf ( n24403 , n24402 );
buf ( n24404 , n24403 );
nand ( n24405 , n24399 , n24404 );
buf ( n24406 , n24405 );
buf ( n24407 , n24406 );
not ( n24408 , n24407 );
or ( n24409 , n24390 , n24408 );
or ( n24410 , n24406 , n24388 );
buf ( n24411 , n860 );
buf ( n24412 , n870 );
xor ( n24413 , n24411 , n24412 );
buf ( n24414 , n24413 );
not ( n24415 , n24414 );
not ( n24416 , n19122 );
or ( n24417 , n24415 , n24416 );
buf ( n24418 , n22573 );
buf ( n24419 , n21727 );
nand ( n24420 , n24418 , n24419 );
buf ( n24421 , n24420 );
nand ( n24422 , n24417 , n24421 );
nand ( n24423 , n24410 , n24422 );
buf ( n24424 , n24423 );
nand ( n24425 , n24409 , n24424 );
buf ( n24426 , n24425 );
or ( n24427 , n24372 , n24426 );
not ( n24428 , n24427 );
xor ( n24429 , n22835 , n22848 );
xnor ( n24430 , n24429 , n22823 );
not ( n24431 , n24430 );
or ( n24432 , n24428 , n24431 );
nand ( n24433 , n24426 , n24372 );
nand ( n24434 , n24432 , n24433 );
buf ( n24435 , n24434 );
xor ( n24436 , n24322 , n24435 );
xor ( n24437 , n22959 , n22976 );
xor ( n24438 , n24437 , n22973 );
buf ( n24439 , n24438 );
and ( n24440 , n24436 , n24439 );
and ( n24441 , n24322 , n24435 );
or ( n24442 , n24440 , n24441 );
buf ( n24443 , n24442 );
buf ( n24444 , n24443 );
and ( n24445 , n24309 , n24444 );
and ( n24446 , n24091 , n24308 );
or ( n24447 , n24445 , n24446 );
buf ( n24448 , n24447 );
buf ( n24449 , n24448 );
xor ( n24450 , n22856 , n22860 );
xor ( n24451 , n24450 , n22870 );
buf ( n24452 , n24451 );
buf ( n24453 , n24452 );
xor ( n24454 , n22894 , n22981 );
xor ( n24455 , n24454 , n22997 );
buf ( n24456 , n24455 );
buf ( n24457 , n24456 );
xor ( n24458 , n24453 , n24457 );
xor ( n24459 , n22878 , n22884 );
xor ( n24460 , n24459 , n22881 );
buf ( n24461 , n24460 );
xor ( n24462 , n22953 , n22923 );
xor ( n24463 , n24462 , n22927 );
buf ( n24464 , n24463 );
buf ( n24465 , n839 );
buf ( n24466 , n892 );
xor ( n24467 , n24465 , n24466 );
buf ( n24468 , n24467 );
not ( n24469 , n24468 );
not ( n24470 , n20599 );
or ( n24471 , n24469 , n24470 );
buf ( n24472 , n23181 );
buf ( n24473 , n24126 );
nand ( n24474 , n24472 , n24473 );
buf ( n24475 , n24474 );
nand ( n24476 , n24471 , n24475 );
buf ( n24477 , n24476 );
buf ( n24478 , n863 );
buf ( n24479 , n869 );
or ( n24480 , n24478 , n24479 );
buf ( n24481 , n870 );
nand ( n24482 , n24480 , n24481 );
buf ( n24483 , n24482 );
buf ( n24484 , n863 );
buf ( n24485 , n869 );
nand ( n24486 , n24484 , n24485 );
buf ( n24487 , n24486 );
and ( n24488 , n24483 , n24487 , n868 );
buf ( n24489 , n24488 );
and ( n24490 , n24477 , n24489 );
buf ( n24491 , n24490 );
not ( n24492 , n24150 );
not ( n24493 , n20325 );
or ( n24494 , n24492 , n24493 );
not ( n24495 , n18847 );
buf ( n24496 , n851 );
buf ( n24497 , n880 );
xor ( n24498 , n24496 , n24497 );
buf ( n24499 , n24498 );
nand ( n24500 , n24495 , n24499 , n22828 );
nand ( n24501 , n24494 , n24500 );
buf ( n24502 , n24501 );
not ( n24503 , n24502 );
buf ( n24504 , n24503 );
not ( n24505 , n24504 );
buf ( n24506 , n843 );
buf ( n24507 , n888 );
xor ( n24508 , n24506 , n24507 );
buf ( n24509 , n24508 );
buf ( n24510 , n24509 );
not ( n24511 , n24510 );
buf ( n24512 , n20357 );
not ( n24513 , n24512 );
or ( n24514 , n24511 , n24513 );
buf ( n24515 , n20363 );
buf ( n24516 , n24099 );
nand ( n24517 , n24515 , n24516 );
buf ( n24518 , n24517 );
buf ( n24519 , n24518 );
nand ( n24520 , n24514 , n24519 );
buf ( n24521 , n24520 );
buf ( n24522 , n24521 );
not ( n24523 , n24522 );
buf ( n24524 , n24523 );
not ( n24525 , n24524 );
or ( n24526 , n24505 , n24525 );
buf ( n24527 , n853 );
buf ( n24528 , n878 );
xor ( n24529 , n24527 , n24528 );
buf ( n24530 , n24529 );
buf ( n24531 , n24530 );
not ( n24532 , n24531 );
buf ( n24533 , n19259 );
not ( n24534 , n24533 );
or ( n24535 , n24532 , n24534 );
buf ( n24536 , n19265 );
buf ( n24537 , n24164 );
nand ( n24538 , n24536 , n24537 );
buf ( n24539 , n24538 );
buf ( n24540 , n24539 );
nand ( n24541 , n24535 , n24540 );
buf ( n24542 , n24541 );
nand ( n24543 , n24526 , n24542 );
buf ( n24544 , n24521 );
buf ( n24545 , n24501 );
nand ( n24546 , n24544 , n24545 );
buf ( n24547 , n24546 );
nand ( n24548 , n24543 , n24547 );
xor ( n24549 , n24491 , n24548 );
buf ( n24550 , n845 );
buf ( n24551 , n886 );
xor ( n24552 , n24550 , n24551 );
buf ( n24553 , n24552 );
buf ( n24554 , n24553 );
not ( n24555 , n24554 );
buf ( n24556 , n20521 );
not ( n24557 , n24556 );
or ( n24558 , n24555 , n24557 );
buf ( n24559 , n20525 );
buf ( n24560 , n24182 );
nand ( n24561 , n24559 , n24560 );
buf ( n24562 , n24561 );
buf ( n24563 , n24562 );
nand ( n24564 , n24558 , n24563 );
buf ( n24565 , n24564 );
not ( n24566 , n24565 );
buf ( n24567 , n855 );
buf ( n24568 , n876 );
xor ( n24569 , n24567 , n24568 );
buf ( n24570 , n24569 );
buf ( n24571 , n24570 );
not ( n24572 , n24571 );
buf ( n24573 , n19077 );
not ( n24574 , n24573 );
or ( n24575 , n24572 , n24574 );
buf ( n24576 , n19082 );
buf ( n24577 , n24226 );
nand ( n24578 , n24576 , n24577 );
buf ( n24579 , n24578 );
buf ( n24580 , n24579 );
nand ( n24581 , n24575 , n24580 );
buf ( n24582 , n24581 );
not ( n24583 , n24582 );
or ( n24584 , n24566 , n24583 );
buf ( n24585 , n24565 );
buf ( n24586 , n24582 );
nor ( n24587 , n24585 , n24586 );
buf ( n24588 , n24587 );
buf ( n24589 , n18977 );
buf ( n24590 , n857 );
buf ( n24591 , n874 );
xor ( n24592 , n24590 , n24591 );
buf ( n24593 , n24592 );
buf ( n24594 , n24593 );
and ( n24595 , n24589 , n24594 );
buf ( n24596 , n20555 );
buf ( n24597 , n24245 );
and ( n24598 , n24596 , n24597 );
nor ( n24599 , n24595 , n24598 );
buf ( n24600 , n24599 );
or ( n24601 , n24588 , n24600 );
nand ( n24602 , n24584 , n24601 );
and ( n24603 , n24549 , n24602 );
and ( n24604 , n24491 , n24548 );
or ( n24605 , n24603 , n24604 );
buf ( n24606 , n24605 );
xor ( n24607 , n24464 , n24606 );
buf ( n24608 , n18944 );
buf ( n24609 , n863 );
nand ( n24610 , n24608 , n24609 );
buf ( n24611 , n24610 );
buf ( n24612 , n24611 );
buf ( n24613 , n24138 );
xor ( n24614 , n24612 , n24613 );
buf ( n24615 , n24111 );
xor ( n24616 , n24614 , n24615 );
buf ( n24617 , n24616 );
buf ( n24618 , n24617 );
not ( n24619 , n24618 );
not ( n24620 , n24351 );
not ( n24621 , n24334 );
not ( n24622 , n24370 );
and ( n24623 , n24621 , n24622 );
and ( n24624 , n24334 , n24370 );
nor ( n24625 , n24623 , n24624 );
not ( n24626 , n24625 );
or ( n24627 , n24620 , n24626 );
or ( n24628 , n24351 , n24625 );
nand ( n24629 , n24627 , n24628 );
buf ( n24630 , n24629 );
not ( n24631 , n24630 );
or ( n24632 , n24619 , n24631 );
buf ( n24633 , n24221 );
buf ( n24634 , n24234 );
xor ( n24635 , n24633 , n24634 );
buf ( n24636 , n24252 );
xnor ( n24637 , n24635 , n24636 );
buf ( n24638 , n24637 );
buf ( n24639 , n24638 );
nand ( n24640 , n24632 , n24639 );
buf ( n24641 , n24640 );
buf ( n24642 , n24641 );
buf ( n24643 , n24629 );
not ( n24644 , n24643 );
buf ( n24645 , n24617 );
not ( n24646 , n24645 );
buf ( n24647 , n24646 );
buf ( n24648 , n24647 );
nand ( n24649 , n24644 , n24648 );
buf ( n24650 , n24649 );
buf ( n24651 , n24650 );
nand ( n24652 , n24642 , n24651 );
buf ( n24653 , n24652 );
buf ( n24654 , n24653 );
and ( n24655 , n24607 , n24654 );
and ( n24656 , n24464 , n24606 );
or ( n24657 , n24655 , n24656 );
buf ( n24658 , n24657 );
buf ( n24659 , n24658 );
xor ( n24660 , n24461 , n24659 );
not ( n24661 , n24255 );
not ( n24662 , n24144 );
or ( n24663 , n24661 , n24662 );
buf ( n24664 , n24254 );
not ( n24665 , n24664 );
buf ( n24666 , n24143 );
nand ( n24667 , n24665 , n24666 );
buf ( n24668 , n24667 );
nand ( n24669 , n24663 , n24668 );
and ( n24670 , n24669 , n24202 );
not ( n24671 , n24669 );
and ( n24672 , n24671 , n24199 );
nor ( n24673 , n24670 , n24672 );
buf ( n24674 , n24673 );
not ( n24675 , n24674 );
buf ( n24676 , n24426 );
buf ( n24677 , n24372 );
xor ( n24678 , n24676 , n24677 );
buf ( n24679 , n24430 );
xnor ( n24680 , n24678 , n24679 );
buf ( n24681 , n24680 );
buf ( n24682 , n24681 );
not ( n24683 , n24682 );
or ( n24684 , n24675 , n24683 );
buf ( n24685 , n837 );
buf ( n24686 , n894 );
xor ( n24687 , n24685 , n24686 );
buf ( n24688 , n24687 );
buf ( n24689 , n24688 );
not ( n24690 , n24689 );
buf ( n24691 , n21297 );
not ( n24692 , n24691 );
or ( n24693 , n24690 , n24692 );
buf ( n24694 , n24209 );
buf ( n24695 , n895 );
nand ( n24696 , n24694 , n24695 );
buf ( n24697 , n24696 );
buf ( n24698 , n24697 );
nand ( n24699 , n24693 , n24698 );
buf ( n24700 , n24699 );
buf ( n24701 , n24700 );
buf ( n24702 , n847 );
buf ( n24703 , n884 );
xor ( n24704 , n24702 , n24703 );
buf ( n24705 , n24704 );
buf ( n24706 , n24705 );
not ( n24707 , n24706 );
buf ( n24708 , n20694 );
not ( n24709 , n24708 );
or ( n24710 , n24707 , n24709 );
buf ( n24711 , n20700 );
buf ( n24712 , n24394 );
nand ( n24713 , n24711 , n24712 );
buf ( n24714 , n24713 );
buf ( n24715 , n24714 );
nand ( n24716 , n24710 , n24715 );
buf ( n24717 , n24716 );
buf ( n24718 , n24717 );
xor ( n24719 , n24701 , n24718 );
xor ( n24720 , n872 , n859 );
buf ( n24721 , n24720 );
not ( n24722 , n24721 );
buf ( n24723 , n19230 );
not ( n24724 , n24723 );
or ( n24725 , n24722 , n24724 );
buf ( n24726 , n19234 );
buf ( n24727 , n24376 );
nand ( n24728 , n24726 , n24727 );
buf ( n24729 , n24728 );
buf ( n24730 , n24729 );
nand ( n24731 , n24725 , n24730 );
buf ( n24732 , n24731 );
buf ( n24733 , n24732 );
and ( n24734 , n24719 , n24733 );
and ( n24735 , n24701 , n24718 );
or ( n24736 , n24734 , n24735 );
buf ( n24737 , n24736 );
buf ( n24738 , n24737 );
buf ( n24739 , n841 );
buf ( n24740 , n890 );
xor ( n24741 , n24739 , n24740 );
buf ( n24742 , n24741 );
buf ( n24743 , n24742 );
not ( n24744 , n24743 );
buf ( n24745 , n21441 );
not ( n24746 , n24745 );
or ( n24747 , n24744 , n24746 );
buf ( n24748 , n20869 );
buf ( n24749 , n24358 );
nand ( n24750 , n24748 , n24749 );
buf ( n24751 , n24750 );
buf ( n24752 , n24751 );
nand ( n24753 , n24747 , n24752 );
buf ( n24754 , n24753 );
buf ( n24755 , n24754 );
not ( n24756 , n24755 );
buf ( n24757 , n863 );
buf ( n24758 , n868 );
xor ( n24759 , n24757 , n24758 );
buf ( n24760 , n24759 );
buf ( n24761 , n24760 );
not ( n24762 , n24761 );
buf ( n24763 , n23893 );
not ( n24764 , n24763 );
or ( n24765 , n24762 , n24764 );
buf ( n24766 , n22916 );
buf ( n24767 , n24339 );
nand ( n24768 , n24766 , n24767 );
buf ( n24769 , n24768 );
buf ( n24770 , n24769 );
nand ( n24771 , n24765 , n24770 );
buf ( n24772 , n24771 );
buf ( n24773 , n24772 );
not ( n24774 , n24773 );
or ( n24775 , n24756 , n24774 );
buf ( n24776 , n24754 );
buf ( n24777 , n24772 );
or ( n24778 , n24776 , n24777 );
buf ( n24779 , n861 );
buf ( n24780 , n870 );
xor ( n24781 , n24779 , n24780 );
buf ( n24782 , n24781 );
buf ( n24783 , n24782 );
not ( n24784 , n24783 );
buf ( n24785 , n19122 );
not ( n24786 , n24785 );
or ( n24787 , n24784 , n24786 );
buf ( n24788 , n21727 );
buf ( n24789 , n24414 );
nand ( n24790 , n24788 , n24789 );
buf ( n24791 , n24790 );
buf ( n24792 , n24791 );
nand ( n24793 , n24787 , n24792 );
buf ( n24794 , n24793 );
buf ( n24795 , n24794 );
nand ( n24796 , n24778 , n24795 );
buf ( n24797 , n24796 );
buf ( n24798 , n24797 );
nand ( n24799 , n24775 , n24798 );
buf ( n24800 , n24799 );
buf ( n24801 , n24800 );
xor ( n24802 , n24738 , n24801 );
xor ( n24803 , n24160 , n24177 );
xor ( n24804 , n24803 , n24195 );
buf ( n24805 , n24804 );
buf ( n24806 , n24805 );
and ( n24807 , n24802 , n24806 );
and ( n24808 , n24738 , n24801 );
or ( n24809 , n24807 , n24808 );
buf ( n24810 , n24809 );
buf ( n24811 , n24810 );
nand ( n24812 , n24684 , n24811 );
buf ( n24813 , n24812 );
buf ( n24814 , n24813 );
buf ( n24815 , n24673 );
not ( n24816 , n24815 );
buf ( n24817 , n24681 );
not ( n24818 , n24817 );
buf ( n24819 , n24818 );
buf ( n24820 , n24819 );
nand ( n24821 , n24816 , n24820 );
buf ( n24822 , n24821 );
buf ( n24823 , n24822 );
nand ( n24824 , n24814 , n24823 );
buf ( n24825 , n24824 );
buf ( n24826 , n24825 );
and ( n24827 , n24660 , n24826 );
and ( n24828 , n24461 , n24659 );
or ( n24829 , n24827 , n24828 );
buf ( n24830 , n24829 );
buf ( n24831 , n24830 );
and ( n24832 , n24458 , n24831 );
and ( n24833 , n24453 , n24457 );
or ( n24834 , n24832 , n24833 );
buf ( n24835 , n24834 );
buf ( n24836 , n24835 );
xor ( n24837 , n24449 , n24836 );
xor ( n24838 , n22042 , n22048 );
xor ( n24839 , n24838 , n22094 );
buf ( n24840 , n24839 );
xor ( n24841 , n22733 , n22736 );
xor ( n24842 , n24841 , n22740 );
buf ( n24843 , n24842 );
buf ( n24844 , n24843 );
xor ( n24845 , n24840 , n24844 );
xor ( n24846 , n22753 , n22875 );
xor ( n24847 , n24846 , n23002 );
buf ( n24848 , n24847 );
buf ( n24849 , n24848 );
xor ( n24850 , n24845 , n24849 );
buf ( n24851 , n24850 );
buf ( n24852 , n24851 );
xor ( n24853 , n24837 , n24852 );
buf ( n24854 , n24853 );
buf ( n24855 , n24854 );
buf ( n24856 , n851 );
buf ( n24857 , n866 );
xor ( n24858 , n24856 , n24857 );
buf ( n24859 , n24858 );
buf ( n24860 , n24859 );
not ( n24861 , n24860 );
buf ( n24862 , n18931 );
not ( n24863 , n24862 );
or ( n24864 , n24861 , n24863 );
buf ( n24865 , n21249 );
buf ( n24866 , n850 );
buf ( n24867 , n866 );
xor ( n24868 , n24866 , n24867 );
buf ( n24869 , n24868 );
buf ( n24870 , n24869 );
nand ( n24871 , n24865 , n24870 );
buf ( n24872 , n24871 );
buf ( n24873 , n24872 );
nand ( n24874 , n24864 , n24873 );
buf ( n24875 , n24874 );
buf ( n24876 , n849 );
buf ( n24877 , n868 );
xor ( n24878 , n24876 , n24877 );
buf ( n24879 , n24878 );
buf ( n24880 , n24879 );
not ( n24881 , n24880 );
buf ( n24882 , n18887 );
not ( n24883 , n24882 );
or ( n24884 , n24881 , n24883 );
buf ( n24885 , n22916 );
buf ( n24886 , n848 );
buf ( n24887 , n868 );
xor ( n24888 , n24886 , n24887 );
buf ( n24889 , n24888 );
buf ( n24890 , n24889 );
nand ( n24891 , n24885 , n24890 );
buf ( n24892 , n24891 );
buf ( n24893 , n24892 );
nand ( n24894 , n24884 , n24893 );
buf ( n24895 , n24894 );
xor ( n24896 , n24875 , n24895 );
buf ( n24897 , n835 );
buf ( n24898 , n882 );
xor ( n24899 , n24897 , n24898 );
buf ( n24900 , n24899 );
buf ( n24901 , n24900 );
not ( n24902 , n24901 );
buf ( n24903 , n19580 );
not ( n24904 , n24903 );
or ( n24905 , n24902 , n24904 );
buf ( n24906 , n19909 );
buf ( n24907 , n834 );
buf ( n24908 , n882 );
xor ( n24909 , n24907 , n24908 );
buf ( n24910 , n24909 );
buf ( n24911 , n24910 );
nand ( n24912 , n24906 , n24911 );
buf ( n24913 , n24912 );
buf ( n24914 , n24913 );
nand ( n24915 , n24905 , n24914 );
buf ( n24916 , n24915 );
not ( n24917 , n24916 );
and ( n24918 , n24896 , n24917 );
not ( n24919 , n24896 );
and ( n24920 , n24919 , n24916 );
nor ( n24921 , n24918 , n24920 );
buf ( n24922 , n847 );
buf ( n24923 , n870 );
xor ( n24924 , n24922 , n24923 );
buf ( n24925 , n24924 );
buf ( n24926 , n24925 );
not ( n24927 , n24926 );
buf ( n24928 , n19122 );
not ( n24929 , n24928 );
or ( n24930 , n24927 , n24929 );
buf ( n24931 , n19131 );
buf ( n24932 , n846 );
buf ( n24933 , n870 );
xor ( n24934 , n24932 , n24933 );
buf ( n24935 , n24934 );
buf ( n24936 , n24935 );
nand ( n24937 , n24931 , n24936 );
buf ( n24938 , n24937 );
buf ( n24939 , n24938 );
nand ( n24940 , n24930 , n24939 );
buf ( n24941 , n24940 );
buf ( n24942 , n24941 );
buf ( n24943 , n845 );
buf ( n24944 , n872 );
xor ( n24945 , n24943 , n24944 );
buf ( n24946 , n24945 );
buf ( n24947 , n24946 );
not ( n24948 , n24947 );
buf ( n24949 , n19230 );
not ( n24950 , n24949 );
or ( n24951 , n24948 , n24950 );
buf ( n24952 , n19235 );
buf ( n24953 , n844 );
buf ( n24954 , n872 );
xor ( n24955 , n24953 , n24954 );
buf ( n24956 , n24955 );
buf ( n24957 , n24956 );
nand ( n24958 , n24952 , n24957 );
buf ( n24959 , n24958 );
buf ( n24960 , n24959 );
nand ( n24961 , n24951 , n24960 );
buf ( n24962 , n24961 );
buf ( n24963 , n24962 );
xor ( n24964 , n24942 , n24963 );
buf ( n24965 , n839 );
buf ( n24966 , n878 );
xor ( n24967 , n24965 , n24966 );
buf ( n24968 , n24967 );
buf ( n24969 , n24968 );
not ( n24970 , n24969 );
buf ( n24971 , n19259 );
not ( n24972 , n24971 );
or ( n24973 , n24970 , n24972 );
buf ( n24974 , n19265 );
buf ( n24975 , n838 );
buf ( n24976 , n878 );
xor ( n24977 , n24975 , n24976 );
buf ( n24978 , n24977 );
buf ( n24979 , n24978 );
nand ( n24980 , n24974 , n24979 );
buf ( n24981 , n24980 );
buf ( n24982 , n24981 );
nand ( n24983 , n24973 , n24982 );
buf ( n24984 , n24983 );
buf ( n24985 , n24984 );
xor ( n24986 , n24964 , n24985 );
buf ( n24987 , n24986 );
not ( n24988 , n24987 );
xor ( n24989 , n24921 , n24988 );
not ( n24990 , n20525 );
not ( n24991 , n24990 );
buf ( n24992 , n20521 );
not ( n24993 , n24992 );
buf ( n24994 , n24993 );
not ( n24995 , n24994 );
or ( n24996 , n24991 , n24995 );
nand ( n24997 , n24996 , n886 );
buf ( n24998 , n837 );
buf ( n24999 , n880 );
xor ( n25000 , n24998 , n24999 );
buf ( n25001 , n25000 );
not ( n25002 , n25001 );
not ( n25003 , n18850 );
or ( n25004 , n25002 , n25003 );
buf ( n25005 , n22271 );
buf ( n25006 , n836 );
buf ( n25007 , n880 );
xor ( n25008 , n25006 , n25007 );
buf ( n25009 , n25008 );
buf ( n25010 , n25009 );
nand ( n25011 , n25005 , n25010 );
buf ( n25012 , n25011 );
nand ( n25013 , n25004 , n25012 );
xor ( n25014 , n24997 , n25013 );
buf ( n25015 , n833 );
buf ( n25016 , n884 );
xor ( n25017 , n25015 , n25016 );
buf ( n25018 , n25017 );
not ( n25019 , n25018 );
buf ( n25020 , n20694 );
buf ( n25021 , n25020 );
buf ( n25022 , n25021 );
not ( n25023 , n25022 );
or ( n25024 , n25019 , n25023 );
buf ( n25025 , n23233 );
buf ( n25026 , n832 );
buf ( n25027 , n884 );
xor ( n25028 , n25026 , n25027 );
buf ( n25029 , n25028 );
buf ( n25030 , n25029 );
nand ( n25031 , n25025 , n25030 );
buf ( n25032 , n25031 );
nand ( n25033 , n25024 , n25032 );
xor ( n25034 , n25014 , n25033 );
xor ( n25035 , n24989 , n25034 );
buf ( n25036 , n854 );
buf ( n25037 , n864 );
and ( n25038 , n25036 , n25037 );
buf ( n25039 , n25038 );
buf ( n25040 , n25039 );
buf ( n25041 , n853 );
buf ( n25042 , n864 );
xor ( n25043 , n25041 , n25042 );
buf ( n25044 , n25043 );
buf ( n25045 , n25044 );
not ( n25046 , n25045 );
buf ( n25047 , n19013 );
not ( n25048 , n25047 );
or ( n25049 , n25046 , n25048 );
buf ( n25050 , n19030 );
buf ( n25051 , n852 );
buf ( n25052 , n864 );
xor ( n25053 , n25051 , n25052 );
buf ( n25054 , n25053 );
buf ( n25055 , n25054 );
nand ( n25056 , n25050 , n25055 );
buf ( n25057 , n25056 );
buf ( n25058 , n25057 );
nand ( n25059 , n25049 , n25058 );
buf ( n25060 , n25059 );
buf ( n25061 , n25060 );
xor ( n25062 , n25040 , n25061 );
buf ( n25063 , n841 );
buf ( n25064 , n876 );
xor ( n25065 , n25063 , n25064 );
buf ( n25066 , n25065 );
buf ( n25067 , n25066 );
not ( n25068 , n25067 );
buf ( n25069 , n19077 );
not ( n25070 , n25069 );
or ( n25071 , n25068 , n25070 );
buf ( n25072 , n20246 );
buf ( n25073 , n840 );
buf ( n25074 , n876 );
xor ( n25075 , n25073 , n25074 );
buf ( n25076 , n25075 );
buf ( n25077 , n25076 );
nand ( n25078 , n25072 , n25077 );
buf ( n25079 , n25078 );
buf ( n25080 , n25079 );
nand ( n25081 , n25071 , n25080 );
buf ( n25082 , n25081 );
buf ( n25083 , n25082 );
xor ( n25084 , n25062 , n25083 );
buf ( n25085 , n25084 );
buf ( n25086 , n25085 );
xor ( n25087 , n874 , n843 );
buf ( n25088 , n25087 );
not ( n25089 , n25088 );
buf ( n25090 , n20549 );
not ( n25091 , n25090 );
or ( n25092 , n25089 , n25091 );
buf ( n25093 , n18987 );
buf ( n25094 , n842 );
buf ( n25095 , n874 );
xor ( n25096 , n25094 , n25095 );
buf ( n25097 , n25096 );
buf ( n25098 , n25097 );
nand ( n25099 , n25093 , n25098 );
buf ( n25100 , n25099 );
buf ( n25101 , n25100 );
nand ( n25102 , n25092 , n25101 );
buf ( n25103 , n25102 );
buf ( n25104 , n25103 );
buf ( n25105 , n834 );
buf ( n25106 , n884 );
xor ( n25107 , n25105 , n25106 );
buf ( n25108 , n25107 );
buf ( n25109 , n25108 );
not ( n25110 , n25109 );
buf ( n25111 , n25022 );
not ( n25112 , n25111 );
or ( n25113 , n25110 , n25112 );
buf ( n25114 , n23233 );
buf ( n25115 , n25018 );
nand ( n25116 , n25114 , n25115 );
buf ( n25117 , n25116 );
buf ( n25118 , n25117 );
nand ( n25119 , n25113 , n25118 );
buf ( n25120 , n25119 );
buf ( n25121 , n25120 );
xor ( n25122 , n25104 , n25121 );
buf ( n25123 , n850 );
buf ( n25124 , n868 );
xor ( n25125 , n25123 , n25124 );
buf ( n25126 , n25125 );
buf ( n25127 , n25126 );
not ( n25128 , n25127 );
buf ( n25129 , n23893 );
not ( n25130 , n25129 );
or ( n25131 , n25128 , n25130 );
buf ( n25132 , n22916 );
buf ( n25133 , n24879 );
nand ( n25134 , n25132 , n25133 );
buf ( n25135 , n25134 );
buf ( n25136 , n25135 );
nand ( n25137 , n25131 , n25136 );
buf ( n25138 , n25137 );
not ( n25139 , n25138 );
buf ( n25140 , n852 );
buf ( n25141 , n866 );
xor ( n25142 , n25140 , n25141 );
buf ( n25143 , n25142 );
buf ( n25144 , n25143 );
not ( n25145 , n25144 );
buf ( n25146 , n18931 );
not ( n25147 , n25146 );
or ( n25148 , n25145 , n25147 );
buf ( n25149 , n18938 );
buf ( n25150 , n24859 );
nand ( n25151 , n25149 , n25150 );
buf ( n25152 , n25151 );
buf ( n25153 , n25152 );
nand ( n25154 , n25148 , n25153 );
buf ( n25155 , n25154 );
not ( n25156 , n25155 );
or ( n25157 , n25139 , n25156 );
buf ( n25158 , n25138 );
buf ( n25159 , n25155 );
nor ( n25160 , n25158 , n25159 );
buf ( n25161 , n25160 );
buf ( n25162 , n840 );
buf ( n25163 , n878 );
xor ( n25164 , n25162 , n25163 );
buf ( n25165 , n25164 );
buf ( n25166 , n25165 );
not ( n25167 , n25166 );
buf ( n25168 , n19259 );
not ( n25169 , n25168 );
or ( n25170 , n25167 , n25169 );
buf ( n25171 , n19265 );
buf ( n25172 , n24968 );
nand ( n25173 , n25171 , n25172 );
buf ( n25174 , n25173 );
buf ( n25175 , n25174 );
nand ( n25176 , n25170 , n25175 );
buf ( n25177 , n25176 );
buf ( n25178 , n25177 );
not ( n25179 , n25178 );
buf ( n25180 , n25179 );
or ( n25181 , n25161 , n25180 );
nand ( n25182 , n25157 , n25181 );
buf ( n25183 , n25182 );
xor ( n25184 , n25122 , n25183 );
buf ( n25185 , n25184 );
buf ( n25186 , n25185 );
xor ( n25187 , n25086 , n25186 );
buf ( n25188 , n25108 );
not ( n25189 , n25188 );
buf ( n25190 , n25022 );
not ( n25191 , n25190 );
or ( n25192 , n25189 , n25191 );
buf ( n25193 , n25117 );
nand ( n25194 , n25192 , n25193 );
buf ( n25195 , n25194 );
buf ( n25196 , n25195 );
not ( n25197 , n25196 );
buf ( n25198 , n25197 );
buf ( n25199 , n25198 );
buf ( n25200 , n851 );
buf ( n25201 , n868 );
xor ( n25202 , n25200 , n25201 );
buf ( n25203 , n25202 );
buf ( n25204 , n25203 );
not ( n25205 , n25204 );
buf ( n25206 , n23893 );
not ( n25207 , n25206 );
or ( n25208 , n25205 , n25207 );
buf ( n25209 , n18892 );
buf ( n25210 , n25126 );
nand ( n25211 , n25209 , n25210 );
buf ( n25212 , n25211 );
buf ( n25213 , n25212 );
nand ( n25214 , n25208 , n25213 );
buf ( n25215 , n25214 );
buf ( n25216 , n25215 );
not ( n25217 , n25216 );
buf ( n25218 , n849 );
buf ( n25219 , n870 );
xor ( n25220 , n25218 , n25219 );
buf ( n25221 , n25220 );
buf ( n25222 , n25221 );
not ( n25223 , n25222 );
buf ( n25224 , n20805 );
not ( n25225 , n25224 );
or ( n25226 , n25223 , n25225 );
buf ( n25227 , n19131 );
buf ( n25228 , n848 );
buf ( n25229 , n870 );
xor ( n25230 , n25228 , n25229 );
buf ( n25231 , n25230 );
buf ( n25232 , n25231 );
nand ( n25233 , n25227 , n25232 );
buf ( n25234 , n25233 );
buf ( n25235 , n25234 );
nand ( n25236 , n25226 , n25235 );
buf ( n25237 , n25236 );
buf ( n25238 , n25237 );
not ( n25239 , n25238 );
or ( n25240 , n25217 , n25239 );
buf ( n25241 , n25237 );
not ( n25242 , n25241 );
buf ( n25243 , n25242 );
buf ( n25244 , n25243 );
not ( n25245 , n25244 );
buf ( n25246 , n25215 );
not ( n25247 , n25246 );
buf ( n25248 , n25247 );
buf ( n25249 , n25248 );
not ( n25250 , n25249 );
or ( n25251 , n25245 , n25250 );
buf ( n25252 , n835 );
buf ( n25253 , n884 );
xor ( n25254 , n25252 , n25253 );
buf ( n25255 , n25254 );
buf ( n25256 , n25255 );
not ( n25257 , n25256 );
buf ( n25258 , n25022 );
not ( n25259 , n25258 );
or ( n25260 , n25257 , n25259 );
buf ( n25261 , n20700 );
buf ( n25262 , n25261 );
buf ( n25263 , n25262 );
buf ( n25264 , n25263 );
buf ( n25265 , n25108 );
nand ( n25266 , n25264 , n25265 );
buf ( n25267 , n25266 );
buf ( n25268 , n25267 );
nand ( n25269 , n25260 , n25268 );
buf ( n25270 , n25269 );
buf ( n25271 , n25270 );
nand ( n25272 , n25251 , n25271 );
buf ( n25273 , n25272 );
buf ( n25274 , n25273 );
nand ( n25275 , n25240 , n25274 );
buf ( n25276 , n25275 );
buf ( n25277 , n25276 );
xor ( n25278 , n25199 , n25277 );
buf ( n25279 , n847 );
buf ( n25280 , n872 );
xor ( n25281 , n25279 , n25280 );
buf ( n25282 , n25281 );
buf ( n25283 , n25282 );
not ( n25284 , n25283 );
not ( n25285 , n20210 );
buf ( n25286 , n25285 );
not ( n25287 , n25286 );
or ( n25288 , n25284 , n25287 );
buf ( n25289 , n19234 );
buf ( n25290 , n846 );
buf ( n25291 , n872 );
xor ( n25292 , n25290 , n25291 );
buf ( n25293 , n25292 );
buf ( n25294 , n25293 );
nand ( n25295 , n25289 , n25294 );
buf ( n25296 , n25295 );
buf ( n25297 , n25296 );
nand ( n25298 , n25288 , n25297 );
buf ( n25299 , n25298 );
buf ( n25300 , n25299 );
buf ( n25301 , n845 );
buf ( n25302 , n874 );
xor ( n25303 , n25301 , n25302 );
buf ( n25304 , n25303 );
buf ( n25305 , n25304 );
not ( n25306 , n25305 );
buf ( n25307 , n18974 );
not ( n25308 , n25307 );
or ( n25309 , n25306 , n25308 );
buf ( n25310 , n21513 );
xor ( n25311 , n874 , n844 );
buf ( n25312 , n25311 );
nand ( n25313 , n25310 , n25312 );
buf ( n25314 , n25313 );
buf ( n25315 , n25314 );
nand ( n25316 , n25309 , n25315 );
buf ( n25317 , n25316 );
buf ( n25318 , n25317 );
xor ( n25319 , n25300 , n25318 );
buf ( n25320 , n839 );
buf ( n25321 , n880 );
xor ( n25322 , n25320 , n25321 );
buf ( n25323 , n25322 );
buf ( n25324 , n25323 );
not ( n25325 , n25324 );
buf ( n25326 , n18850 );
not ( n25327 , n25326 );
or ( n25328 , n25325 , n25327 );
buf ( n25329 , n23917 );
buf ( n25330 , n838 );
buf ( n25331 , n880 );
xor ( n25332 , n25330 , n25331 );
buf ( n25333 , n25332 );
buf ( n25334 , n25333 );
nand ( n25335 , n25329 , n25334 );
buf ( n25336 , n25335 );
buf ( n25337 , n25336 );
nand ( n25338 , n25328 , n25337 );
buf ( n25339 , n25338 );
buf ( n25340 , n25339 );
and ( n25341 , n25319 , n25340 );
and ( n25342 , n25300 , n25318 );
or ( n25343 , n25341 , n25342 );
buf ( n25344 , n25343 );
buf ( n25345 , n25344 );
and ( n25346 , n25278 , n25345 );
and ( n25347 , n25199 , n25277 );
or ( n25348 , n25346 , n25347 );
buf ( n25349 , n25348 );
buf ( n25350 , n25349 );
xor ( n25351 , n25187 , n25350 );
buf ( n25352 , n25351 );
xor ( n25353 , n25035 , n25352 );
buf ( n25354 , n856 );
buf ( n25355 , n864 );
and ( n25356 , n25354 , n25355 );
buf ( n25357 , n25356 );
buf ( n25358 , n25357 );
buf ( n25359 , n843 );
buf ( n25360 , n876 );
xor ( n25361 , n25359 , n25360 );
buf ( n25362 , n25361 );
buf ( n25363 , n25362 );
not ( n25364 , n25363 );
buf ( n25365 , n19153 );
not ( n25366 , n25365 );
or ( n25367 , n25364 , n25366 );
buf ( n25368 , n19082 );
buf ( n25369 , n842 );
buf ( n25370 , n876 );
xor ( n25371 , n25369 , n25370 );
buf ( n25372 , n25371 );
buf ( n25373 , n25372 );
nand ( n25374 , n25368 , n25373 );
buf ( n25375 , n25374 );
buf ( n25376 , n25375 );
nand ( n25377 , n25367 , n25376 );
buf ( n25378 , n25377 );
buf ( n25379 , n25378 );
xor ( n25380 , n25358 , n25379 );
buf ( n25381 , n23983 );
not ( n25382 , n25381 );
buf ( n25383 , n20521 );
not ( n25384 , n25383 );
or ( n25385 , n25382 , n25384 );
buf ( n25386 , n20525 );
buf ( n25387 , n833 );
buf ( n25388 , n886 );
xor ( n25389 , n25387 , n25388 );
buf ( n25390 , n25389 );
buf ( n25391 , n25390 );
nand ( n25392 , n25386 , n25391 );
buf ( n25393 , n25392 );
buf ( n25394 , n25393 );
nand ( n25395 , n25385 , n25394 );
buf ( n25396 , n25395 );
buf ( n25397 , n25396 );
and ( n25398 , n25380 , n25397 );
and ( n25399 , n25358 , n25379 );
or ( n25400 , n25398 , n25399 );
buf ( n25401 , n25400 );
buf ( n25402 , n25401 );
buf ( n25403 , n23922 );
not ( n25404 , n25403 );
buf ( n25405 , n20642 );
not ( n25406 , n25405 );
or ( n25407 , n25404 , n25406 );
buf ( n25408 , n20325 );
buf ( n25409 , n25323 );
nand ( n25410 , n25408 , n25409 );
buf ( n25411 , n25410 );
buf ( n25412 , n25411 );
nand ( n25413 , n25407 , n25412 );
buf ( n25414 , n25413 );
buf ( n25415 , n25414 );
buf ( n25416 , n23901 );
not ( n25417 , n25416 );
buf ( n25418 , n23893 );
not ( n25419 , n25418 );
or ( n25420 , n25417 , n25419 );
buf ( n25421 , n18892 );
buf ( n25422 , n25203 );
nand ( n25423 , n25421 , n25422 );
buf ( n25424 , n25423 );
buf ( n25425 , n25424 );
nand ( n25426 , n25420 , n25425 );
buf ( n25427 , n25426 );
buf ( n25428 , n25427 );
or ( n25429 , n25415 , n25428 );
buf ( n25430 , n23950 );
not ( n25431 , n25430 );
buf ( n25432 , n19122 );
not ( n25433 , n25432 );
or ( n25434 , n25431 , n25433 );
buf ( n25435 , n21727 );
buf ( n25436 , n25221 );
nand ( n25437 , n25435 , n25436 );
buf ( n25438 , n25437 );
buf ( n25439 , n25438 );
nand ( n25440 , n25434 , n25439 );
buf ( n25441 , n25440 );
buf ( n25442 , n25441 );
nand ( n25443 , n25429 , n25442 );
buf ( n25444 , n25443 );
buf ( n25445 , n25444 );
buf ( n25446 , n25427 );
buf ( n25447 , n25414 );
nand ( n25448 , n25446 , n25447 );
buf ( n25449 , n25448 );
buf ( n25450 , n25449 );
nand ( n25451 , n25445 , n25450 );
buf ( n25452 , n25451 );
buf ( n25453 , n25452 );
buf ( n25454 , n25285 );
buf ( n25455 , n23966 );
and ( n25456 , n25454 , n25455 );
buf ( n25457 , n19234 );
buf ( n25458 , n25282 );
and ( n25459 , n25457 , n25458 );
nor ( n25460 , n25456 , n25459 );
buf ( n25461 , n25460 );
buf ( n25462 , n25461 );
not ( n25463 , n25462 );
buf ( n25464 , n25463 );
buf ( n25465 , n25464 );
not ( n25466 , n25465 );
buf ( n25467 , n23654 );
not ( n25468 , n25467 );
buf ( n25469 , n19580 );
not ( n25470 , n25469 );
or ( n25471 , n25468 , n25470 );
buf ( n25472 , n837 );
buf ( n25473 , n882 );
xor ( n25474 , n25472 , n25473 );
buf ( n25475 , n25474 );
buf ( n25476 , n25475 );
buf ( n25477 , n19909 );
nand ( n25478 , n25476 , n25477 );
buf ( n25479 , n25478 );
buf ( n25480 , n25479 );
nand ( n25481 , n25471 , n25480 );
buf ( n25482 , n25481 );
buf ( n25483 , n25482 );
not ( n25484 , n25483 );
or ( n25485 , n25466 , n25484 );
not ( n25486 , n25482 );
buf ( n25487 , n25486 );
not ( n25488 , n25487 );
buf ( n25489 , n25461 );
not ( n25490 , n25489 );
or ( n25491 , n25488 , n25490 );
buf ( n25492 , n23638 );
not ( n25493 , n25492 );
buf ( n25494 , n18974 );
not ( n25495 , n25494 );
or ( n25496 , n25493 , n25495 );
buf ( n25497 , n20555 );
buf ( n25498 , n25304 );
nand ( n25499 , n25497 , n25498 );
buf ( n25500 , n25499 );
buf ( n25501 , n25500 );
nand ( n25502 , n25496 , n25501 );
buf ( n25503 , n25502 );
buf ( n25504 , n25503 );
nand ( n25505 , n25491 , n25504 );
buf ( n25506 , n25505 );
buf ( n25507 , n25506 );
nand ( n25508 , n25485 , n25507 );
buf ( n25509 , n25508 );
buf ( n25510 , n25509 );
xor ( n25511 , n25453 , n25510 );
not ( n25512 , n20363 );
not ( n25513 , n888 );
or ( n25514 , n25512 , n25513 );
nand ( n25515 , n23848 , n22303 );
nand ( n25516 , n25514 , n25515 );
buf ( n25517 , n25516 );
not ( n25518 , n25517 );
buf ( n25519 , n25518 );
buf ( n25520 , n25519 );
not ( n25521 , n25520 );
buf ( n25522 , n23881 );
not ( n25523 , n25522 );
buf ( n25524 , n18931 );
not ( n25525 , n25524 );
or ( n25526 , n25523 , n25525 );
buf ( n25527 , n21249 );
buf ( n25528 , n853 );
buf ( n25529 , n866 );
xor ( n25530 , n25528 , n25529 );
buf ( n25531 , n25530 );
buf ( n25532 , n25531 );
nand ( n25533 , n25527 , n25532 );
buf ( n25534 , n25533 );
buf ( n25535 , n25534 );
nand ( n25536 , n25526 , n25535 );
buf ( n25537 , n25536 );
buf ( n25538 , n25537 );
not ( n25539 , n25538 );
buf ( n25540 , n25539 );
buf ( n25541 , n25540 );
not ( n25542 , n25541 );
or ( n25543 , n25521 , n25542 );
buf ( n25544 , n23827 );
not ( n25545 , n25544 );
buf ( n25546 , n19479 );
not ( n25547 , n25546 );
or ( n25548 , n25545 , n25547 );
buf ( n25549 , n19265 );
buf ( n25550 , n841 );
buf ( n25551 , n878 );
xor ( n25552 , n25550 , n25551 );
buf ( n25553 , n25552 );
buf ( n25554 , n25553 );
nand ( n25555 , n25549 , n25554 );
buf ( n25556 , n25555 );
buf ( n25557 , n25556 );
nand ( n25558 , n25548 , n25557 );
buf ( n25559 , n25558 );
buf ( n25560 , n25559 );
nand ( n25561 , n25543 , n25560 );
buf ( n25562 , n25561 );
buf ( n25563 , n25562 );
buf ( n25564 , n25516 );
buf ( n25565 , n25537 );
nand ( n25566 , n25564 , n25565 );
buf ( n25567 , n25566 );
buf ( n25568 , n25567 );
nand ( n25569 , n25563 , n25568 );
buf ( n25570 , n25569 );
buf ( n25571 , n25570 );
and ( n25572 , n25511 , n25571 );
and ( n25573 , n25453 , n25510 );
or ( n25574 , n25572 , n25573 );
buf ( n25575 , n25574 );
buf ( n25576 , n25575 );
xor ( n25577 , n25402 , n25576 );
xor ( n25578 , n25199 , n25277 );
xor ( n25579 , n25578 , n25345 );
buf ( n25580 , n25579 );
buf ( n25581 , n25580 );
and ( n25582 , n25577 , n25581 );
and ( n25583 , n25402 , n25576 );
or ( n25584 , n25582 , n25583 );
buf ( n25585 , n25584 );
xor ( n25586 , n25353 , n25585 );
buf ( n25587 , n25586 );
buf ( n25588 , n25553 );
not ( n25589 , n25588 );
buf ( n25590 , n19259 );
not ( n25591 , n25590 );
or ( n25592 , n25589 , n25591 );
buf ( n25593 , n19265 );
buf ( n25594 , n25165 );
nand ( n25595 , n25593 , n25594 );
buf ( n25596 , n25595 );
buf ( n25597 , n25596 );
nand ( n25598 , n25592 , n25597 );
buf ( n25599 , n25598 );
buf ( n25600 , n25599 );
not ( n25601 , n25600 );
buf ( n25602 , n25531 );
not ( n25603 , n25602 );
buf ( n25604 , n18931 );
not ( n25605 , n25604 );
or ( n25606 , n25603 , n25605 );
buf ( n25607 , n21249 );
buf ( n25608 , n25143 );
nand ( n25609 , n25607 , n25608 );
buf ( n25610 , n25609 );
buf ( n25611 , n25610 );
nand ( n25612 , n25606 , n25611 );
buf ( n25613 , n25612 );
buf ( n25614 , n25613 );
not ( n25615 , n25614 );
buf ( n25616 , n25615 );
buf ( n25617 , n25616 );
not ( n25618 , n25617 );
or ( n25619 , n25601 , n25618 );
buf ( n25620 , n25599 );
not ( n25621 , n25620 );
buf ( n25622 , n25613 );
nand ( n25623 , n25621 , n25622 );
buf ( n25624 , n25623 );
buf ( n25625 , n25624 );
nand ( n25626 , n25619 , n25625 );
buf ( n25627 , n25626 );
buf ( n25628 , n25627 );
buf ( n25629 , n855 );
buf ( n25630 , n864 );
xor ( n25631 , n25629 , n25630 );
buf ( n25632 , n25631 );
buf ( n25633 , n25632 );
not ( n25634 , n25633 );
buf ( n25635 , n19013 );
not ( n25636 , n25635 );
or ( n25637 , n25634 , n25636 );
buf ( n25638 , n19030 );
buf ( n25639 , n854 );
buf ( n25640 , n864 );
xor ( n25641 , n25639 , n25640 );
buf ( n25642 , n25641 );
buf ( n25643 , n25642 );
nand ( n25644 , n25638 , n25643 );
buf ( n25645 , n25644 );
buf ( n25646 , n25645 );
nand ( n25647 , n25637 , n25646 );
buf ( n25648 , n25647 );
buf ( n25649 , n25648 );
not ( n25650 , n25649 );
buf ( n25651 , n25650 );
buf ( n25652 , n25651 );
and ( n25653 , n25628 , n25652 );
not ( n25654 , n25628 );
buf ( n25655 , n25648 );
and ( n25656 , n25654 , n25655 );
nor ( n25657 , n25653 , n25656 );
buf ( n25658 , n25657 );
buf ( n25659 , n25658 );
not ( n25660 , n25659 );
buf ( n25661 , n25660 );
not ( n25662 , n25661 );
xor ( n25663 , n25358 , n25379 );
xor ( n25664 , n25663 , n25397 );
buf ( n25665 , n25664 );
not ( n25666 , n25665 );
or ( n25667 , n25662 , n25666 );
buf ( n25668 , n25661 );
buf ( n25669 , n25665 );
or ( n25670 , n25668 , n25669 );
xor ( n25671 , n25237 , n25248 );
xnor ( n25672 , n25671 , n25270 );
buf ( n25673 , n25672 );
nand ( n25674 , n25670 , n25673 );
buf ( n25675 , n25674 );
nand ( n25676 , n25667 , n25675 );
buf ( n25677 , n25676 );
buf ( n25678 , n857 );
buf ( n25679 , n864 );
and ( n25680 , n25678 , n25679 );
buf ( n25681 , n25680 );
buf ( n25682 , n25681 );
buf ( n25683 , n23809 );
not ( n25684 , n25683 );
buf ( n25685 , n19013 );
not ( n25686 , n25685 );
or ( n25687 , n25684 , n25686 );
buf ( n25688 , n19030 );
buf ( n25689 , n25632 );
nand ( n25690 , n25688 , n25689 );
buf ( n25691 , n25690 );
buf ( n25692 , n25691 );
nand ( n25693 , n25687 , n25692 );
buf ( n25694 , n25693 );
buf ( n25695 , n25694 );
xor ( n25696 , n25682 , n25695 );
buf ( n25697 , n23865 );
not ( n25698 , n25697 );
buf ( n25699 , n25022 );
not ( n25700 , n25699 );
or ( n25701 , n25698 , n25700 );
buf ( n25702 , n25263 );
buf ( n25703 , n25255 );
nand ( n25704 , n25702 , n25703 );
buf ( n25705 , n25704 );
buf ( n25706 , n25705 );
nand ( n25707 , n25701 , n25706 );
buf ( n25708 , n25707 );
buf ( n25709 , n25708 );
and ( n25710 , n25696 , n25709 );
and ( n25711 , n25682 , n25695 );
or ( n25712 , n25710 , n25711 );
buf ( n25713 , n25712 );
buf ( n25714 , n25713 );
xor ( n25715 , n25300 , n25318 );
xor ( n25716 , n25715 , n25340 );
buf ( n25717 , n25716 );
buf ( n25718 , n25717 );
xor ( n25719 , n25714 , n25718 );
not ( n25720 , n20358 );
not ( n25721 , n25720 );
buf ( n25722 , n20363 );
not ( n25723 , n25722 );
buf ( n25724 , n25723 );
not ( n25725 , n25724 );
or ( n25726 , n25721 , n25725 );
nand ( n25727 , n25726 , n888 );
buf ( n25728 , n25727 );
buf ( n25729 , n25390 );
not ( n25730 , n25729 );
buf ( n25731 , n20521 );
not ( n25732 , n25731 );
or ( n25733 , n25730 , n25732 );
buf ( n25734 , n20525 );
buf ( n25735 , n832 );
buf ( n25736 , n886 );
xor ( n25737 , n25735 , n25736 );
buf ( n25738 , n25737 );
buf ( n25739 , n25738 );
nand ( n25740 , n25734 , n25739 );
buf ( n25741 , n25740 );
buf ( n25742 , n25741 );
nand ( n25743 , n25733 , n25742 );
buf ( n25744 , n25743 );
buf ( n25745 , n25744 );
xor ( n25746 , n25728 , n25745 );
buf ( n25747 , n25475 );
not ( n25748 , n25747 );
buf ( n25749 , n19580 );
not ( n25750 , n25749 );
or ( n25751 , n25748 , n25750 );
buf ( n25752 , n19910 );
buf ( n25753 , n836 );
buf ( n25754 , n882 );
xor ( n25755 , n25753 , n25754 );
buf ( n25756 , n25755 );
buf ( n25757 , n25756 );
nand ( n25758 , n25752 , n25757 );
buf ( n25759 , n25758 );
buf ( n25760 , n25759 );
nand ( n25761 , n25751 , n25760 );
buf ( n25762 , n25761 );
buf ( n25763 , n25762 );
xor ( n25764 , n25746 , n25763 );
buf ( n25765 , n25764 );
buf ( n25766 , n25765 );
and ( n25767 , n25719 , n25766 );
and ( n25768 , n25714 , n25718 );
or ( n25769 , n25767 , n25768 );
buf ( n25770 , n25769 );
buf ( n25771 , n25770 );
xor ( n25772 , n25677 , n25771 );
buf ( n25773 , n25616 );
not ( n25774 , n25773 );
buf ( n25775 , n25651 );
not ( n25776 , n25775 );
or ( n25777 , n25774 , n25776 );
buf ( n25778 , n25599 );
nand ( n25779 , n25777 , n25778 );
buf ( n25780 , n25779 );
buf ( n25781 , n25780 );
buf ( n25782 , n25648 );
buf ( n25783 , n25613 );
nand ( n25784 , n25782 , n25783 );
buf ( n25785 , n25784 );
buf ( n25786 , n25785 );
nand ( n25787 , n25781 , n25786 );
buf ( n25788 , n25787 );
buf ( n25789 , n25788 );
buf ( n25790 , n855 );
buf ( n25791 , n864 );
and ( n25792 , n25790 , n25791 );
buf ( n25793 , n25792 );
buf ( n25794 , n25793 );
buf ( n25795 , n25311 );
not ( n25796 , n25795 );
buf ( n25797 , n20549 );
not ( n25798 , n25797 );
or ( n25799 , n25796 , n25798 );
buf ( n25800 , n21513 );
buf ( n25801 , n25087 );
nand ( n25802 , n25800 , n25801 );
buf ( n25803 , n25802 );
buf ( n25804 , n25803 );
nand ( n25805 , n25799 , n25804 );
buf ( n25806 , n25805 );
buf ( n25807 , n25806 );
xor ( n25808 , n25794 , n25807 );
buf ( n25809 , n25756 );
not ( n25810 , n25809 );
buf ( n25811 , n19580 );
not ( n25812 , n25811 );
or ( n25813 , n25810 , n25812 );
buf ( n25814 , n19910 );
buf ( n25815 , n24900 );
nand ( n25816 , n25814 , n25815 );
buf ( n25817 , n25816 );
buf ( n25818 , n25817 );
nand ( n25819 , n25813 , n25818 );
buf ( n25820 , n25819 );
buf ( n25821 , n25820 );
xor ( n25822 , n25808 , n25821 );
buf ( n25823 , n25822 );
buf ( n25824 , n25823 );
xor ( n25825 , n25789 , n25824 );
xor ( n25826 , n25728 , n25745 );
and ( n25827 , n25826 , n25763 );
and ( n25828 , n25728 , n25745 );
or ( n25829 , n25827 , n25828 );
buf ( n25830 , n25829 );
buf ( n25831 , n25830 );
xor ( n25832 , n25825 , n25831 );
buf ( n25833 , n25832 );
buf ( n25834 , n25833 );
xor ( n25835 , n25772 , n25834 );
buf ( n25836 , n25835 );
buf ( n25837 , n25836 );
xor ( n25838 , n25714 , n25718 );
xor ( n25839 , n25838 , n25766 );
buf ( n25840 , n25839 );
buf ( n25841 , n25840 );
xor ( n25842 , n23799 , n23816 );
and ( n25843 , n25842 , n23834 );
and ( n25844 , n23799 , n23816 );
or ( n25845 , n25843 , n25844 );
buf ( n25846 , n25845 );
buf ( n25847 , n25846 );
xor ( n25848 , n25682 , n25695 );
xor ( n25849 , n25848 , n25709 );
buf ( n25850 , n25849 );
buf ( n25851 , n25850 );
xor ( n25852 , n25847 , n25851 );
and ( n25853 , n25503 , n25486 );
not ( n25854 , n25503 );
and ( n25855 , n25854 , n25482 );
or ( n25856 , n25853 , n25855 );
and ( n25857 , n25856 , n25464 );
not ( n25858 , n25856 );
and ( n25859 , n25858 , n25461 );
nor ( n25860 , n25857 , n25859 );
buf ( n25861 , n25860 );
and ( n25862 , n25852 , n25861 );
and ( n25863 , n25847 , n25851 );
or ( n25864 , n25862 , n25863 );
buf ( n25865 , n25864 );
buf ( n25866 , n25865 );
xor ( n25867 , n25841 , n25866 );
xor ( n25868 , n25658 , n25672 );
not ( n25869 , n25665 );
xor ( n25870 , n25868 , n25869 );
buf ( n25871 , n25870 );
and ( n25872 , n25867 , n25871 );
and ( n25873 , n25841 , n25866 );
or ( n25874 , n25872 , n25873 );
buf ( n25875 , n25874 );
buf ( n25876 , n25875 );
xor ( n25877 , n25837 , n25876 );
xnor ( n25878 , n25427 , n25414 );
buf ( n25879 , n25878 );
buf ( n25880 , n25441 );
buf ( n25881 , n25880 );
buf ( n25882 , n25881 );
buf ( n25883 , n25882 );
not ( n25884 , n25883 );
buf ( n25885 , n25884 );
buf ( n25886 , n25885 );
and ( n25887 , n25879 , n25886 );
not ( n25888 , n25879 );
buf ( n25889 , n25882 );
and ( n25890 , n25888 , n25889 );
nor ( n25891 , n25887 , n25890 );
buf ( n25892 , n25891 );
buf ( n25893 , n25892 );
xnor ( n25894 , n25540 , n25516 );
xor ( n25895 , n25559 , n25894 );
buf ( n25896 , n25895 );
xor ( n25897 , n25893 , n25896 );
buf ( n25898 , n23670 );
not ( n25899 , n25898 );
buf ( n25900 , n19153 );
not ( n25901 , n25900 );
or ( n25902 , n25899 , n25901 );
buf ( n25903 , n19082 );
buf ( n25904 , n25362 );
nand ( n25905 , n25903 , n25904 );
buf ( n25906 , n25905 );
buf ( n25907 , n25906 );
nand ( n25908 , n25902 , n25907 );
buf ( n25909 , n25908 );
buf ( n25910 , n25909 );
buf ( n25911 , n25396 );
not ( n25912 , n25911 );
buf ( n25913 , n25912 );
buf ( n25914 , n25913 );
xor ( n25915 , n25910 , n25914 );
buf ( n25916 , n23887 );
buf ( n25917 , n23907 );
or ( n25918 , n25916 , n25917 );
buf ( n25919 , n23928 );
nand ( n25920 , n25918 , n25919 );
buf ( n25921 , n25920 );
buf ( n25922 , n25921 );
buf ( n25923 , n23887 );
buf ( n25924 , n23907 );
nand ( n25925 , n25923 , n25924 );
buf ( n25926 , n25925 );
buf ( n25927 , n25926 );
nand ( n25928 , n25922 , n25927 );
buf ( n25929 , n25928 );
buf ( n25930 , n25929 );
xor ( n25931 , n25915 , n25930 );
buf ( n25932 , n25931 );
buf ( n25933 , n25932 );
and ( n25934 , n25897 , n25933 );
and ( n25935 , n25893 , n25896 );
or ( n25936 , n25934 , n25935 );
buf ( n25937 , n25936 );
buf ( n25938 , n25937 );
xor ( n25939 , n23483 , n23498 );
and ( n25940 , n25939 , n23542 );
and ( n25941 , n23483 , n23498 );
or ( n25942 , n25940 , n25941 );
buf ( n25943 , n25942 );
buf ( n25944 , n25943 );
not ( n25945 , n23580 );
not ( n25946 , n23622 );
or ( n25947 , n25945 , n25946 );
not ( n25948 , n23626 );
not ( n25949 , n23623 );
or ( n25950 , n25948 , n25949 );
nand ( n25951 , n25950 , n23677 );
nand ( n25952 , n25947 , n25951 );
buf ( n25953 , n25952 );
xor ( n25954 , n25944 , n25953 );
not ( n25955 , n23842 );
not ( n25956 , n23852 );
or ( n25957 , n25955 , n25956 );
not ( n25958 , n23841 );
and ( n25959 , n23843 , n23851 , n890 );
not ( n25960 , n25959 );
or ( n25961 , n25958 , n25960 );
nand ( n25962 , n25961 , n23869 );
nand ( n25963 , n25957 , n25962 );
buf ( n25964 , n25963 );
or ( n25965 , n23989 , n23972 );
nand ( n25966 , n25965 , n23956 );
buf ( n25967 , n23989 );
buf ( n25968 , n23972 );
nand ( n25969 , n25967 , n25968 );
buf ( n25970 , n25969 );
nand ( n25971 , n25966 , n25970 );
buf ( n25972 , n25971 );
xor ( n25973 , n25964 , n25972 );
not ( n25974 , n23644 );
nand ( n25975 , n25974 , n23661 );
nand ( n25976 , n23675 , n25975 );
not ( n25977 , n23661 );
nand ( n25978 , n25977 , n23644 );
nand ( n25979 , n25976 , n25978 );
buf ( n25980 , n25979 );
xor ( n25981 , n25973 , n25980 );
buf ( n25982 , n25981 );
buf ( n25983 , n25982 );
and ( n25984 , n25954 , n25983 );
and ( n25985 , n25944 , n25953 );
or ( n25986 , n25984 , n25985 );
buf ( n25987 , n25986 );
buf ( n25988 , n25987 );
xor ( n25989 , n25938 , n25988 );
xor ( n25990 , n25910 , n25914 );
and ( n25991 , n25990 , n25930 );
and ( n25992 , n25910 , n25914 );
or ( n25993 , n25991 , n25992 );
buf ( n25994 , n25993 );
buf ( n25995 , n25994 );
xor ( n25996 , n25964 , n25972 );
and ( n25997 , n25996 , n25980 );
and ( n25998 , n25964 , n25972 );
or ( n25999 , n25997 , n25998 );
buf ( n26000 , n25999 );
buf ( n26001 , n26000 );
xor ( n26002 , n25995 , n26001 );
xor ( n26003 , n25453 , n25510 );
xor ( n26004 , n26003 , n25571 );
buf ( n26005 , n26004 );
buf ( n26006 , n26005 );
xor ( n26007 , n26002 , n26006 );
buf ( n26008 , n26007 );
buf ( n26009 , n26008 );
and ( n26010 , n25989 , n26009 );
and ( n26011 , n25938 , n25988 );
or ( n26012 , n26010 , n26011 );
buf ( n26013 , n26012 );
buf ( n26014 , n26013 );
and ( n26015 , n25877 , n26014 );
and ( n26016 , n25837 , n25876 );
or ( n26017 , n26015 , n26016 );
buf ( n26018 , n26017 );
buf ( n26019 , n26018 );
xor ( n26020 , n25587 , n26019 );
xor ( n26021 , n25677 , n25771 );
and ( n26022 , n26021 , n25834 );
and ( n26023 , n25677 , n25771 );
or ( n26024 , n26022 , n26023 );
buf ( n26025 , n26024 );
buf ( n26026 , n26025 );
xor ( n26027 , n25789 , n25824 );
and ( n26028 , n26027 , n25831 );
and ( n26029 , n25789 , n25824 );
or ( n26030 , n26028 , n26029 );
buf ( n26031 , n26030 );
buf ( n26032 , n26031 );
buf ( n26033 , n25372 );
not ( n26034 , n26033 );
buf ( n26035 , n19153 );
not ( n26036 , n26035 );
or ( n26037 , n26034 , n26036 );
buf ( n26038 , n20246 );
buf ( n26039 , n25066 );
nand ( n26040 , n26038 , n26039 );
buf ( n26041 , n26040 );
buf ( n26042 , n26041 );
nand ( n26043 , n26037 , n26042 );
buf ( n26044 , n26043 );
buf ( n26045 , n25642 );
not ( n26046 , n26045 );
buf ( n26047 , n20302 );
not ( n26048 , n26047 );
or ( n26049 , n26046 , n26048 );
buf ( n26050 , n19027 );
buf ( n26051 , n25044 );
nand ( n26052 , n26050 , n26051 );
buf ( n26053 , n26052 );
buf ( n26054 , n26053 );
nand ( n26055 , n26049 , n26054 );
buf ( n26056 , n26055 );
or ( n26057 , n26044 , n26056 );
buf ( n26058 , n25738 );
not ( n26059 , n26058 );
buf ( n26060 , n20521 );
not ( n26061 , n26060 );
or ( n26062 , n26059 , n26061 );
buf ( n26063 , n20525 );
buf ( n26064 , n886 );
nand ( n26065 , n26063 , n26064 );
buf ( n26066 , n26065 );
buf ( n26067 , n26066 );
nand ( n26068 , n26062 , n26067 );
buf ( n26069 , n26068 );
nand ( n26070 , n26057 , n26069 );
buf ( n26071 , n25372 );
not ( n26072 , n26071 );
buf ( n26073 , n19077 );
not ( n26074 , n26073 );
or ( n26075 , n26072 , n26074 );
buf ( n26076 , n26041 );
nand ( n26077 , n26075 , n26076 );
buf ( n26078 , n26077 );
buf ( n26079 , n26078 );
buf ( n26080 , n26056 );
nand ( n26081 , n26079 , n26080 );
buf ( n26082 , n26081 );
nand ( n26083 , n26070 , n26082 );
buf ( n26084 , n26083 );
xor ( n26085 , n25794 , n25807 );
and ( n26086 , n26085 , n25821 );
and ( n26087 , n25794 , n25807 );
or ( n26088 , n26086 , n26087 );
buf ( n26089 , n26088 );
buf ( n26090 , n26089 );
xor ( n26091 , n26084 , n26090 );
buf ( n26092 , n25333 );
not ( n26093 , n26092 );
buf ( n26094 , n19614 );
not ( n26095 , n26094 );
or ( n26096 , n26093 , n26095 );
buf ( n26097 , n18860 );
buf ( n26098 , n25001 );
nand ( n26099 , n26097 , n26098 );
buf ( n26100 , n26099 );
buf ( n26101 , n26100 );
nand ( n26102 , n26096 , n26101 );
buf ( n26103 , n26102 );
buf ( n26104 , n25293 );
not ( n26105 , n26104 );
buf ( n26106 , n19230 );
not ( n26107 , n26106 );
or ( n26108 , n26105 , n26107 );
buf ( n26109 , n19235 );
buf ( n26110 , n24946 );
nand ( n26111 , n26109 , n26110 );
buf ( n26112 , n26111 );
buf ( n26113 , n26112 );
nand ( n26114 , n26108 , n26113 );
buf ( n26115 , n26114 );
xor ( n26116 , n26103 , n26115 );
buf ( n26117 , n25231 );
not ( n26118 , n26117 );
buf ( n26119 , n19125 );
not ( n26120 , n26119 );
or ( n26121 , n26118 , n26120 );
buf ( n26122 , n19134 );
buf ( n26123 , n24925 );
nand ( n26124 , n26122 , n26123 );
buf ( n26125 , n26124 );
buf ( n26126 , n26125 );
nand ( n26127 , n26121 , n26126 );
buf ( n26128 , n26127 );
and ( n26129 , n26116 , n26128 );
and ( n26130 , n26103 , n26115 );
or ( n26131 , n26129 , n26130 );
buf ( n26132 , n26131 );
xor ( n26133 , n26091 , n26132 );
buf ( n26134 , n26133 );
buf ( n26135 , n26134 );
xor ( n26136 , n26032 , n26135 );
xor ( n26137 , n26069 , n26078 );
buf ( n26138 , n26137 );
buf ( n26139 , n26056 );
xor ( n26140 , n26138 , n26139 );
buf ( n26141 , n26140 );
buf ( n26142 , n26141 );
xor ( n26143 , n25155 , n25138 );
and ( n26144 , n26143 , n25177 );
not ( n26145 , n26143 );
and ( n26146 , n26145 , n25180 );
nor ( n26147 , n26144 , n26146 );
buf ( n26148 , n26147 );
xor ( n26149 , n26142 , n26148 );
xor ( n26150 , n26103 , n26115 );
xor ( n26151 , n26150 , n26128 );
buf ( n26152 , n26151 );
and ( n26153 , n26149 , n26152 );
and ( n26154 , n26142 , n26148 );
or ( n26155 , n26153 , n26154 );
buf ( n26156 , n26155 );
buf ( n26157 , n26156 );
xor ( n26158 , n26136 , n26157 );
buf ( n26159 , n26158 );
buf ( n26160 , n26159 );
xor ( n26161 , n26026 , n26160 );
xor ( n26162 , n26142 , n26148 );
xor ( n26163 , n26162 , n26152 );
buf ( n26164 , n26163 );
xor ( n26165 , n25402 , n25576 );
xor ( n26166 , n26165 , n25581 );
buf ( n26167 , n26166 );
nand ( n26168 , n26164 , n26167 );
xor ( n26169 , n25995 , n26001 );
and ( n26170 , n26169 , n26006 );
and ( n26171 , n25995 , n26001 );
or ( n26172 , n26170 , n26171 );
buf ( n26173 , n26172 );
nand ( n26174 , n26164 , n26173 );
nand ( n26175 , n26167 , n26173 );
nand ( n26176 , n26168 , n26174 , n26175 );
buf ( n26177 , n26176 );
xor ( n26178 , n26161 , n26177 );
buf ( n26179 , n26178 );
buf ( n26180 , n26179 );
xor ( n26181 , n26020 , n26180 );
buf ( n26182 , n26181 );
buf ( n26183 , n26182 );
xor ( n26184 , n19455 , n19473 );
and ( n26185 , n26184 , n19493 );
and ( n26186 , n19455 , n19473 );
or ( n26187 , n26185 , n26186 );
buf ( n26188 , n26187 );
buf ( n26189 , n26188 );
xor ( n26190 , n19299 , n19347 );
and ( n26191 , n26190 , n19395 );
and ( n26192 , n19299 , n19347 );
or ( n26193 , n26191 , n26192 );
buf ( n26194 , n26193 );
buf ( n26195 , n26194 );
xor ( n26196 , n26189 , n26195 );
buf ( n26197 , n19489 );
xor ( n26198 , n19406 , n19420 );
and ( n26199 , n26198 , n19435 );
and ( n26200 , n19406 , n19420 );
or ( n26201 , n26199 , n26200 );
buf ( n26202 , n26201 );
buf ( n26203 , n26202 );
xor ( n26204 , n26197 , n26203 );
xor ( n26205 , n19511 , n19525 );
and ( n26206 , n26205 , n19540 );
and ( n26207 , n19511 , n19525 );
or ( n26208 , n26206 , n26207 );
buf ( n26209 , n26208 );
buf ( n26210 , n26209 );
xor ( n26211 , n26204 , n26210 );
buf ( n26212 , n26211 );
buf ( n26213 , n26212 );
xor ( n26214 , n26196 , n26213 );
buf ( n26215 , n26214 );
buf ( n26216 , n26215 );
xor ( n26217 , n19438 , n19496 );
and ( n26218 , n26217 , n19543 );
and ( n26219 , n19438 , n19496 );
or ( n26220 , n26218 , n26219 );
buf ( n26221 , n26220 );
buf ( n26222 , n26221 );
buf ( n26223 , n846 );
buf ( n26224 , n864 );
and ( n26225 , n26223 , n26224 );
buf ( n26226 , n26225 );
buf ( n26227 , n26226 );
buf ( n26228 , n19413 );
not ( n26229 , n26228 );
buf ( n26230 , n19330 );
not ( n26231 , n26230 );
or ( n26232 , n26229 , n26231 );
buf ( n26233 , n19030 );
buf ( n26234 , n864 );
buf ( n26235 , n844 );
xor ( n26236 , n26234 , n26235 );
buf ( n26237 , n26236 );
buf ( n26238 , n26237 );
nand ( n26239 , n26233 , n26238 );
buf ( n26240 , n26239 );
buf ( n26241 , n26240 );
nand ( n26242 , n26232 , n26241 );
buf ( n26243 , n26242 );
buf ( n26244 , n26243 );
xor ( n26245 , n26227 , n26244 );
buf ( n26246 , n19504 );
not ( n26247 , n26246 );
buf ( n26248 , n19125 );
not ( n26249 , n26248 );
or ( n26250 , n26247 , n26249 );
buf ( n26251 , n19134 );
buf ( n26252 , n838 );
buf ( n26253 , n870 );
xor ( n26254 , n26252 , n26253 );
buf ( n26255 , n26254 );
buf ( n26256 , n26255 );
nand ( n26257 , n26251 , n26256 );
buf ( n26258 , n26257 );
buf ( n26259 , n26258 );
nand ( n26260 , n26250 , n26259 );
buf ( n26261 , n26260 );
buf ( n26262 , n26261 );
xor ( n26263 , n26245 , n26262 );
buf ( n26264 , n26263 );
buf ( n26265 , n26264 );
buf ( n26266 , n19448 );
not ( n26267 , n26266 );
buf ( n26268 , n18931 );
not ( n26269 , n26268 );
or ( n26270 , n26267 , n26269 );
buf ( n26271 , n18944 );
buf ( n26272 , n842 );
buf ( n26273 , n866 );
xor ( n26274 , n26272 , n26273 );
buf ( n26275 , n26274 );
buf ( n26276 , n26275 );
nand ( n26277 , n26271 , n26276 );
buf ( n26278 , n26277 );
buf ( n26279 , n26278 );
nand ( n26280 , n26270 , n26279 );
buf ( n26281 , n26280 );
buf ( n26282 , n26281 );
buf ( n26283 , n19518 );
not ( n26284 , n26283 );
buf ( n26285 , n18977 );
not ( n26286 , n26285 );
or ( n26287 , n26284 , n26286 );
buf ( n26288 , n18987 );
buf ( n26289 , n834 );
buf ( n26290 , n874 );
xor ( n26291 , n26289 , n26290 );
buf ( n26292 , n26291 );
buf ( n26293 , n26292 );
nand ( n26294 , n26288 , n26293 );
buf ( n26295 , n26294 );
buf ( n26296 , n26295 );
nand ( n26297 , n26287 , n26296 );
buf ( n26298 , n26297 );
buf ( n26299 , n26298 );
xor ( n26300 , n26282 , n26299 );
buf ( n26301 , n19466 );
not ( n26302 , n26301 );
buf ( n26303 , n18887 );
not ( n26304 , n26303 );
or ( n26305 , n26302 , n26304 );
buf ( n26306 , n18898 );
buf ( n26307 , n840 );
buf ( n26308 , n868 );
xor ( n26309 , n26307 , n26308 );
buf ( n26310 , n26309 );
buf ( n26311 , n26310 );
nand ( n26312 , n26306 , n26311 );
buf ( n26313 , n26312 );
buf ( n26314 , n26313 );
nand ( n26315 , n26305 , n26314 );
buf ( n26316 , n26315 );
buf ( n26317 , n26316 );
xor ( n26318 , n26300 , n26317 );
buf ( n26319 , n26318 );
buf ( n26320 , n26319 );
xor ( n26321 , n26265 , n26320 );
buf ( n26322 , n19428 );
not ( n26323 , n26322 );
buf ( n26324 , n19230 );
not ( n26325 , n26324 );
or ( n26326 , n26323 , n26325 );
buf ( n26327 , n19235 );
xor ( n26328 , n872 , n836 );
buf ( n26329 , n26328 );
nand ( n26330 , n26327 , n26329 );
buf ( n26331 , n26330 );
buf ( n26332 , n26331 );
nand ( n26333 , n26326 , n26332 );
buf ( n26334 , n26333 );
buf ( n26335 , n19533 );
not ( n26336 , n26335 );
buf ( n26337 , n19153 );
not ( n26338 , n26337 );
or ( n26339 , n26336 , n26338 );
buf ( n26340 , n19085 );
xor ( n26341 , n876 , n832 );
buf ( n26342 , n26341 );
nand ( n26343 , n26340 , n26342 );
buf ( n26344 , n26343 );
buf ( n26345 , n26344 );
nand ( n26346 , n26339 , n26345 );
buf ( n26347 , n26346 );
xor ( n26348 , n26334 , n26347 );
buf ( n26349 , n19479 );
buf ( n26350 , n19265 );
or ( n26351 , n26349 , n26350 );
buf ( n26352 , n878 );
nand ( n26353 , n26351 , n26352 );
buf ( n26354 , n26353 );
xor ( n26355 , n26348 , n26354 );
buf ( n26356 , n26355 );
xor ( n26357 , n26321 , n26356 );
buf ( n26358 , n26357 );
buf ( n26359 , n26358 );
xor ( n26360 , n26222 , n26359 );
xor ( n26361 , n19056 , n19283 );
and ( n26362 , n26361 , n19398 );
and ( n26363 , n19056 , n19283 );
or ( n26364 , n26362 , n26363 );
buf ( n26365 , n26364 );
buf ( n26366 , n26365 );
xor ( n26367 , n26360 , n26366 );
buf ( n26368 , n26367 );
buf ( n26369 , n26368 );
xor ( n26370 , n26216 , n26369 );
xor ( n26371 , n19546 , n19564 );
and ( n26372 , n26371 , n19777 );
and ( n26373 , n19546 , n19564 );
or ( n26374 , n26372 , n26373 );
buf ( n26375 , n26374 );
buf ( n26376 , n26375 );
xor ( n26377 , n26370 , n26376 );
buf ( n26378 , n26377 );
buf ( n26379 , n26378 );
xor ( n26380 , n25587 , n26019 );
and ( n26381 , n26380 , n26180 );
and ( n26382 , n25587 , n26019 );
or ( n26383 , n26381 , n26382 );
buf ( n26384 , n26383 );
buf ( n26385 , n26384 );
buf ( n26386 , n856 );
buf ( n26387 , n886 );
xor ( n26388 , n26386 , n26387 );
buf ( n26389 , n26388 );
not ( n26390 , n26389 );
not ( n26391 , n20521 );
or ( n26392 , n26390 , n26391 );
buf ( n26393 , n855 );
buf ( n26394 , n886 );
xor ( n26395 , n26393 , n26394 );
buf ( n26396 , n26395 );
nand ( n26397 , n20525 , n26396 );
nand ( n26398 , n26392 , n26397 );
buf ( n26399 , n862 );
buf ( n26400 , n880 );
xor ( n26401 , n26399 , n26400 );
buf ( n26402 , n26401 );
buf ( n26403 , n26402 );
not ( n26404 , n26403 );
buf ( n26405 , n19614 );
not ( n26406 , n26405 );
or ( n26407 , n26404 , n26406 );
buf ( n26408 , n18860 );
buf ( n26409 , n861 );
buf ( n26410 , n880 );
xor ( n26411 , n26409 , n26410 );
buf ( n26412 , n26411 );
buf ( n26413 , n26412 );
nand ( n26414 , n26408 , n26413 );
buf ( n26415 , n26414 );
buf ( n26416 , n26415 );
nand ( n26417 , n26407 , n26416 );
buf ( n26418 , n26417 );
xor ( n26419 , n26398 , n26418 );
buf ( n26420 , n854 );
buf ( n26421 , n888 );
xor ( n26422 , n26420 , n26421 );
buf ( n26423 , n26422 );
buf ( n26424 , n26423 );
not ( n26425 , n26424 );
buf ( n26426 , n20358 );
not ( n26427 , n26426 );
or ( n26428 , n26425 , n26427 );
buf ( n26429 , n20363 );
buf ( n26430 , n853 );
buf ( n26431 , n888 );
xor ( n26432 , n26430 , n26431 );
buf ( n26433 , n26432 );
buf ( n26434 , n26433 );
nand ( n26435 , n26429 , n26434 );
buf ( n26436 , n26435 );
buf ( n26437 , n26436 );
nand ( n26438 , n26428 , n26437 );
buf ( n26439 , n26438 );
xor ( n26440 , n26419 , n26439 );
buf ( n26441 , n850 );
buf ( n26442 , n892 );
xor ( n26443 , n26441 , n26442 );
buf ( n26444 , n26443 );
buf ( n26445 , n26444 );
not ( n26446 , n26445 );
buf ( n26447 , n23175 );
not ( n26448 , n26447 );
or ( n26449 , n26446 , n26448 );
buf ( n26450 , n22818 );
buf ( n26451 , n849 );
buf ( n26452 , n892 );
xor ( n26453 , n26451 , n26452 );
buf ( n26454 , n26453 );
buf ( n26455 , n26454 );
nand ( n26456 , n26450 , n26455 );
buf ( n26457 , n26456 );
buf ( n26458 , n26457 );
nand ( n26459 , n26449 , n26458 );
buf ( n26460 , n26459 );
not ( n26461 , n21297 );
buf ( n26462 , n848 );
buf ( n26463 , n894 );
xor ( n26464 , n26462 , n26463 );
buf ( n26465 , n26464 );
not ( n26466 , n26465 );
or ( n26467 , n26461 , n26466 );
buf ( n26468 , n847 );
buf ( n26469 , n894 );
xor ( n26470 , n26468 , n26469 );
buf ( n26471 , n26470 );
buf ( n26472 , n26471 );
buf ( n26473 , n895 );
nand ( n26474 , n26472 , n26473 );
buf ( n26475 , n26474 );
nand ( n26476 , n26467 , n26475 );
not ( n26477 , n26476 );
nand ( n26478 , n863 , n19265 );
and ( n26479 , n26477 , n26478 );
not ( n26480 , n26477 );
nand ( n26481 , n19265 , n863 );
not ( n26482 , n26481 );
and ( n26483 , n26480 , n26482 );
nor ( n26484 , n26479 , n26483 );
xor ( n26485 , n26460 , n26484 );
buf ( n26486 , n26485 );
buf ( n26487 , n852 );
buf ( n26488 , n890 );
xor ( n26489 , n26487 , n26488 );
buf ( n26490 , n26489 );
buf ( n26491 , n26490 );
not ( n26492 , n26491 );
buf ( n26493 , n21441 );
not ( n26494 , n26493 );
or ( n26495 , n26492 , n26494 );
buf ( n26496 , n20869 );
buf ( n26497 , n851 );
buf ( n26498 , n890 );
xor ( n26499 , n26497 , n26498 );
buf ( n26500 , n26499 );
buf ( n26501 , n26500 );
nand ( n26502 , n26496 , n26501 );
buf ( n26503 , n26502 );
buf ( n26504 , n26503 );
nand ( n26505 , n26495 , n26504 );
buf ( n26506 , n26505 );
buf ( n26507 , n858 );
buf ( n26508 , n884 );
xor ( n26509 , n26507 , n26508 );
buf ( n26510 , n26509 );
buf ( n26511 , n26510 );
not ( n26512 , n26511 );
buf ( n26513 , n25022 );
not ( n26514 , n26513 );
or ( n26515 , n26512 , n26514 );
buf ( n26516 , n23233 );
buf ( n26517 , n857 );
buf ( n26518 , n884 );
xor ( n26519 , n26517 , n26518 );
buf ( n26520 , n26519 );
buf ( n26521 , n26520 );
nand ( n26522 , n26516 , n26521 );
buf ( n26523 , n26522 );
buf ( n26524 , n26523 );
nand ( n26525 , n26515 , n26524 );
buf ( n26526 , n26525 );
xor ( n26527 , n26506 , n26526 );
buf ( n26528 , n860 );
buf ( n26529 , n882 );
xor ( n26530 , n26528 , n26529 );
buf ( n26531 , n26530 );
buf ( n26532 , n26531 );
not ( n26533 , n26532 );
buf ( n26534 , n19580 );
buf ( n26535 , n26534 );
not ( n26536 , n26535 );
or ( n26537 , n26533 , n26536 );
not ( n26538 , n19569 );
buf ( n26539 , n26538 );
buf ( n26540 , n859 );
buf ( n26541 , n882 );
xor ( n26542 , n26540 , n26541 );
buf ( n26543 , n26542 );
buf ( n26544 , n26543 );
nand ( n26545 , n26539 , n26544 );
buf ( n26546 , n26545 );
buf ( n26547 , n26546 );
nand ( n26548 , n26537 , n26547 );
buf ( n26549 , n26548 );
xor ( n26550 , n26527 , n26549 );
nand ( n26551 , n26440 , n26486 , n26550 );
not ( n26552 , n26486 );
not ( n26553 , n26550 );
nand ( n26554 , n26552 , n26553 );
not ( n26555 , n26554 );
nand ( n26556 , n26555 , n26440 );
not ( n26557 , n26440 );
not ( n26558 , n26550 );
nor ( n26559 , n26558 , n26486 );
nand ( n26560 , n26557 , n26559 );
nand ( n26561 , n26557 , n26486 , n26553 );
nand ( n26562 , n26551 , n26556 , n26560 , n26561 );
buf ( n26563 , n26562 );
buf ( n26564 , n851 );
buf ( n26565 , n894 );
xor ( n26566 , n26564 , n26565 );
buf ( n26567 , n26566 );
buf ( n26568 , n26567 );
not ( n26569 , n26568 );
buf ( n26570 , n23288 );
not ( n26571 , n26570 );
or ( n26572 , n26569 , n26571 );
buf ( n26573 , n850 );
buf ( n26574 , n894 );
xor ( n26575 , n26573 , n26574 );
buf ( n26576 , n26575 );
buf ( n26577 , n26576 );
buf ( n26578 , n895 );
nand ( n26579 , n26577 , n26578 );
buf ( n26580 , n26579 );
buf ( n26581 , n26580 );
nand ( n26582 , n26572 , n26581 );
buf ( n26583 , n26582 );
buf ( n26584 , n26583 );
buf ( n26585 , n863 );
buf ( n26586 , n883 );
or ( n26587 , n26585 , n26586 );
buf ( n26588 , n884 );
nand ( n26589 , n26587 , n26588 );
buf ( n26590 , n26589 );
buf ( n26591 , n863 );
buf ( n26592 , n883 );
nand ( n26593 , n26591 , n26592 );
buf ( n26594 , n26593 );
and ( n26595 , n26590 , n26594 , n882 );
buf ( n26596 , n26595 );
and ( n26597 , n26584 , n26596 );
buf ( n26598 , n26597 );
buf ( n26599 , n26598 );
xor ( n26600 , n882 , n862 );
buf ( n26601 , n26600 );
not ( n26602 , n26601 );
buf ( n26603 , n19580 );
not ( n26604 , n26603 );
or ( n26605 , n26602 , n26604 );
buf ( n26606 , n19910 );
buf ( n26607 , n861 );
buf ( n26608 , n882 );
xor ( n26609 , n26607 , n26608 );
buf ( n26610 , n26609 );
buf ( n26611 , n26610 );
nand ( n26612 , n26606 , n26611 );
buf ( n26613 , n26612 );
buf ( n26614 , n26613 );
nand ( n26615 , n26605 , n26614 );
buf ( n26616 , n26615 );
buf ( n26617 , n26616 );
xor ( n26618 , n26599 , n26617 );
xor ( n26619 , n884 , n860 );
buf ( n26620 , n26619 );
not ( n26621 , n26620 );
buf ( n26622 , n25022 );
not ( n26623 , n26622 );
or ( n26624 , n26621 , n26623 );
buf ( n26625 , n25263 );
buf ( n26626 , n859 );
buf ( n26627 , n884 );
xor ( n26628 , n26626 , n26627 );
buf ( n26629 , n26628 );
buf ( n26630 , n26629 );
nand ( n26631 , n26625 , n26630 );
buf ( n26632 , n26631 );
buf ( n26633 , n26632 );
nand ( n26634 , n26624 , n26633 );
buf ( n26635 , n26634 );
buf ( n26636 , n26635 );
and ( n26637 , n26618 , n26636 );
and ( n26638 , n26599 , n26617 );
or ( n26639 , n26637 , n26638 );
buf ( n26640 , n26639 );
buf ( n26641 , n26640 );
buf ( n26642 , n26610 );
not ( n26643 , n26642 );
buf ( n26644 , n26534 );
not ( n26645 , n26644 );
or ( n26646 , n26643 , n26645 );
buf ( n26647 , n19910 );
buf ( n26648 , n26531 );
nand ( n26649 , n26647 , n26648 );
buf ( n26650 , n26649 );
buf ( n26651 , n26650 );
nand ( n26652 , n26646 , n26651 );
buf ( n26653 , n26652 );
buf ( n26654 , n26653 );
buf ( n26655 , n863 );
buf ( n26656 , n881 );
or ( n26657 , n26655 , n26656 );
buf ( n26658 , n882 );
nand ( n26659 , n26657 , n26658 );
buf ( n26660 , n26659 );
buf ( n26661 , n26660 );
buf ( n26662 , n863 );
buf ( n26663 , n881 );
nand ( n26664 , n26662 , n26663 );
buf ( n26665 , n26664 );
buf ( n26666 , n26665 );
buf ( n26667 , n880 );
and ( n26668 , n26661 , n26666 , n26667 );
buf ( n26669 , n26668 );
buf ( n26670 , n26669 );
buf ( n26671 , n849 );
buf ( n26672 , n894 );
xor ( n26673 , n26671 , n26672 );
buf ( n26674 , n26673 );
buf ( n26675 , n26674 );
not ( n26676 , n26675 );
buf ( n26677 , n21297 );
not ( n26678 , n26677 );
or ( n26679 , n26676 , n26678 );
buf ( n26680 , n26465 );
buf ( n26681 , n895 );
nand ( n26682 , n26680 , n26681 );
buf ( n26683 , n26682 );
buf ( n26684 , n26683 );
nand ( n26685 , n26679 , n26684 );
buf ( n26686 , n26685 );
buf ( n26687 , n26686 );
xor ( n26688 , n26670 , n26687 );
buf ( n26689 , n26688 );
buf ( n26690 , n26689 );
xor ( n26691 , n26654 , n26690 );
buf ( n26692 , n20325 );
buf ( n26693 , n863 );
and ( n26694 , n26692 , n26693 );
buf ( n26695 , n26694 );
buf ( n26696 , n26695 );
buf ( n26697 , n26576 );
not ( n26698 , n26697 );
buf ( n26699 , n21297 );
not ( n26700 , n26699 );
or ( n26701 , n26698 , n26700 );
buf ( n26702 , n26674 );
buf ( n26703 , n895 );
nand ( n26704 , n26702 , n26703 );
buf ( n26705 , n26704 );
buf ( n26706 , n26705 );
nand ( n26707 , n26701 , n26706 );
buf ( n26708 , n26707 );
buf ( n26709 , n26708 );
xor ( n26710 , n26696 , n26709 );
buf ( n26711 , n852 );
buf ( n26712 , n892 );
xor ( n26713 , n26711 , n26712 );
buf ( n26714 , n26713 );
buf ( n26715 , n26714 );
not ( n26716 , n26715 );
buf ( n26717 , n23175 );
not ( n26718 , n26717 );
or ( n26719 , n26716 , n26718 );
buf ( n26720 , n22818 );
buf ( n26721 , n851 );
buf ( n26722 , n892 );
xor ( n26723 , n26721 , n26722 );
buf ( n26724 , n26723 );
buf ( n26725 , n26724 );
nand ( n26726 , n26720 , n26725 );
buf ( n26727 , n26726 );
buf ( n26728 , n26727 );
nand ( n26729 , n26719 , n26728 );
buf ( n26730 , n26729 );
buf ( n26731 , n26730 );
and ( n26732 , n26710 , n26731 );
and ( n26733 , n26696 , n26709 );
or ( n26734 , n26732 , n26733 );
buf ( n26735 , n26734 );
buf ( n26736 , n26735 );
xor ( n26737 , n26691 , n26736 );
buf ( n26738 , n26737 );
buf ( n26739 , n26738 );
xor ( n26740 , n26641 , n26739 );
xor ( n26741 , n26696 , n26709 );
xor ( n26742 , n26741 , n26731 );
buf ( n26743 , n26742 );
buf ( n26744 , n26743 );
buf ( n26745 , n857 );
buf ( n26746 , n888 );
xor ( n26747 , n26745 , n26746 );
buf ( n26748 , n26747 );
buf ( n26749 , n26748 );
not ( n26750 , n26749 );
buf ( n26751 , n20358 );
not ( n26752 , n26751 );
or ( n26753 , n26750 , n26752 );
buf ( n26754 , n20363 );
buf ( n26755 , n856 );
buf ( n26756 , n888 );
xor ( n26757 , n26755 , n26756 );
buf ( n26758 , n26757 );
buf ( n26759 , n26758 );
nand ( n26760 , n26754 , n26759 );
buf ( n26761 , n26760 );
buf ( n26762 , n26761 );
nand ( n26763 , n26753 , n26762 );
buf ( n26764 , n26763 );
buf ( n26765 , n26764 );
not ( n26766 , n26765 );
buf ( n26767 , n859 );
buf ( n26768 , n886 );
xor ( n26769 , n26767 , n26768 );
buf ( n26770 , n26769 );
buf ( n26771 , n26770 );
not ( n26772 , n26771 );
buf ( n26773 , n20521 );
not ( n26774 , n26773 );
or ( n26775 , n26772 , n26774 );
buf ( n26776 , n20525 );
buf ( n26777 , n858 );
buf ( n26778 , n886 );
xor ( n26779 , n26777 , n26778 );
buf ( n26780 , n26779 );
buf ( n26781 , n26780 );
nand ( n26782 , n26776 , n26781 );
buf ( n26783 , n26782 );
buf ( n26784 , n26783 );
nand ( n26785 , n26775 , n26784 );
buf ( n26786 , n26785 );
buf ( n26787 , n26786 );
not ( n26788 , n26787 );
or ( n26789 , n26766 , n26788 );
buf ( n26790 , n26786 );
buf ( n26791 , n26764 );
or ( n26792 , n26790 , n26791 );
xor ( n26793 , n892 , n853 );
buf ( n26794 , n26793 );
not ( n26795 , n26794 );
buf ( n26796 , n23175 );
not ( n26797 , n26796 );
or ( n26798 , n26795 , n26797 );
buf ( n26799 , n23181 );
buf ( n26800 , n26714 );
nand ( n26801 , n26799 , n26800 );
buf ( n26802 , n26801 );
buf ( n26803 , n26802 );
nand ( n26804 , n26798 , n26803 );
buf ( n26805 , n26804 );
buf ( n26806 , n26805 );
nand ( n26807 , n26792 , n26806 );
buf ( n26808 , n26807 );
buf ( n26809 , n26808 );
nand ( n26810 , n26789 , n26809 );
buf ( n26811 , n26810 );
buf ( n26812 , n26811 );
xor ( n26813 , n26744 , n26812 );
xor ( n26814 , n882 , n863 );
buf ( n26815 , n26814 );
not ( n26816 , n26815 );
buf ( n26817 , n19580 );
not ( n26818 , n26817 );
or ( n26819 , n26816 , n26818 );
buf ( n26820 , n19910 );
buf ( n26821 , n26600 );
nand ( n26822 , n26820 , n26821 );
buf ( n26823 , n26822 );
buf ( n26824 , n26823 );
nand ( n26825 , n26819 , n26824 );
buf ( n26826 , n26825 );
buf ( n26827 , n26826 );
buf ( n26828 , n855 );
buf ( n26829 , n890 );
xor ( n26830 , n26828 , n26829 );
buf ( n26831 , n26830 );
buf ( n26832 , n26831 );
not ( n26833 , n26832 );
buf ( n26834 , n21441 );
not ( n26835 , n26834 );
or ( n26836 , n26833 , n26835 );
buf ( n26837 , n20869 );
xor ( n26838 , n890 , n854 );
buf ( n26839 , n26838 );
nand ( n26840 , n26837 , n26839 );
buf ( n26841 , n26840 );
buf ( n26842 , n26841 );
nand ( n26843 , n26836 , n26842 );
buf ( n26844 , n26843 );
buf ( n26845 , n26844 );
xor ( n26846 , n26827 , n26845 );
xor ( n26847 , n884 , n861 );
buf ( n26848 , n26847 );
not ( n26849 , n26848 );
buf ( n26850 , n25022 );
not ( n26851 , n26850 );
or ( n26852 , n26849 , n26851 );
buf ( n26853 , n25263 );
buf ( n26854 , n26619 );
nand ( n26855 , n26853 , n26854 );
buf ( n26856 , n26855 );
buf ( n26857 , n26856 );
nand ( n26858 , n26852 , n26857 );
buf ( n26859 , n26858 );
buf ( n26860 , n26859 );
and ( n26861 , n26846 , n26860 );
and ( n26862 , n26827 , n26845 );
or ( n26863 , n26861 , n26862 );
buf ( n26864 , n26863 );
buf ( n26865 , n26864 );
and ( n26866 , n26813 , n26865 );
and ( n26867 , n26744 , n26812 );
or ( n26868 , n26866 , n26867 );
buf ( n26869 , n26868 );
buf ( n26870 , n26869 );
and ( n26871 , n26740 , n26870 );
and ( n26872 , n26641 , n26739 );
or ( n26873 , n26871 , n26872 );
buf ( n26874 , n26873 );
buf ( n26875 , n26874 );
xor ( n26876 , n26563 , n26875 );
xor ( n26877 , n26654 , n26690 );
and ( n26878 , n26877 , n26736 );
and ( n26879 , n26654 , n26690 );
or ( n26880 , n26878 , n26879 );
buf ( n26881 , n26880 );
buf ( n26882 , n26881 );
and ( n26883 , n26670 , n26687 );
buf ( n26884 , n26883 );
buf ( n26885 , n26884 );
buf ( n26886 , n855 );
buf ( n26887 , n888 );
xor ( n26888 , n26886 , n26887 );
buf ( n26889 , n26888 );
buf ( n26890 , n26889 );
not ( n26891 , n26890 );
buf ( n26892 , n23144 );
not ( n26893 , n26892 );
or ( n26894 , n26891 , n26893 );
buf ( n26895 , n20363 );
buf ( n26896 , n26423 );
nand ( n26897 , n26895 , n26896 );
buf ( n26898 , n26897 );
buf ( n26899 , n26898 );
nand ( n26900 , n26894 , n26899 );
buf ( n26901 , n26900 );
not ( n26902 , n26724 );
not ( n26903 , n23175 );
or ( n26904 , n26902 , n26903 );
buf ( n26905 , n22818 );
buf ( n26906 , n26444 );
nand ( n26907 , n26905 , n26906 );
buf ( n26908 , n26907 );
nand ( n26909 , n26904 , n26908 );
or ( n26910 , n26901 , n26909 );
buf ( n26911 , n863 );
buf ( n26912 , n880 );
xor ( n26913 , n26911 , n26912 );
buf ( n26914 , n26913 );
buf ( n26915 , n26914 );
not ( n26916 , n26915 );
buf ( n26917 , n19614 );
not ( n26918 , n26917 );
or ( n26919 , n26916 , n26918 );
buf ( n26920 , n18860 );
buf ( n26921 , n26402 );
nand ( n26922 , n26920 , n26921 );
buf ( n26923 , n26922 );
buf ( n26924 , n26923 );
nand ( n26925 , n26919 , n26924 );
buf ( n26926 , n26925 );
nand ( n26927 , n26910 , n26926 );
buf ( n26928 , n26927 );
nand ( n26929 , n26909 , n26901 );
buf ( n26930 , n26929 );
nand ( n26931 , n26928 , n26930 );
buf ( n26932 , n26931 );
buf ( n26933 , n26932 );
xor ( n26934 , n26885 , n26933 );
buf ( n26935 , n857 );
buf ( n26936 , n886 );
xor ( n26937 , n26935 , n26936 );
buf ( n26938 , n26937 );
buf ( n26939 , n26938 );
not ( n26940 , n26939 );
buf ( n26941 , n23027 );
not ( n26942 , n26941 );
or ( n26943 , n26940 , n26942 );
buf ( n26944 , n20525 );
buf ( n26945 , n26389 );
nand ( n26946 , n26944 , n26945 );
buf ( n26947 , n26946 );
buf ( n26948 , n26947 );
nand ( n26949 , n26943 , n26948 );
buf ( n26950 , n26949 );
buf ( n26951 , n26950 );
xor ( n26952 , n890 , n853 );
buf ( n26953 , n26952 );
not ( n26954 , n26953 );
buf ( n26955 , n21441 );
not ( n26956 , n26955 );
or ( n26957 , n26954 , n26956 );
buf ( n26958 , n20869 );
buf ( n26959 , n26490 );
nand ( n26960 , n26958 , n26959 );
buf ( n26961 , n26960 );
buf ( n26962 , n26961 );
nand ( n26963 , n26957 , n26962 );
buf ( n26964 , n26963 );
buf ( n26965 , n26964 );
or ( n26966 , n26951 , n26965 );
buf ( n26967 , n26629 );
not ( n26968 , n26967 );
buf ( n26969 , n25022 );
not ( n26970 , n26969 );
or ( n26971 , n26968 , n26970 );
buf ( n26972 , n25263 );
buf ( n26973 , n26510 );
nand ( n26974 , n26972 , n26973 );
buf ( n26975 , n26974 );
buf ( n26976 , n26975 );
nand ( n26977 , n26971 , n26976 );
buf ( n26978 , n26977 );
buf ( n26979 , n26978 );
nand ( n26980 , n26966 , n26979 );
buf ( n26981 , n26980 );
buf ( n26982 , n26981 );
buf ( n26983 , n26950 );
buf ( n26984 , n26964 );
nand ( n26985 , n26983 , n26984 );
buf ( n26986 , n26985 );
buf ( n26987 , n26986 );
nand ( n26988 , n26982 , n26987 );
buf ( n26989 , n26988 );
buf ( n26990 , n26989 );
xor ( n26991 , n26934 , n26990 );
buf ( n26992 , n26991 );
buf ( n26993 , n26992 );
xor ( n26994 , n26882 , n26993 );
buf ( n26995 , n26838 );
not ( n26996 , n26995 );
buf ( n26997 , n21441 );
not ( n26998 , n26997 );
or ( n26999 , n26996 , n26998 );
buf ( n27000 , n20869 );
buf ( n27001 , n26952 );
nand ( n27002 , n27000 , n27001 );
buf ( n27003 , n27002 );
buf ( n27004 , n27003 );
nand ( n27005 , n26999 , n27004 );
buf ( n27006 , n27005 );
not ( n27007 , n27006 );
buf ( n27008 , n26758 );
not ( n27009 , n27008 );
buf ( n27010 , n23144 );
not ( n27011 , n27010 );
or ( n27012 , n27009 , n27011 );
buf ( n27013 , n20363 );
buf ( n27014 , n26889 );
nand ( n27015 , n27013 , n27014 );
buf ( n27016 , n27015 );
buf ( n27017 , n27016 );
nand ( n27018 , n27012 , n27017 );
buf ( n27019 , n27018 );
not ( n27020 , n27019 );
nand ( n27021 , n27007 , n27020 );
not ( n27022 , n27021 );
buf ( n27023 , n23320 );
buf ( n27024 , n26938 );
nand ( n27025 , n27023 , n27024 );
buf ( n27026 , n27025 );
nand ( n27027 , n20521 , n26780 );
nand ( n27028 , n27026 , n27027 );
not ( n27029 , n27028 );
or ( n27030 , n27022 , n27029 );
buf ( n27031 , n27006 );
buf ( n27032 , n27019 );
nand ( n27033 , n27031 , n27032 );
buf ( n27034 , n27033 );
nand ( n27035 , n27030 , n27034 );
buf ( n27036 , n27035 );
xor ( n27037 , n26901 , n26926 );
xor ( n27038 , n27037 , n26909 );
buf ( n27039 , n27038 );
xor ( n27040 , n27036 , n27039 );
xor ( n27041 , n26964 , n26950 );
xor ( n27042 , n27041 , n26978 );
buf ( n27043 , n27042 );
and ( n27044 , n27040 , n27043 );
and ( n27045 , n27036 , n27039 );
or ( n27046 , n27044 , n27045 );
buf ( n27047 , n27046 );
buf ( n27048 , n27047 );
xor ( n27049 , n26994 , n27048 );
buf ( n27050 , n27049 );
buf ( n27051 , n27050 );
xor ( n27052 , n26876 , n27051 );
buf ( n27053 , n27052 );
buf ( n27054 , n27053 );
xor ( n27055 , n27036 , n27039 );
xor ( n27056 , n27055 , n27043 );
buf ( n27057 , n27056 );
buf ( n27058 , n27057 );
xor ( n27059 , n26599 , n26617 );
xor ( n27060 , n27059 , n26636 );
buf ( n27061 , n27060 );
buf ( n27062 , n27061 );
xor ( n27063 , n27028 , n27007 );
not ( n27064 , n27020 );
xnor ( n27065 , n27063 , n27064 );
buf ( n27066 , n27065 );
xor ( n27067 , n27062 , n27066 );
buf ( n27068 , n26583 );
buf ( n27069 , n26595 );
xor ( n27070 , n27068 , n27069 );
buf ( n27071 , n27070 );
buf ( n27072 , n27071 );
buf ( n27073 , n26538 );
buf ( n27074 , n863 );
and ( n27075 , n27073 , n27074 );
buf ( n27076 , n27075 );
buf ( n27077 , n27076 );
not ( n27078 , n23144 );
xor ( n27079 , n888 , n858 );
not ( n27080 , n27079 );
or ( n27081 , n27078 , n27080 );
buf ( n27082 , n20363 );
buf ( n27083 , n26748 );
nand ( n27084 , n27082 , n27083 );
buf ( n27085 , n27084 );
nand ( n27086 , n27081 , n27085 );
buf ( n27087 , n27086 );
xor ( n27088 , n27077 , n27087 );
buf ( n27089 , n854 );
buf ( n27090 , n892 );
xor ( n27091 , n27089 , n27090 );
buf ( n27092 , n27091 );
buf ( n27093 , n27092 );
not ( n27094 , n27093 );
buf ( n27095 , n23175 );
not ( n27096 , n27095 );
or ( n27097 , n27094 , n27096 );
buf ( n27098 , n23181 );
buf ( n27099 , n26793 );
nand ( n27100 , n27098 , n27099 );
buf ( n27101 , n27100 );
buf ( n27102 , n27101 );
nand ( n27103 , n27097 , n27102 );
buf ( n27104 , n27103 );
buf ( n27105 , n27104 );
and ( n27106 , n27088 , n27105 );
and ( n27107 , n27077 , n27087 );
or ( n27108 , n27106 , n27107 );
buf ( n27109 , n27108 );
buf ( n27110 , n27109 );
xor ( n27111 , n27072 , n27110 );
buf ( n27112 , n852 );
buf ( n27113 , n894 );
xor ( n27114 , n27112 , n27113 );
buf ( n27115 , n27114 );
buf ( n27116 , n27115 );
not ( n27117 , n27116 );
buf ( n27118 , n23288 );
not ( n27119 , n27118 );
or ( n27120 , n27117 , n27119 );
buf ( n27121 , n26567 );
buf ( n27122 , n895 );
nand ( n27123 , n27121 , n27122 );
buf ( n27124 , n27123 );
buf ( n27125 , n27124 );
nand ( n27126 , n27120 , n27125 );
buf ( n27127 , n27126 );
buf ( n27128 , n27127 );
buf ( n27129 , n860 );
buf ( n27130 , n886 );
xor ( n27131 , n27129 , n27130 );
buf ( n27132 , n27131 );
buf ( n27133 , n27132 );
not ( n27134 , n27133 );
buf ( n27135 , n20521 );
not ( n27136 , n27135 );
or ( n27137 , n27134 , n27136 );
buf ( n27138 , n20525 );
buf ( n27139 , n26770 );
nand ( n27140 , n27138 , n27139 );
buf ( n27141 , n27140 );
buf ( n27142 , n27141 );
nand ( n27143 , n27137 , n27142 );
buf ( n27144 , n27143 );
buf ( n27145 , n27144 );
xor ( n27146 , n27128 , n27145 );
xor ( n27147 , n884 , n862 );
buf ( n27148 , n27147 );
not ( n27149 , n27148 );
buf ( n27150 , n25022 );
not ( n27151 , n27150 );
or ( n27152 , n27149 , n27151 );
buf ( n27153 , n25263 );
buf ( n27154 , n26847 );
nand ( n27155 , n27153 , n27154 );
buf ( n27156 , n27155 );
buf ( n27157 , n27156 );
nand ( n27158 , n27152 , n27157 );
buf ( n27159 , n27158 );
buf ( n27160 , n27159 );
and ( n27161 , n27146 , n27160 );
and ( n27162 , n27128 , n27145 );
or ( n27163 , n27161 , n27162 );
buf ( n27164 , n27163 );
buf ( n27165 , n27164 );
and ( n27166 , n27111 , n27165 );
and ( n27167 , n27072 , n27110 );
or ( n27168 , n27166 , n27167 );
buf ( n27169 , n27168 );
buf ( n27170 , n27169 );
and ( n27171 , n27067 , n27170 );
and ( n27172 , n27062 , n27066 );
or ( n27173 , n27171 , n27172 );
buf ( n27174 , n27173 );
buf ( n27175 , n27174 );
xor ( n27176 , n27058 , n27175 );
xor ( n27177 , n26641 , n26739 );
xor ( n27178 , n27177 , n26870 );
buf ( n27179 , n27178 );
buf ( n27180 , n27179 );
xor ( n27181 , n27176 , n27180 );
buf ( n27182 , n27181 );
buf ( n27183 , n27182 );
buf ( n27184 , n23076 );
not ( n27185 , n27184 );
buf ( n27186 , n21441 );
not ( n27187 , n27186 );
or ( n27188 , n27185 , n27187 );
buf ( n27189 , n20869 );
xor ( n27190 , n890 , n856 );
buf ( n27191 , n27190 );
nand ( n27192 , n27189 , n27191 );
buf ( n27193 , n27192 );
buf ( n27194 , n27193 );
nand ( n27195 , n27188 , n27194 );
buf ( n27196 , n27195 );
xor ( n27197 , n884 , n863 );
buf ( n27198 , n27197 );
not ( n27199 , n27198 );
buf ( n27200 , n25022 );
not ( n27201 , n27200 );
or ( n27202 , n27199 , n27201 );
buf ( n27203 , n25263 );
buf ( n27204 , n27147 );
nand ( n27205 , n27203 , n27204 );
buf ( n27206 , n27205 );
buf ( n27207 , n27206 );
nand ( n27208 , n27202 , n27207 );
buf ( n27209 , n27208 );
xor ( n27210 , n27196 , n27209 );
buf ( n27211 , n27210 );
buf ( n27212 , n863 );
buf ( n27213 , n885 );
or ( n27214 , n27212 , n27213 );
buf ( n27215 , n886 );
nand ( n27216 , n27214 , n27215 );
buf ( n27217 , n27216 );
buf ( n27218 , n27217 );
buf ( n27219 , n863 );
buf ( n27220 , n885 );
nand ( n27221 , n27219 , n27220 );
buf ( n27222 , n27221 );
buf ( n27223 , n27222 );
buf ( n27224 , n884 );
nand ( n27225 , n27218 , n27223 , n27224 );
buf ( n27226 , n27225 );
buf ( n27227 , n27226 );
not ( n27228 , n27227 );
buf ( n27229 , n23274 );
not ( n27230 , n27229 );
buf ( n27231 , n23175 );
not ( n27232 , n27231 );
or ( n27233 , n27230 , n27232 );
buf ( n27234 , n23181 );
buf ( n27235 , n27092 );
nand ( n27236 , n27234 , n27235 );
buf ( n27237 , n27236 );
buf ( n27238 , n27237 );
nand ( n27239 , n27233 , n27238 );
buf ( n27240 , n27239 );
buf ( n27241 , n27240 );
not ( n27242 , n27241 );
or ( n27243 , n27228 , n27242 );
buf ( n27244 , n27240 );
buf ( n27245 , n27226 );
or ( n27246 , n27244 , n27245 );
nand ( n27247 , n27243 , n27246 );
buf ( n27248 , n27247 );
buf ( n27249 , n27248 );
xor ( n27250 , n27211 , n27249 );
buf ( n27251 , n27250 );
buf ( n27252 , n27251 );
xor ( n27253 , n23242 , n23263 );
and ( n27254 , n27253 , n23281 );
and ( n27255 , n23242 , n23263 );
or ( n27256 , n27254 , n27255 );
buf ( n27257 , n27256 );
buf ( n27258 , n27257 );
buf ( n27259 , n23082 );
buf ( n27260 , n23061 );
or ( n27261 , n27259 , n27260 );
buf ( n27262 , n23041 );
nand ( n27263 , n27261 , n27262 );
buf ( n27264 , n27263 );
buf ( n27265 , n27264 );
buf ( n27266 , n23082 );
buf ( n27267 , n23061 );
nand ( n27268 , n27266 , n27267 );
buf ( n27269 , n27268 );
buf ( n27270 , n27269 );
nand ( n27271 , n27265 , n27270 );
buf ( n27272 , n27271 );
buf ( n27273 , n27272 );
xor ( n27274 , n27258 , n27273 );
buf ( n27275 , n23054 );
not ( n27276 , n27275 );
buf ( n27277 , n21297 );
not ( n27278 , n27277 );
or ( n27279 , n27276 , n27278 );
buf ( n27280 , n27115 );
buf ( n27281 , n895 );
nand ( n27282 , n27280 , n27281 );
buf ( n27283 , n27282 );
buf ( n27284 , n27283 );
nand ( n27285 , n27279 , n27284 );
buf ( n27286 , n27285 );
buf ( n27287 , n27286 );
buf ( n27288 , n23035 );
not ( n27289 , n27288 );
buf ( n27290 , n20521 );
not ( n27291 , n27290 );
or ( n27292 , n27289 , n27291 );
buf ( n27293 , n20525 );
buf ( n27294 , n27132 );
nand ( n27295 , n27293 , n27294 );
buf ( n27296 , n27295 );
buf ( n27297 , n27296 );
nand ( n27298 , n27292 , n27297 );
buf ( n27299 , n27298 );
buf ( n27300 , n27299 );
xor ( n27301 , n27287 , n27300 );
buf ( n27302 , n23256 );
not ( n27303 , n27302 );
buf ( n27304 , n23144 );
not ( n27305 , n27304 );
or ( n27306 , n27303 , n27305 );
buf ( n27307 , n27079 );
buf ( n27308 , n20363 );
nand ( n27309 , n27307 , n27308 );
buf ( n27310 , n27309 );
buf ( n27311 , n27310 );
nand ( n27312 , n27306 , n27311 );
buf ( n27313 , n27312 );
buf ( n27314 , n27313 );
xor ( n27315 , n27301 , n27314 );
buf ( n27316 , n27315 );
buf ( n27317 , n27316 );
xor ( n27318 , n27274 , n27317 );
buf ( n27319 , n27318 );
buf ( n27320 , n27319 );
xor ( n27321 , n27252 , n27320 );
xor ( n27322 , n23230 , n23284 );
and ( n27323 , n27322 , n23333 );
and ( n27324 , n23230 , n23284 );
or ( n27325 , n27323 , n27324 );
buf ( n27326 , n27325 );
buf ( n27327 , n27326 );
xor ( n27328 , n27321 , n27327 );
buf ( n27329 , n27328 );
buf ( n27330 , n27329 );
buf ( n27331 , n859 );
buf ( n27332 , n892 );
xor ( n27333 , n27331 , n27332 );
buf ( n27334 , n27333 );
not ( n27335 , n27334 );
not ( n27336 , n23175 );
or ( n27337 , n27335 , n27336 );
buf ( n27338 , n23181 );
buf ( n27339 , n858 );
buf ( n27340 , n892 );
xor ( n27341 , n27339 , n27340 );
buf ( n27342 , n27341 );
buf ( n27343 , n27342 );
nand ( n27344 , n27338 , n27343 );
buf ( n27345 , n27344 );
nand ( n27346 , n27337 , n27345 );
buf ( n27347 , n861 );
buf ( n27348 , n890 );
xor ( n27349 , n27347 , n27348 );
buf ( n27350 , n27349 );
not ( n27351 , n27350 );
not ( n27352 , n21441 );
or ( n27353 , n27351 , n27352 );
buf ( n27354 , n20869 );
buf ( n27355 , n860 );
buf ( n27356 , n890 );
xor ( n27357 , n27355 , n27356 );
buf ( n27358 , n27357 );
buf ( n27359 , n27358 );
nand ( n27360 , n27354 , n27359 );
buf ( n27361 , n27360 );
nand ( n27362 , n27353 , n27361 );
xor ( n27363 , n27346 , n27362 );
buf ( n27364 , n863 );
buf ( n27365 , n888 );
xor ( n27366 , n27364 , n27365 );
buf ( n27367 , n27366 );
not ( n27368 , n27367 );
not ( n27369 , n23144 );
or ( n27370 , n27368 , n27369 );
buf ( n27371 , n20363 );
buf ( n27372 , n27371 );
buf ( n27373 , n23139 );
nand ( n27374 , n27372 , n27373 );
buf ( n27375 , n27374 );
nand ( n27376 , n27370 , n27375 );
and ( n27377 , n27363 , n27376 );
and ( n27378 , n27346 , n27362 );
or ( n27379 , n27377 , n27378 );
buf ( n27380 , n23158 );
buf ( n27381 , n23109 );
not ( n27382 , n27381 );
buf ( n27383 , n23124 );
not ( n27384 , n27383 );
or ( n27385 , n27382 , n27384 );
buf ( n27386 , n23124 );
buf ( n27387 , n23109 );
or ( n27388 , n27386 , n27387 );
nand ( n27389 , n27385 , n27388 );
buf ( n27390 , n27389 );
buf ( n27391 , n27390 );
xor ( n27392 , n27380 , n27391 );
buf ( n27393 , n27392 );
not ( n27394 , n27393 );
xor ( n27395 , n27379 , n27394 );
buf ( n27396 , n27358 );
not ( n27397 , n27396 );
buf ( n27398 , n21441 );
not ( n27399 , n27398 );
or ( n27400 , n27397 , n27399 );
buf ( n27401 , n20869 );
buf ( n27402 , n23088 );
nand ( n27403 , n27401 , n27402 );
buf ( n27404 , n27403 );
buf ( n27405 , n27404 );
nand ( n27406 , n27400 , n27405 );
buf ( n27407 , n27406 );
buf ( n27408 , n27342 );
not ( n27409 , n27408 );
buf ( n27410 , n23175 );
not ( n27411 , n27410 );
or ( n27412 , n27409 , n27411 );
buf ( n27413 , n23181 );
buf ( n27414 , n23170 );
nand ( n27415 , n27413 , n27414 );
buf ( n27416 , n27415 );
buf ( n27417 , n27416 );
nand ( n27418 , n27412 , n27417 );
buf ( n27419 , n27418 );
xor ( n27420 , n27407 , n27419 );
buf ( n27421 , n857 );
buf ( n27422 , n894 );
xor ( n27423 , n27421 , n27422 );
buf ( n27424 , n27423 );
buf ( n27425 , n27424 );
not ( n27426 , n27425 );
buf ( n27427 , n23288 );
not ( n27428 , n27427 );
or ( n27429 , n27426 , n27428 );
buf ( n27430 , n23116 );
buf ( n27431 , n895 );
nand ( n27432 , n27430 , n27431 );
buf ( n27433 , n27432 );
buf ( n27434 , n27433 );
nand ( n27435 , n27429 , n27434 );
buf ( n27436 , n27435 );
buf ( n27437 , n27436 );
buf ( n27438 , n863 );
buf ( n27439 , n889 );
or ( n27440 , n27438 , n27439 );
buf ( n27441 , n890 );
nand ( n27442 , n27440 , n27441 );
buf ( n27443 , n27442 );
buf ( n27444 , n27443 );
buf ( n27445 , n863 );
buf ( n27446 , n889 );
nand ( n27447 , n27445 , n27446 );
buf ( n27448 , n27447 );
buf ( n27449 , n27448 );
buf ( n27450 , n888 );
nand ( n27451 , n27444 , n27449 , n27450 );
buf ( n27452 , n27451 );
buf ( n27453 , n27452 );
not ( n27454 , n27453 );
buf ( n27455 , n27454 );
buf ( n27456 , n27455 );
nand ( n27457 , n27437 , n27456 );
buf ( n27458 , n27457 );
buf ( n27459 , n27458 );
not ( n27460 , n27459 );
buf ( n27461 , n27460 );
and ( n27462 , n27420 , n27461 );
not ( n27463 , n27420 );
and ( n27464 , n27463 , n27458 );
or ( n27465 , n27462 , n27464 );
xnor ( n27466 , n27395 , n27465 );
not ( n27467 , n27466 );
buf ( n27468 , n27467 );
buf ( n27469 , n863 );
buf ( n27470 , n893 );
or ( n27471 , n27469 , n27470 );
buf ( n27472 , n894 );
nand ( n27473 , n27471 , n27472 );
buf ( n27474 , n27473 );
buf ( n27475 , n27474 );
buf ( n27476 , n863 );
buf ( n27477 , n893 );
nand ( n27478 , n27476 , n27477 );
buf ( n27479 , n27478 );
buf ( n27480 , n27479 );
buf ( n27481 , n892 );
and ( n27482 , n27475 , n27480 , n27481 );
buf ( n27483 , n27482 );
buf ( n27484 , n27483 );
buf ( n27485 , n861 );
buf ( n27486 , n894 );
xor ( n27487 , n27485 , n27486 );
buf ( n27488 , n27487 );
buf ( n27489 , n27488 );
not ( n27490 , n27489 );
buf ( n27491 , n21297 );
not ( n27492 , n27491 );
or ( n27493 , n27490 , n27492 );
buf ( n27494 , n860 );
buf ( n27495 , n894 );
xor ( n27496 , n27494 , n27495 );
buf ( n27497 , n27496 );
buf ( n27498 , n27497 );
buf ( n27499 , n895 );
nand ( n27500 , n27498 , n27499 );
buf ( n27501 , n27500 );
buf ( n27502 , n27501 );
nand ( n27503 , n27493 , n27502 );
buf ( n27504 , n27503 );
buf ( n27505 , n27504 );
xor ( n27506 , n27484 , n27505 );
buf ( n27507 , n27506 );
buf ( n27508 , n27507 );
xor ( n27509 , n24449 , n24836 );
and ( n27510 , n27509 , n24852 );
and ( n27511 , n24449 , n24836 );
or ( n27512 , n27510 , n27511 );
buf ( n27513 , n27512 );
buf ( n27514 , n27513 );
xor ( n27515 , n27072 , n27110 );
xor ( n27516 , n27515 , n27165 );
buf ( n27517 , n27516 );
buf ( n27518 , n27517 );
xor ( n27519 , n27077 , n27087 );
xor ( n27520 , n27519 , n27105 );
buf ( n27521 , n27520 );
buf ( n27522 , n27521 );
xor ( n27523 , n27128 , n27145 );
xor ( n27524 , n27523 , n27160 );
buf ( n27525 , n27524 );
buf ( n27526 , n27525 );
xor ( n27527 , n27522 , n27526 );
buf ( n27528 , n27209 );
buf ( n27529 , n27196 );
or ( n27530 , n27528 , n27529 );
buf ( n27531 , n27530 );
not ( n27532 , n27531 );
not ( n27533 , n27248 );
or ( n27534 , n27532 , n27533 );
buf ( n27535 , n27196 );
buf ( n27536 , n27209 );
nand ( n27537 , n27535 , n27536 );
buf ( n27538 , n27537 );
nand ( n27539 , n27534 , n27538 );
buf ( n27540 , n27539 );
and ( n27541 , n27527 , n27540 );
and ( n27542 , n27522 , n27526 );
or ( n27543 , n27541 , n27542 );
buf ( n27544 , n27543 );
buf ( n27545 , n27544 );
xor ( n27546 , n27518 , n27545 );
buf ( n27547 , n26805 );
buf ( n27548 , n27547 );
not ( n27549 , n27548 );
xnor ( n27550 , n26786 , n26764 );
buf ( n27551 , n27550 );
not ( n27552 , n27551 );
or ( n27553 , n27549 , n27552 );
buf ( n27554 , n27550 );
buf ( n27555 , n27547 );
or ( n27556 , n27554 , n27555 );
nand ( n27557 , n27553 , n27556 );
buf ( n27558 , n27557 );
buf ( n27559 , n27558 );
xor ( n27560 , n26827 , n26845 );
xor ( n27561 , n27560 , n26860 );
buf ( n27562 , n27561 );
buf ( n27563 , n27562 );
xor ( n27564 , n27559 , n27563 );
buf ( n27565 , n27190 );
not ( n27566 , n27565 );
buf ( n27567 , n21441 );
not ( n27568 , n27567 );
or ( n27569 , n27566 , n27568 );
buf ( n27570 , n20869 );
buf ( n27571 , n27570 );
buf ( n27572 , n26831 );
nand ( n27573 , n27571 , n27572 );
buf ( n27574 , n27573 );
buf ( n27575 , n27574 );
nand ( n27576 , n27569 , n27575 );
buf ( n27577 , n27576 );
buf ( n27578 , n27577 );
buf ( n27579 , n27240 );
not ( n27580 , n27579 );
buf ( n27581 , n27226 );
nor ( n27582 , n27580 , n27581 );
buf ( n27583 , n27582 );
buf ( n27584 , n27583 );
xor ( n27585 , n27578 , n27584 );
xor ( n27586 , n27287 , n27300 );
and ( n27587 , n27586 , n27314 );
and ( n27588 , n27287 , n27300 );
or ( n27589 , n27587 , n27588 );
buf ( n27590 , n27589 );
buf ( n27591 , n27590 );
and ( n27592 , n27585 , n27591 );
and ( n27593 , n27578 , n27584 );
or ( n27594 , n27592 , n27593 );
buf ( n27595 , n27594 );
buf ( n27596 , n27595 );
xor ( n27597 , n27564 , n27596 );
buf ( n27598 , n27597 );
buf ( n27599 , n27598 );
xor ( n27600 , n27546 , n27599 );
buf ( n27601 , n27600 );
buf ( n27602 , n27601 );
buf ( n27603 , n863 );
buf ( n27604 , n877 );
or ( n27605 , n27603 , n27604 );
buf ( n27606 , n878 );
nand ( n27607 , n27605 , n27606 );
buf ( n27608 , n27607 );
buf ( n27609 , n27608 );
buf ( n27610 , n863 );
buf ( n27611 , n877 );
nand ( n27612 , n27610 , n27611 );
buf ( n27613 , n27612 );
buf ( n27614 , n27613 );
buf ( n27615 , n876 );
nand ( n27616 , n27609 , n27614 , n27615 );
buf ( n27617 , n27616 );
buf ( n27618 , n27617 );
not ( n27619 , n27618 );
xor ( n27620 , n894 , n845 );
buf ( n27621 , n27620 );
not ( n27622 , n27621 );
buf ( n27623 , n20132 );
not ( n27624 , n27623 );
or ( n27625 , n27622 , n27624 );
xor ( n27626 , n894 , n844 );
buf ( n27627 , n27626 );
buf ( n27628 , n895 );
nand ( n27629 , n27627 , n27628 );
buf ( n27630 , n27629 );
buf ( n27631 , n27630 );
nand ( n27632 , n27625 , n27631 );
buf ( n27633 , n27632 );
buf ( n27634 , n27633 );
nand ( n27635 , n27619 , n27634 );
buf ( n27636 , n27635 );
buf ( n27637 , n27636 );
not ( n27638 , n27637 );
buf ( n27639 , n856 );
buf ( n27640 , n882 );
xor ( n27641 , n27639 , n27640 );
buf ( n27642 , n27641 );
buf ( n27643 , n27642 );
not ( n27644 , n27643 );
buf ( n27645 , n19580 );
not ( n27646 , n27645 );
or ( n27647 , n27644 , n27646 );
buf ( n27648 , n26538 );
xor ( n27649 , n882 , n855 );
buf ( n27650 , n27649 );
nand ( n27651 , n27648 , n27650 );
buf ( n27652 , n27651 );
buf ( n27653 , n27652 );
nand ( n27654 , n27647 , n27653 );
buf ( n27655 , n27654 );
buf ( n27656 , n27655 );
nor ( n27657 , n27638 , n27656 );
buf ( n27658 , n27657 );
buf ( n27659 , n27658 );
not ( n27660 , n27659 );
buf ( n27661 , n27636 );
not ( n27662 , n27661 );
buf ( n27663 , n27655 );
nand ( n27664 , n27662 , n27663 );
buf ( n27665 , n27664 );
buf ( n27666 , n27665 );
nand ( n27667 , n27660 , n27666 );
buf ( n27668 , n27667 );
buf ( n27669 , n27668 );
buf ( n27670 , n854 );
buf ( n27671 , n884 );
xor ( n27672 , n27670 , n27671 );
buf ( n27673 , n27672 );
buf ( n27674 , n27673 );
not ( n27675 , n27674 );
buf ( n27676 , n25022 );
not ( n27677 , n27676 );
or ( n27678 , n27675 , n27677 );
buf ( n27679 , n25263 );
buf ( n27680 , n853 );
buf ( n27681 , n884 );
xor ( n27682 , n27680 , n27681 );
buf ( n27683 , n27682 );
buf ( n27684 , n27683 );
nand ( n27685 , n27679 , n27684 );
buf ( n27686 , n27685 );
buf ( n27687 , n27686 );
nand ( n27688 , n27678 , n27687 );
buf ( n27689 , n27688 );
buf ( n27690 , n27689 );
not ( n27691 , n27690 );
buf ( n27692 , n27691 );
and ( n27693 , n27669 , n27692 );
not ( n27694 , n27669 );
buf ( n27695 , n27690 );
and ( n27696 , n27694 , n27695 );
nor ( n27697 , n27693 , n27696 );
buf ( n27698 , n27697 );
buf ( n27699 , n27698 );
buf ( n27700 , n27617 );
not ( n27701 , n27700 );
buf ( n27702 , n27633 );
not ( n27703 , n27702 );
or ( n27704 , n27701 , n27703 );
buf ( n27705 , n27633 );
buf ( n27706 , n27617 );
or ( n27707 , n27705 , n27706 );
nand ( n27708 , n27704 , n27707 );
buf ( n27709 , n27708 );
buf ( n27710 , n27709 );
buf ( n27711 , n846 );
buf ( n27712 , n894 );
xor ( n27713 , n27711 , n27712 );
buf ( n27714 , n27713 );
buf ( n27715 , n27714 );
not ( n27716 , n27715 );
buf ( n27717 , n21297 );
not ( n27718 , n27717 );
or ( n27719 , n27716 , n27718 );
buf ( n27720 , n27620 );
buf ( n27721 , n895 );
nand ( n27722 , n27720 , n27721 );
buf ( n27723 , n27722 );
buf ( n27724 , n27723 );
nand ( n27725 , n27719 , n27724 );
buf ( n27726 , n27725 );
buf ( n27727 , n27726 );
buf ( n27728 , n19082 );
buf ( n27729 , n863 );
and ( n27730 , n27728 , n27729 );
buf ( n27731 , n27730 );
buf ( n27732 , n27731 );
xor ( n27733 , n27727 , n27732 );
buf ( n27734 , n23144 );
not ( n27735 , n27734 );
buf ( n27736 , n27735 );
buf ( n27737 , n27736 );
buf ( n27738 , n852 );
buf ( n27739 , n888 );
xnor ( n27740 , n27738 , n27739 );
buf ( n27741 , n27740 );
buf ( n27742 , n27741 );
or ( n27743 , n27737 , n27742 );
buf ( n27744 , n25724 );
buf ( n27745 , n851 );
buf ( n27746 , n888 );
xor ( n27747 , n27745 , n27746 );
buf ( n27748 , n27747 );
buf ( n27749 , n27748 );
not ( n27750 , n27749 );
buf ( n27751 , n27750 );
buf ( n27752 , n27751 );
or ( n27753 , n27744 , n27752 );
nand ( n27754 , n27743 , n27753 );
buf ( n27755 , n27754 );
buf ( n27756 , n27755 );
and ( n27757 , n27733 , n27756 );
and ( n27758 , n27727 , n27732 );
or ( n27759 , n27757 , n27758 );
buf ( n27760 , n27759 );
buf ( n27761 , n27760 );
xor ( n27762 , n27710 , n27761 );
xor ( n27763 , n892 , n848 );
buf ( n27764 , n27763 );
not ( n27765 , n27764 );
buf ( n27766 , n23175 );
not ( n27767 , n27766 );
or ( n27768 , n27765 , n27767 );
buf ( n27769 , n22818 );
xor ( n27770 , n892 , n847 );
buf ( n27771 , n27770 );
nand ( n27772 , n27769 , n27771 );
buf ( n27773 , n27772 );
buf ( n27774 , n27773 );
nand ( n27775 , n27768 , n27774 );
buf ( n27776 , n27775 );
buf ( n27777 , n27776 );
buf ( n27778 , n859 );
buf ( n27779 , n880 );
xor ( n27780 , n27778 , n27779 );
buf ( n27781 , n27780 );
buf ( n27782 , n27781 );
not ( n27783 , n27782 );
buf ( n27784 , n18860 );
not ( n27785 , n27784 );
or ( n27786 , n27783 , n27785 );
buf ( n27787 , n18850 );
buf ( n27788 , n860 );
buf ( n27789 , n880 );
xor ( n27790 , n27788 , n27789 );
buf ( n27791 , n27790 );
buf ( n27792 , n27791 );
nand ( n27793 , n27787 , n27792 );
buf ( n27794 , n27793 );
buf ( n27795 , n27794 );
nand ( n27796 , n27786 , n27795 );
buf ( n27797 , n27796 );
buf ( n27798 , n27797 );
xor ( n27799 , n27777 , n27798 );
buf ( n27800 , n862 );
buf ( n27801 , n878 );
xor ( n27802 , n27800 , n27801 );
buf ( n27803 , n27802 );
buf ( n27804 , n27803 );
not ( n27805 , n27804 );
buf ( n27806 , n19259 );
not ( n27807 , n27806 );
or ( n27808 , n27805 , n27807 );
buf ( n27809 , n19265 );
buf ( n27810 , n861 );
buf ( n27811 , n878 );
xor ( n27812 , n27810 , n27811 );
buf ( n27813 , n27812 );
buf ( n27814 , n27813 );
nand ( n27815 , n27809 , n27814 );
buf ( n27816 , n27815 );
buf ( n27817 , n27816 );
nand ( n27818 , n27808 , n27817 );
buf ( n27819 , n27818 );
buf ( n27820 , n27819 );
and ( n27821 , n27799 , n27820 );
and ( n27822 , n27777 , n27798 );
or ( n27823 , n27821 , n27822 );
buf ( n27824 , n27823 );
buf ( n27825 , n27824 );
and ( n27826 , n27762 , n27825 );
and ( n27827 , n27710 , n27761 );
or ( n27828 , n27826 , n27827 );
buf ( n27829 , n27828 );
buf ( n27830 , n27829 );
xor ( n27831 , n27699 , n27830 );
not ( n27832 , n27748 );
not ( n27833 , n20358 );
or ( n27834 , n27832 , n27833 );
buf ( n27835 , n850 );
buf ( n27836 , n888 );
xor ( n27837 , n27835 , n27836 );
buf ( n27838 , n27837 );
nand ( n27839 , n20363 , n27838 );
nand ( n27840 , n27834 , n27839 );
buf ( n27841 , n27781 );
not ( n27842 , n27841 );
buf ( n27843 , n18850 );
not ( n27844 , n27843 );
or ( n27845 , n27842 , n27844 );
buf ( n27846 , n22271 );
buf ( n27847 , n858 );
buf ( n27848 , n880 );
xor ( n27849 , n27847 , n27848 );
buf ( n27850 , n27849 );
buf ( n27851 , n27850 );
nand ( n27852 , n27846 , n27851 );
buf ( n27853 , n27852 );
buf ( n27854 , n27853 );
nand ( n27855 , n27845 , n27854 );
buf ( n27856 , n27855 );
xor ( n27857 , n27840 , n27856 );
buf ( n27858 , n27813 );
not ( n27859 , n27858 );
buf ( n27860 , n19259 );
not ( n27861 , n27860 );
or ( n27862 , n27859 , n27861 );
buf ( n27863 , n19265 );
buf ( n27864 , n860 );
buf ( n27865 , n878 );
xor ( n27866 , n27864 , n27865 );
buf ( n27867 , n27866 );
buf ( n27868 , n27867 );
nand ( n27869 , n27863 , n27868 );
buf ( n27870 , n27869 );
buf ( n27871 , n27870 );
nand ( n27872 , n27862 , n27871 );
buf ( n27873 , n27872 );
xor ( n27874 , n27857 , n27873 );
buf ( n27875 , n27874 );
buf ( n27876 , n850 );
buf ( n27877 , n890 );
xor ( n27878 , n27876 , n27877 );
buf ( n27879 , n27878 );
buf ( n27880 , n27879 );
not ( n27881 , n27880 );
buf ( n27882 , n21441 );
not ( n27883 , n27882 );
or ( n27884 , n27881 , n27883 );
buf ( n27885 , n20869 );
buf ( n27886 , n849 );
buf ( n27887 , n890 );
xor ( n27888 , n27886 , n27887 );
buf ( n27889 , n27888 );
buf ( n27890 , n27889 );
nand ( n27891 , n27885 , n27890 );
buf ( n27892 , n27891 );
buf ( n27893 , n27892 );
nand ( n27894 , n27884 , n27893 );
buf ( n27895 , n27894 );
not ( n27896 , n27895 );
buf ( n27897 , n854 );
buf ( n27898 , n886 );
xor ( n27899 , n27897 , n27898 );
buf ( n27900 , n27899 );
buf ( n27901 , n27900 );
not ( n27902 , n27901 );
buf ( n27903 , n20521 );
not ( n27904 , n27903 );
or ( n27905 , n27902 , n27904 );
buf ( n27906 , n23320 );
buf ( n27907 , n853 );
buf ( n27908 , n886 );
xor ( n27909 , n27907 , n27908 );
buf ( n27910 , n27909 );
buf ( n27911 , n27910 );
nand ( n27912 , n27906 , n27911 );
buf ( n27913 , n27912 );
buf ( n27914 , n27913 );
nand ( n27915 , n27905 , n27914 );
buf ( n27916 , n27915 );
not ( n27917 , n27916 );
or ( n27918 , n27896 , n27917 );
or ( n27919 , n27895 , n27916 );
buf ( n27920 , n856 );
buf ( n27921 , n884 );
xor ( n27922 , n27920 , n27921 );
buf ( n27923 , n27922 );
buf ( n27924 , n27923 );
not ( n27925 , n27924 );
buf ( n27926 , n25022 );
not ( n27927 , n27926 );
or ( n27928 , n27925 , n27927 );
buf ( n27929 , n23233 );
buf ( n27930 , n855 );
buf ( n27931 , n884 );
xor ( n27932 , n27930 , n27931 );
buf ( n27933 , n27932 );
buf ( n27934 , n27933 );
nand ( n27935 , n27929 , n27934 );
buf ( n27936 , n27935 );
buf ( n27937 , n27936 );
nand ( n27938 , n27928 , n27937 );
buf ( n27939 , n27938 );
nand ( n27940 , n27919 , n27939 );
nand ( n27941 , n27918 , n27940 );
buf ( n27942 , n27941 );
or ( n27943 , n27875 , n27942 );
not ( n27944 , n27889 );
not ( n27945 , n21441 );
or ( n27946 , n27944 , n27945 );
buf ( n27947 , n20869 );
buf ( n27948 , n848 );
buf ( n27949 , n890 );
xor ( n27950 , n27948 , n27949 );
buf ( n27951 , n27950 );
buf ( n27952 , n27951 );
nand ( n27953 , n27947 , n27952 );
buf ( n27954 , n27953 );
nand ( n27955 , n27946 , n27954 );
buf ( n27956 , n27955 );
buf ( n27957 , n857 );
buf ( n27958 , n882 );
xor ( n27959 , n27957 , n27958 );
buf ( n27960 , n27959 );
not ( n27961 , n27960 );
not ( n27962 , n19580 );
or ( n27963 , n27961 , n27962 );
buf ( n27964 , n26538 );
buf ( n27965 , n27642 );
nand ( n27966 , n27964 , n27965 );
buf ( n27967 , n27966 );
nand ( n27968 , n27963 , n27967 );
buf ( n27969 , n27968 );
xor ( n27970 , n27956 , n27969 );
buf ( n27971 , n27970 );
buf ( n27972 , n27971 );
buf ( n27973 , n27933 );
not ( n27974 , n27973 );
buf ( n27975 , n25022 );
not ( n27976 , n27975 );
or ( n27977 , n27974 , n27976 );
buf ( n27978 , n23233 );
buf ( n27979 , n27673 );
nand ( n27980 , n27978 , n27979 );
buf ( n27981 , n27980 );
buf ( n27982 , n27981 );
nand ( n27983 , n27977 , n27982 );
buf ( n27984 , n27983 );
buf ( n27985 , n27984 );
xor ( n27986 , n27972 , n27985 );
buf ( n27987 , n27986 );
buf ( n27988 , n27987 );
nand ( n27989 , n27943 , n27988 );
buf ( n27990 , n27989 );
buf ( n27991 , n27990 );
buf ( n27992 , n27941 );
buf ( n27993 , n27874 );
nand ( n27994 , n27992 , n27993 );
buf ( n27995 , n27994 );
buf ( n27996 , n27995 );
nand ( n27997 , n27991 , n27996 );
buf ( n27998 , n27997 );
buf ( n27999 , n27998 );
and ( n28000 , n27831 , n27999 );
and ( n28001 , n27699 , n27830 );
or ( n28002 , n28000 , n28001 );
buf ( n28003 , n28002 );
buf ( n28004 , n28003 );
buf ( n28005 , n20555 );
buf ( n28006 , n863 );
and ( n28007 , n28005 , n28006 );
buf ( n28008 , n28007 );
buf ( n28009 , n28008 );
buf ( n28010 , n27626 );
not ( n28011 , n28010 );
buf ( n28012 , n23288 );
not ( n28013 , n28012 );
or ( n28014 , n28011 , n28013 );
buf ( n28015 , n843 );
buf ( n28016 , n894 );
xor ( n28017 , n28015 , n28016 );
buf ( n28018 , n28017 );
buf ( n28019 , n28018 );
buf ( n28020 , n895 );
nand ( n28021 , n28019 , n28020 );
buf ( n28022 , n28021 );
buf ( n28023 , n28022 );
nand ( n28024 , n28014 , n28023 );
buf ( n28025 , n28024 );
buf ( n28026 , n28025 );
xor ( n28027 , n28009 , n28026 );
buf ( n28028 , n27838 );
not ( n28029 , n28028 );
buf ( n28030 , n20358 );
not ( n28031 , n28030 );
or ( n28032 , n28029 , n28031 );
buf ( n28033 , n20363 );
buf ( n28034 , n849 );
buf ( n28035 , n888 );
xor ( n28036 , n28034 , n28035 );
buf ( n28037 , n28036 );
buf ( n28038 , n28037 );
nand ( n28039 , n28033 , n28038 );
buf ( n28040 , n28039 );
buf ( n28041 , n28040 );
nand ( n28042 , n28032 , n28041 );
buf ( n28043 , n28042 );
buf ( n28044 , n28043 );
xor ( n28045 , n28027 , n28044 );
buf ( n28046 , n28045 );
buf ( n28047 , n28046 );
buf ( n28048 , n27951 );
not ( n28049 , n28048 );
buf ( n28050 , n21441 );
not ( n28051 , n28050 );
or ( n28052 , n28049 , n28051 );
buf ( n28053 , n20869 );
buf ( n28054 , n847 );
buf ( n28055 , n890 );
xor ( n28056 , n28054 , n28055 );
buf ( n28057 , n28056 );
buf ( n28058 , n28057 );
nand ( n28059 , n28053 , n28058 );
buf ( n28060 , n28059 );
buf ( n28061 , n28060 );
nand ( n28062 , n28052 , n28061 );
buf ( n28063 , n28062 );
buf ( n28064 , n28063 );
buf ( n28065 , n862 );
buf ( n28066 , n876 );
xor ( n28067 , n28065 , n28066 );
buf ( n28068 , n28067 );
buf ( n28069 , n28068 );
not ( n28070 , n28069 );
buf ( n28071 , n19153 );
not ( n28072 , n28071 );
or ( n28073 , n28070 , n28072 );
buf ( n28074 , n19082 );
buf ( n28075 , n861 );
buf ( n28076 , n876 );
xor ( n28077 , n28075 , n28076 );
buf ( n28078 , n28077 );
buf ( n28079 , n28078 );
nand ( n28080 , n28074 , n28079 );
buf ( n28081 , n28080 );
buf ( n28082 , n28081 );
nand ( n28083 , n28073 , n28082 );
buf ( n28084 , n28083 );
buf ( n28085 , n28084 );
xor ( n28086 , n28064 , n28085 );
xor ( n28087 , n886 , n852 );
buf ( n28088 , n28087 );
not ( n28089 , n28088 );
buf ( n28090 , n23027 );
not ( n28091 , n28090 );
or ( n28092 , n28089 , n28091 );
buf ( n28093 , n20525 );
buf ( n28094 , n851 );
buf ( n28095 , n886 );
xor ( n28096 , n28094 , n28095 );
buf ( n28097 , n28096 );
buf ( n28098 , n28097 );
nand ( n28099 , n28093 , n28098 );
buf ( n28100 , n28099 );
buf ( n28101 , n28100 );
nand ( n28102 , n28092 , n28101 );
buf ( n28103 , n28102 );
buf ( n28104 , n28103 );
xor ( n28105 , n28086 , n28104 );
buf ( n28106 , n28105 );
buf ( n28107 , n28106 );
xor ( n28108 , n28047 , n28107 );
buf ( n28109 , n27867 );
not ( n28110 , n28109 );
buf ( n28111 , n19259 );
not ( n28112 , n28111 );
or ( n28113 , n28110 , n28112 );
buf ( n28114 , n19265 );
buf ( n28115 , n859 );
buf ( n28116 , n878 );
xor ( n28117 , n28115 , n28116 );
buf ( n28118 , n28117 );
buf ( n28119 , n28118 );
nand ( n28120 , n28114 , n28119 );
buf ( n28121 , n28120 );
buf ( n28122 , n28121 );
nand ( n28123 , n28113 , n28122 );
buf ( n28124 , n28123 );
buf ( n28125 , n28124 );
not ( n28126 , n28125 );
buf ( n28127 , n27850 );
not ( n28128 , n28127 );
buf ( n28129 , n18850 );
not ( n28130 , n28129 );
or ( n28131 , n28128 , n28130 );
buf ( n28132 , n23917 );
buf ( n28133 , n857 );
buf ( n28134 , n880 );
xor ( n28135 , n28133 , n28134 );
buf ( n28136 , n28135 );
buf ( n28137 , n28136 );
nand ( n28138 , n28132 , n28137 );
buf ( n28139 , n28138 );
buf ( n28140 , n28139 );
nand ( n28141 , n28131 , n28140 );
buf ( n28142 , n28141 );
buf ( n28143 , n28142 );
not ( n28144 , n28143 );
buf ( n28145 , n28144 );
buf ( n28146 , n28145 );
not ( n28147 , n28146 );
or ( n28148 , n28126 , n28147 );
buf ( n28149 , n28124 );
buf ( n28150 , n28145 );
or ( n28151 , n28149 , n28150 );
nand ( n28152 , n28148 , n28151 );
buf ( n28153 , n28152 );
buf ( n28154 , n28153 );
buf ( n28155 , n846 );
buf ( n28156 , n892 );
xor ( n28157 , n28155 , n28156 );
buf ( n28158 , n28157 );
buf ( n28159 , n28158 );
not ( n28160 , n28159 );
buf ( n28161 , n23175 );
not ( n28162 , n28161 );
or ( n28163 , n28160 , n28162 );
buf ( n28164 , n22818 );
buf ( n28165 , n845 );
buf ( n28166 , n892 );
xor ( n28167 , n28165 , n28166 );
buf ( n28168 , n28167 );
buf ( n28169 , n28168 );
nand ( n28170 , n28164 , n28169 );
buf ( n28171 , n28170 );
buf ( n28172 , n28171 );
nand ( n28173 , n28163 , n28172 );
buf ( n28174 , n28173 );
buf ( n28175 , n28174 );
and ( n28176 , n28154 , n28175 );
not ( n28177 , n28154 );
buf ( n28178 , n28174 );
not ( n28179 , n28178 );
buf ( n28180 , n28179 );
buf ( n28181 , n28180 );
and ( n28182 , n28177 , n28181 );
nor ( n28183 , n28176 , n28182 );
buf ( n28184 , n28183 );
buf ( n28185 , n28184 );
xor ( n28186 , n28108 , n28185 );
buf ( n28187 , n28186 );
not ( n28188 , n28187 );
not ( n28189 , n27955 );
not ( n28190 , n27968 );
or ( n28191 , n28189 , n28190 );
or ( n28192 , n27955 , n27968 );
not ( n28193 , n27933 );
not ( n28194 , n25022 );
or ( n28195 , n28193 , n28194 );
nand ( n28196 , n28195 , n27981 );
nand ( n28197 , n28192 , n28196 );
nand ( n28198 , n28191 , n28197 );
buf ( n28199 , n28198 );
xor ( n28200 , n27840 , n27856 );
and ( n28201 , n28200 , n27873 );
and ( n28202 , n27840 , n27856 );
or ( n28203 , n28201 , n28202 );
buf ( n28204 , n28203 );
xor ( n28205 , n28199 , n28204 );
buf ( n28206 , n28205 );
buf ( n28207 , n28206 );
buf ( n28208 , n27910 );
not ( n28209 , n28208 );
buf ( n28210 , n20521 );
not ( n28211 , n28210 );
or ( n28212 , n28209 , n28211 );
buf ( n28213 , n20525 );
buf ( n28214 , n28087 );
nand ( n28215 , n28213 , n28214 );
buf ( n28216 , n28215 );
buf ( n28217 , n28216 );
nand ( n28218 , n28212 , n28217 );
buf ( n28219 , n28218 );
not ( n28220 , n28219 );
buf ( n28221 , n27770 );
not ( n28222 , n28221 );
buf ( n28223 , n23175 );
not ( n28224 , n28223 );
or ( n28225 , n28222 , n28224 );
buf ( n28226 , n22818 );
buf ( n28227 , n28158 );
nand ( n28228 , n28226 , n28227 );
buf ( n28229 , n28228 );
buf ( n28230 , n28229 );
nand ( n28231 , n28225 , n28230 );
buf ( n28232 , n28231 );
not ( n28233 , n28232 );
or ( n28234 , n28220 , n28233 );
buf ( n28235 , n28219 );
buf ( n28236 , n28232 );
or ( n28237 , n28235 , n28236 );
buf ( n28238 , n863 );
buf ( n28239 , n876 );
xor ( n28240 , n28238 , n28239 );
buf ( n28241 , n28240 );
buf ( n28242 , n28241 );
not ( n28243 , n28242 );
buf ( n28244 , n19077 );
not ( n28245 , n28244 );
or ( n28246 , n28243 , n28245 );
buf ( n28247 , n19082 );
buf ( n28248 , n28068 );
nand ( n28249 , n28247 , n28248 );
buf ( n28250 , n28249 );
buf ( n28251 , n28250 );
nand ( n28252 , n28246 , n28251 );
buf ( n28253 , n28252 );
buf ( n28254 , n28253 );
nand ( n28255 , n28237 , n28254 );
buf ( n28256 , n28255 );
nand ( n28257 , n28234 , n28256 );
buf ( n28258 , n28257 );
not ( n28259 , n28258 );
buf ( n28260 , n28259 );
buf ( n28261 , n28260 );
and ( n28262 , n28207 , n28261 );
not ( n28263 , n28207 );
buf ( n28264 , n28257 );
and ( n28265 , n28263 , n28264 );
nor ( n28266 , n28262 , n28265 );
buf ( n28267 , n28266 );
nand ( n28268 , n28188 , n28267 );
not ( n28269 , n28268 );
xor ( n28270 , n27699 , n27830 );
xor ( n28271 , n28270 , n27999 );
buf ( n28272 , n28271 );
not ( n28273 , n28272 );
or ( n28274 , n28269 , n28273 );
buf ( n28275 , n28267 );
not ( n28276 , n28275 );
buf ( n28277 , n28187 );
nand ( n28278 , n28276 , n28277 );
buf ( n28279 , n28278 );
nand ( n28280 , n28274 , n28279 );
buf ( n28281 , n28280 );
xor ( n28282 , n28004 , n28281 );
xor ( n28283 , n28047 , n28107 );
and ( n28284 , n28283 , n28185 );
and ( n28285 , n28047 , n28107 );
or ( n28286 , n28284 , n28285 );
buf ( n28287 , n28286 );
buf ( n28288 , n28287 );
buf ( n28289 , n27658 );
not ( n28290 , n27689 );
buf ( n28291 , n28290 );
or ( n28292 , n28289 , n28291 );
buf ( n28293 , n27665 );
nand ( n28294 , n28292 , n28293 );
buf ( n28295 , n28294 );
buf ( n28296 , n28295 );
buf ( n28297 , n28078 );
not ( n28298 , n28297 );
buf ( n28299 , n19153 );
not ( n28300 , n28299 );
or ( n28301 , n28298 , n28300 );
buf ( n28302 , n20246 );
buf ( n28303 , n860 );
buf ( n28304 , n876 );
xor ( n28305 , n28303 , n28304 );
buf ( n28306 , n28305 );
buf ( n28307 , n28306 );
nand ( n28308 , n28302 , n28307 );
buf ( n28309 , n28308 );
buf ( n28310 , n28309 );
nand ( n28311 , n28301 , n28310 );
buf ( n28312 , n28311 );
buf ( n28313 , n28312 );
not ( n28314 , n28313 );
buf ( n28315 , n28314 );
not ( n28316 , n28097 );
not ( n28317 , n20521 );
or ( n28318 , n28316 , n28317 );
buf ( n28319 , n850 );
buf ( n28320 , n886 );
xor ( n28321 , n28319 , n28320 );
buf ( n28322 , n28321 );
nand ( n28323 , n28322 , n20525 );
nand ( n28324 , n28318 , n28323 );
xor ( n28325 , n28315 , n28324 );
buf ( n28326 , n863 );
buf ( n28327 , n874 );
xor ( n28328 , n28326 , n28327 );
buf ( n28329 , n28328 );
buf ( n28330 , n28329 );
not ( n28331 , n28330 );
buf ( n28332 , n20549 );
not ( n28333 , n28332 );
or ( n28334 , n28331 , n28333 );
buf ( n28335 , n18987 );
xor ( n28336 , n874 , n862 );
buf ( n28337 , n28336 );
nand ( n28338 , n28335 , n28337 );
buf ( n28339 , n28338 );
buf ( n28340 , n28339 );
nand ( n28341 , n28334 , n28340 );
buf ( n28342 , n28341 );
not ( n28343 , n28342 );
xor ( n28344 , n28325 , n28343 );
buf ( n28345 , n28344 );
xor ( n28346 , n28296 , n28345 );
buf ( n28347 , n28136 );
not ( n28348 , n28347 );
buf ( n28349 , n18850 );
not ( n28350 , n28349 );
or ( n28351 , n28348 , n28350 );
buf ( n28352 , n856 );
buf ( n28353 , n880 );
xor ( n28354 , n28352 , n28353 );
buf ( n28355 , n28354 );
buf ( n28356 , n28355 );
buf ( n28357 , n20325 );
nand ( n28358 , n28356 , n28357 );
buf ( n28359 , n28358 );
buf ( n28360 , n28359 );
nand ( n28361 , n28351 , n28360 );
buf ( n28362 , n28361 );
buf ( n28363 , n28362 );
not ( n28364 , n28363 );
buf ( n28365 , n28364 );
buf ( n28366 , n28037 );
not ( n28367 , n28366 );
buf ( n28368 , n20358 );
not ( n28369 , n28368 );
or ( n28370 , n28367 , n28369 );
buf ( n28371 , n20363 );
buf ( n28372 , n848 );
buf ( n28373 , n888 );
xor ( n28374 , n28372 , n28373 );
buf ( n28375 , n28374 );
buf ( n28376 , n28375 );
nand ( n28377 , n28371 , n28376 );
buf ( n28378 , n28377 );
buf ( n28379 , n28378 );
nand ( n28380 , n28370 , n28379 );
buf ( n28381 , n28380 );
xor ( n28382 , n28365 , n28381 );
buf ( n28383 , n28118 );
not ( n28384 , n28383 );
buf ( n28385 , n19259 );
not ( n28386 , n28385 );
or ( n28387 , n28384 , n28386 );
buf ( n28388 , n19265 );
buf ( n28389 , n858 );
buf ( n28390 , n878 );
xor ( n28391 , n28389 , n28390 );
buf ( n28392 , n28391 );
buf ( n28393 , n28392 );
nand ( n28394 , n28388 , n28393 );
buf ( n28395 , n28394 );
buf ( n28396 , n28395 );
nand ( n28397 , n28387 , n28396 );
buf ( n28398 , n28397 );
xnor ( n28399 , n28382 , n28398 );
buf ( n28400 , n28399 );
xor ( n28401 , n28346 , n28400 );
buf ( n28402 , n28401 );
buf ( n28403 , n28402 );
xor ( n28404 , n28288 , n28403 );
buf ( n28405 , n28203 );
not ( n28406 , n28405 );
buf ( n28407 , n28198 );
not ( n28408 , n28407 );
or ( n28409 , n28406 , n28408 );
buf ( n28410 , n28203 );
buf ( n28411 , n28198 );
or ( n28412 , n28410 , n28411 );
buf ( n28413 , n28257 );
nand ( n28414 , n28412 , n28413 );
buf ( n28415 , n28414 );
buf ( n28416 , n28415 );
nand ( n28417 , n28409 , n28416 );
buf ( n28418 , n28417 );
buf ( n28419 , n28418 );
buf ( n28420 , n27649 );
not ( n28421 , n28420 );
buf ( n28422 , n26534 );
not ( n28423 , n28422 );
or ( n28424 , n28421 , n28423 );
buf ( n28425 , n19910 );
buf ( n28426 , n854 );
buf ( n28427 , n882 );
xor ( n28428 , n28426 , n28427 );
buf ( n28429 , n28428 );
buf ( n28430 , n28429 );
nand ( n28431 , n28425 , n28430 );
buf ( n28432 , n28431 );
buf ( n28433 , n28432 );
nand ( n28434 , n28424 , n28433 );
buf ( n28435 , n28434 );
buf ( n28436 , n28435 );
buf ( n28437 , n863 );
buf ( n28438 , n875 );
or ( n28439 , n28437 , n28438 );
buf ( n28440 , n876 );
nand ( n28441 , n28439 , n28440 );
buf ( n28442 , n28441 );
buf ( n28443 , n28442 );
buf ( n28444 , n863 );
buf ( n28445 , n875 );
nand ( n28446 , n28444 , n28445 );
buf ( n28447 , n28446 );
buf ( n28448 , n28447 );
buf ( n28449 , n874 );
and ( n28450 , n28443 , n28448 , n28449 );
buf ( n28451 , n28450 );
buf ( n28452 , n28451 );
buf ( n28453 , n28168 );
not ( n28454 , n28453 );
buf ( n28455 , n23175 );
not ( n28456 , n28455 );
or ( n28457 , n28454 , n28456 );
buf ( n28458 , n22818 );
buf ( n28459 , n844 );
buf ( n28460 , n892 );
xor ( n28461 , n28459 , n28460 );
buf ( n28462 , n28461 );
buf ( n28463 , n28462 );
nand ( n28464 , n28458 , n28463 );
buf ( n28465 , n28464 );
buf ( n28466 , n28465 );
nand ( n28467 , n28457 , n28466 );
buf ( n28468 , n28467 );
buf ( n28469 , n28468 );
xor ( n28470 , n28452 , n28469 );
buf ( n28471 , n28470 );
buf ( n28472 , n28471 );
xor ( n28473 , n28436 , n28472 );
not ( n28474 , n28142 );
not ( n28475 , n28174 );
or ( n28476 , n28474 , n28475 );
not ( n28477 , n28180 );
not ( n28478 , n28145 );
or ( n28479 , n28477 , n28478 );
nand ( n28480 , n28479 , n28124 );
nand ( n28481 , n28476 , n28480 );
buf ( n28482 , n28481 );
xor ( n28483 , n28473 , n28482 );
buf ( n28484 , n28483 );
buf ( n28485 , n28484 );
xor ( n28486 , n28419 , n28485 );
xor ( n28487 , n28009 , n28026 );
and ( n28488 , n28487 , n28044 );
and ( n28489 , n28009 , n28026 );
or ( n28490 , n28488 , n28489 );
buf ( n28491 , n28490 );
buf ( n28492 , n28491 );
xor ( n28493 , n28064 , n28085 );
and ( n28494 , n28493 , n28104 );
and ( n28495 , n28064 , n28085 );
or ( n28496 , n28494 , n28495 );
buf ( n28497 , n28496 );
buf ( n28498 , n28497 );
xor ( n28499 , n28492 , n28498 );
buf ( n28500 , n28018 );
not ( n28501 , n28500 );
buf ( n28502 , n21297 );
not ( n28503 , n28502 );
or ( n28504 , n28501 , n28503 );
buf ( n28505 , n842 );
buf ( n28506 , n894 );
xor ( n28507 , n28505 , n28506 );
buf ( n28508 , n28507 );
buf ( n28509 , n28508 );
buf ( n28510 , n895 );
nand ( n28511 , n28509 , n28510 );
buf ( n28512 , n28511 );
buf ( n28513 , n28512 );
nand ( n28514 , n28504 , n28513 );
buf ( n28515 , n28514 );
buf ( n28516 , n28515 );
buf ( n28517 , n28057 );
not ( n28518 , n28517 );
buf ( n28519 , n21441 );
not ( n28520 , n28519 );
or ( n28521 , n28518 , n28520 );
buf ( n28522 , n20869 );
buf ( n28523 , n846 );
buf ( n28524 , n890 );
xor ( n28525 , n28523 , n28524 );
buf ( n28526 , n28525 );
buf ( n28527 , n28526 );
nand ( n28528 , n28522 , n28527 );
buf ( n28529 , n28528 );
buf ( n28530 , n28529 );
nand ( n28531 , n28521 , n28530 );
buf ( n28532 , n28531 );
buf ( n28533 , n28532 );
xor ( n28534 , n28516 , n28533 );
buf ( n28535 , n27683 );
not ( n28536 , n28535 );
buf ( n28537 , n25022 );
not ( n28538 , n28537 );
or ( n28539 , n28536 , n28538 );
buf ( n28540 , n23233 );
buf ( n28541 , n852 );
buf ( n28542 , n884 );
xor ( n28543 , n28541 , n28542 );
buf ( n28544 , n28543 );
buf ( n28545 , n28544 );
nand ( n28546 , n28540 , n28545 );
buf ( n28547 , n28546 );
buf ( n28548 , n28547 );
nand ( n28549 , n28539 , n28548 );
buf ( n28550 , n28549 );
buf ( n28551 , n28550 );
xor ( n28552 , n28534 , n28551 );
buf ( n28553 , n28552 );
buf ( n28554 , n28553 );
xor ( n28555 , n28499 , n28554 );
buf ( n28556 , n28555 );
buf ( n28557 , n28556 );
xor ( n28558 , n28486 , n28557 );
buf ( n28559 , n28558 );
buf ( n28560 , n28559 );
xor ( n28561 , n28404 , n28560 );
buf ( n28562 , n28561 );
buf ( n28563 , n28562 );
and ( n28564 , n28282 , n28563 );
and ( n28565 , n28004 , n28281 );
or ( n28566 , n28564 , n28565 );
buf ( n28567 , n28566 );
buf ( n28568 , n28567 );
buf ( n28569 , n863 );
buf ( n28570 , n879 );
or ( n28571 , n28569 , n28570 );
buf ( n28572 , n880 );
nand ( n28573 , n28571 , n28572 );
buf ( n28574 , n28573 );
buf ( n28575 , n28574 );
buf ( n28576 , n863 );
buf ( n28577 , n879 );
nand ( n28578 , n28576 , n28577 );
buf ( n28579 , n28578 );
buf ( n28580 , n28579 );
buf ( n28581 , n878 );
and ( n28582 , n28575 , n28580 , n28581 );
buf ( n28583 , n28582 );
buf ( n28584 , n28583 );
buf ( n28585 , n26471 );
not ( n28586 , n28585 );
buf ( n28587 , n22776 );
not ( n28588 , n28587 );
or ( n28589 , n28586 , n28588 );
buf ( n28590 , n27714 );
buf ( n28591 , n895 );
nand ( n28592 , n28590 , n28591 );
buf ( n28593 , n28592 );
buf ( n28594 , n28593 );
nand ( n28595 , n28589 , n28594 );
buf ( n28596 , n28595 );
buf ( n28597 , n28596 );
and ( n28598 , n28584 , n28597 );
buf ( n28599 , n28598 );
buf ( n28600 , n28599 );
not ( n28601 , n28600 );
xor ( n28602 , n882 , n858 );
buf ( n28603 , n28602 );
not ( n28604 , n28603 );
buf ( n28605 , n19580 );
not ( n28606 , n28605 );
or ( n28607 , n28604 , n28606 );
buf ( n28608 , n26538 );
buf ( n28609 , n27960 );
nand ( n28610 , n28608 , n28609 );
buf ( n28611 , n28610 );
buf ( n28612 , n28611 );
nand ( n28613 , n28607 , n28612 );
buf ( n28614 , n28613 );
not ( n28615 , n28614 );
buf ( n28616 , n28615 );
nand ( n28617 , n28601 , n28616 );
buf ( n28618 , n28617 );
buf ( n28619 , n28618 );
not ( n28620 , n28619 );
buf ( n28621 , n26433 );
not ( n28622 , n28621 );
buf ( n28623 , n23144 );
not ( n28624 , n28623 );
or ( n28625 , n28622 , n28624 );
buf ( n28626 , n27741 );
not ( n28627 , n28626 );
buf ( n28628 , n20363 );
nand ( n28629 , n28627 , n28628 );
buf ( n28630 , n28629 );
buf ( n28631 , n28630 );
nand ( n28632 , n28625 , n28631 );
buf ( n28633 , n28632 );
buf ( n28634 , n28633 );
not ( n28635 , n28634 );
buf ( n28636 , n26412 );
not ( n28637 , n28636 );
buf ( n28638 , n19614 );
not ( n28639 , n28638 );
or ( n28640 , n28637 , n28639 );
buf ( n28641 , n22271 );
buf ( n28642 , n27791 );
nand ( n28643 , n28641 , n28642 );
buf ( n28644 , n28643 );
buf ( n28645 , n28644 );
nand ( n28646 , n28640 , n28645 );
buf ( n28647 , n28646 );
buf ( n28648 , n28647 );
not ( n28649 , n28648 );
or ( n28650 , n28635 , n28649 );
buf ( n28651 , n28647 );
buf ( n28652 , n28633 );
or ( n28653 , n28651 , n28652 );
buf ( n28654 , n863 );
buf ( n28655 , n878 );
xor ( n28656 , n28654 , n28655 );
buf ( n28657 , n28656 );
buf ( n28658 , n28657 );
not ( n28659 , n28658 );
buf ( n28660 , n19479 );
not ( n28661 , n28660 );
or ( n28662 , n28659 , n28661 );
buf ( n28663 , n19265 );
buf ( n28664 , n27803 );
nand ( n28665 , n28663 , n28664 );
buf ( n28666 , n28665 );
buf ( n28667 , n28666 );
nand ( n28668 , n28662 , n28667 );
buf ( n28669 , n28668 );
buf ( n28670 , n28669 );
nand ( n28671 , n28653 , n28670 );
buf ( n28672 , n28671 );
buf ( n28673 , n28672 );
nand ( n28674 , n28650 , n28673 );
buf ( n28675 , n28674 );
buf ( n28676 , n28675 );
not ( n28677 , n28676 );
or ( n28678 , n28620 , n28677 );
buf ( n28679 , n28614 );
buf ( n28680 , n28599 );
nand ( n28681 , n28679 , n28680 );
buf ( n28682 , n28681 );
buf ( n28683 , n28682 );
nand ( n28684 , n28678 , n28683 );
buf ( n28685 , n28684 );
buf ( n28686 , n28685 );
xor ( n28687 , n27710 , n27761 );
xor ( n28688 , n28687 , n27825 );
buf ( n28689 , n28688 );
buf ( n28690 , n28689 );
xor ( n28691 , n28686 , n28690 );
buf ( n28692 , n28253 );
buf ( n28693 , n28219 );
xor ( n28694 , n28692 , n28693 );
buf ( n28695 , n28694 );
buf ( n28696 , n28695 );
buf ( n28697 , n28232 );
xor ( n28698 , n28696 , n28697 );
buf ( n28699 , n28698 );
buf ( n28700 , n28699 );
and ( n28701 , n28691 , n28700 );
and ( n28702 , n28686 , n28690 );
or ( n28703 , n28701 , n28702 );
buf ( n28704 , n28703 );
buf ( n28705 , n28704 );
buf ( n28706 , n26543 );
not ( n28707 , n28706 );
buf ( n28708 , n19580 );
not ( n28709 , n28708 );
or ( n28710 , n28707 , n28709 );
buf ( n28711 , n26538 );
buf ( n28712 , n28602 );
nand ( n28713 , n28711 , n28712 );
buf ( n28714 , n28713 );
buf ( n28715 , n28714 );
nand ( n28716 , n28710 , n28715 );
buf ( n28717 , n28716 );
buf ( n28718 , n28717 );
xor ( n28719 , n28584 , n28597 );
buf ( n28720 , n28719 );
buf ( n28721 , n28720 );
or ( n28722 , n28718 , n28721 );
buf ( n28723 , n26520 );
not ( n28724 , n28723 );
buf ( n28725 , n25022 );
not ( n28726 , n28725 );
or ( n28727 , n28724 , n28726 );
buf ( n28728 , n23233 );
buf ( n28729 , n27923 );
nand ( n28730 , n28728 , n28729 );
buf ( n28731 , n28730 );
buf ( n28732 , n28731 );
nand ( n28733 , n28727 , n28732 );
buf ( n28734 , n28733 );
buf ( n28735 , n28734 );
nand ( n28736 , n28722 , n28735 );
buf ( n28737 , n28736 );
buf ( n28738 , n28737 );
buf ( n28739 , n28720 );
buf ( n28740 , n28717 );
nand ( n28741 , n28739 , n28740 );
buf ( n28742 , n28741 );
buf ( n28743 , n28742 );
nand ( n28744 , n28738 , n28743 );
buf ( n28745 , n28744 );
buf ( n28746 , n28745 );
xor ( n28747 , n27777 , n27798 );
xor ( n28748 , n28747 , n27820 );
buf ( n28749 , n28748 );
buf ( n28750 , n28749 );
xor ( n28751 , n28746 , n28750 );
buf ( n28752 , n28599 );
buf ( n28753 , n28615 );
xor ( n28754 , n28752 , n28753 );
buf ( n28755 , n28754 );
buf ( n28756 , n28755 );
not ( n28757 , n28756 );
buf ( n28758 , n28675 );
not ( n28759 , n28758 );
or ( n28760 , n28757 , n28759 );
buf ( n28761 , n28675 );
buf ( n28762 , n28755 );
or ( n28763 , n28761 , n28762 );
nand ( n28764 , n28760 , n28763 );
buf ( n28765 , n28764 );
buf ( n28766 , n28765 );
and ( n28767 , n28751 , n28766 );
and ( n28768 , n28746 , n28750 );
or ( n28769 , n28767 , n28768 );
buf ( n28770 , n28769 );
buf ( n28771 , n28770 );
not ( n28772 , n28771 );
buf ( n28773 , n28772 );
buf ( n28774 , n28773 );
not ( n28775 , n28774 );
buf ( n28776 , n28775 );
buf ( n28777 , n28776 );
not ( n28778 , n28777 );
xor ( n28779 , n27727 , n27732 );
xor ( n28780 , n28779 , n27756 );
buf ( n28781 , n28780 );
buf ( n28782 , n28781 );
buf ( n28783 , n26454 );
not ( n28784 , n28783 );
buf ( n28785 , n23175 );
not ( n28786 , n28785 );
or ( n28787 , n28784 , n28786 );
buf ( n28788 , n22818 );
buf ( n28789 , n27763 );
nand ( n28790 , n28788 , n28789 );
buf ( n28791 , n28790 );
buf ( n28792 , n28791 );
nand ( n28793 , n28787 , n28792 );
buf ( n28794 , n28793 );
not ( n28795 , n28794 );
buf ( n28796 , n28795 );
not ( n28797 , n28796 );
buf ( n28798 , n26500 );
not ( n28799 , n28798 );
buf ( n28800 , n21441 );
not ( n28801 , n28800 );
or ( n28802 , n28799 , n28801 );
buf ( n28803 , n20869 );
buf ( n28804 , n27879 );
nand ( n28805 , n28803 , n28804 );
buf ( n28806 , n28805 );
buf ( n28807 , n28806 );
nand ( n28808 , n28802 , n28807 );
buf ( n28809 , n28808 );
buf ( n28810 , n28809 );
not ( n28811 , n28810 );
buf ( n28812 , n28811 );
buf ( n28813 , n28812 );
not ( n28814 , n28813 );
or ( n28815 , n28797 , n28814 );
buf ( n28816 , n26396 );
not ( n28817 , n28816 );
buf ( n28818 , n23027 );
not ( n28819 , n28818 );
or ( n28820 , n28817 , n28819 );
buf ( n28821 , n20525 );
buf ( n28822 , n27900 );
nand ( n28823 , n28821 , n28822 );
buf ( n28824 , n28823 );
buf ( n28825 , n28824 );
nand ( n28826 , n28820 , n28825 );
buf ( n28827 , n28826 );
buf ( n28828 , n28827 );
nand ( n28829 , n28815 , n28828 );
buf ( n28830 , n28829 );
buf ( n28831 , n28830 );
buf ( n28832 , n28809 );
not ( n28833 , n28795 );
buf ( n28834 , n28833 );
nand ( n28835 , n28832 , n28834 );
buf ( n28836 , n28835 );
buf ( n28837 , n28836 );
nand ( n28838 , n28831 , n28837 );
buf ( n28839 , n28838 );
buf ( n28840 , n28839 );
xor ( n28841 , n28782 , n28840 );
buf ( n28842 , n27939 );
not ( n28843 , n28842 );
buf ( n28844 , n28843 );
buf ( n28845 , n28844 );
not ( n28846 , n28845 );
xor ( n28847 , n27895 , n27916 );
buf ( n28848 , n28847 );
not ( n28849 , n28848 );
or ( n28850 , n28846 , n28849 );
buf ( n28851 , n28847 );
buf ( n28852 , n28844 );
or ( n28853 , n28851 , n28852 );
nand ( n28854 , n28850 , n28853 );
buf ( n28855 , n28854 );
buf ( n28856 , n28855 );
and ( n28857 , n28841 , n28856 );
and ( n28858 , n28782 , n28840 );
or ( n28859 , n28857 , n28858 );
buf ( n28860 , n28859 );
buf ( n28861 , n28860 );
not ( n28862 , n28861 );
or ( n28863 , n28778 , n28862 );
buf ( n28864 , n28860 );
buf ( n28865 , n28776 );
or ( n28866 , n28864 , n28865 );
xor ( n28867 , n27941 , n27987 );
xor ( n28868 , n28867 , n27874 );
buf ( n28869 , n28868 );
nand ( n28870 , n28866 , n28869 );
buf ( n28871 , n28870 );
buf ( n28872 , n28871 );
nand ( n28873 , n28863 , n28872 );
buf ( n28874 , n28873 );
buf ( n28875 , n28874 );
xor ( n28876 , n28705 , n28875 );
buf ( n28877 , n28187 );
not ( n28878 , n28877 );
buf ( n28879 , n28267 );
not ( n28880 , n28879 );
and ( n28881 , n28878 , n28880 );
buf ( n28882 , n28187 );
buf ( n28883 , n28267 );
and ( n28884 , n28882 , n28883 );
nor ( n28885 , n28881 , n28884 );
buf ( n28886 , n28885 );
buf ( n28887 , n28886 );
not ( n28888 , n28887 );
buf ( n28889 , n28272 );
not ( n28890 , n28889 );
or ( n28891 , n28888 , n28890 );
buf ( n28892 , n28886 );
buf ( n28893 , n28272 );
or ( n28894 , n28892 , n28893 );
nand ( n28895 , n28891 , n28894 );
buf ( n28896 , n28895 );
buf ( n28897 , n28896 );
xor ( n28898 , n28876 , n28897 );
buf ( n28899 , n28898 );
buf ( n28900 , n28899 );
xor ( n28901 , n28686 , n28690 );
xor ( n28902 , n28901 , n28700 );
buf ( n28903 , n28902 );
buf ( n28904 , n28903 );
not ( n28905 , n26478 );
nand ( n28906 , n28905 , n26476 );
not ( n28907 , n26477 );
not ( n28908 , n26481 );
or ( n28909 , n28907 , n28908 );
nand ( n28910 , n28909 , n26460 );
nand ( n28911 , n28906 , n28910 );
xor ( n28912 , n26506 , n26526 );
and ( n28913 , n28912 , n26549 );
and ( n28914 , n26506 , n26526 );
or ( n28915 , n28913 , n28914 );
xor ( n28916 , n28911 , n28915 );
buf ( n28917 , n26398 );
not ( n28918 , n28917 );
buf ( n28919 , n26418 );
not ( n28920 , n28919 );
or ( n28921 , n28918 , n28920 );
buf ( n28922 , n26398 );
buf ( n28923 , n26418 );
or ( n28924 , n28922 , n28923 );
buf ( n28925 , n26439 );
nand ( n28926 , n28924 , n28925 );
buf ( n28927 , n28926 );
buf ( n28928 , n28927 );
nand ( n28929 , n28921 , n28928 );
buf ( n28930 , n28929 );
and ( n28931 , n28916 , n28930 );
and ( n28932 , n28911 , n28915 );
or ( n28933 , n28931 , n28932 );
buf ( n28934 , n28933 );
xor ( n28935 , n28782 , n28840 );
xor ( n28936 , n28935 , n28856 );
buf ( n28937 , n28936 );
buf ( n28938 , n28937 );
xor ( n28939 , n28934 , n28938 );
buf ( n28940 , n28734 );
not ( n28941 , n28940 );
xor ( n28942 , n28717 , n28720 );
not ( n28943 , n28942 );
or ( n28944 , n28941 , n28943 );
or ( n28945 , n28942 , n28940 );
nand ( n28946 , n28944 , n28945 );
buf ( n28947 , n28946 );
not ( n28948 , n28947 );
xor ( n28949 , n28647 , n28633 );
xnor ( n28950 , n28949 , n28669 );
buf ( n28951 , n28950 );
not ( n28952 , n28951 );
or ( n28953 , n28948 , n28952 );
xor ( n28954 , n28812 , n28827 );
xnor ( n28955 , n28954 , n28833 );
buf ( n28956 , n28955 );
nand ( n28957 , n28953 , n28956 );
buf ( n28958 , n28957 );
buf ( n28959 , n28958 );
buf ( n28960 , n28950 );
not ( n28961 , n28960 );
not ( n28962 , n28946 );
buf ( n28963 , n28962 );
nand ( n28964 , n28961 , n28963 );
buf ( n28965 , n28964 );
buf ( n28966 , n28965 );
nand ( n28967 , n28959 , n28966 );
buf ( n28968 , n28967 );
buf ( n28969 , n28968 );
and ( n28970 , n28939 , n28969 );
and ( n28971 , n28934 , n28938 );
or ( n28972 , n28970 , n28971 );
buf ( n28973 , n28972 );
buf ( n28974 , n28973 );
xor ( n28975 , n28904 , n28974 );
xor ( n28976 , n28773 , n28860 );
buf ( n28977 , n28868 );
not ( n28978 , n28977 );
buf ( n28979 , n28978 );
and ( n28980 , n28976 , n28979 );
not ( n28981 , n28976 );
and ( n28982 , n28981 , n28868 );
nor ( n28983 , n28980 , n28982 );
buf ( n28984 , n28983 );
and ( n28985 , n28975 , n28984 );
and ( n28986 , n28904 , n28974 );
or ( n28987 , n28985 , n28986 );
buf ( n28988 , n28987 );
buf ( n28989 , n28988 );
buf ( n28990 , n23238 );
not ( n28991 , n28990 );
buf ( n28992 , n22776 );
not ( n28993 , n28992 );
or ( n28994 , n28991 , n28993 );
buf ( n28995 , n862 );
buf ( n28996 , n894 );
xor ( n28997 , n28995 , n28996 );
buf ( n28998 , n28997 );
buf ( n28999 , n28998 );
buf ( n29000 , n895 );
nand ( n29001 , n28999 , n29000 );
buf ( n29002 , n29001 );
buf ( n29003 , n29002 );
nand ( n29004 , n28994 , n29003 );
buf ( n29005 , n29004 );
buf ( n29006 , n29005 );
buf ( n29007 , n9989 );
xor ( n29008 , n866 , n839 );
buf ( n29009 , n29008 );
not ( n29010 , n29009 );
buf ( n29011 , n18931 );
not ( n29012 , n29011 );
or ( n29013 , n29010 , n29012 );
buf ( n29014 , n18944 );
buf ( n29015 , n838 );
buf ( n29016 , n866 );
xor ( n29017 , n29015 , n29016 );
buf ( n29018 , n29017 );
buf ( n29019 , n29018 );
nand ( n29020 , n29014 , n29019 );
buf ( n29021 , n29020 );
buf ( n29022 , n29021 );
nand ( n29023 , n29013 , n29022 );
buf ( n29024 , n29023 );
buf ( n29025 , n29024 );
buf ( n29026 , n835 );
buf ( n29027 , n870 );
xor ( n29028 , n29026 , n29027 );
buf ( n29029 , n29028 );
buf ( n29030 , n29029 );
not ( n29031 , n29030 );
buf ( n29032 , n19125 );
not ( n29033 , n29032 );
or ( n29034 , n29031 , n29033 );
buf ( n29035 , n19134 );
buf ( n29036 , n834 );
buf ( n29037 , n870 );
xor ( n29038 , n29036 , n29037 );
buf ( n29039 , n29038 );
buf ( n29040 , n29039 );
nand ( n29041 , n29035 , n29040 );
buf ( n29042 , n29041 );
buf ( n29043 , n29042 );
nand ( n29044 , n29034 , n29043 );
buf ( n29045 , n29044 );
buf ( n29046 , n29045 );
xor ( n29047 , n29025 , n29046 );
buf ( n29048 , n864 );
buf ( n29049 , n841 );
xor ( n29050 , n29048 , n29049 );
buf ( n29051 , n29050 );
buf ( n29052 , n29051 );
not ( n29053 , n29052 );
buf ( n29054 , n19330 );
not ( n29055 , n29054 );
or ( n29056 , n29053 , n29055 );
buf ( n29057 , n19030 );
buf ( n29058 , n864 );
buf ( n29059 , n840 );
xor ( n29060 , n29058 , n29059 );
buf ( n29061 , n29060 );
buf ( n29062 , n29061 );
nand ( n29063 , n29057 , n29062 );
buf ( n29064 , n29063 );
buf ( n29065 , n29064 );
nand ( n29066 , n29056 , n29065 );
buf ( n29067 , n29066 );
buf ( n29068 , n29067 );
and ( n29069 , n29047 , n29068 );
and ( n29070 , n29025 , n29046 );
or ( n29071 , n29069 , n29070 );
buf ( n29072 , n29071 );
buf ( n29073 , n29072 );
xor ( n29074 , n868 , n837 );
buf ( n29075 , n29074 );
not ( n29076 , n29075 );
buf ( n29077 , n18887 );
not ( n29078 , n29077 );
or ( n29079 , n29076 , n29078 );
buf ( n29080 , n18898 );
buf ( n29081 , n836 );
buf ( n29082 , n868 );
xor ( n29083 , n29081 , n29082 );
buf ( n29084 , n29083 );
buf ( n29085 , n29084 );
nand ( n29086 , n29080 , n29085 );
buf ( n29087 , n29086 );
buf ( n29088 , n29087 );
nand ( n29089 , n29079 , n29088 );
buf ( n29090 , n29089 );
buf ( n29091 , n29090 );
buf ( n29092 , n18984 );
not ( n29093 , n29092 );
buf ( n29094 , n18977 );
not ( n29095 , n29094 );
buf ( n29096 , n29095 );
buf ( n29097 , n29096 );
not ( n29098 , n29097 );
or ( n29099 , n29093 , n29098 );
buf ( n29100 , n874 );
nand ( n29101 , n29099 , n29100 );
buf ( n29102 , n29101 );
buf ( n29103 , n29102 );
xor ( n29104 , n29091 , n29103 );
buf ( n29105 , n833 );
buf ( n29106 , n872 );
xor ( n29107 , n29105 , n29106 );
buf ( n29108 , n29107 );
buf ( n29109 , n29108 );
not ( n29110 , n29109 );
buf ( n29111 , n19230 );
not ( n29112 , n29111 );
or ( n29113 , n29110 , n29112 );
buf ( n29114 , n19235 );
buf ( n29115 , n832 );
buf ( n29116 , n872 );
xor ( n29117 , n29115 , n29116 );
buf ( n29118 , n29117 );
buf ( n29119 , n29118 );
nand ( n29120 , n29114 , n29119 );
buf ( n29121 , n29120 );
buf ( n29122 , n29121 );
nand ( n29123 , n29113 , n29122 );
buf ( n29124 , n29123 );
buf ( n29125 , n29124 );
and ( n29126 , n29104 , n29125 );
and ( n29127 , n29091 , n29103 );
or ( n29128 , n29126 , n29127 );
buf ( n29129 , n29128 );
buf ( n29130 , n29129 );
xor ( n29131 , n29073 , n29130 );
buf ( n29132 , n29018 );
not ( n29133 , n29132 );
buf ( n29134 , n18931 );
not ( n29135 , n29134 );
buf ( n29136 , n29135 );
buf ( n29137 , n29136 );
not ( n29138 , n29137 );
buf ( n29139 , n29138 );
buf ( n29140 , n29139 );
not ( n29141 , n29140 );
or ( n29142 , n29133 , n29141 );
buf ( n29143 , n18944 );
buf ( n29144 , n837 );
buf ( n29145 , n866 );
xor ( n29146 , n29144 , n29145 );
buf ( n29147 , n29146 );
buf ( n29148 , n29147 );
nand ( n29149 , n29143 , n29148 );
buf ( n29150 , n29149 );
buf ( n29151 , n29150 );
nand ( n29152 , n29142 , n29151 );
buf ( n29153 , n29152 );
buf ( n29154 , n29118 );
not ( n29155 , n29154 );
buf ( n29156 , n19230 );
not ( n29157 , n29156 );
or ( n29158 , n29155 , n29157 );
buf ( n29159 , n19234 );
buf ( n29160 , n872 );
nand ( n29161 , n29159 , n29160 );
buf ( n29162 , n29161 );
buf ( n29163 , n29162 );
nand ( n29164 , n29158 , n29163 );
buf ( n29165 , n29164 );
xnor ( n29166 , n29153 , n29165 );
buf ( n29167 , n29166 );
buf ( n29168 , n29061 );
not ( n29169 , n29168 );
buf ( n29170 , n19330 );
not ( n29171 , n29170 );
or ( n29172 , n29169 , n29171 );
buf ( n29173 , n19030 );
buf ( n29174 , n864 );
buf ( n29175 , n839 );
xor ( n29176 , n29174 , n29175 );
buf ( n29177 , n29176 );
buf ( n29178 , n29177 );
nand ( n29179 , n29173 , n29178 );
buf ( n29180 , n29179 );
buf ( n29181 , n29180 );
nand ( n29182 , n29172 , n29181 );
buf ( n29183 , n29182 );
buf ( n29184 , n29183 );
xnor ( n29185 , n29167 , n29184 );
buf ( n29186 , n29185 );
buf ( n29187 , n29186 );
xor ( n29188 , n29131 , n29187 );
buf ( n29189 , n29188 );
buf ( n29190 , n29189 );
and ( n29191 , n29048 , n29049 );
buf ( n29192 , n29191 );
buf ( n29193 , n29192 );
buf ( n29194 , n29084 );
not ( n29195 , n29194 );
buf ( n29196 , n18887 );
not ( n29197 , n29196 );
or ( n29198 , n29195 , n29197 );
buf ( n29199 , n18898 );
buf ( n29200 , n835 );
buf ( n29201 , n868 );
xor ( n29202 , n29200 , n29201 );
buf ( n29203 , n29202 );
buf ( n29204 , n29203 );
nand ( n29205 , n29199 , n29204 );
buf ( n29206 , n29205 );
buf ( n29207 , n29206 );
nand ( n29208 , n29198 , n29207 );
buf ( n29209 , n29208 );
buf ( n29210 , n29209 );
xor ( n29211 , n29193 , n29210 );
buf ( n29212 , n29039 );
not ( n29213 , n29212 );
buf ( n29214 , n19125 );
not ( n29215 , n29214 );
or ( n29216 , n29213 , n29215 );
buf ( n29217 , n19134 );
buf ( n29218 , n870 );
buf ( n29219 , n833 );
xor ( n29220 , n29218 , n29219 );
buf ( n29221 , n29220 );
buf ( n29222 , n29221 );
nand ( n29223 , n29217 , n29222 );
buf ( n29224 , n29223 );
buf ( n29225 , n29224 );
nand ( n29226 , n29216 , n29225 );
buf ( n29227 , n29226 );
buf ( n29228 , n29227 );
not ( n29229 , n29228 );
buf ( n29230 , n29229 );
buf ( n29231 , n29230 );
xor ( n29232 , n29211 , n29231 );
buf ( n29233 , n29232 );
buf ( n29234 , n29233 );
buf ( n29235 , n864 );
buf ( n29236 , n842 );
and ( n29237 , n29235 , n29236 );
buf ( n29238 , n29237 );
buf ( n29239 , n29238 );
buf ( n29240 , n832 );
buf ( n29241 , n874 );
xor ( n29242 , n29240 , n29241 );
buf ( n29243 , n29242 );
buf ( n29244 , n29243 );
not ( n29245 , n29244 );
buf ( n29246 , n18977 );
not ( n29247 , n29246 );
or ( n29248 , n29245 , n29247 );
buf ( n29249 , n18987 );
buf ( n29250 , n874 );
nand ( n29251 , n29249 , n29250 );
buf ( n29252 , n29251 );
buf ( n29253 , n29252 );
nand ( n29254 , n29248 , n29253 );
buf ( n29255 , n29254 );
buf ( n29256 , n29255 );
xor ( n29257 , n29239 , n29256 );
xor ( n29258 , n866 , n840 );
buf ( n29259 , n29258 );
not ( n29260 , n29259 );
buf ( n29261 , n18931 );
not ( n29262 , n29261 );
or ( n29263 , n29260 , n29262 );
buf ( n29264 , n18944 );
buf ( n29265 , n29008 );
nand ( n29266 , n29264 , n29265 );
buf ( n29267 , n29266 );
buf ( n29268 , n29267 );
nand ( n29269 , n29263 , n29268 );
buf ( n29270 , n29269 );
buf ( n29271 , n29270 );
xor ( n29272 , n868 , n838 );
buf ( n29273 , n29272 );
not ( n29274 , n29273 );
buf ( n29275 , n18887 );
not ( n29276 , n29275 );
or ( n29277 , n29274 , n29276 );
buf ( n29278 , n18898 );
buf ( n29279 , n29074 );
nand ( n29280 , n29278 , n29279 );
buf ( n29281 , n29280 );
buf ( n29282 , n29281 );
nand ( n29283 , n29277 , n29282 );
buf ( n29284 , n29283 );
buf ( n29285 , n29284 );
nand ( n29286 , n29271 , n29285 );
buf ( n29287 , n29286 );
buf ( n29288 , n29287 );
buf ( n29289 , n29270 );
buf ( n29290 , n29284 );
or ( n29291 , n29289 , n29290 );
buf ( n29292 , n834 );
buf ( n29293 , n872 );
xor ( n29294 , n29292 , n29293 );
buf ( n29295 , n29294 );
buf ( n29296 , n29295 );
not ( n29297 , n29296 );
buf ( n29298 , n19230 );
not ( n29299 , n29298 );
or ( n29300 , n29297 , n29299 );
buf ( n29301 , n19235 );
buf ( n29302 , n29108 );
nand ( n29303 , n29301 , n29302 );
buf ( n29304 , n29303 );
buf ( n29305 , n29304 );
nand ( n29306 , n29300 , n29305 );
buf ( n29307 , n29306 );
buf ( n29308 , n29307 );
nand ( n29309 , n29291 , n29308 );
buf ( n29310 , n29309 );
buf ( n29311 , n29310 );
nand ( n29312 , n29288 , n29311 );
buf ( n29313 , n29312 );
buf ( n29314 , n29313 );
and ( n29315 , n29257 , n29314 );
and ( n29316 , n29239 , n29256 );
or ( n29317 , n29315 , n29316 );
buf ( n29318 , n29317 );
buf ( n29319 , n29318 );
xor ( n29320 , n29234 , n29319 );
buf ( n29321 , n843 );
buf ( n29322 , n864 );
and ( n29323 , n29321 , n29322 );
buf ( n29324 , n29323 );
buf ( n29325 , n29324 );
xor ( n29326 , n29235 , n29236 );
buf ( n29327 , n29326 );
buf ( n29328 , n29327 );
not ( n29329 , n29328 );
buf ( n29330 , n19330 );
not ( n29331 , n29330 );
or ( n29332 , n29329 , n29331 );
buf ( n29333 , n19030 );
buf ( n29334 , n29051 );
nand ( n29335 , n29333 , n29334 );
buf ( n29336 , n29335 );
buf ( n29337 , n29336 );
nand ( n29338 , n29332 , n29337 );
buf ( n29339 , n29338 );
buf ( n29340 , n29339 );
xor ( n29341 , n29325 , n29340 );
buf ( n29342 , n836 );
buf ( n29343 , n870 );
xor ( n29344 , n29342 , n29343 );
buf ( n29345 , n29344 );
buf ( n29346 , n29345 );
not ( n29347 , n29346 );
buf ( n29348 , n19125 );
not ( n29349 , n29348 );
or ( n29350 , n29347 , n29349 );
buf ( n29351 , n19134 );
buf ( n29352 , n29029 );
nand ( n29353 , n29351 , n29352 );
buf ( n29354 , n29353 );
buf ( n29355 , n29354 );
nand ( n29356 , n29350 , n29355 );
buf ( n29357 , n29356 );
buf ( n29358 , n29357 );
and ( n29359 , n29341 , n29358 );
and ( n29360 , n29325 , n29340 );
or ( n29361 , n29359 , n29360 );
buf ( n29362 , n29361 );
buf ( n29363 , n29362 );
xor ( n29364 , n29091 , n29103 );
xor ( n29365 , n29364 , n29125 );
buf ( n29366 , n29365 );
buf ( n29367 , n29366 );
xor ( n29368 , n29363 , n29367 );
xor ( n29369 , n29025 , n29046 );
xor ( n29370 , n29369 , n29068 );
buf ( n29371 , n29370 );
buf ( n29372 , n29371 );
and ( n29373 , n29368 , n29372 );
and ( n29374 , n29363 , n29367 );
or ( n29375 , n29373 , n29374 );
buf ( n29376 , n29375 );
buf ( n29377 , n29376 );
xor ( n29378 , n29320 , n29377 );
buf ( n29379 , n29378 );
buf ( n29380 , n29379 );
xor ( n29381 , n29190 , n29380 );
xor ( n29382 , n29239 , n29256 );
xor ( n29383 , n29382 , n29314 );
buf ( n29384 , n29383 );
buf ( n29385 , n29384 );
buf ( n29386 , n29255 );
not ( n29387 , n29386 );
buf ( n29388 , n29387 );
buf ( n29389 , n29388 );
buf ( n29390 , n839 );
buf ( n29391 , n868 );
xor ( n29392 , n29390 , n29391 );
buf ( n29393 , n29392 );
buf ( n29394 , n29393 );
not ( n29395 , n29394 );
buf ( n29396 , n18887 );
not ( n29397 , n29396 );
or ( n29398 , n29395 , n29397 );
buf ( n29399 , n18898 );
buf ( n29400 , n29272 );
nand ( n29401 , n29399 , n29400 );
buf ( n29402 , n29401 );
buf ( n29403 , n29402 );
nand ( n29404 , n29398 , n29403 );
buf ( n29405 , n29404 );
buf ( n29406 , n29405 );
and ( n29407 , n26234 , n26235 );
buf ( n29408 , n29407 );
buf ( n29409 , n29408 );
or ( n29410 , n29406 , n29409 );
buf ( n29411 , n835 );
buf ( n29412 , n872 );
xor ( n29413 , n29411 , n29412 );
buf ( n29414 , n29413 );
buf ( n29415 , n29414 );
not ( n29416 , n29415 );
buf ( n29417 , n19230 );
not ( n29418 , n29417 );
or ( n29419 , n29416 , n29418 );
buf ( n29420 , n19235 );
buf ( n29421 , n29295 );
nand ( n29422 , n29420 , n29421 );
buf ( n29423 , n29422 );
buf ( n29424 , n29423 );
nand ( n29425 , n29419 , n29424 );
buf ( n29426 , n29425 );
buf ( n29427 , n29426 );
nand ( n29428 , n29410 , n29427 );
buf ( n29429 , n29428 );
buf ( n29430 , n29429 );
buf ( n29431 , n29405 );
buf ( n29432 , n29408 );
nand ( n29433 , n29431 , n29432 );
buf ( n29434 , n29433 );
buf ( n29435 , n29434 );
nand ( n29436 , n29430 , n29435 );
buf ( n29437 , n29436 );
buf ( n29438 , n29437 );
xor ( n29439 , n29389 , n29438 );
buf ( n29440 , n837 );
buf ( n29441 , n870 );
xor ( n29442 , n29440 , n29441 );
buf ( n29443 , n29442 );
buf ( n29444 , n29443 );
not ( n29445 , n29444 );
buf ( n29446 , n19125 );
not ( n29447 , n29446 );
or ( n29448 , n29445 , n29447 );
buf ( n29449 , n19134 );
buf ( n29450 , n29345 );
nand ( n29451 , n29449 , n29450 );
buf ( n29452 , n29451 );
buf ( n29453 , n29452 );
nand ( n29454 , n29448 , n29453 );
buf ( n29455 , n29454 );
buf ( n29456 , n29455 );
or ( n29457 , n19085 , n19153 );
nand ( n29458 , n29457 , n876 );
buf ( n29459 , n29458 );
xor ( n29460 , n29456 , n29459 );
buf ( n29461 , n833 );
buf ( n29462 , n874 );
xor ( n29463 , n29461 , n29462 );
buf ( n29464 , n29463 );
buf ( n29465 , n29464 );
not ( n29466 , n29465 );
buf ( n29467 , n18977 );
not ( n29468 , n29467 );
or ( n29469 , n29466 , n29468 );
buf ( n29470 , n18987 );
buf ( n29471 , n29243 );
nand ( n29472 , n29470 , n29471 );
buf ( n29473 , n29472 );
buf ( n29474 , n29473 );
nand ( n29475 , n29469 , n29474 );
buf ( n29476 , n29475 );
buf ( n29477 , n29476 );
and ( n29478 , n29460 , n29477 );
and ( n29479 , n29456 , n29459 );
or ( n29480 , n29478 , n29479 );
buf ( n29481 , n29480 );
buf ( n29482 , n29481 );
and ( n29483 , n29439 , n29482 );
and ( n29484 , n29389 , n29438 );
or ( n29485 , n29483 , n29484 );
buf ( n29486 , n29485 );
buf ( n29487 , n29486 );
xor ( n29488 , n29385 , n29487 );
buf ( n29489 , n843 );
buf ( n29490 , n864 );
xor ( n29491 , n29489 , n29490 );
buf ( n29492 , n29491 );
buf ( n29493 , n29492 );
not ( n29494 , n29493 );
buf ( n29495 , n19330 );
not ( n29496 , n29495 );
or ( n29497 , n29494 , n29496 );
buf ( n29498 , n19030 );
buf ( n29499 , n29327 );
nand ( n29500 , n29498 , n29499 );
buf ( n29501 , n29500 );
buf ( n29502 , n29501 );
nand ( n29503 , n29497 , n29502 );
buf ( n29504 , n29503 );
buf ( n29505 , n29504 );
buf ( n29506 , n841 );
buf ( n29507 , n866 );
xor ( n29508 , n29506 , n29507 );
buf ( n29509 , n29508 );
buf ( n29510 , n29509 );
not ( n29511 , n29510 );
buf ( n29512 , n18931 );
not ( n29513 , n29512 );
or ( n29514 , n29511 , n29513 );
buf ( n29515 , n18944 );
buf ( n29516 , n29258 );
nand ( n29517 , n29515 , n29516 );
buf ( n29518 , n29517 );
buf ( n29519 , n29518 );
nand ( n29520 , n29514 , n29519 );
buf ( n29521 , n29520 );
buf ( n29522 , n29521 );
or ( n29523 , n29505 , n29522 );
buf ( n29524 , n26341 );
not ( n29525 , n29524 );
buf ( n29526 , n19153 );
not ( n29527 , n29526 );
or ( n29528 , n29525 , n29527 );
buf ( n29529 , n19085 );
buf ( n29530 , n876 );
nand ( n29531 , n29529 , n29530 );
buf ( n29532 , n29531 );
buf ( n29533 , n29532 );
nand ( n29534 , n29528 , n29533 );
buf ( n29535 , n29534 );
buf ( n29536 , n29535 );
nand ( n29537 , n29523 , n29536 );
buf ( n29538 , n29537 );
buf ( n29539 , n29538 );
buf ( n29540 , n29504 );
buf ( n29541 , n29521 );
nand ( n29542 , n29540 , n29541 );
buf ( n29543 , n29542 );
buf ( n29544 , n29543 );
nand ( n29545 , n29539 , n29544 );
buf ( n29546 , n29545 );
buf ( n29547 , n29546 );
xor ( n29548 , n29325 , n29340 );
xor ( n29549 , n29548 , n29358 );
buf ( n29550 , n29549 );
buf ( n29551 , n29550 );
xor ( n29552 , n29547 , n29551 );
xor ( n29553 , n29270 , n29307 );
buf ( n29554 , n29553 );
buf ( n29555 , n29284 );
xor ( n29556 , n29554 , n29555 );
buf ( n29557 , n29556 );
buf ( n29558 , n29557 );
and ( n29559 , n29552 , n29558 );
and ( n29560 , n29547 , n29551 );
or ( n29561 , n29559 , n29560 );
buf ( n29562 , n29561 );
buf ( n29563 , n29562 );
and ( n29564 , n29488 , n29563 );
and ( n29565 , n29385 , n29487 );
or ( n29566 , n29564 , n29565 );
buf ( n29567 , n29566 );
buf ( n29568 , n29567 );
xor ( n29569 , n29381 , n29568 );
buf ( n29570 , n29569 );
buf ( n29571 , n29570 );
and ( n29572 , n28452 , n28469 );
buf ( n29573 , n29572 );
buf ( n29574 , n29573 );
buf ( n29575 , n28312 );
not ( n29576 , n29575 );
buf ( n29577 , n28324 );
not ( n29578 , n29577 );
or ( n29579 , n29576 , n29578 );
buf ( n29580 , n28315 );
not ( n29581 , n29580 );
buf ( n29582 , n28324 );
not ( n29583 , n29582 );
buf ( n29584 , n29583 );
buf ( n29585 , n29584 );
not ( n29586 , n29585 );
or ( n29587 , n29581 , n29586 );
buf ( n29588 , n28342 );
nand ( n29589 , n29587 , n29588 );
buf ( n29590 , n29589 );
buf ( n29591 , n29590 );
nand ( n29592 , n29579 , n29591 );
buf ( n29593 , n29592 );
buf ( n29594 , n29593 );
xor ( n29595 , n29574 , n29594 );
xor ( n29596 , n28516 , n28533 );
and ( n29597 , n29596 , n28551 );
and ( n29598 , n28516 , n28533 );
or ( n29599 , n29597 , n29598 );
buf ( n29600 , n29599 );
buf ( n29601 , n29600 );
xor ( n29602 , n29595 , n29601 );
buf ( n29603 , n29602 );
buf ( n29604 , n29603 );
xor ( n29605 , n28492 , n28498 );
and ( n29606 , n29605 , n28554 );
and ( n29607 , n28492 , n28498 );
or ( n29608 , n29606 , n29607 );
buf ( n29609 , n29608 );
buf ( n29610 , n29609 );
xor ( n29611 , n29604 , n29610 );
xor ( n29612 , n28296 , n28345 );
and ( n29613 , n29612 , n28400 );
and ( n29614 , n28296 , n28345 );
or ( n29615 , n29613 , n29614 );
buf ( n29616 , n29615 );
buf ( n29617 , n29616 );
xor ( n29618 , n29611 , n29617 );
buf ( n29619 , n29618 );
buf ( n29620 , n29619 );
buf ( n29621 , n28365 );
not ( n29622 , n29621 );
buf ( n29623 , n28381 );
not ( n29624 , n29623 );
buf ( n29625 , n29624 );
buf ( n29626 , n29625 );
not ( n29627 , n29626 );
or ( n29628 , n29622 , n29627 );
buf ( n29629 , n28398 );
nand ( n29630 , n29628 , n29629 );
buf ( n29631 , n29630 );
buf ( n29632 , n29631 );
buf ( n29633 , n28381 );
buf ( n29634 , n28362 );
nand ( n29635 , n29633 , n29634 );
buf ( n29636 , n29635 );
buf ( n29637 , n29636 );
nand ( n29638 , n29632 , n29637 );
buf ( n29639 , n29638 );
buf ( n29640 , n29639 );
buf ( n29641 , n28526 );
not ( n29642 , n29641 );
buf ( n29643 , n21441 );
not ( n29644 , n29643 );
or ( n29645 , n29642 , n29644 );
buf ( n29646 , n20869 );
buf ( n29647 , n845 );
buf ( n29648 , n890 );
xor ( n29649 , n29647 , n29648 );
buf ( n29650 , n29649 );
buf ( n29651 , n29650 );
nand ( n29652 , n29646 , n29651 );
buf ( n29653 , n29652 );
buf ( n29654 , n29653 );
nand ( n29655 , n29645 , n29654 );
buf ( n29656 , n29655 );
buf ( n29657 , n29656 );
buf ( n29658 , n28544 );
not ( n29659 , n29658 );
buf ( n29660 , n20694 );
not ( n29661 , n29660 );
or ( n29662 , n29659 , n29661 );
buf ( n29663 , n20700 );
buf ( n29664 , n851 );
buf ( n29665 , n884 );
xor ( n29666 , n29664 , n29665 );
buf ( n29667 , n29666 );
buf ( n29668 , n29667 );
nand ( n29669 , n29663 , n29668 );
buf ( n29670 , n29669 );
buf ( n29671 , n29670 );
nand ( n29672 , n29662 , n29671 );
buf ( n29673 , n29672 );
buf ( n29674 , n29673 );
xor ( n29675 , n29657 , n29674 );
buf ( n29676 , n28429 );
not ( n29677 , n29676 );
buf ( n29678 , n19580 );
not ( n29679 , n29678 );
or ( n29680 , n29677 , n29679 );
buf ( n29681 , n19910 );
buf ( n29682 , n853 );
buf ( n29683 , n882 );
xor ( n29684 , n29682 , n29683 );
buf ( n29685 , n29684 );
buf ( n29686 , n29685 );
nand ( n29687 , n29681 , n29686 );
buf ( n29688 , n29687 );
buf ( n29689 , n29688 );
nand ( n29690 , n29680 , n29689 );
buf ( n29691 , n29690 );
buf ( n29692 , n29691 );
xor ( n29693 , n29675 , n29692 );
buf ( n29694 , n29693 );
buf ( n29695 , n29694 );
xor ( n29696 , n29640 , n29695 );
buf ( n29697 , n28322 );
not ( n29698 , n29697 );
buf ( n29699 , n21817 );
not ( n29700 , n29699 );
or ( n29701 , n29698 , n29700 );
buf ( n29702 , n20525 );
buf ( n29703 , n849 );
buf ( n29704 , n886 );
xor ( n29705 , n29703 , n29704 );
buf ( n29706 , n29705 );
buf ( n29707 , n29706 );
nand ( n29708 , n29702 , n29707 );
buf ( n29709 , n29708 );
buf ( n29710 , n29709 );
nand ( n29711 , n29701 , n29710 );
buf ( n29712 , n29711 );
not ( n29713 , n28355 );
not ( n29714 , n18850 );
or ( n29715 , n29713 , n29714 );
buf ( n29716 , n20325 );
buf ( n29717 , n855 );
buf ( n29718 , n880 );
xor ( n29719 , n29717 , n29718 );
buf ( n29720 , n29719 );
buf ( n29721 , n29720 );
nand ( n29722 , n29716 , n29721 );
buf ( n29723 , n29722 );
nand ( n29724 , n29715 , n29723 );
xor ( n29725 , n29712 , n29724 );
buf ( n29726 , n28392 );
not ( n29727 , n29726 );
buf ( n29728 , n19259 );
not ( n29729 , n29728 );
or ( n29730 , n29727 , n29729 );
buf ( n29731 , n19265 );
buf ( n29732 , n857 );
buf ( n29733 , n878 );
xor ( n29734 , n29732 , n29733 );
buf ( n29735 , n29734 );
buf ( n29736 , n29735 );
nand ( n29737 , n29731 , n29736 );
buf ( n29738 , n29737 );
buf ( n29739 , n29738 );
nand ( n29740 , n29730 , n29739 );
buf ( n29741 , n29740 );
xor ( n29742 , n29725 , n29741 );
buf ( n29743 , n29742 );
xor ( n29744 , n29696 , n29743 );
buf ( n29745 , n29744 );
buf ( n29746 , n29745 );
and ( n29747 , n19221 , n863 );
buf ( n29748 , n29747 );
buf ( n29749 , n28375 );
not ( n29750 , n29749 );
buf ( n29751 , n20358 );
not ( n29752 , n29751 );
or ( n29753 , n29750 , n29752 );
buf ( n29754 , n847 );
buf ( n29755 , n888 );
xor ( n29756 , n29754 , n29755 );
buf ( n29757 , n29756 );
buf ( n29758 , n29757 );
buf ( n29759 , n20363 );
nand ( n29760 , n29758 , n29759 );
buf ( n29761 , n29760 );
buf ( n29762 , n29761 );
nand ( n29763 , n29753 , n29762 );
buf ( n29764 , n29763 );
buf ( n29765 , n29764 );
xor ( n29766 , n29748 , n29765 );
buf ( n29767 , n28462 );
not ( n29768 , n29767 );
buf ( n29769 , n20599 );
not ( n29770 , n29769 );
or ( n29771 , n29768 , n29770 );
buf ( n29772 , n22818 );
buf ( n29773 , n843 );
buf ( n29774 , n892 );
xor ( n29775 , n29773 , n29774 );
buf ( n29776 , n29775 );
buf ( n29777 , n29776 );
nand ( n29778 , n29772 , n29777 );
buf ( n29779 , n29778 );
buf ( n29780 , n29779 );
nand ( n29781 , n29771 , n29780 );
buf ( n29782 , n29781 );
buf ( n29783 , n29782 );
xor ( n29784 , n29766 , n29783 );
buf ( n29785 , n29784 );
buf ( n29786 , n29785 );
buf ( n29787 , n28508 );
not ( n29788 , n29787 );
buf ( n29789 , n22776 );
not ( n29790 , n29789 );
or ( n29791 , n29788 , n29790 );
buf ( n29792 , n841 );
buf ( n29793 , n894 );
xor ( n29794 , n29792 , n29793 );
buf ( n29795 , n29794 );
buf ( n29796 , n29795 );
buf ( n29797 , n895 );
nand ( n29798 , n29796 , n29797 );
buf ( n29799 , n29798 );
buf ( n29800 , n29799 );
nand ( n29801 , n29791 , n29800 );
buf ( n29802 , n29801 );
buf ( n29803 , n29802 );
buf ( n29804 , n28306 );
not ( n29805 , n29804 );
buf ( n29806 , n19153 );
not ( n29807 , n29806 );
or ( n29808 , n29805 , n29807 );
buf ( n29809 , n20246 );
buf ( n29810 , n859 );
buf ( n29811 , n876 );
xor ( n29812 , n29810 , n29811 );
buf ( n29813 , n29812 );
buf ( n29814 , n29813 );
nand ( n29815 , n29809 , n29814 );
buf ( n29816 , n29815 );
buf ( n29817 , n29816 );
nand ( n29818 , n29808 , n29817 );
buf ( n29819 , n29818 );
buf ( n29820 , n29819 );
xor ( n29821 , n29803 , n29820 );
buf ( n29822 , n28336 );
not ( n29823 , n29822 );
buf ( n29824 , n18974 );
not ( n29825 , n29824 );
or ( n29826 , n29823 , n29825 );
buf ( n29827 , n20555 );
buf ( n29828 , n861 );
buf ( n29829 , n874 );
xor ( n29830 , n29828 , n29829 );
buf ( n29831 , n29830 );
buf ( n29832 , n29831 );
nand ( n29833 , n29827 , n29832 );
buf ( n29834 , n29833 );
buf ( n29835 , n29834 );
nand ( n29836 , n29826 , n29835 );
buf ( n29837 , n29836 );
buf ( n29838 , n29837 );
xor ( n29839 , n29821 , n29838 );
buf ( n29840 , n29839 );
buf ( n29841 , n29840 );
xor ( n29842 , n29786 , n29841 );
xor ( n29843 , n28436 , n28472 );
and ( n29844 , n29843 , n28482 );
and ( n29845 , n28436 , n28472 );
or ( n29846 , n29844 , n29845 );
buf ( n29847 , n29846 );
buf ( n29848 , n29847 );
xor ( n29849 , n29842 , n29848 );
buf ( n29850 , n29849 );
buf ( n29851 , n29850 );
xor ( n29852 , n29746 , n29851 );
xor ( n29853 , n28419 , n28485 );
and ( n29854 , n29853 , n28557 );
and ( n29855 , n28419 , n28485 );
or ( n29856 , n29854 , n29855 );
buf ( n29857 , n29856 );
buf ( n29858 , n29857 );
xor ( n29859 , n29852 , n29858 );
buf ( n29860 , n29859 );
buf ( n29861 , n29860 );
xor ( n29862 , n29620 , n29861 );
xor ( n29863 , n28288 , n28403 );
and ( n29864 , n29863 , n28560 );
and ( n29865 , n28288 , n28403 );
or ( n29866 , n29864 , n29865 );
buf ( n29867 , n29866 );
buf ( n29868 , n29867 );
and ( n29869 , n29862 , n29868 );
and ( n29870 , n29620 , n29861 );
or ( n29871 , n29869 , n29870 );
buf ( n29872 , n29871 );
buf ( n29873 , n29872 );
not ( n29874 , n18553 );
not ( n29875 , n831 );
or ( n29876 , n29874 , n29875 );
buf ( n29877 , n888 );
buf ( n29878 , n9799 );
xor ( n29879 , n29877 , n29878 );
buf ( n29880 , n9821 );
xor ( n29881 , n29879 , n29880 );
buf ( n29882 , n29881 );
buf ( n29883 , n29882 );
buf ( n29884 , n889 );
buf ( n29885 , n9912 );
xor ( n29886 , n29884 , n29885 );
buf ( n29887 , n9916 );
and ( n29888 , n29886 , n29887 );
and ( n29889 , n29884 , n29885 );
or ( n29890 , n29888 , n29889 );
buf ( n29891 , n29890 );
buf ( n29892 , n29891 );
nor ( n29893 , n29883 , n29892 );
buf ( n29894 , n29893 );
buf ( n29895 , n29894 );
not ( n29896 , n29895 );
buf ( n29897 , n29896 );
buf ( n29898 , n29897 );
buf ( n29899 , n891 );
buf ( n29900 , n10050 );
xor ( n29901 , n29899 , n29900 );
buf ( n29902 , n10054 );
xor ( n29903 , n29901 , n29902 );
buf ( n29904 , n29903 );
buf ( n29905 , n29904 );
buf ( n29906 , n892 );
buf ( n29907 , n10088 );
xor ( n29908 , n29906 , n29907 );
buf ( n29909 , n10115 );
and ( n29910 , n29908 , n29909 );
and ( n29911 , n29906 , n29907 );
or ( n29912 , n29910 , n29911 );
buf ( n29913 , n29912 );
buf ( n29914 , n29913 );
nor ( n29915 , n29905 , n29914 );
buf ( n29916 , n29915 );
buf ( n29917 , n29916 );
buf ( n29918 , n890 );
not ( n29919 , n29918 );
not ( n29920 , n9984 );
buf ( n29921 , n29920 );
not ( n29922 , n29921 );
or ( n29923 , n29919 , n29922 );
buf ( n29924 , n890 );
not ( n29925 , n29924 );
buf ( n29926 , n9984 );
nand ( n29927 , n29925 , n29926 );
buf ( n29928 , n29927 );
buf ( n29929 , n29928 );
nand ( n29930 , n29923 , n29929 );
buf ( n29931 , n29930 );
buf ( n29932 , n29931 );
buf ( n29933 , n29007 );
and ( n29934 , n29932 , n29933 );
not ( n29935 , n29932 );
buf ( n29936 , n29007 );
not ( n29937 , n29936 );
buf ( n29938 , n29937 );
buf ( n29939 , n29938 );
and ( n29940 , n29935 , n29939 );
nor ( n29941 , n29934 , n29940 );
buf ( n29942 , n29941 );
buf ( n29943 , n29942 );
xor ( n29944 , n29899 , n29900 );
and ( n29945 , n29944 , n29902 );
and ( n29946 , n29899 , n29900 );
or ( n29947 , n29945 , n29946 );
buf ( n29948 , n29947 );
buf ( n29949 , n29948 );
nor ( n29950 , n29943 , n29949 );
buf ( n29951 , n29950 );
buf ( n29952 , n29951 );
nor ( n29953 , n29917 , n29952 );
buf ( n29954 , n29953 );
buf ( n29955 , n893 );
buf ( n29956 , n10180 );
xor ( n29957 , n29955 , n29956 );
buf ( n29958 , n10174 );
xor ( n29959 , n29957 , n29958 );
buf ( n29960 , n29959 );
buf ( n29961 , n29960 );
and ( n29962 , n1185 , n1190 );
buf ( n29963 , n29962 );
buf ( n29964 , n29963 );
nand ( n29965 , n29961 , n29964 );
buf ( n29966 , n29965 );
buf ( n29967 , n29966 );
not ( n29968 , n29967 );
buf ( n29969 , n29968 );
buf ( n29970 , n29960 );
not ( n29971 , n29970 );
buf ( n29972 , n29971 );
buf ( n29973 , n29972 );
buf ( n29974 , n29963 );
not ( n29975 , n29974 );
buf ( n29976 , n29975 );
buf ( n29977 , n29976 );
and ( n29978 , n29973 , n29977 );
buf ( n29979 , n1176 );
buf ( n29980 , n1193 );
nand ( n29981 , n29979 , n29980 );
buf ( n29982 , n29981 );
buf ( n29983 , n29982 );
buf ( n29984 , n1184 );
and ( n29985 , n29983 , n29984 );
buf ( n29986 , n1175 );
buf ( n29987 , n1192 );
and ( n29988 , n29986 , n29987 );
buf ( n29989 , n29988 );
buf ( n29990 , n29989 );
nor ( n29991 , n29985 , n29990 );
buf ( n29992 , n29991 );
buf ( n29993 , n29992 );
nor ( n29994 , n29978 , n29993 );
buf ( n29995 , n29994 );
or ( n29996 , n29969 , n29995 );
xor ( n29997 , n29906 , n29907 );
xor ( n29998 , n29997 , n29909 );
buf ( n29999 , n29998 );
buf ( n30000 , n29999 );
not ( n30001 , n30000 );
buf ( n30002 , n30001 );
buf ( n30003 , n30002 );
xor ( n30004 , n29955 , n29956 );
and ( n30005 , n30004 , n29958 );
and ( n30006 , n29955 , n29956 );
or ( n30007 , n30005 , n30006 );
buf ( n30008 , n30007 );
buf ( n30009 , n30008 );
not ( n30010 , n30009 );
buf ( n30011 , n30010 );
buf ( n30012 , n30011 );
nand ( n30013 , n30003 , n30012 );
buf ( n30014 , n30013 );
nand ( n30015 , n29996 , n30014 );
buf ( n30016 , n30011 );
not ( n30017 , n30016 );
buf ( n30018 , n29999 );
nand ( n30019 , n30017 , n30018 );
buf ( n30020 , n30019 );
nand ( n30021 , n30015 , n30020 );
nand ( n30022 , n29954 , n30021 );
not ( n30023 , n30022 );
buf ( n30024 , n30023 );
xor ( n30025 , n29884 , n29885 );
xor ( n30026 , n30025 , n29887 );
buf ( n30027 , n30026 );
buf ( n30028 , n30027 );
buf ( n30029 , n9984 );
not ( n30030 , n30029 );
buf ( n30031 , n29007 );
not ( n30032 , n30031 );
or ( n30033 , n30030 , n30032 );
buf ( n30034 , n29007 );
buf ( n30035 , n9984 );
or ( n30036 , n30034 , n30035 );
buf ( n30037 , n890 );
nand ( n30038 , n30036 , n30037 );
buf ( n30039 , n30038 );
buf ( n30040 , n30039 );
nand ( n30041 , n30033 , n30040 );
buf ( n30042 , n30041 );
buf ( n30043 , n30042 );
nor ( n30044 , n30028 , n30043 );
buf ( n30045 , n30044 );
buf ( n30046 , n30045 );
not ( n30047 , n30046 );
buf ( n30048 , n30047 );
buf ( n30049 , n30048 );
nand ( n30050 , n29898 , n30024 , n30049 );
buf ( n30051 , n30050 );
buf ( n30052 , n30051 );
buf ( n30053 , n29897 );
buf ( n30054 , n29942 );
buf ( n30055 , n29948 );
nor ( n30056 , n30054 , n30055 );
buf ( n30057 , n30056 );
buf ( n30058 , n30057 );
buf ( n30059 , n29904 );
buf ( n30060 , n29913 );
nand ( n30061 , n30059 , n30060 );
buf ( n30062 , n30061 );
buf ( n30063 , n30062 );
or ( n30064 , n30058 , n30063 );
buf ( n30065 , n29942 );
buf ( n30066 , n29948 );
nand ( n30067 , n30065 , n30066 );
buf ( n30068 , n30067 );
buf ( n30069 , n30068 );
nand ( n30070 , n30064 , n30069 );
buf ( n30071 , n30070 );
buf ( n30072 , n30071 );
buf ( n30073 , n30048 );
nand ( n30074 , n30053 , n30072 , n30073 );
buf ( n30075 , n30074 );
buf ( n30076 , n30075 );
buf ( n30077 , n29894 );
not ( n30078 , n30077 );
buf ( n30079 , n30027 );
buf ( n30080 , n30042 );
nand ( n30081 , n30079 , n30080 );
buf ( n30082 , n30081 );
buf ( n30083 , n30082 );
not ( n30084 , n30083 );
and ( n30085 , n30078 , n30084 );
buf ( n30086 , n29882 );
buf ( n30087 , n29891 );
and ( n30088 , n30086 , n30087 );
buf ( n30089 , n30088 );
buf ( n30090 , n30089 );
nor ( n30091 , n30085 , n30090 );
buf ( n30092 , n30091 );
buf ( n30093 , n30092 );
nand ( n30094 , n30052 , n30076 , n30093 );
buf ( n30095 , n30094 );
buf ( n30096 , n30095 );
not ( n30097 , n30096 );
buf ( n30098 , n30097 );
buf ( n30099 , n30098 );
not ( n30100 , n30099 );
buf ( n30101 , n30100 );
buf ( n30102 , n30101 );
not ( n30103 , n30102 );
buf ( n30104 , n884 );
buf ( n30105 , n9354 );
xor ( n30106 , n30104 , n30105 );
buf ( n30107 , n9359 );
xor ( n30108 , n30106 , n30107 );
buf ( n30109 , n30108 );
buf ( n30110 , n30109 );
buf ( n30111 , n885 );
buf ( n30112 , n9489 );
xor ( n30113 , n30111 , n30112 );
buf ( n30114 , n9497 );
and ( n30115 , n30113 , n30114 );
and ( n30116 , n30111 , n30112 );
or ( n30117 , n30115 , n30116 );
buf ( n30118 , n30117 );
buf ( n30119 , n30118 );
nor ( n30120 , n30110 , n30119 );
buf ( n30121 , n30120 );
buf ( n30122 , n30121 );
not ( n30123 , n30122 );
buf ( n30124 , n30123 );
buf ( n30125 , n30124 );
xor ( n30126 , n30111 , n30112 );
xor ( n30127 , n30126 , n30114 );
buf ( n30128 , n30127 );
buf ( n30129 , n30128 );
buf ( n30130 , n886 );
buf ( n30131 , n9614 );
xor ( n30132 , n30130 , n30131 );
buf ( n30133 , n9619 );
and ( n30134 , n30132 , n30133 );
and ( n30135 , n30130 , n30131 );
or ( n30136 , n30134 , n30135 );
buf ( n30137 , n30136 );
buf ( n30138 , n30137 );
or ( n30139 , n30129 , n30138 );
buf ( n30140 , n30139 );
buf ( n30141 , n30140 );
buf ( n30142 , n887 );
buf ( n30143 , n9720 );
xor ( n30144 , n30142 , n30143 );
buf ( n30145 , n9725 );
xor ( n30146 , n30144 , n30145 );
buf ( n30147 , n30146 );
not ( n30148 , n30147 );
xor ( n30149 , n29877 , n29878 );
and ( n30150 , n30149 , n29880 );
and ( n30151 , n29877 , n29878 );
or ( n30152 , n30150 , n30151 );
buf ( n30153 , n30152 );
not ( n30154 , n30153 );
and ( n30155 , n30148 , n30154 );
xor ( n30156 , n30130 , n30131 );
xor ( n30157 , n30156 , n30133 );
buf ( n30158 , n30157 );
buf ( n30159 , n30158 );
xor ( n30160 , n30142 , n30143 );
and ( n30161 , n30160 , n30145 );
and ( n30162 , n30142 , n30143 );
or ( n30163 , n30161 , n30162 );
buf ( n30164 , n30163 );
buf ( n30165 , n30164 );
nor ( n30166 , n30159 , n30165 );
buf ( n30167 , n30166 );
nor ( n30168 , n30155 , n30167 );
buf ( n30169 , n30168 );
and ( n30170 , n30125 , n30141 , n30169 );
buf ( n30171 , n30170 );
buf ( n30172 , n30171 );
not ( n30173 , n30172 );
or ( n30174 , n30103 , n30173 );
buf ( n30175 , n30167 );
buf ( n30176 , n30147 );
buf ( n30177 , n30153 );
nand ( n30178 , n30176 , n30177 );
buf ( n30179 , n30178 );
buf ( n30180 , n30179 );
or ( n30181 , n30175 , n30180 );
buf ( n30182 , n30158 );
buf ( n30183 , n30164 );
nand ( n30184 , n30182 , n30183 );
buf ( n30185 , n30184 );
buf ( n30186 , n30185 );
nand ( n30187 , n30181 , n30186 );
buf ( n30188 , n30187 );
buf ( n30189 , n30188 );
not ( n30190 , n30189 );
buf ( n30191 , n30121 );
buf ( n30192 , n30128 );
buf ( n30193 , n30137 );
nor ( n30194 , n30192 , n30193 );
buf ( n30195 , n30194 );
buf ( n30196 , n30195 );
nor ( n30197 , n30191 , n30196 );
buf ( n30198 , n30197 );
buf ( n30199 , n30198 );
not ( n30200 , n30199 );
or ( n30201 , n30190 , n30200 );
buf ( n30202 , n30121 );
not ( n30203 , n30202 );
buf ( n30204 , n30128 );
buf ( n30205 , n30137 );
nand ( n30206 , n30204 , n30205 );
buf ( n30207 , n30206 );
buf ( n30208 , n30207 );
not ( n30209 , n30208 );
and ( n30210 , n30203 , n30209 );
buf ( n30211 , n30109 );
buf ( n30212 , n30118 );
and ( n30213 , n30211 , n30212 );
buf ( n30214 , n30213 );
buf ( n30215 , n30214 );
nor ( n30216 , n30210 , n30215 );
buf ( n30217 , n30216 );
buf ( n30218 , n30217 );
nand ( n30219 , n30201 , n30218 );
buf ( n30220 , n30219 );
buf ( n30221 , n30220 );
not ( n30222 , n30221 );
buf ( n30223 , n30222 );
buf ( n30224 , n30223 );
nand ( n30225 , n30174 , n30224 );
buf ( n30226 , n30225 );
buf ( n30227 , n883 );
buf ( n30228 , n9248 );
xor ( n30229 , n30227 , n30228 );
buf ( n30230 , n9253 );
xor ( n30231 , n30229 , n30230 );
buf ( n30232 , n30231 );
buf ( n30233 , n30232 );
xor ( n30234 , n30104 , n30105 );
and ( n30235 , n30234 , n30107 );
and ( n30236 , n30104 , n30105 );
or ( n30237 , n30235 , n30236 );
buf ( n30238 , n30237 );
buf ( n30239 , n30238 );
nor ( n30240 , n30233 , n30239 );
buf ( n30241 , n30240 );
buf ( n30242 , n30241 );
not ( n30243 , n30242 );
buf ( n30244 , n30243 );
buf ( n30245 , n30244 );
buf ( n30246 , n30232 );
buf ( n30247 , n30238 );
nand ( n30248 , n30246 , n30247 );
buf ( n30249 , n30248 );
buf ( n30250 , n30249 );
buf ( n30251 , n30250 );
buf ( n30252 , n30251 );
buf ( n30253 , n30252 );
nand ( n30254 , n30245 , n30253 );
buf ( n30255 , n30254 );
xnor ( n30256 , n30226 , n30255 );
nand ( n30257 , n30256 , n1152 );
nand ( n30258 , n29876 , n30257 );
buf ( n30259 , n30258 );
or ( n30260 , n30147 , n30153 );
not ( n30261 , n30260 );
nor ( n30262 , n30261 , n30167 , n30195 );
buf ( n30263 , n30262 );
not ( n30264 , n30263 );
buf ( n30265 , n30095 );
buf ( n30266 , n30265 );
buf ( n30267 , n30266 );
buf ( n30268 , n30267 );
not ( n30269 , n30268 );
or ( n30270 , n30264 , n30269 );
buf ( n30271 , n30188 );
not ( n30272 , n30271 );
buf ( n30273 , n30140 );
not ( n30274 , n30273 );
or ( n30275 , n30272 , n30274 );
buf ( n30276 , n30207 );
nand ( n30277 , n30275 , n30276 );
buf ( n30278 , n30277 );
buf ( n30279 , n30278 );
not ( n30280 , n30279 );
buf ( n30281 , n30280 );
buf ( n30282 , n30281 );
nand ( n30283 , n30270 , n30282 );
buf ( n30284 , n30283 );
buf ( n30285 , n30284 );
buf ( n30286 , n30124 );
not ( n30287 , n30286 );
buf ( n30288 , n30214 );
nor ( n30289 , n30287 , n30288 );
buf ( n30290 , n30289 );
buf ( n30291 , n30290 );
and ( n30292 , n30285 , n30291 );
not ( n30293 , n30285 );
buf ( n30294 , n30290 );
not ( n30295 , n30294 );
buf ( n30296 , n30295 );
buf ( n30297 , n30296 );
and ( n30298 , n30293 , n30297 );
nor ( n30299 , n30292 , n30298 );
buf ( n30300 , n30299 );
nand ( n30301 , n30300 , n1152 );
buf ( n30302 , n10279 );
buf ( n30303 , n9840 );
not ( n30304 , n30303 );
buf ( n30305 , n30304 );
buf ( n30306 , n30305 );
or ( n30307 , n9734 , n9730 );
buf ( n30308 , n30307 );
nand ( n30309 , n30306 , n30308 );
buf ( n30310 , n30309 );
buf ( n30311 , n30310 );
nor ( n30312 , n30302 , n30311 );
buf ( n30313 , n30312 );
buf ( n30314 , n30313 );
not ( n30315 , n30314 );
buf ( n30316 , n10249 );
buf ( n30317 , n30316 );
buf ( n30318 , n30317 );
buf ( n30319 , n30318 );
not ( n30320 , n30319 );
or ( n30321 , n30315 , n30320 );
buf ( n30322 , n9630 );
not ( n30323 , n30322 );
buf ( n30324 , n10270 );
not ( n30325 , n30324 );
or ( n30326 , n30323 , n30325 );
buf ( n30327 , n10288 );
nand ( n30328 , n30326 , n30327 );
buf ( n30329 , n30328 );
buf ( n30330 , n30329 );
not ( n30331 , n30330 );
buf ( n30332 , n30331 );
buf ( n30333 , n30332 );
nand ( n30334 , n30321 , n30333 );
buf ( n30335 , n30334 );
buf ( n30336 , n30335 );
not ( n30337 , n9516 );
nor ( n30338 , n30337 , n10297 );
buf ( n30339 , n30338 );
and ( n30340 , n30336 , n30339 );
not ( n30341 , n30336 );
buf ( n30342 , n30338 );
not ( n30343 , n30342 );
buf ( n30344 , n30343 );
buf ( n30345 , n30344 );
and ( n30346 , n30341 , n30345 );
nor ( n30347 , n30340 , n30346 );
buf ( n30348 , n30347 );
nand ( n30349 , n30348 , n831 );
nand ( n30350 , n30301 , n30349 );
buf ( n30351 , n30350 );
not ( n30352 , n831 );
and ( n30353 , n30305 , n10261 );
buf ( n30354 , n30353 );
not ( n30355 , n30354 );
buf ( n30356 , n10252 );
not ( n30357 , n30356 );
or ( n30358 , n30355 , n30357 );
buf ( n30359 , n30318 );
not ( n30360 , n30359 );
buf ( n30361 , n30360 );
buf ( n30362 , n30361 );
buf ( n30363 , n30353 );
or ( n30364 , n30362 , n30363 );
nand ( n30365 , n30358 , n30364 );
buf ( n30366 , n30365 );
not ( n30367 , n30366 );
or ( n30368 , n30352 , n30367 );
buf ( n30369 , n30260 );
buf ( n30370 , n30179 );
and ( n30371 , n30369 , n30370 );
buf ( n30372 , n30371 );
and ( n30373 , n30372 , n30098 );
not ( n30374 , n30372 );
and ( n30375 , n30374 , n30267 );
or ( n30376 , n30373 , n30375 );
nand ( n30377 , n30376 , n1152 );
nand ( n30378 , n30368 , n30377 );
buf ( n30379 , n30378 );
buf ( n30380 , n9997 );
buf ( n30381 , n30380 );
buf ( n30382 , n30381 );
buf ( n30383 , n30382 );
buf ( n30384 , n10143 );
buf ( n30385 , n10135 );
nand ( n30386 , n30384 , n30385 );
buf ( n30387 , n30386 );
buf ( n30388 , n30387 );
buf ( n30389 , n10239 );
not ( n30390 , n30389 );
buf ( n30391 , n30390 );
buf ( n30392 , n30391 );
not ( n30393 , n30392 );
buf ( n30394 , n10143 );
buf ( n30395 , n10160 );
buf ( n30396 , n30395 );
buf ( n30397 , n30396 );
buf ( n30398 , n30397 );
nand ( n30399 , n30393 , n30394 , n30398 );
buf ( n30400 , n30399 );
buf ( n30401 , n30400 );
nand ( n30402 , n30383 , n30388 , n30401 );
buf ( n30403 , n30402 );
buf ( n30404 , n30403 );
not ( n30405 , n30404 );
buf ( n30406 , n10006 );
not ( n30407 , n30406 );
buf ( n30408 , n9924 );
nand ( n30409 , n30407 , n30408 );
buf ( n30410 , n30409 );
buf ( n30411 , n30410 );
not ( n30412 , n30411 );
or ( n30413 , n30405 , n30412 );
buf ( n30414 , n30403 );
buf ( n30415 , n30410 );
or ( n30416 , n30414 , n30415 );
nand ( n30417 , n30413 , n30416 );
buf ( n30418 , n30417 );
and ( n30419 , n831 , n30418 );
not ( n30420 , n831 );
buf ( n30421 , n30089 );
not ( n30422 , n30421 );
buf ( n30423 , n29897 );
nand ( n30424 , n30422 , n30423 );
buf ( n30425 , n30424 );
buf ( n30426 , n30425 );
not ( n30427 , n30426 );
buf ( n30428 , n30082 );
buf ( n30429 , n30027 );
buf ( n30430 , n30042 );
nor ( n30431 , n30429 , n30430 );
buf ( n30432 , n30431 );
buf ( n30433 , n30432 );
not ( n30434 , n30433 );
buf ( n30435 , n29954 );
buf ( n30436 , n30435 );
buf ( n30437 , n30436 );
buf ( n30438 , n30437 );
not ( n30439 , n30021 );
not ( n30440 , n30439 );
buf ( n30441 , n30440 );
nand ( n30442 , n30434 , n30438 , n30441 );
buf ( n30443 , n30442 );
buf ( n30444 , n30443 );
buf ( n30445 , n30071 );
buf ( n30446 , n30432 );
not ( n30447 , n30446 );
buf ( n30448 , n30447 );
buf ( n30449 , n30448 );
nand ( n30450 , n30445 , n30449 );
buf ( n30451 , n30450 );
buf ( n30452 , n30451 );
nand ( n30453 , n30428 , n30444 , n30452 );
buf ( n30454 , n30453 );
buf ( n30455 , n30454 );
not ( n30456 , n30455 );
or ( n30457 , n30427 , n30456 );
buf ( n30458 , n30454 );
buf ( n30459 , n30425 );
or ( n30460 , n30458 , n30459 );
nand ( n30461 , n30457 , n30460 );
buf ( n30462 , n30461 );
and ( n30463 , n30420 , n30462 );
nor ( n30464 , n30419 , n30463 );
not ( n30465 , n30464 );
buf ( n30466 , n30168 );
not ( n30467 , n30466 );
buf ( n30468 , n30095 );
not ( n30469 , n30468 );
or ( n30470 , n30467 , n30469 );
buf ( n30471 , n30188 );
not ( n30472 , n30471 );
buf ( n30473 , n30472 );
buf ( n30474 , n30473 );
nand ( n30475 , n30470 , n30474 );
buf ( n30476 , n30475 );
buf ( n30477 , n30476 );
buf ( n30478 , n30140 );
buf ( n30479 , n30207 );
nand ( n30480 , n30478 , n30479 );
buf ( n30481 , n30480 );
buf ( n30482 , n30481 );
not ( n30483 , n30482 );
buf ( n30484 , n30483 );
buf ( n30485 , n30484 );
and ( n30486 , n30477 , n30485 );
not ( n30487 , n30477 );
buf ( n30488 , n30481 );
and ( n30489 , n30487 , n30488 );
nor ( n30490 , n30486 , n30489 );
buf ( n30491 , n30490 );
and ( n30492 , n1152 , n30491 );
not ( n30493 , n1152 );
buf ( n30494 , n9843 );
not ( n30495 , n30494 );
buf ( n30496 , n10249 );
not ( n30497 , n30496 );
or ( n30498 , n30495 , n30497 );
buf ( n30499 , n10270 );
not ( n30500 , n30499 );
buf ( n30501 , n30500 );
buf ( n30502 , n30501 );
nand ( n30503 , n30498 , n30502 );
buf ( n30504 , n30503 );
buf ( n30505 , n30504 );
buf ( n30506 , n9537 );
not ( n30507 , n30506 );
buf ( n30508 , n9627 );
not ( n30509 , n30508 );
or ( n30510 , n30507 , n30509 );
buf ( n30511 , n10288 );
nand ( n30512 , n30510 , n30511 );
buf ( n30513 , n30512 );
buf ( n30514 , n30513 );
not ( n30515 , n30514 );
buf ( n30516 , n30515 );
buf ( n30517 , n30516 );
and ( n30518 , n30505 , n30517 );
not ( n30519 , n30505 );
buf ( n30520 , n30513 );
and ( n30521 , n30519 , n30520 );
nor ( n30522 , n30518 , n30521 );
buf ( n30523 , n30522 );
and ( n30524 , n30493 , n30523 );
nor ( n30525 , n30492 , n30524 );
not ( n30526 , n1152 );
buf ( n30527 , n30260 );
not ( n30528 , n30527 );
buf ( n30529 , n30095 );
not ( n30530 , n30529 );
or ( n30531 , n30528 , n30530 );
buf ( n30532 , n30179 );
nand ( n30533 , n30531 , n30532 );
buf ( n30534 , n30533 );
buf ( n30535 , n30534 );
buf ( n30536 , n30167 );
not ( n30537 , n30536 );
buf ( n30538 , n30185 );
nand ( n30539 , n30537 , n30538 );
buf ( n30540 , n30539 );
buf ( n30541 , n30540 );
not ( n30542 , n30541 );
buf ( n30543 , n30542 );
buf ( n30544 , n30543 );
and ( n30545 , n30535 , n30544 );
not ( n30546 , n30535 );
buf ( n30547 , n30540 );
and ( n30548 , n30546 , n30547 );
nor ( n30549 , n30545 , n30548 );
buf ( n30550 , n30549 );
not ( n30551 , n30550 );
or ( n30552 , n30526 , n30551 );
buf ( n30553 , n30305 );
not ( n30554 , n30553 );
buf ( n30555 , n10249 );
not ( n30556 , n30555 );
or ( n30557 , n30554 , n30556 );
buf ( n30558 , n10261 );
nand ( n30559 , n30557 , n30558 );
buf ( n30560 , n30559 );
buf ( n30561 , n30560 );
buf ( n30562 , n30307 );
buf ( n30563 , n10267 );
nand ( n30564 , n30562 , n30563 );
buf ( n30565 , n30564 );
buf ( n30566 , n30565 );
not ( n30567 , n30566 );
buf ( n30568 , n30567 );
buf ( n30569 , n30568 );
and ( n30570 , n30561 , n30569 );
not ( n30571 , n30561 );
buf ( n30572 , n30565 );
and ( n30573 , n30571 , n30572 );
nor ( n30574 , n30570 , n30573 );
buf ( n30575 , n30574 );
nand ( n30576 , n30575 , n831 );
nand ( n30577 , n30552 , n30576 );
not ( n30578 , n831 );
buf ( n30579 , n10229 );
buf ( n30580 , n10238 );
nand ( n30581 , n30579 , n30580 );
buf ( n30582 , n30581 );
buf ( n30583 , n30582 );
buf ( n30584 , n10213 );
not ( n30585 , n30584 );
buf ( n30586 , n30585 );
buf ( n30587 , n30586 );
and ( n30588 , n30583 , n30587 );
not ( n30589 , n30583 );
buf ( n30590 , n10213 );
and ( n30591 , n30589 , n30590 );
nor ( n30592 , n30588 , n30591 );
buf ( n30593 , n30592 );
not ( n30594 , n30593 );
or ( n30595 , n30578 , n30594 );
buf ( n30596 , n30014 );
buf ( n30597 , n30020 );
nand ( n30598 , n30596 , n30597 );
buf ( n30599 , n30598 );
buf ( n30600 , n30599 );
buf ( n30601 , n29995 );
not ( n30602 , n30601 );
buf ( n30603 , n29966 );
nand ( n30604 , n30602 , n30603 );
buf ( n30605 , n30604 );
buf ( n30606 , n30605 );
xnor ( n30607 , n30600 , n30606 );
buf ( n30608 , n30607 );
nand ( n30609 , n30608 , n1152 );
nand ( n30610 , n30595 , n30609 );
not ( n30611 , n831 );
buf ( n30612 , n10189 );
not ( n30613 , n30612 );
buf ( n30614 , n10210 );
nand ( n30615 , n30613 , n30614 );
buf ( n30616 , n30615 );
xor ( n30617 , n30616 , n10201 );
not ( n30618 , n30617 );
or ( n30619 , n30611 , n30618 );
buf ( n30620 , n29992 );
buf ( n30621 , n29976 );
not ( n30622 , n30621 );
buf ( n30623 , n29972 );
not ( n30624 , n30623 );
or ( n30625 , n30622 , n30624 );
buf ( n30626 , n29966 );
nand ( n30627 , n30625 , n30626 );
buf ( n30628 , n30627 );
buf ( n30629 , n30628 );
xor ( n30630 , n30620 , n30629 );
buf ( n30631 , n30630 );
nand ( n30632 , n30631 , n1152 );
nand ( n30633 , n30619 , n30632 );
not ( n30634 , n831 );
buf ( n30635 , n8884 );
not ( n30636 , n30635 );
buf ( n30637 , n8414 );
nor ( n30638 , n30636 , n30637 );
buf ( n30639 , n30638 );
buf ( n30640 , n30639 );
not ( n30641 , n30640 );
buf ( n30642 , n18807 );
not ( n30643 , n30642 );
or ( n30644 , n30641 , n30643 );
buf ( n30645 , n18812 );
buf ( n30646 , n18820 );
and ( n30647 , n30645 , n30646 );
buf ( n30648 , n8788 );
nor ( n30649 , n30647 , n30648 );
buf ( n30650 , n30649 );
buf ( n30651 , n30650 );
nand ( n30652 , n30644 , n30651 );
buf ( n30653 , n30652 );
buf ( n30654 , n30653 );
buf ( n30655 , n8777 );
not ( n30656 , n30655 );
buf ( n30657 , n8794 );
nor ( n30658 , n30656 , n30657 );
buf ( n30659 , n30658 );
buf ( n30660 , n30659 );
and ( n30661 , n30654 , n30660 );
not ( n30662 , n30654 );
buf ( n30663 , n30659 );
not ( n30664 , n30663 );
buf ( n30665 , n30664 );
buf ( n30666 , n30665 );
and ( n30667 , n30662 , n30666 );
nor ( n30668 , n30661 , n30667 );
buf ( n30669 , n30668 );
not ( n30670 , n30669 );
or ( n30671 , n30634 , n30670 );
buf ( n30672 , n878 );
buf ( n30673 , n8401 );
xor ( n30674 , n30672 , n30673 );
buf ( n30675 , n8406 );
xor ( n30676 , n30674 , n30675 );
buf ( n30677 , n30676 );
not ( n30678 , n30677 );
buf ( n30679 , n879 );
buf ( n30680 , n8737 );
xor ( n30681 , n30679 , n30680 );
buf ( n30682 , n8742 );
and ( n30683 , n30681 , n30682 );
and ( n30684 , n30679 , n30680 );
or ( n30685 , n30683 , n30684 );
buf ( n30686 , n30685 );
not ( n30687 , n30686 );
and ( n30688 , n30678 , n30687 );
buf ( n30689 , n880 );
buf ( n30690 , n8706 );
xor ( n30691 , n30689 , n30690 );
buf ( n30692 , n8725 );
and ( n30693 , n30691 , n30692 );
and ( n30694 , n30689 , n30690 );
or ( n30695 , n30693 , n30694 );
buf ( n30696 , n30695 );
xor ( n30697 , n30679 , n30680 );
xor ( n30698 , n30697 , n30682 );
buf ( n30699 , n30698 );
nor ( n30700 , n30696 , n30699 );
nor ( n30701 , n30688 , n30700 );
buf ( n30702 , n877 );
buf ( n30703 , n8159 );
xor ( n30704 , n30702 , n30703 );
buf ( n30705 , n8163 );
xor ( n30706 , n30704 , n30705 );
buf ( n30707 , n30706 );
buf ( n30708 , n30707 );
xor ( n30709 , n30672 , n30673 );
and ( n30710 , n30709 , n30675 );
and ( n30711 , n30672 , n30673 );
or ( n30712 , n30710 , n30711 );
buf ( n30713 , n30712 );
buf ( n30714 , n30713 );
nor ( n30715 , n30708 , n30714 );
buf ( n30716 , n30715 );
buf ( n30717 , n30716 );
not ( n30718 , n30717 );
buf ( n30719 , n30718 );
and ( n30720 , n30701 , n30719 );
buf ( n30721 , n30720 );
not ( n30722 , n30721 );
buf ( n30723 , n881 );
buf ( n30724 , n8978 );
xor ( n30725 , n30723 , n30724 );
buf ( n30726 , n8983 );
and ( n30727 , n30725 , n30726 );
and ( n30728 , n30723 , n30724 );
or ( n30729 , n30727 , n30728 );
buf ( n30730 , n30729 );
buf ( n30731 , n30730 );
not ( n30732 , n30731 );
xor ( n30733 , n30689 , n30690 );
xor ( n30734 , n30733 , n30692 );
buf ( n30735 , n30734 );
buf ( n30736 , n30735 );
not ( n30737 , n30736 );
buf ( n30738 , n30737 );
buf ( n30739 , n30738 );
nand ( n30740 , n30732 , n30739 );
buf ( n30741 , n30740 );
buf ( n30742 , n30741 );
buf ( n30743 , n30241 );
xor ( n30744 , n30227 , n30228 );
and ( n30745 , n30744 , n30230 );
and ( n30746 , n30227 , n30228 );
or ( n30747 , n30745 , n30746 );
buf ( n30748 , n30747 );
buf ( n30749 , n30748 );
buf ( n30750 , n882 );
buf ( n30751 , n9123 );
xor ( n30752 , n30750 , n30751 );
buf ( n30753 , n9128 );
xor ( n30754 , n30752 , n30753 );
buf ( n30755 , n30754 );
buf ( n30756 , n30755 );
nor ( n30757 , n30749 , n30756 );
buf ( n30758 , n30757 );
buf ( n30759 , n30758 );
nor ( n30760 , n30743 , n30759 );
buf ( n30761 , n30760 );
buf ( n30762 , n30761 );
xor ( n30763 , n30723 , n30724 );
xor ( n30764 , n30763 , n30726 );
buf ( n30765 , n30764 );
buf ( n30766 , n30765 );
xor ( n30767 , n30750 , n30751 );
and ( n30768 , n30767 , n30753 );
and ( n30769 , n30750 , n30751 );
or ( n30770 , n30768 , n30769 );
buf ( n30771 , n30770 );
buf ( n30772 , n30771 );
nor ( n30773 , n30766 , n30772 );
buf ( n30774 , n30773 );
buf ( n30775 , n30774 );
not ( n30776 , n30775 );
buf ( n30777 , n30776 );
buf ( n30778 , n30777 );
and ( n30779 , n30742 , n30762 , n30778 );
buf ( n30780 , n30779 );
buf ( n30781 , n30780 );
not ( n30782 , n30781 );
buf ( n30783 , n30226 );
not ( n30784 , n30783 );
or ( n30785 , n30782 , n30784 );
buf ( n30786 , n30755 );
buf ( n30787 , n30748 );
nor ( n30788 , n30786 , n30787 );
buf ( n30789 , n30788 );
buf ( n30790 , n30789 );
buf ( n30791 , n30249 );
or ( n30792 , n30790 , n30791 );
buf ( n30793 , n30755 );
buf ( n30794 , n30748 );
nand ( n30795 , n30793 , n30794 );
buf ( n30796 , n30795 );
buf ( n30797 , n30796 );
nand ( n30798 , n30792 , n30797 );
buf ( n30799 , n30798 );
buf ( n30800 , n30799 );
not ( n30801 , n30800 );
buf ( n30802 , n30730 );
buf ( n30803 , n30735 );
nor ( n30804 , n30802 , n30803 );
buf ( n30805 , n30804 );
buf ( n30806 , n30805 );
buf ( n30807 , n30774 );
nor ( n30808 , n30806 , n30807 );
buf ( n30809 , n30808 );
buf ( n30810 , n30809 );
not ( n30811 , n30810 );
or ( n30812 , n30801 , n30811 );
buf ( n30813 , n30741 );
buf ( n30814 , n30765 );
buf ( n30815 , n30771 );
and ( n30816 , n30814 , n30815 );
buf ( n30817 , n30816 );
buf ( n30818 , n30817 );
and ( n30819 , n30813 , n30818 );
buf ( n30820 , n30730 );
not ( n30821 , n30820 );
buf ( n30822 , n30738 );
nor ( n30823 , n30821 , n30822 );
buf ( n30824 , n30823 );
buf ( n30825 , n30824 );
nor ( n30826 , n30819 , n30825 );
buf ( n30827 , n30826 );
buf ( n30828 , n30827 );
nand ( n30829 , n30812 , n30828 );
buf ( n30830 , n30829 );
buf ( n30831 , n30830 );
not ( n30832 , n30831 );
buf ( n30833 , n30832 );
buf ( n30834 , n30833 );
nand ( n30835 , n30785 , n30834 );
buf ( n30836 , n30835 );
buf ( n30837 , n30836 );
not ( n30838 , n30837 );
or ( n30839 , n30722 , n30838 );
buf ( n30840 , n30696 );
buf ( n30841 , n30699 );
nand ( n30842 , n30840 , n30841 );
buf ( n30843 , n30842 );
buf ( n30844 , n30677 );
buf ( n30845 , n30686 );
nand ( n30846 , n30844 , n30845 );
buf ( n30847 , n30846 );
and ( n30848 , n30843 , n30847 );
buf ( n30849 , n30677 );
not ( n30850 , n30849 );
buf ( n30851 , n30850 );
buf ( n30852 , n30851 );
buf ( n30853 , n30686 );
not ( n30854 , n30853 );
buf ( n30855 , n30854 );
buf ( n30856 , n30855 );
nand ( n30857 , n30852 , n30856 );
buf ( n30858 , n30857 );
not ( n30859 , n30858 );
nor ( n30860 , n30848 , n30859 );
buf ( n30861 , n30860 );
and ( n30862 , n30719 , n30861 );
buf ( n30863 , n30707 );
not ( n30864 , n30863 );
buf ( n30865 , n30864 );
buf ( n30866 , n30865 );
buf ( n30867 , n30713 );
not ( n30868 , n30867 );
buf ( n30869 , n30868 );
buf ( n30870 , n30869 );
nor ( n30871 , n30866 , n30870 );
buf ( n30872 , n30871 );
buf ( n30873 , n30872 );
buf ( n30874 , n30873 );
buf ( n30875 , n30874 );
nor ( n30876 , n30862 , n30875 );
buf ( n30877 , n30876 );
nand ( n30878 , n30839 , n30877 );
buf ( n30879 , n30878 );
buf ( n30880 , n30879 );
xor ( n30881 , n30702 , n30703 );
and ( n30882 , n30881 , n30705 );
and ( n30883 , n30702 , n30703 );
or ( n30884 , n30882 , n30883 );
buf ( n30885 , n30884 );
buf ( n30886 , n30885 );
not ( n30887 , n30886 );
buf ( n30888 , n876 );
buf ( n30889 , n7947 );
xor ( n30890 , n30888 , n30889 );
buf ( n30891 , n7951 );
xor ( n30892 , n30890 , n30891 );
buf ( n30893 , n30892 );
buf ( n30894 , n30893 );
not ( n30895 , n30894 );
buf ( n30896 , n30895 );
buf ( n30897 , n30896 );
nand ( n30898 , n30887 , n30897 );
buf ( n30899 , n30898 );
buf ( n30900 , n30899 );
not ( n30901 , n30900 );
buf ( n30902 , n30901 );
buf ( n30903 , n30902 );
not ( n30904 , n30903 );
buf ( n30905 , n30904 );
buf ( n30906 , n30905 );
buf ( n30907 , n30893 );
buf ( n30908 , n30885 );
buf ( n30909 , n30908 );
buf ( n30910 , n30909 );
buf ( n30911 , n30910 );
nand ( n30912 , n30907 , n30911 );
buf ( n30913 , n30912 );
buf ( n30914 , n30913 );
and ( n30915 , n30906 , n30914 );
buf ( n30916 , n30915 );
buf ( n30917 , n30916 );
and ( n30918 , n30880 , n30917 );
not ( n30919 , n30880 );
buf ( n30920 , n30916 );
not ( n30921 , n30920 );
buf ( n30922 , n30921 );
buf ( n30923 , n30922 );
and ( n30924 , n30919 , n30923 );
nor ( n30925 , n30918 , n30924 );
buf ( n30926 , n30925 );
nand ( n30927 , n30926 , n1152 );
nand ( n30928 , n30671 , n30927 );
buf ( n30929 , n30928 );
not ( n30930 , n831 );
buf ( n30931 , n8883 );
not ( n30932 , n30931 );
buf ( n30933 , n30932 );
buf ( n30934 , n30933 );
buf ( n30935 , n8748 );
nand ( n30936 , n30934 , n30935 );
buf ( n30937 , n30936 );
buf ( n30938 , n30937 );
not ( n30939 , n30938 );
buf ( n30940 , n18807 );
not ( n30941 , n30940 );
buf ( n30942 , n30941 );
buf ( n30943 , n30942 );
not ( n30944 , n30943 );
buf ( n30945 , n30944 );
buf ( n30946 , n30945 );
not ( n30947 , n30946 );
or ( n30948 , n30939 , n30947 );
buf ( n30949 , n30942 );
not ( n30950 , n30949 );
buf ( n30951 , n30950 );
buf ( n30952 , n30951 );
buf ( n30953 , n30937 );
or ( n30954 , n30952 , n30953 );
nand ( n30955 , n30948 , n30954 );
buf ( n30956 , n30955 );
not ( n30957 , n30956 );
or ( n30958 , n30930 , n30957 );
not ( n30959 , n30700 );
and ( n30960 , n30843 , n30959 );
xor ( n30961 , n30960 , n30836 );
nand ( n30962 , n30961 , n1152 );
nand ( n30963 , n30958 , n30962 );
buf ( n30964 , n30963 );
nand ( n30965 , n15271 , n14941 );
buf ( n30966 , n30965 );
buf ( n30967 , n15634 );
buf ( n30968 , n15332 );
xor ( n30969 , n30967 , n30968 );
buf ( n30970 , n30969 );
buf ( n30971 , n30970 );
not ( n30972 , n30971 );
buf ( n30973 , n30972 );
buf ( n30974 , n30973 );
nand ( n30975 , n30966 , n30974 );
buf ( n30976 , n30975 );
buf ( n30977 , n30976 );
not ( n30978 , n30977 );
buf ( n30979 , n14126 );
buf ( n30980 , n14121 );
nand ( n30981 , n30979 , n30980 );
buf ( n30982 , n30981 );
buf ( n30983 , n30982 );
not ( n30984 , n30983 );
buf ( n30985 , n30984 );
not ( n30986 , n30985 );
buf ( n30987 , n14510 );
buf ( n30988 , n14500 );
xor ( n30989 , n30987 , n30988 );
buf ( n30990 , n30989 );
not ( n30991 , n30990 );
and ( n30992 , n30986 , n30991 );
buf ( n30993 , n14126 );
not ( n30994 , n30993 );
buf ( n30995 , n14528 );
not ( n30996 , n30995 );
or ( n30997 , n30994 , n30996 );
buf ( n30998 , n14534 );
buf ( n30999 , n14121 );
nand ( n31000 , n30998 , n30999 );
buf ( n31001 , n31000 );
buf ( n31002 , n31001 );
nand ( n31003 , n30997 , n31002 );
buf ( n31004 , n31003 );
buf ( n31005 , n31004 );
and ( n31006 , n13276 , n13658 );
buf ( n31007 , n31006 );
nor ( n31008 , n31005 , n31007 );
buf ( n31009 , n31008 );
nor ( n31010 , n30992 , n31009 );
and ( n31011 , n30987 , n30988 );
buf ( n31012 , n31011 );
buf ( n31013 , n31012 );
not ( n31014 , n31013 );
buf ( n31015 , n31014 );
buf ( n31016 , n31015 );
xnor ( n31017 , n15290 , n15284 );
buf ( n31018 , n31017 );
nand ( n31019 , n31016 , n31018 );
buf ( n31020 , n31019 );
buf ( n31021 , n15284 );
buf ( n31022 , n15290 );
nand ( n31023 , n31021 , n31022 );
buf ( n31024 , n31023 );
buf ( n31025 , n31024 );
xnor ( n31026 , n14941 , n15271 );
buf ( n31027 , n31026 );
nand ( n31028 , n31025 , n31027 );
buf ( n31029 , n31028 );
nand ( n31030 , n31020 , n31029 );
not ( n31031 , n31030 );
nand ( n31032 , n31010 , n31031 );
not ( n31033 , n31032 );
buf ( n31034 , n31033 );
not ( n31035 , n31034 );
buf ( n31036 , n31035 );
buf ( n31037 , n31036 );
nor ( n31038 , n30978 , n31037 );
buf ( n31039 , n31038 );
buf ( n31040 , n864 );
buf ( n31041 , n3320 );
xor ( n31042 , n31040 , n31041 );
buf ( n31043 , n3783 );
and ( n31044 , n31042 , n31043 );
and ( n31045 , n31040 , n31041 );
or ( n31046 , n31044 , n31045 );
buf ( n31047 , n31046 );
buf ( n31048 , n31047 );
buf ( n31049 , n3794 );
not ( n31050 , n31049 );
buf ( n31051 , n4328 );
not ( n31052 , n31051 );
or ( n31053 , n31050 , n31052 );
buf ( n31054 , n4325 );
buf ( n31055 , n4335 );
nand ( n31056 , n31054 , n31055 );
buf ( n31057 , n31056 );
buf ( n31058 , n31057 );
nand ( n31059 , n31053 , n31058 );
buf ( n31060 , n31059 );
buf ( n31061 , n31060 );
nor ( n31062 , n31048 , n31061 );
buf ( n31063 , n31062 );
not ( n31064 , n13719 );
not ( n31065 , n13739 );
or ( n31066 , n31064 , n31065 );
buf ( n31067 , n13713 );
buf ( n31068 , n13746 );
nand ( n31069 , n31067 , n31068 );
buf ( n31070 , n31069 );
nand ( n31071 , n31066 , n31070 );
buf ( n31072 , n31071 );
buf ( n31073 , n4325 );
buf ( n31074 , n3794 );
and ( n31075 , n31073 , n31074 );
buf ( n31076 , n31075 );
buf ( n31077 , n31076 );
nor ( n31078 , n31072 , n31077 );
buf ( n31079 , n31078 );
nor ( n31080 , n31063 , n31079 );
buf ( n31081 , n13706 );
not ( n31082 , n31081 );
buf ( n31083 , n13687 );
not ( n31084 , n31083 );
or ( n31085 , n31082 , n31084 );
buf ( n31086 , n13688 );
buf ( n31087 , n13709 );
nand ( n31088 , n31086 , n31087 );
buf ( n31089 , n31088 );
buf ( n31090 , n31089 );
nand ( n31091 , n31085 , n31090 );
buf ( n31092 , n31091 );
not ( n31093 , n31092 );
and ( n31094 , n13713 , n13719 );
not ( n31095 , n31094 );
and ( n31096 , n31093 , n31095 );
not ( n31097 , n12715 );
buf ( n31098 , n31097 );
not ( n31099 , n31098 );
buf ( n31100 , n12802 );
not ( n31101 , n31100 );
or ( n31102 , n31099 , n31101 );
not ( n31103 , n12802 );
nand ( n31104 , n31103 , n12715 );
buf ( n31105 , n31104 );
nand ( n31106 , n31102 , n31105 );
buf ( n31107 , n31106 );
buf ( n31108 , n31107 );
and ( n31109 , n13688 , n13706 );
buf ( n31110 , n31109 );
nor ( n31111 , n31108 , n31110 );
buf ( n31112 , n31111 );
nor ( n31113 , n31096 , n31112 );
nand ( n31114 , n31080 , n31113 );
not ( n31115 , n31114 );
and ( n31116 , n12396 , n12574 );
buf ( n31117 , n31116 );
not ( n31118 , n31117 );
buf ( n31119 , n12815 );
not ( n31120 , n31119 );
buf ( n31121 , n13230 );
not ( n31122 , n31121 );
or ( n31123 , n31120 , n31122 );
buf ( n31124 , n13236 );
buf ( n31125 , n13229 );
nand ( n31126 , n31124 , n31125 );
buf ( n31127 , n31126 );
buf ( n31128 , n31127 );
nand ( n31129 , n31123 , n31128 );
buf ( n31130 , n31129 );
buf ( n31131 , n31130 );
not ( n31132 , n31131 );
buf ( n31133 , n31132 );
buf ( n31134 , n31133 );
nand ( n31135 , n31118 , n31134 );
buf ( n31136 , n31135 );
buf ( n31137 , n31136 );
buf ( n31138 , n13199 );
not ( n31139 , n31138 );
buf ( n31140 , n13215 );
not ( n31141 , n31140 );
or ( n31142 , n31139 , n31141 );
buf ( n31143 , n13273 );
nand ( n31144 , n31142 , n31143 );
buf ( n31145 , n31144 );
not ( n31146 , n31145 );
not ( n31147 , n13661 );
or ( n31148 , n31146 , n31147 );
buf ( n31149 , n13658 );
buf ( n31150 , n13277 );
nand ( n31151 , n31149 , n31150 );
buf ( n31152 , n31151 );
nand ( n31153 , n31148 , n31152 );
buf ( n31154 , n13229 );
buf ( n31155 , n12815 );
and ( n31156 , n31154 , n31155 );
buf ( n31157 , n31156 );
nor ( n31158 , n31153 , n31157 );
buf ( n31159 , n12700 );
buf ( n31160 , n12704 );
xor ( n31161 , n31159 , n31160 );
buf ( n31162 , n31161 );
buf ( n31163 , n12715 );
buf ( n31164 , n12802 );
and ( n31165 , n31163 , n31164 );
buf ( n31166 , n31165 );
nor ( n31167 , n31162 , n31166 );
nor ( n31168 , n31158 , n31167 );
buf ( n31169 , n31168 );
and ( n31170 , n31159 , n31160 );
buf ( n31171 , n31170 );
not ( n31172 , n31171 );
xnor ( n31173 , n12396 , n12574 );
nand ( n31174 , n31172 , n31173 );
buf ( n31175 , n31174 );
nand ( n31176 , n31137 , n31169 , n31175 );
buf ( n31177 , n31176 );
buf ( n31178 , n31177 );
not ( n31179 , n31178 );
buf ( n31180 , n31179 );
nand ( n31181 , n31115 , n31180 );
not ( n31182 , n31181 );
and ( n31183 , n31039 , n31182 );
buf ( n31184 , n31183 );
not ( n31185 , n31184 );
buf ( n31186 , n870 );
buf ( n31187 , n6313 );
xor ( n31188 , n31186 , n31187 );
buf ( n31189 , n6318 );
xor ( n31190 , n31188 , n31189 );
buf ( n31191 , n31190 );
buf ( n31192 , n31191 );
buf ( n31193 , n871 );
buf ( n31194 , n6757 );
xor ( n31195 , n31193 , n31194 );
buf ( n31196 , n6762 );
and ( n31197 , n31195 , n31196 );
and ( n31198 , n31193 , n31194 );
or ( n31199 , n31197 , n31198 );
buf ( n31200 , n31199 );
buf ( n31201 , n31200 );
nor ( n31202 , n31192 , n31201 );
buf ( n31203 , n31202 );
buf ( n31204 , n31203 );
xor ( n31205 , n31193 , n31194 );
xor ( n31206 , n31205 , n31196 );
buf ( n31207 , n31206 );
buf ( n31208 , n31207 );
buf ( n31209 , n872 );
buf ( n31210 , n6841 );
xor ( n31211 , n31209 , n31210 );
buf ( n31212 , n6846 );
and ( n31213 , n31211 , n31212 );
and ( n31214 , n31209 , n31210 );
or ( n31215 , n31213 , n31214 );
buf ( n31216 , n31215 );
buf ( n31217 , n31216 );
nor ( n31218 , n31208 , n31217 );
buf ( n31219 , n31218 );
buf ( n31220 , n31219 );
nor ( n31221 , n31204 , n31220 );
buf ( n31222 , n31221 );
buf ( n31223 , n31222 );
not ( n31224 , n31223 );
buf ( n31225 , n31224 );
buf ( n31226 , n31225 );
not ( n31227 , n31226 );
buf ( n31228 , n31227 );
buf ( n31229 , n867 );
buf ( n31230 , n5492 );
xor ( n31231 , n31229 , n31230 );
buf ( n31232 , n5487 );
and ( n31233 , n31231 , n31232 );
and ( n31234 , n31229 , n31230 );
or ( n31235 , n31233 , n31234 );
buf ( n31236 , n31235 );
buf ( n31237 , n31236 );
not ( n31238 , n31237 );
buf ( n31239 , n866 );
buf ( n31240 , n5139 );
xor ( n31241 , n31239 , n31240 );
buf ( n31242 , n5168 );
xor ( n31243 , n31241 , n31242 );
buf ( n31244 , n31243 );
buf ( n31245 , n31244 );
not ( n31246 , n31245 );
buf ( n31247 , n31246 );
buf ( n31248 , n31247 );
nand ( n31249 , n31238 , n31248 );
buf ( n31250 , n31249 );
buf ( n31251 , n31250 );
buf ( n31252 , n868 );
buf ( n31253 , n5860 );
xor ( n31254 , n31252 , n31253 );
buf ( n31255 , n5865 );
and ( n31256 , n31254 , n31255 );
and ( n31257 , n31252 , n31253 );
or ( n31258 , n31256 , n31257 );
buf ( n31259 , n31258 );
buf ( n31260 , n31259 );
not ( n31261 , n31260 );
xor ( n31262 , n31229 , n31230 );
xor ( n31263 , n31262 , n31232 );
buf ( n31264 , n31263 );
buf ( n31265 , n31264 );
not ( n31266 , n31265 );
buf ( n31267 , n31266 );
buf ( n31268 , n31267 );
nand ( n31269 , n31261 , n31268 );
buf ( n31270 , n31269 );
buf ( n31271 , n31270 );
and ( n31272 , n31251 , n31271 );
buf ( n31273 , n31272 );
buf ( n31274 , n30902 );
not ( n31275 , n31274 );
buf ( n31276 , n30719 );
buf ( n31277 , n30701 );
nand ( n31278 , n31275 , n31276 , n31277 );
buf ( n31279 , n31278 );
buf ( n31280 , n31279 );
not ( n31281 , n31280 );
buf ( n31282 , n31281 );
and ( n31283 , n31228 , n31273 , n31282 );
xor ( n31284 , n31252 , n31253 );
xor ( n31285 , n31284 , n31255 );
buf ( n31286 , n31285 );
buf ( n31287 , n31286 );
buf ( n31288 , n869 );
buf ( n31289 , n6188 );
xor ( n31290 , n31288 , n31289 );
buf ( n31291 , n6193 );
and ( n31292 , n31290 , n31291 );
and ( n31293 , n31288 , n31289 );
or ( n31294 , n31292 , n31293 );
buf ( n31295 , n31294 );
buf ( n31296 , n31295 );
nor ( n31297 , n31287 , n31296 );
buf ( n31298 , n31297 );
buf ( n31299 , n31298 );
xor ( n31300 , n31288 , n31289 );
xor ( n31301 , n31300 , n31291 );
buf ( n31302 , n31301 );
buf ( n31303 , n31302 );
xor ( n31304 , n31186 , n31187 );
and ( n31305 , n31304 , n31189 );
and ( n31306 , n31186 , n31187 );
or ( n31307 , n31305 , n31306 );
buf ( n31308 , n31307 );
buf ( n31309 , n31308 );
nor ( n31310 , n31303 , n31309 );
buf ( n31311 , n31310 );
buf ( n31312 , n31311 );
nor ( n31313 , n31299 , n31312 );
buf ( n31314 , n31313 );
buf ( n31315 , n31314 );
buf ( n31316 , n31315 );
buf ( n31317 , n31316 );
buf ( n31318 , n30836 );
buf ( n31319 , n31318 );
buf ( n31320 , n31319 );
buf ( n31321 , n873 );
buf ( n31322 , n7128 );
xor ( n31323 , n31321 , n31322 );
buf ( n31324 , n7133 );
and ( n31325 , n31323 , n31324 );
and ( n31326 , n31321 , n31322 );
or ( n31327 , n31325 , n31326 );
buf ( n31328 , n31327 );
buf ( n31329 , n31328 );
xor ( n31330 , n31209 , n31210 );
xor ( n31331 , n31330 , n31212 );
buf ( n31332 , n31331 );
buf ( n31333 , n31332 );
nor ( n31334 , n31329 , n31333 );
buf ( n31335 , n31334 );
buf ( n31336 , n31335 );
buf ( n31337 , n874 );
buf ( n31338 , n7446 );
xor ( n31339 , n31337 , n31338 );
buf ( n31340 , n7451 );
and ( n31341 , n31339 , n31340 );
and ( n31342 , n31337 , n31338 );
or ( n31343 , n31341 , n31342 );
buf ( n31344 , n31343 );
buf ( n31345 , n31344 );
xor ( n31346 , n31321 , n31322 );
xor ( n31347 , n31346 , n31324 );
buf ( n31348 , n31347 );
buf ( n31349 , n31348 );
nor ( n31350 , n31345 , n31349 );
buf ( n31351 , n31350 );
buf ( n31352 , n31351 );
nor ( n31353 , n31336 , n31352 );
buf ( n31354 , n31353 );
buf ( n31355 , n31354 );
buf ( n31356 , n875 );
buf ( n31357 , n7712 );
xor ( n31358 , n31356 , n31357 );
buf ( n31359 , n7716 );
and ( n31360 , n31358 , n31359 );
and ( n31361 , n31356 , n31357 );
or ( n31362 , n31360 , n31361 );
buf ( n31363 , n31362 );
not ( n31364 , n31363 );
not ( n31365 , n31364 );
xor ( n31366 , n31337 , n31338 );
xor ( n31367 , n31366 , n31340 );
buf ( n31368 , n31367 );
buf ( n31369 , n31368 );
not ( n31370 , n31369 );
buf ( n31371 , n31370 );
not ( n31372 , n31371 );
or ( n31373 , n31365 , n31372 );
xor ( n31374 , n31356 , n31357 );
xor ( n31375 , n31374 , n31359 );
buf ( n31376 , n31375 );
buf ( n31377 , n31376 );
not ( n31378 , n31377 );
buf ( n31379 , n31378 );
xor ( n31380 , n30888 , n30889 );
and ( n31381 , n31380 , n30891 );
and ( n31382 , n30888 , n30889 );
or ( n31383 , n31381 , n31382 );
buf ( n31384 , n31383 );
buf ( n31385 , n31384 );
not ( n31386 , n31385 );
buf ( n31387 , n31386 );
nand ( n31388 , n31379 , n31387 );
nand ( n31389 , n31373 , n31388 );
not ( n31390 , n31389 );
buf ( n31391 , n31390 );
nand ( n31392 , n31355 , n31391 );
buf ( n31393 , n31392 );
buf ( n31394 , n31393 );
not ( n31395 , n31394 );
buf ( n31396 , n31395 );
and ( n31397 , n31317 , n31320 , n31396 );
buf ( n31398 , n865 );
buf ( n31399 , n4842 );
xor ( n31400 , n31398 , n31399 );
buf ( n31401 , n4365 );
and ( n31402 , n31400 , n31401 );
and ( n31403 , n31398 , n31399 );
or ( n31404 , n31402 , n31403 );
buf ( n31405 , n31404 );
buf ( n31406 , n31405 );
xor ( n31407 , n31040 , n31041 );
xor ( n31408 , n31407 , n31043 );
buf ( n31409 , n31408 );
buf ( n31410 , n31409 );
nor ( n31411 , n31406 , n31410 );
buf ( n31412 , n31411 );
xor ( n31413 , n31398 , n31399 );
xor ( n31414 , n31413 , n31401 );
buf ( n31415 , n31414 );
xor ( n31416 , n31239 , n31240 );
and ( n31417 , n31416 , n31242 );
and ( n31418 , n31239 , n31240 );
or ( n31419 , n31417 , n31418 );
buf ( n31420 , n31419 );
nor ( n31421 , n31415 , n31420 );
nor ( n31422 , n31412 , n31421 );
buf ( n31423 , n31422 );
buf ( n31424 , n31423 );
buf ( n31425 , n31424 );
nand ( n31426 , n31283 , n31397 , n31425 );
buf ( n31427 , n31412 );
not ( n31428 , n31427 );
buf ( n31429 , n31428 );
buf ( n31430 , n31298 );
buf ( n31431 , n31430 );
buf ( n31432 , n31431 );
buf ( n31433 , n31432 );
not ( n31434 , n31433 );
buf ( n31435 , n31434 );
or ( n31436 , n31415 , n31420 );
and ( n31437 , n31429 , n31435 , n31436 );
buf ( n31438 , n31298 );
not ( n31439 , n31438 );
buf ( n31440 , n31302 );
buf ( n31441 , n31308 );
nand ( n31442 , n31440 , n31441 );
buf ( n31443 , n31442 );
buf ( n31444 , n31443 );
not ( n31445 , n31444 );
and ( n31446 , n31439 , n31445 );
buf ( n31447 , n31286 );
buf ( n31448 , n31295 );
and ( n31449 , n31447 , n31448 );
buf ( n31450 , n31449 );
buf ( n31451 , n31450 );
nor ( n31452 , n31446 , n31451 );
buf ( n31453 , n31452 );
buf ( n31454 , n31453 );
not ( n31455 , n31454 );
buf ( n31456 , n31455 );
buf ( n31457 , n31456 );
not ( n31458 , n31457 );
buf ( n31459 , n31354 );
not ( n31460 , n31459 );
buf ( n31461 , n31376 );
buf ( n31462 , n31384 );
nand ( n31463 , n31461 , n31462 );
buf ( n31464 , n31463 );
buf ( n31465 , n31464 );
not ( n31466 , n31465 );
buf ( n31467 , n31466 );
buf ( n31468 , n31467 );
not ( n31469 , n31468 );
nand ( n31470 , n31371 , n31364 );
buf ( n31471 , n31470 );
not ( n31472 , n31471 );
or ( n31473 , n31469 , n31472 );
buf ( n31474 , n31371 );
not ( n31475 , n31474 );
buf ( n31476 , n31363 );
nand ( n31477 , n31475 , n31476 );
buf ( n31478 , n31477 );
buf ( n31479 , n31478 );
nand ( n31480 , n31473 , n31479 );
buf ( n31481 , n31480 );
buf ( n31482 , n31481 );
not ( n31483 , n31482 );
or ( n31484 , n31460 , n31483 );
buf ( n31485 , n31335 );
not ( n31486 , n31485 );
buf ( n31487 , n31486 );
buf ( n31488 , n31487 );
buf ( n31489 , n31348 );
buf ( n31490 , n31344 );
and ( n31491 , n31489 , n31490 );
buf ( n31492 , n31491 );
buf ( n31493 , n31492 );
and ( n31494 , n31488 , n31493 );
buf ( n31495 , n31332 );
buf ( n31496 , n31328 );
nand ( n31497 , n31495 , n31496 );
buf ( n31498 , n31497 );
buf ( n31499 , n31498 );
not ( n31500 , n31499 );
buf ( n31501 , n31500 );
buf ( n31502 , n31501 );
nor ( n31503 , n31494 , n31502 );
buf ( n31504 , n31503 );
buf ( n31505 , n31504 );
nand ( n31506 , n31484 , n31505 );
buf ( n31507 , n31506 );
buf ( n31508 , n31507 );
buf ( n31509 , n31207 );
buf ( n31510 , n31216 );
nand ( n31511 , n31509 , n31510 );
buf ( n31512 , n31511 );
buf ( n31513 , n31512 );
not ( n31514 , n31513 );
buf ( n31515 , n31514 );
buf ( n31516 , n31515 );
not ( n31517 , n31516 );
buf ( n31518 , n31203 );
not ( n31519 , n31518 );
buf ( n31520 , n31519 );
buf ( n31521 , n31520 );
not ( n31522 , n31521 );
or ( n31523 , n31517 , n31522 );
buf ( n31524 , n31191 );
buf ( n31525 , n31524 );
buf ( n31526 , n31525 );
buf ( n31527 , n31526 );
buf ( n31528 , n31200 );
nand ( n31529 , n31527 , n31528 );
buf ( n31530 , n31529 );
buf ( n31531 , n31530 );
nand ( n31532 , n31523 , n31531 );
buf ( n31533 , n31532 );
buf ( n31534 , n31533 );
nor ( n31535 , n31508 , n31534 );
buf ( n31536 , n31535 );
buf ( n31537 , n31536 );
buf ( n31538 , n31396 );
nor ( n31539 , n30902 , n30716 );
not ( n31540 , n31539 );
not ( n31541 , n30860 );
or ( n31542 , n31540 , n31541 );
not ( n31543 , n30872 );
not ( n31544 , n30899 );
or ( n31545 , n31543 , n31544 );
nand ( n31546 , n31545 , n30913 );
not ( n31547 , n31546 );
nand ( n31548 , n31542 , n31547 );
buf ( n31549 , n31548 );
nand ( n31550 , n31538 , n31549 );
buf ( n31551 , n31550 );
buf ( n31552 , n31551 );
nand ( n31553 , n31458 , n31537 , n31552 );
buf ( n31554 , n31553 );
buf ( n31555 , n31456 );
not ( n31556 , n31555 );
buf ( n31557 , n31533 );
buf ( n31558 , n31228 );
nor ( n31559 , n31557 , n31558 );
buf ( n31560 , n31559 );
buf ( n31561 , n31560 );
nand ( n31562 , n31556 , n31561 );
buf ( n31563 , n31562 );
buf ( n31564 , n31450 );
not ( n31565 , n31564 );
buf ( n31566 , n31565 );
buf ( n31567 , n31566 );
buf ( n31568 , n31311 );
nand ( n31569 , n31567 , n31568 );
buf ( n31570 , n31569 );
buf ( n31571 , n31570 );
buf ( n31572 , n31250 );
not ( n31573 , n31572 );
buf ( n31574 , n31573 );
buf ( n31575 , n31574 );
buf ( n31576 , n31270 );
not ( n31577 , n31576 );
buf ( n31578 , n31577 );
buf ( n31579 , n31578 );
nor ( n31580 , n31575 , n31579 );
buf ( n31581 , n31580 );
buf ( n31582 , n31581 );
and ( n31583 , n31571 , n31582 );
buf ( n31584 , n31583 );
nand ( n31585 , n31437 , n31554 , n31563 , n31584 );
not ( n31586 , n31422 );
buf ( n31587 , n31236 );
not ( n31588 , n31587 );
buf ( n31589 , n31247 );
nand ( n31590 , n31588 , n31589 );
buf ( n31591 , n31590 );
buf ( n31592 , n31591 );
not ( n31593 , n31592 );
buf ( n31594 , n31264 );
buf ( n31595 , n31259 );
nand ( n31596 , n31594 , n31595 );
buf ( n31597 , n31596 );
buf ( n31598 , n31597 );
not ( n31599 , n31598 );
buf ( n31600 , n31599 );
buf ( n31601 , n31600 );
not ( n31602 , n31601 );
or ( n31603 , n31593 , n31602 );
buf ( n31604 , n31236 );
buf ( n31605 , n31244 );
buf ( n31606 , n31605 );
buf ( n31607 , n31606 );
buf ( n31608 , n31607 );
nand ( n31609 , n31604 , n31608 );
buf ( n31610 , n31609 );
buf ( n31611 , n31610 );
nand ( n31612 , n31603 , n31611 );
buf ( n31613 , n31612 );
not ( n31614 , n31613 );
or ( n31615 , n31586 , n31614 );
buf ( n31616 , n31415 );
buf ( n31617 , n31420 );
nand ( n31618 , n31616 , n31617 );
buf ( n31619 , n31618 );
not ( n31620 , n31619 );
not ( n31621 , n31412 );
and ( n31622 , n31620 , n31621 );
buf ( n31623 , n31409 );
buf ( n31624 , n31623 );
buf ( n31625 , n31624 );
and ( n31626 , n31625 , n31405 );
nor ( n31627 , n31622 , n31626 );
nand ( n31628 , n31615 , n31627 );
not ( n31629 , n31628 );
nand ( n31630 , n31426 , n31585 , n31629 );
not ( n31631 , n31630 );
not ( n31632 , n31631 );
buf ( n31633 , n31632 );
not ( n31634 , n31633 );
or ( n31635 , n31185 , n31634 );
buf ( n31636 , n31039 );
not ( n31637 , n31636 );
buf ( n31638 , n31107 );
buf ( n31639 , n31109 );
nand ( n31640 , n31638 , n31639 );
buf ( n31641 , n31640 );
buf ( n31642 , n31641 );
buf ( n31643 , n31092 );
buf ( n31644 , n31094 );
nand ( n31645 , n31643 , n31644 );
buf ( n31646 , n31645 );
buf ( n31647 , n31646 );
and ( n31648 , n31642 , n31647 );
buf ( n31649 , n31648 );
buf ( n31650 , n31649 );
not ( n31651 , n31650 );
nand ( n31652 , n31071 , n31076 );
nand ( n31653 , n31060 , n31071 , n31047 );
nand ( n31654 , n31652 , n31653 );
nand ( n31655 , n31095 , n31093 );
nand ( n31656 , n31654 , n31655 );
buf ( n31657 , n31656 );
not ( n31658 , n31657 );
or ( n31659 , n31651 , n31658 );
buf ( n31660 , n31177 );
buf ( n31661 , n31107 );
buf ( n31662 , n31109 );
nor ( n31663 , n31661 , n31662 );
buf ( n31664 , n31663 );
buf ( n31665 , n31664 );
nor ( n31666 , n31660 , n31665 );
buf ( n31667 , n31666 );
buf ( n31668 , n31667 );
nand ( n31669 , n31659 , n31668 );
buf ( n31670 , n31669 );
buf ( n31671 , n31158 );
buf ( n31672 , n31671 );
buf ( n31673 , n31672 );
buf ( n31674 , n31673 );
buf ( n31675 , n31130 );
buf ( n31676 , n31116 );
nand ( n31677 , n31675 , n31676 );
buf ( n31678 , n31677 );
buf ( n31679 , n31678 );
or ( n31680 , n31674 , n31679 );
buf ( n31681 , n31153 );
buf ( n31682 , n31681 );
buf ( n31683 , n31682 );
buf ( n31684 , n31683 );
buf ( n31685 , n31157 );
buf ( n31686 , n31685 );
buf ( n31687 , n31686 );
buf ( n31688 , n31687 );
nand ( n31689 , n31684 , n31688 );
buf ( n31690 , n31689 );
buf ( n31691 , n31690 );
nand ( n31692 , n31680 , n31691 );
buf ( n31693 , n31692 );
not ( n31694 , n31693 );
buf ( n31695 , n31162 );
buf ( n31696 , n31166 );
and ( n31697 , n31695 , n31696 );
buf ( n31698 , n31697 );
buf ( n31699 , n31698 );
not ( n31700 , n31699 );
buf ( n31701 , n31174 );
not ( n31702 , n31701 );
or ( n31703 , n31700 , n31702 );
buf ( n31704 , n31173 );
not ( n31705 , n31704 );
buf ( n31706 , n31171 );
nand ( n31707 , n31705 , n31706 );
buf ( n31708 , n31707 );
buf ( n31709 , n31708 );
nand ( n31710 , n31703 , n31709 );
buf ( n31711 , n31710 );
not ( n31712 , n31116 );
not ( n31713 , n31130 );
and ( n31714 , n31712 , n31713 );
nor ( n31715 , n31714 , n31673 );
nand ( n31716 , n31711 , n31715 );
nand ( n31717 , n31694 , n31716 );
buf ( n31718 , n31717 );
not ( n31719 , n31718 );
buf ( n31720 , n31719 );
nand ( n31721 , n31670 , n31720 );
buf ( n31722 , n31721 );
not ( n31723 , n31722 );
or ( n31724 , n31637 , n31723 );
buf ( n31725 , n30976 );
not ( n31726 , n31725 );
not ( n31727 , n30990 );
nand ( n31728 , n31727 , n30982 );
buf ( n31729 , n31728 );
not ( n31730 , n31729 );
buf ( n31731 , n31004 );
buf ( n31732 , n31006 );
and ( n31733 , n31731 , n31732 );
buf ( n31734 , n31733 );
buf ( n31735 , n31734 );
not ( n31736 , n31735 );
or ( n31737 , n31730 , n31736 );
buf ( n31738 , n30985 );
buf ( n31739 , n30990 );
nand ( n31740 , n31738 , n31739 );
buf ( n31741 , n31740 );
buf ( n31742 , n31741 );
nand ( n31743 , n31737 , n31742 );
buf ( n31744 , n31743 );
buf ( n31745 , n31744 );
buf ( n31746 , n31031 );
nand ( n31747 , n31745 , n31746 );
buf ( n31748 , n31747 );
buf ( n31749 , n31748 );
not ( n31750 , n31029 );
buf ( n31751 , n31015 );
buf ( n31752 , n31017 );
nor ( n31753 , n31751 , n31752 );
buf ( n31754 , n31753 );
not ( n31755 , n31754 );
or ( n31756 , n31750 , n31755 );
or ( n31757 , n31026 , n31024 );
nand ( n31758 , n31756 , n31757 );
not ( n31759 , n31758 );
buf ( n31760 , n31759 );
nand ( n31761 , n31749 , n31760 );
buf ( n31762 , n31761 );
buf ( n31763 , n31762 );
not ( n31764 , n31763 );
or ( n31765 , n31726 , n31764 );
nor ( n31766 , n30965 , n30973 );
buf ( n31767 , n31766 );
not ( n31768 , n31767 );
buf ( n31769 , n31768 );
buf ( n31770 , n31769 );
nand ( n31771 , n31765 , n31770 );
buf ( n31772 , n31771 );
buf ( n31773 , n31772 );
not ( n31774 , n31773 );
buf ( n31775 , n31774 );
buf ( n31776 , n31775 );
nand ( n31777 , n31724 , n31776 );
buf ( n31778 , n31777 );
buf ( n31779 , n31778 );
not ( n31780 , n31779 );
buf ( n31781 , n31780 );
buf ( n31782 , n31781 );
nand ( n31783 , n31635 , n31782 );
buf ( n31784 , n31783 );
buf ( n31785 , n31784 );
not ( n31786 , n15923 );
not ( n31787 , n15650 );
or ( n31788 , n31786 , n31787 );
buf ( n31789 , n15930 );
buf ( n31790 , n15920 );
nand ( n31791 , n31789 , n31790 );
buf ( n31792 , n31791 );
nand ( n31793 , n31788 , n31792 );
and ( n31794 , n30967 , n30968 );
buf ( n31795 , n31794 );
or ( n31796 , n31793 , n31795 );
buf ( n31797 , n31796 );
nand ( n31798 , n31795 , n31793 );
buf ( n31799 , n31798 );
nand ( n31800 , n31797 , n31799 );
buf ( n31801 , n31800 );
buf ( n31802 , n31801 );
not ( n31803 , n31802 );
buf ( n31804 , n31803 );
buf ( n31805 , n31804 );
and ( n31806 , n31785 , n31805 );
not ( n31807 , n31785 );
buf ( n31808 , n31801 );
and ( n31809 , n31807 , n31808 );
nor ( n31810 , n31806 , n31809 );
buf ( n31811 , n31810 );
and ( n31812 , n1152 , n31811 );
not ( n31813 , n1152 );
and ( n31814 , n31813 , n16776 );
nor ( n31815 , n31812 , n31814 );
nand ( n31816 , n18421 , n831 );
buf ( n31817 , n31630 );
nor ( n31818 , n31181 , n31036 );
and ( n31819 , n31817 , n31818 );
buf ( n31820 , n31033 );
not ( n31821 , n31820 );
buf ( n31822 , n31721 );
not ( n31823 , n31822 );
or ( n31824 , n31821 , n31823 );
buf ( n31825 , n31762 );
not ( n31826 , n31825 );
buf ( n31827 , n31826 );
buf ( n31828 , n31827 );
nand ( n31829 , n31824 , n31828 );
buf ( n31830 , n31829 );
nor ( n31831 , n31819 , n31830 );
buf ( n31832 , n31831 );
buf ( n31833 , n30976 );
buf ( n31834 , n31769 );
nand ( n31835 , n31833 , n31834 );
buf ( n31836 , n31835 );
not ( n31837 , n31836 );
nand ( n31838 , n31837 , n1152 );
buf ( n31839 , n31838 );
and ( n31840 , n31832 , n31839 );
not ( n31841 , n31832 );
nand ( n31842 , n31836 , n1152 );
buf ( n31843 , n31842 );
and ( n31844 , n31841 , n31843 );
or ( n31845 , n31840 , n31844 );
buf ( n31846 , n31845 );
nand ( n31847 , n31816 , n31846 );
buf ( n31848 , n8894 );
not ( n31849 , n31848 );
buf ( n31850 , n10359 );
not ( n31851 , n31850 );
or ( n31852 , n31849 , n31851 );
not ( n31853 , n8427 );
not ( n31854 , n8772 );
or ( n31855 , n31853 , n31854 );
nand ( n31856 , n31855 , n8797 );
buf ( n31857 , n31856 );
not ( n31858 , n31857 );
buf ( n31859 , n31858 );
buf ( n31860 , n31859 );
nand ( n31861 , n31852 , n31860 );
buf ( n31862 , n31861 );
nand ( n31863 , n18430 , n18434 );
not ( n31864 , n31863 );
and ( n31865 , n31862 , n31864 );
not ( n31866 , n31862 );
and ( n31867 , n31866 , n31863 );
nor ( n31868 , n31865 , n31867 );
nand ( n31869 , n31868 , n831 );
buf ( n31870 , n31282 );
not ( n31871 , n31870 );
buf ( n31872 , n30780 );
not ( n31873 , n31872 );
buf ( n31874 , n30226 );
not ( n31875 , n31874 );
or ( n31876 , n31873 , n31875 );
buf ( n31877 , n30833 );
nand ( n31878 , n31876 , n31877 );
buf ( n31879 , n31878 );
buf ( n31880 , n31879 );
not ( n31881 , n31880 );
or ( n31882 , n31871 , n31881 );
buf ( n31883 , n31548 );
not ( n31884 , n31883 );
buf ( n31885 , n31884 );
buf ( n31886 , n31885 );
nand ( n31887 , n31882 , n31886 );
buf ( n31888 , n31887 );
buf ( n31889 , n31888 );
buf ( n31890 , n31388 );
buf ( n31891 , n31890 );
buf ( n31892 , n31891 );
buf ( n31893 , n31892 );
buf ( n31894 , n31464 );
buf ( n31895 , n31894 );
buf ( n31896 , n31895 );
buf ( n31897 , n31896 );
nand ( n31898 , n31893 , n31897 );
buf ( n31899 , n31898 );
buf ( n31900 , n31899 );
not ( n31901 , n31900 );
buf ( n31902 , n31901 );
buf ( n31903 , n31902 );
and ( n31904 , n31889 , n31903 );
not ( n31905 , n31889 );
buf ( n31906 , n31899 );
and ( n31907 , n31905 , n31906 );
nor ( n31908 , n31904 , n31907 );
buf ( n31909 , n31908 );
nand ( n31910 , n31909 , n1152 );
nand ( n31911 , n31869 , n31910 );
not ( n31912 , n1152 );
not ( n31913 , n30959 );
not ( n31914 , n31879 );
or ( n31915 , n31913 , n31914 );
nand ( n31916 , n31915 , n30843 );
buf ( n31917 , n31916 );
buf ( n31918 , n30858 );
buf ( n31919 , n30847 );
nand ( n31920 , n31918 , n31919 );
buf ( n31921 , n31920 );
buf ( n31922 , n31921 );
not ( n31923 , n31922 );
buf ( n31924 , n31923 );
buf ( n31925 , n31924 );
and ( n31926 , n31917 , n31925 );
not ( n31927 , n31917 );
buf ( n31928 , n31921 );
and ( n31929 , n31927 , n31928 );
nor ( n31930 , n31926 , n31929 );
buf ( n31931 , n31930 );
not ( n31932 , n31931 );
or ( n31933 , n31912 , n31932 );
buf ( n31934 , n30933 );
not ( n31935 , n31934 );
buf ( n31936 , n18807 );
not ( n31937 , n31936 );
or ( n31938 , n31935 , n31937 );
buf ( n31939 , n8748 );
nand ( n31940 , n31938 , n31939 );
buf ( n31941 , n31940 );
buf ( n31942 , n31941 );
buf ( n31943 , n8766 );
buf ( n31944 , n8762 );
nand ( n31945 , n31943 , n31944 );
buf ( n31946 , n31945 );
buf ( n31947 , n31946 );
not ( n31948 , n31947 );
buf ( n31949 , n31948 );
buf ( n31950 , n31949 );
and ( n31951 , n31942 , n31950 );
not ( n31952 , n31942 );
buf ( n31953 , n31946 );
and ( n31954 , n31952 , n31953 );
nor ( n31955 , n31951 , n31954 );
buf ( n31956 , n31955 );
nand ( n31957 , n31956 , n831 );
nand ( n31958 , n31933 , n31957 );
buf ( n31959 , n31115 );
not ( n31960 , n31959 );
buf ( n31961 , n31426 );
buf ( n31962 , n31585 );
buf ( n31963 , n31629 );
nand ( n31964 , n31961 , n31962 , n31963 );
buf ( n31965 , n31964 );
buf ( n31966 , n31965 );
buf ( n31967 , n31966 );
buf ( n31968 , n31967 );
buf ( n31969 , n31968 );
not ( n31970 , n31969 );
or ( n31971 , n31960 , n31970 );
and ( n31972 , n31093 , n31095 );
nor ( n31973 , n31972 , n31112 );
not ( n31974 , n31973 );
not ( n31975 , n31654 );
or ( n31976 , n31974 , n31975 );
not ( n31977 , n31646 );
not ( n31978 , n31664 );
and ( n31979 , n31977 , n31978 );
not ( n31980 , n31641 );
nor ( n31981 , n31979 , n31980 );
nand ( n31982 , n31976 , n31981 );
buf ( n31983 , n31982 );
not ( n31984 , n31983 );
buf ( n31985 , n31984 );
buf ( n31986 , n31985 );
nand ( n31987 , n31971 , n31986 );
buf ( n31988 , n31987 );
buf ( n31989 , n31988 );
buf ( n31990 , n31167 );
not ( n31991 , n31990 );
buf ( n31992 , n31698 );
buf ( n31993 , n31992 );
not ( n31994 , n31993 );
buf ( n31995 , n31994 );
nand ( n31996 , n31991 , n31995 );
buf ( n31997 , n31996 );
not ( n31998 , n31997 );
buf ( n31999 , n31998 );
buf ( n32000 , n31999 );
and ( n32001 , n31989 , n32000 );
not ( n32002 , n31989 );
buf ( n32003 , n31996 );
and ( n32004 , n32002 , n32003 );
nor ( n32005 , n32001 , n32004 );
buf ( n32006 , n32005 );
nand ( n32007 , n32006 , n1152 );
or ( n32008 , n10070 , n10120 );
buf ( n32009 , n32008 );
not ( n32010 , n32009 );
buf ( n32011 , n10239 );
not ( n32012 , n32011 );
or ( n32013 , n32010 , n32012 );
buf ( n32014 , n10123 );
nand ( n32015 , n32013 , n32014 );
buf ( n32016 , n32015 );
buf ( n32017 , n32016 );
buf ( n32018 , n10132 );
buf ( n32019 , n10066 );
not ( n32020 , n32019 );
buf ( n32021 , n32020 );
buf ( n32022 , n32021 );
nand ( n32023 , n32018 , n32022 );
buf ( n32024 , n32023 );
buf ( n32025 , n32024 );
not ( n32026 , n32025 );
buf ( n32027 , n32026 );
buf ( n32028 , n32027 );
and ( n32029 , n32017 , n32028 );
not ( n32030 , n32017 );
buf ( n32031 , n32024 );
and ( n32032 , n32030 , n32031 );
nor ( n32033 , n32029 , n32032 );
buf ( n32034 , n32033 );
nand ( n32035 , n32034 , n831 );
nand ( n32036 , n18801 , n831 );
buf ( n32037 , n30439 );
buf ( n32038 , n29916 );
not ( n32039 , n32038 );
buf ( n32040 , n32039 );
buf ( n32041 , n32040 );
buf ( n32042 , n30062 );
nand ( n32043 , n32041 , n32042 );
buf ( n32044 , n32043 );
buf ( n32045 , n32044 );
and ( n32046 , n32037 , n32045 );
not ( n32047 , n32037 );
buf ( n32048 , n32044 );
not ( n32049 , n32048 );
buf ( n32050 , n32049 );
buf ( n32051 , n32050 );
and ( n32052 , n32047 , n32051 );
nor ( n32053 , n32046 , n32052 );
buf ( n32054 , n32053 );
nand ( n32055 , n32054 , n1152 );
nand ( n32056 , n16709 , n831 );
nand ( n32057 , n18641 , n831 );
not ( n32058 , n30701 );
not ( n32059 , n31879 );
or ( n32060 , n32058 , n32059 );
not ( n32061 , n30861 );
nand ( n32062 , n32060 , n32061 );
buf ( n32063 , n32062 );
buf ( n32064 , n30875 );
not ( n32065 , n32064 );
buf ( n32066 , n30719 );
nand ( n32067 , n32065 , n32066 );
buf ( n32068 , n32067 );
buf ( n32069 , n32068 );
not ( n32070 , n32069 );
buf ( n32071 , n32070 );
buf ( n32072 , n32071 );
and ( n32073 , n32063 , n32072 );
not ( n32074 , n32063 );
buf ( n32075 , n32068 );
and ( n32076 , n32074 , n32075 );
nor ( n32077 , n32073 , n32076 );
buf ( n32078 , n32077 );
nand ( n32079 , n32078 , n1152 );
not ( n32080 , n31721 );
buf ( n32081 , n31314 );
not ( n32082 , n32081 );
buf ( n32083 , n31533 );
not ( n32084 , n32083 );
or ( n32085 , n32082 , n32084 );
buf ( n32086 , n31453 );
nand ( n32087 , n32085 , n32086 );
buf ( n32088 , n32087 );
buf ( n32089 , n32088 );
buf ( n32090 , n32089 );
buf ( n32091 , n32090 );
nor ( n32092 , n31628 , n32091 );
not ( n32093 , n32092 );
or ( n32094 , n31507 , n31396 );
buf ( n32095 , n31314 );
buf ( n32096 , n31222 );
and ( n32097 , n32095 , n32096 );
buf ( n32098 , n32097 );
buf ( n32099 , n32098 );
buf ( n32100 , n32099 );
buf ( n32101 , n32100 );
buf ( n32102 , n31320 );
buf ( n32103 , n31282 );
nand ( n32104 , n32102 , n32103 );
buf ( n32105 , n32104 );
buf ( n32106 , n32105 );
buf ( n32107 , n31507 );
not ( n32108 , n32107 );
buf ( n32109 , n32108 );
buf ( n32110 , n32109 );
buf ( n32111 , n31885 );
nand ( n32112 , n32106 , n32110 , n32111 );
buf ( n32113 , n32112 );
nand ( n32114 , n32094 , n32101 , n32113 );
not ( n32115 , n32114 );
or ( n32116 , n32093 , n32115 );
nand ( n32117 , n31436 , n31429 );
not ( n32118 , n32117 );
buf ( n32119 , n31581 );
nand ( n32120 , n32118 , n32119 );
and ( n32121 , n32120 , n31629 );
nor ( n32122 , n32121 , n31181 );
nand ( n32123 , n32116 , n32122 );
nand ( n32124 , n32080 , n32123 );
buf ( n32125 , n32124 );
buf ( n32126 , n31009 );
not ( n32127 , n32126 );
buf ( n32128 , n32127 );
buf ( n32129 , n32128 );
buf ( n32130 , n31734 );
not ( n32131 , n32130 );
buf ( n32132 , n32131 );
buf ( n32133 , n32132 );
nand ( n32134 , n32129 , n32133 );
buf ( n32135 , n32134 );
buf ( n32136 , n32135 );
xnor ( n32137 , n32125 , n32136 );
buf ( n32138 , n32137 );
nand ( n32139 , n32138 , n1152 );
buf ( n32140 , n31174 );
not ( n32141 , n32140 );
nor ( n32142 , n32141 , n31990 );
buf ( n32143 , n32142 );
buf ( n32144 , n31136 );
buf ( n32145 , n32144 );
buf ( n32146 , n32145 );
buf ( n32147 , n32146 );
nand ( n32148 , n32143 , n32147 );
buf ( n32149 , n32148 );
buf ( n32150 , n32149 );
buf ( n32151 , n31114 );
nor ( n32152 , n32150 , n32151 );
buf ( n32153 , n32152 );
buf ( n32154 , n32153 );
not ( n32155 , n32154 );
buf ( n32156 , n31632 );
not ( n32157 , n32156 );
or ( n32158 , n32155 , n32157 );
buf ( n32159 , n31982 );
not ( n32160 , n32159 );
not ( n32161 , n32149 );
buf ( n32162 , n32161 );
not ( n32163 , n32162 );
or ( n32164 , n32160 , n32163 );
buf ( n32165 , n32146 );
not ( n32166 , n32165 );
buf ( n32167 , n31711 );
buf ( n32168 , n32167 );
buf ( n32169 , n32168 );
buf ( n32170 , n32169 );
not ( n32171 , n32170 );
or ( n32172 , n32166 , n32171 );
buf ( n32173 , n31678 );
nand ( n32174 , n32172 , n32173 );
buf ( n32175 , n32174 );
buf ( n32176 , n32175 );
not ( n32177 , n32176 );
buf ( n32178 , n32177 );
buf ( n32179 , n32178 );
nand ( n32180 , n32164 , n32179 );
buf ( n32181 , n32180 );
buf ( n32182 , n32181 );
not ( n32183 , n32182 );
buf ( n32184 , n32183 );
buf ( n32185 , n32184 );
nand ( n32186 , n32158 , n32185 );
buf ( n32187 , n32186 );
buf ( n32188 , n32187 );
buf ( n32189 , n31673 );
not ( n32190 , n32189 );
buf ( n32191 , n31690 );
nand ( n32192 , n32190 , n32191 );
buf ( n32193 , n32192 );
buf ( n32194 , n32193 );
not ( n32195 , n32194 );
buf ( n32196 , n32195 );
buf ( n32197 , n32196 );
and ( n32198 , n32188 , n32197 );
not ( n32199 , n32188 );
buf ( n32200 , n32193 );
and ( n32201 , n32199 , n32200 );
nor ( n32202 , n32198 , n32201 );
buf ( n32203 , n32202 );
nand ( n32204 , n32203 , n1152 );
xor ( n32205 , n19715 , n19760 );
xor ( n32206 , n32205 , n19772 );
buf ( n32207 , n32206 );
buf ( n32208 , n19797 );
buf ( n32209 , n844 );
buf ( n32210 , n870 );
xor ( n32211 , n32209 , n32210 );
buf ( n32212 , n32211 );
buf ( n32213 , n32212 );
not ( n32214 , n32213 );
buf ( n32215 , n19125 );
not ( n32216 , n32215 );
or ( n32217 , n32214 , n32216 );
buf ( n32218 , n19134 );
buf ( n32219 , n19802 );
nand ( n32220 , n32218 , n32219 );
buf ( n32221 , n32220 );
buf ( n32222 , n32221 );
nand ( n32223 , n32217 , n32222 );
buf ( n32224 , n32223 );
buf ( n32225 , n32224 );
xor ( n32226 , n32208 , n32225 );
buf ( n32227 , n851 );
buf ( n32228 , n864 );
xor ( n32229 , n32227 , n32228 );
buf ( n32230 , n32229 );
buf ( n32231 , n32230 );
not ( n32232 , n32231 );
buf ( n32233 , n19013 );
not ( n32234 , n32233 );
or ( n32235 , n32232 , n32234 );
buf ( n32236 , n19030 );
buf ( n32237 , n19968 );
nand ( n32238 , n32236 , n32237 );
buf ( n32239 , n32238 );
buf ( n32240 , n32239 );
nand ( n32241 , n32235 , n32240 );
buf ( n32242 , n32241 );
buf ( n32243 , n32242 );
not ( n32244 , n32243 );
buf ( n32245 , n835 );
buf ( n32246 , n880 );
xor ( n32247 , n32245 , n32246 );
buf ( n32248 , n32247 );
buf ( n32249 , n32248 );
not ( n32250 , n32249 );
buf ( n32251 , n18850 );
not ( n32252 , n32251 );
or ( n32253 , n32250 , n32252 );
buf ( n32254 , n18860 );
buf ( n32255 , n19790 );
nand ( n32256 , n32254 , n32255 );
buf ( n32257 , n32256 );
buf ( n32258 , n32257 );
nand ( n32259 , n32253 , n32258 );
buf ( n32260 , n32259 );
buf ( n32261 , n32260 );
not ( n32262 , n32261 );
or ( n32263 , n32244 , n32262 );
buf ( n32264 , n32260 );
buf ( n32265 , n32242 );
or ( n32266 , n32264 , n32265 );
buf ( n32267 , n849 );
buf ( n32268 , n866 );
xor ( n32269 , n32267 , n32268 );
buf ( n32270 , n32269 );
buf ( n32271 , n32270 );
not ( n32272 , n32271 );
buf ( n32273 , n18931 );
not ( n32274 , n32273 );
or ( n32275 , n32272 , n32274 );
buf ( n32276 , n18944 );
buf ( n32277 , n19846 );
nand ( n32278 , n32276 , n32277 );
buf ( n32279 , n32278 );
buf ( n32280 , n32279 );
nand ( n32281 , n32275 , n32280 );
buf ( n32282 , n32281 );
buf ( n32283 , n32282 );
nand ( n32284 , n32266 , n32283 );
buf ( n32285 , n32284 );
buf ( n32286 , n32285 );
nand ( n32287 , n32263 , n32286 );
buf ( n32288 , n32287 );
buf ( n32289 , n32288 );
and ( n32290 , n32226 , n32289 );
and ( n32291 , n32208 , n32225 );
or ( n32292 , n32290 , n32291 );
buf ( n32293 , n32292 );
buf ( n32294 , n32293 );
xor ( n32295 , n19801 , n19815 );
xor ( n32296 , n32295 , n19833 );
buf ( n32297 , n32296 );
buf ( n32298 , n32297 );
xor ( n32299 , n32294 , n32298 );
buf ( n32300 , n852 );
buf ( n32301 , n864 );
and ( n32302 , n32300 , n32301 );
buf ( n32303 , n32302 );
buf ( n32304 , n32303 );
buf ( n32305 , n843 );
buf ( n32306 , n872 );
xor ( n32307 , n32305 , n32306 );
buf ( n32308 , n32307 );
buf ( n32309 , n32308 );
not ( n32310 , n32309 );
buf ( n32311 , n19230 );
not ( n32312 , n32311 );
or ( n32313 , n32310 , n32312 );
buf ( n32314 , n19235 );
buf ( n32315 , n19922 );
nand ( n32316 , n32314 , n32315 );
buf ( n32317 , n32316 );
buf ( n32318 , n32317 );
nand ( n32319 , n32313 , n32318 );
buf ( n32320 , n32319 );
buf ( n32321 , n32320 );
xor ( n32322 , n32304 , n32321 );
buf ( n32323 , n841 );
buf ( n32324 , n874 );
xor ( n32325 , n32323 , n32324 );
buf ( n32326 , n32325 );
buf ( n32327 , n32326 );
not ( n32328 , n32327 );
buf ( n32329 , n18977 );
not ( n32330 , n32329 );
or ( n32331 , n32328 , n32330 );
buf ( n32332 , n18987 );
buf ( n32333 , n19986 );
nand ( n32334 , n32332 , n32333 );
buf ( n32335 , n32334 );
buf ( n32336 , n32335 );
nand ( n32337 , n32331 , n32336 );
buf ( n32338 , n32337 );
buf ( n32339 , n32338 );
and ( n32340 , n32322 , n32339 );
and ( n32341 , n32304 , n32321 );
or ( n32342 , n32340 , n32341 );
buf ( n32343 , n32342 );
buf ( n32344 , n32343 );
buf ( n32345 , n847 );
buf ( n32346 , n868 );
xor ( n32347 , n32345 , n32346 );
buf ( n32348 , n32347 );
buf ( n32349 , n32348 );
not ( n32350 , n32349 );
buf ( n32351 , n18887 );
not ( n32352 , n32351 );
or ( n32353 , n32350 , n32352 );
buf ( n32354 , n18892 );
buf ( n32355 , n19860 );
nand ( n32356 , n32354 , n32355 );
buf ( n32357 , n32356 );
buf ( n32358 , n32357 );
nand ( n32359 , n32353 , n32358 );
buf ( n32360 , n32359 );
buf ( n32361 , n32360 );
buf ( n32362 , n839 );
buf ( n32363 , n876 );
xor ( n32364 , n32362 , n32363 );
buf ( n32365 , n32364 );
buf ( n32366 , n32365 );
not ( n32367 , n32366 );
buf ( n32368 , n19077 );
not ( n32369 , n32368 );
or ( n32370 , n32367 , n32369 );
buf ( n32371 , n19085 );
buf ( n32372 , n19875 );
nand ( n32373 , n32371 , n32372 );
buf ( n32374 , n32373 );
buf ( n32375 , n32374 );
nand ( n32376 , n32370 , n32375 );
buf ( n32377 , n32376 );
buf ( n32378 , n32377 );
xor ( n32379 , n32361 , n32378 );
buf ( n32380 , n845 );
buf ( n32381 , n870 );
xor ( n32382 , n32380 , n32381 );
buf ( n32383 , n32382 );
buf ( n32384 , n32383 );
not ( n32385 , n32384 );
buf ( n32386 , n19125 );
not ( n32387 , n32386 );
or ( n32388 , n32385 , n32387 );
buf ( n32389 , n19134 );
buf ( n32390 , n32212 );
nand ( n32391 , n32389 , n32390 );
buf ( n32392 , n32391 );
buf ( n32393 , n32392 );
nand ( n32394 , n32388 , n32393 );
buf ( n32395 , n32394 );
buf ( n32396 , n32395 );
and ( n32397 , n32379 , n32396 );
and ( n32398 , n32361 , n32378 );
or ( n32399 , n32397 , n32398 );
buf ( n32400 , n32399 );
buf ( n32401 , n32400 );
xor ( n32402 , n32344 , n32401 );
buf ( n32403 , n25022 );
buf ( n32404 , n25263 );
or ( n32405 , n32403 , n32404 );
buf ( n32406 , n884 );
nand ( n32407 , n32405 , n32406 );
buf ( n32408 , n32407 );
buf ( n32409 , n32408 );
xor ( n32410 , n882 , n833 );
buf ( n32411 , n32410 );
not ( n32412 , n32411 );
buf ( n32413 , n26534 );
not ( n32414 , n32413 );
or ( n32415 , n32412 , n32414 );
buf ( n32416 , n19910 );
buf ( n32417 , n19897 );
nand ( n32418 , n32416 , n32417 );
buf ( n32419 , n32418 );
buf ( n32420 , n32419 );
nand ( n32421 , n32415 , n32420 );
buf ( n32422 , n32421 );
buf ( n32423 , n32422 );
xor ( n32424 , n32409 , n32423 );
buf ( n32425 , n837 );
buf ( n32426 , n878 );
xor ( n32427 , n32425 , n32426 );
buf ( n32428 , n32427 );
buf ( n32429 , n32428 );
not ( n32430 , n32429 );
buf ( n32431 , n19479 );
not ( n32432 , n32431 );
or ( n32433 , n32430 , n32432 );
buf ( n32434 , n19265 );
buf ( n32435 , n19940 );
nand ( n32436 , n32434 , n32435 );
buf ( n32437 , n32436 );
buf ( n32438 , n32437 );
nand ( n32439 , n32433 , n32438 );
buf ( n32440 , n32439 );
buf ( n32441 , n32440 );
and ( n32442 , n32424 , n32441 );
and ( n32443 , n32409 , n32423 );
or ( n32444 , n32442 , n32443 );
buf ( n32445 , n32444 );
buf ( n32446 , n32445 );
and ( n32447 , n32402 , n32446 );
and ( n32448 , n32344 , n32401 );
or ( n32449 , n32447 , n32448 );
buf ( n32450 , n32449 );
buf ( n32451 , n32450 );
and ( n32452 , n32299 , n32451 );
and ( n32453 , n32294 , n32298 );
or ( n32454 , n32452 , n32453 );
buf ( n32455 , n32454 );
xor ( n32456 , n19838 , n19841 );
xor ( n32457 , n32456 , n20009 );
buf ( n32458 , n32457 );
xor ( n32459 , n32455 , n32458 );
xor ( n32460 , n19918 , n19935 );
xor ( n32461 , n32460 , n19953 );
buf ( n32462 , n32461 );
buf ( n32463 , n32462 );
xor ( n32464 , n19859 , n19873 );
xor ( n32465 , n32464 , n19888 );
buf ( n32466 , n32465 );
buf ( n32467 , n32466 );
or ( n32468 , n32463 , n32467 );
xor ( n32469 , n19964 , n19981 );
xor ( n32470 , n32469 , n19999 );
buf ( n32471 , n32470 );
buf ( n32472 , n32471 );
nand ( n32473 , n32468 , n32472 );
buf ( n32474 , n32473 );
buf ( n32475 , n32474 );
buf ( n32476 , n32462 );
buf ( n32477 , n32466 );
nand ( n32478 , n32476 , n32477 );
buf ( n32479 , n32478 );
buf ( n32480 , n32479 );
nand ( n32481 , n32475 , n32480 );
buf ( n32482 , n32481 );
buf ( n32483 , n32482 );
xor ( n32484 , n19893 , n19958 );
xor ( n32485 , n32484 , n20004 );
buf ( n32486 , n32485 );
buf ( n32487 , n32486 );
xor ( n32488 , n32483 , n32487 );
xor ( n32489 , n20017 , n20020 );
xor ( n32490 , n32489 , n20041 );
buf ( n32491 , n32490 );
and ( n32492 , n32488 , n32491 );
and ( n32493 , n32483 , n32487 );
or ( n32494 , n32492 , n32493 );
buf ( n32495 , n32494 );
and ( n32496 , n32459 , n32495 );
and ( n32497 , n32455 , n32458 );
or ( n32498 , n32496 , n32497 );
xor ( n32499 , n32207 , n32498 );
xor ( n32500 , n19785 , n20014 );
xor ( n32501 , n32500 , n20088 );
buf ( n32502 , n32501 );
and ( n32503 , n32499 , n32502 );
and ( n32504 , n32207 , n32498 );
or ( n32505 , n32503 , n32504 );
not ( n32506 , n32505 );
not ( n32507 , n20095 );
nand ( n32508 , n32506 , n32507 );
xor ( n32509 , n19401 , n19780 );
and ( n32510 , n32509 , n20093 );
and ( n32511 , n19401 , n19780 );
or ( n32512 , n32510 , n32511 );
buf ( n32513 , n32512 );
not ( n32514 , n32513 );
not ( n32515 , n26378 );
nand ( n32516 , n32514 , n32515 );
nand ( n32517 , n32508 , n32516 );
xor ( n32518 , n26216 , n26369 );
and ( n32519 , n32518 , n26376 );
and ( n32520 , n26216 , n26369 );
or ( n32521 , n32519 , n32520 );
buf ( n32522 , n32521 );
not ( n32523 , n32522 );
xor ( n32524 , n26189 , n26195 );
and ( n32525 , n32524 , n26213 );
and ( n32526 , n26189 , n26195 );
or ( n32527 , n32525 , n32526 );
buf ( n32528 , n32527 );
buf ( n32529 , n32528 );
xor ( n32530 , n26227 , n26244 );
and ( n32531 , n32530 , n26262 );
and ( n32532 , n26227 , n26244 );
or ( n32533 , n32531 , n32532 );
buf ( n32534 , n32533 );
buf ( n32535 , n32534 );
xor ( n32536 , n26282 , n26299 );
and ( n32537 , n32536 , n26317 );
and ( n32538 , n26282 , n26299 );
or ( n32539 , n32537 , n32538 );
buf ( n32540 , n32539 );
buf ( n32541 , n32540 );
xor ( n32542 , n32535 , n32541 );
buf ( n32543 , n26275 );
not ( n32544 , n32543 );
buf ( n32545 , n18931 );
not ( n32546 , n32545 );
or ( n32547 , n32544 , n32546 );
buf ( n32548 , n18944 );
buf ( n32549 , n29509 );
nand ( n32550 , n32548 , n32549 );
buf ( n32551 , n32550 );
buf ( n32552 , n32551 );
nand ( n32553 , n32547 , n32552 );
buf ( n32554 , n32553 );
buf ( n32555 , n32554 );
buf ( n32556 , n26328 );
not ( n32557 , n32556 );
buf ( n32558 , n19230 );
not ( n32559 , n32558 );
or ( n32560 , n32557 , n32559 );
buf ( n32561 , n19235 );
buf ( n32562 , n29414 );
nand ( n32563 , n32561 , n32562 );
buf ( n32564 , n32563 );
buf ( n32565 , n32564 );
nand ( n32566 , n32560 , n32565 );
buf ( n32567 , n32566 );
buf ( n32568 , n32567 );
xor ( n32569 , n32555 , n32568 );
buf ( n32570 , n26310 );
not ( n32571 , n32570 );
buf ( n32572 , n18887 );
not ( n32573 , n32572 );
or ( n32574 , n32571 , n32573 );
buf ( n32575 , n18898 );
buf ( n32576 , n29393 );
nand ( n32577 , n32575 , n32576 );
buf ( n32578 , n32577 );
buf ( n32579 , n32578 );
nand ( n32580 , n32574 , n32579 );
buf ( n32581 , n32580 );
buf ( n32582 , n32581 );
xor ( n32583 , n32569 , n32582 );
buf ( n32584 , n32583 );
buf ( n32585 , n32584 );
xor ( n32586 , n32542 , n32585 );
buf ( n32587 , n32586 );
buf ( n32588 , n32587 );
xor ( n32589 , n26265 , n26320 );
and ( n32590 , n32589 , n26356 );
and ( n32591 , n26265 , n26320 );
or ( n32592 , n32590 , n32591 );
buf ( n32593 , n32592 );
buf ( n32594 , n32593 );
xor ( n32595 , n32588 , n32594 );
buf ( n32596 , n845 );
buf ( n32597 , n864 );
and ( n32598 , n32596 , n32597 );
buf ( n32599 , n32598 );
buf ( n32600 , n32599 );
buf ( n32601 , n26255 );
not ( n32602 , n32601 );
buf ( n32603 , n19125 );
not ( n32604 , n32603 );
or ( n32605 , n32602 , n32604 );
buf ( n32606 , n19134 );
buf ( n32607 , n29443 );
nand ( n32608 , n32606 , n32607 );
buf ( n32609 , n32608 );
buf ( n32610 , n32609 );
nand ( n32611 , n32605 , n32610 );
buf ( n32612 , n32611 );
buf ( n32613 , n32612 );
xor ( n32614 , n32600 , n32613 );
buf ( n32615 , n26292 );
not ( n32616 , n32615 );
buf ( n32617 , n18977 );
not ( n32618 , n32617 );
or ( n32619 , n32616 , n32618 );
buf ( n32620 , n18987 );
buf ( n32621 , n29464 );
nand ( n32622 , n32620 , n32621 );
buf ( n32623 , n32622 );
buf ( n32624 , n32623 );
nand ( n32625 , n32619 , n32624 );
buf ( n32626 , n32625 );
buf ( n32627 , n32626 );
xor ( n32628 , n32614 , n32627 );
buf ( n32629 , n32628 );
buf ( n32630 , n32629 );
buf ( n32631 , n29535 );
not ( n32632 , n32631 );
buf ( n32633 , n32632 );
buf ( n32634 , n32633 );
buf ( n32635 , n26237 );
not ( n32636 , n32635 );
buf ( n32637 , n19330 );
not ( n32638 , n32637 );
or ( n32639 , n32636 , n32638 );
buf ( n32640 , n19030 );
buf ( n32641 , n29492 );
nand ( n32642 , n32640 , n32641 );
buf ( n32643 , n32642 );
buf ( n32644 , n32643 );
nand ( n32645 , n32639 , n32644 );
buf ( n32646 , n32645 );
buf ( n32647 , n32646 );
xor ( n32648 , n32634 , n32647 );
buf ( n32649 , n26347 );
buf ( n32650 , n26334 );
or ( n32651 , n32649 , n32650 );
buf ( n32652 , n26354 );
nand ( n32653 , n32651 , n32652 );
buf ( n32654 , n32653 );
buf ( n32655 , n32654 );
buf ( n32656 , n26347 );
buf ( n32657 , n26334 );
nand ( n32658 , n32656 , n32657 );
buf ( n32659 , n32658 );
buf ( n32660 , n32659 );
nand ( n32661 , n32655 , n32660 );
buf ( n32662 , n32661 );
buf ( n32663 , n32662 );
xor ( n32664 , n32648 , n32663 );
buf ( n32665 , n32664 );
buf ( n32666 , n32665 );
xor ( n32667 , n32630 , n32666 );
xor ( n32668 , n26197 , n26203 );
and ( n32669 , n32668 , n26210 );
and ( n32670 , n26197 , n26203 );
or ( n32671 , n32669 , n32670 );
buf ( n32672 , n32671 );
buf ( n32673 , n32672 );
xor ( n32674 , n32667 , n32673 );
buf ( n32675 , n32674 );
buf ( n32676 , n32675 );
xor ( n32677 , n32595 , n32676 );
buf ( n32678 , n32677 );
buf ( n32679 , n32678 );
xor ( n32680 , n32529 , n32679 );
xor ( n32681 , n26222 , n26359 );
and ( n32682 , n32681 , n26366 );
and ( n32683 , n26222 , n26359 );
or ( n32684 , n32682 , n32683 );
buf ( n32685 , n32684 );
buf ( n32686 , n32685 );
xor ( n32687 , n32680 , n32686 );
buf ( n32688 , n32687 );
not ( n32689 , n32688 );
nand ( n32690 , n32523 , n32689 );
buf ( n32691 , n29405 );
buf ( n32692 , n29408 );
xor ( n32693 , n32691 , n32692 );
buf ( n32694 , n32693 );
buf ( n32695 , n32694 );
buf ( n32696 , n29426 );
xor ( n32697 , n32695 , n32696 );
buf ( n32698 , n32697 );
buf ( n32699 , n32698 );
xor ( n32700 , n29504 , n29521 );
buf ( n32701 , n32700 );
buf ( n32702 , n29535 );
and ( n32703 , n32701 , n32702 );
not ( n32704 , n32701 );
buf ( n32705 , n32633 );
and ( n32706 , n32704 , n32705 );
nor ( n32707 , n32703 , n32706 );
buf ( n32708 , n32707 );
buf ( n32709 , n32708 );
xor ( n32710 , n32699 , n32709 );
xor ( n32711 , n32634 , n32647 );
and ( n32712 , n32711 , n32663 );
and ( n32713 , n32634 , n32647 );
or ( n32714 , n32712 , n32713 );
buf ( n32715 , n32714 );
buf ( n32716 , n32715 );
xor ( n32717 , n32710 , n32716 );
buf ( n32718 , n32717 );
buf ( n32719 , n32718 );
xor ( n32720 , n32535 , n32541 );
and ( n32721 , n32720 , n32585 );
and ( n32722 , n32535 , n32541 );
or ( n32723 , n32721 , n32722 );
buf ( n32724 , n32723 );
buf ( n32725 , n32724 );
xor ( n32726 , n32600 , n32613 );
and ( n32727 , n32726 , n32627 );
and ( n32728 , n32600 , n32613 );
or ( n32729 , n32727 , n32728 );
buf ( n32730 , n32729 );
buf ( n32731 , n32730 );
xor ( n32732 , n32555 , n32568 );
and ( n32733 , n32732 , n32582 );
and ( n32734 , n32555 , n32568 );
or ( n32735 , n32733 , n32734 );
buf ( n32736 , n32735 );
buf ( n32737 , n32736 );
xor ( n32738 , n32731 , n32737 );
xor ( n32739 , n29456 , n29459 );
xor ( n32740 , n32739 , n29477 );
buf ( n32741 , n32740 );
buf ( n32742 , n32741 );
xor ( n32743 , n32738 , n32742 );
buf ( n32744 , n32743 );
buf ( n32745 , n32744 );
xor ( n32746 , n32725 , n32745 );
xor ( n32747 , n32630 , n32666 );
and ( n32748 , n32747 , n32673 );
and ( n32749 , n32630 , n32666 );
or ( n32750 , n32748 , n32749 );
buf ( n32751 , n32750 );
buf ( n32752 , n32751 );
xor ( n32753 , n32746 , n32752 );
buf ( n32754 , n32753 );
buf ( n32755 , n32754 );
xor ( n32756 , n32719 , n32755 );
xor ( n32757 , n32588 , n32594 );
and ( n32758 , n32757 , n32676 );
and ( n32759 , n32588 , n32594 );
or ( n32760 , n32758 , n32759 );
buf ( n32761 , n32760 );
buf ( n32762 , n32761 );
xor ( n32763 , n32756 , n32762 );
buf ( n32764 , n32763 );
not ( n32765 , n32764 );
xor ( n32766 , n32529 , n32679 );
and ( n32767 , n32766 , n32686 );
and ( n32768 , n32529 , n32679 );
or ( n32769 , n32767 , n32768 );
buf ( n32770 , n32769 );
not ( n32771 , n32770 );
nand ( n32772 , n32765 , n32771 );
nand ( n32773 , n32690 , n32772 );
nor ( n32774 , n32517 , n32773 );
not ( n32775 , n32774 );
xor ( n32776 , n32699 , n32709 );
and ( n32777 , n32776 , n32716 );
and ( n32778 , n32699 , n32709 );
or ( n32779 , n32777 , n32778 );
buf ( n32780 , n32779 );
buf ( n32781 , n32780 );
xor ( n32782 , n29389 , n29438 );
xor ( n32783 , n32782 , n29482 );
buf ( n32784 , n32783 );
buf ( n32785 , n32784 );
xor ( n32786 , n32731 , n32737 );
and ( n32787 , n32786 , n32742 );
and ( n32788 , n32731 , n32737 );
or ( n32789 , n32787 , n32788 );
buf ( n32790 , n32789 );
buf ( n32791 , n32790 );
xor ( n32792 , n32785 , n32791 );
xor ( n32793 , n29547 , n29551 );
xor ( n32794 , n32793 , n29558 );
buf ( n32795 , n32794 );
buf ( n32796 , n32795 );
xor ( n32797 , n32792 , n32796 );
buf ( n32798 , n32797 );
buf ( n32799 , n32798 );
xor ( n32800 , n32781 , n32799 );
xor ( n32801 , n32725 , n32745 );
and ( n32802 , n32801 , n32752 );
and ( n32803 , n32725 , n32745 );
or ( n32804 , n32802 , n32803 );
buf ( n32805 , n32804 );
buf ( n32806 , n32805 );
and ( n32807 , n32800 , n32806 );
and ( n32808 , n32781 , n32799 );
or ( n32809 , n32807 , n32808 );
buf ( n32810 , n32809 );
xor ( n32811 , n29363 , n29367 );
xor ( n32812 , n32811 , n29372 );
buf ( n32813 , n32812 );
buf ( n32814 , n32813 );
xor ( n32815 , n29385 , n29487 );
xor ( n32816 , n32815 , n29563 );
buf ( n32817 , n32816 );
buf ( n32818 , n32817 );
xor ( n32819 , n32814 , n32818 );
xor ( n32820 , n32785 , n32791 );
and ( n32821 , n32820 , n32796 );
and ( n32822 , n32785 , n32791 );
or ( n32823 , n32821 , n32822 );
buf ( n32824 , n32823 );
buf ( n32825 , n32824 );
xor ( n32826 , n32819 , n32825 );
buf ( n32827 , n32826 );
or ( n32828 , n32810 , n32827 );
xor ( n32829 , n32781 , n32799 );
xor ( n32830 , n32829 , n32806 );
buf ( n32831 , n32830 );
xor ( n32832 , n32719 , n32755 );
and ( n32833 , n32832 , n32762 );
and ( n32834 , n32719 , n32755 );
or ( n32835 , n32833 , n32834 );
buf ( n32836 , n32835 );
or ( n32837 , n32831 , n32836 );
nand ( n32838 , n32828 , n32837 );
nor ( n32839 , n32775 , n32838 );
not ( n32840 , n32839 );
xor ( n32841 , n32304 , n32321 );
xor ( n32842 , n32841 , n32339 );
buf ( n32843 , n32842 );
buf ( n32844 , n32843 );
not ( n32845 , n32844 );
buf ( n32846 , n32845 );
buf ( n32847 , n32846 );
not ( n32848 , n32847 );
xor ( n32849 , n32242 , n32282 );
xnor ( n32850 , n32849 , n32260 );
buf ( n32851 , n32850 );
not ( n32852 , n32851 );
or ( n32853 , n32848 , n32852 );
buf ( n32854 , n24869 );
not ( n32855 , n32854 );
buf ( n32856 , n18931 );
not ( n32857 , n32856 );
or ( n32858 , n32855 , n32857 );
buf ( n32859 , n18944 );
buf ( n32860 , n32270 );
nand ( n32861 , n32859 , n32860 );
buf ( n32862 , n32861 );
buf ( n32863 , n32862 );
nand ( n32864 , n32858 , n32863 );
buf ( n32865 , n32864 );
buf ( n32866 , n32865 );
buf ( n32867 , n25054 );
not ( n32868 , n32867 );
buf ( n32869 , n19013 );
not ( n32870 , n32869 );
or ( n32871 , n32868 , n32870 );
buf ( n32872 , n19030 );
buf ( n32873 , n32230 );
nand ( n32874 , n32872 , n32873 );
buf ( n32875 , n32874 );
buf ( n32876 , n32875 );
nand ( n32877 , n32871 , n32876 );
buf ( n32878 , n32877 );
buf ( n32879 , n32878 );
xor ( n32880 , n32866 , n32879 );
buf ( n32881 , n25076 );
not ( n32882 , n32881 );
buf ( n32883 , n19153 );
not ( n32884 , n32883 );
or ( n32885 , n32882 , n32884 );
buf ( n32886 , n20246 );
buf ( n32887 , n32886 );
buf ( n32888 , n32365 );
nand ( n32889 , n32887 , n32888 );
buf ( n32890 , n32889 );
buf ( n32891 , n32890 );
nand ( n32892 , n32885 , n32891 );
buf ( n32893 , n32892 );
buf ( n32894 , n32893 );
and ( n32895 , n32880 , n32894 );
and ( n32896 , n32866 , n32879 );
or ( n32897 , n32895 , n32896 );
buf ( n32898 , n32897 );
buf ( n32899 , n32898 );
nand ( n32900 , n32853 , n32899 );
buf ( n32901 , n32900 );
buf ( n32902 , n32901 );
not ( n32903 , n32850 );
nand ( n32904 , n32903 , n32843 );
buf ( n32905 , n32904 );
nand ( n32906 , n32902 , n32905 );
buf ( n32907 , n32906 );
buf ( n32908 , n32907 );
buf ( n32909 , n24956 );
not ( n32910 , n32909 );
buf ( n32911 , n25285 );
not ( n32912 , n32911 );
or ( n32913 , n32910 , n32912 );
buf ( n32914 , n19234 );
buf ( n32915 , n32308 );
nand ( n32916 , n32914 , n32915 );
buf ( n32917 , n32916 );
buf ( n32918 , n32917 );
nand ( n32919 , n32913 , n32918 );
buf ( n32920 , n32919 );
buf ( n32921 , n32920 );
buf ( n32922 , n25097 );
not ( n32923 , n32922 );
buf ( n32924 , n18977 );
not ( n32925 , n32924 );
or ( n32926 , n32923 , n32925 );
buf ( n32927 , n18987 );
buf ( n32928 , n32326 );
nand ( n32929 , n32927 , n32928 );
buf ( n32930 , n32929 );
buf ( n32931 , n32930 );
nand ( n32932 , n32926 , n32931 );
buf ( n32933 , n32932 );
buf ( n32934 , n32933 );
xor ( n32935 , n32921 , n32934 );
buf ( n32936 , n24910 );
not ( n32937 , n32936 );
buf ( n32938 , n19580 );
not ( n32939 , n32938 );
or ( n32940 , n32937 , n32939 );
buf ( n32941 , n26538 );
buf ( n32942 , n32410 );
nand ( n32943 , n32941 , n32942 );
buf ( n32944 , n32943 );
buf ( n32945 , n32944 );
nand ( n32946 , n32940 , n32945 );
buf ( n32947 , n32946 );
buf ( n32948 , n32947 );
not ( n32949 , n32948 );
buf ( n32950 , n32949 );
buf ( n32951 , n32950 );
and ( n32952 , n32935 , n32951 );
and ( n32953 , n32921 , n32934 );
or ( n32954 , n32952 , n32953 );
buf ( n32955 , n32954 );
buf ( n32956 , n32955 );
xor ( n32957 , n32361 , n32378 );
xor ( n32958 , n32957 , n32396 );
buf ( n32959 , n32958 );
buf ( n32960 , n32959 );
xor ( n32961 , n32956 , n32960 );
xor ( n32962 , n32409 , n32423 );
xor ( n32963 , n32962 , n32441 );
buf ( n32964 , n32963 );
buf ( n32965 , n32964 );
and ( n32966 , n32961 , n32965 );
and ( n32967 , n32956 , n32960 );
or ( n32968 , n32966 , n32967 );
buf ( n32969 , n32968 );
buf ( n32970 , n32969 );
xor ( n32971 , n32908 , n32970 );
xor ( n32972 , n32466 , n32462 );
buf ( n32973 , n32972 );
buf ( n32974 , n32471 );
xor ( n32975 , n32973 , n32974 );
buf ( n32976 , n32975 );
buf ( n32977 , n32976 );
xor ( n32978 , n32971 , n32977 );
buf ( n32979 , n32978 );
buf ( n32980 , n32979 );
xor ( n32981 , n25104 , n25121 );
and ( n32982 , n32981 , n25183 );
and ( n32983 , n25104 , n25121 );
or ( n32984 , n32982 , n32983 );
buf ( n32985 , n32984 );
buf ( n32986 , n32985 );
not ( n32987 , n24875 );
not ( n32988 , n24916 );
or ( n32989 , n32987 , n32988 );
buf ( n32990 , n24916 );
buf ( n32991 , n24875 );
nor ( n32992 , n32990 , n32991 );
buf ( n32993 , n32992 );
buf ( n32994 , n24895 );
not ( n32995 , n32994 );
buf ( n32996 , n32995 );
or ( n32997 , n32993 , n32996 );
nand ( n32998 , n32989 , n32997 );
buf ( n32999 , n32998 );
buf ( n33000 , n25013 );
not ( n33001 , n33000 );
buf ( n33002 , n24997 );
not ( n33003 , n33002 );
or ( n33004 , n33001 , n33003 );
not ( n33005 , n24997 );
not ( n33006 , n33005 );
not ( n33007 , n25013 );
not ( n33008 , n33007 );
or ( n33009 , n33006 , n33008 );
nand ( n33010 , n33009 , n25033 );
buf ( n33011 , n33010 );
nand ( n33012 , n33004 , n33011 );
buf ( n33013 , n33012 );
buf ( n33014 , n33013 );
xor ( n33015 , n32999 , n33014 );
xor ( n33016 , n25040 , n25061 );
and ( n33017 , n33016 , n25083 );
and ( n33018 , n25040 , n25061 );
or ( n33019 , n33017 , n33018 );
buf ( n33020 , n33019 );
buf ( n33021 , n33020 );
xor ( n33022 , n33015 , n33021 );
buf ( n33023 , n33022 );
buf ( n33024 , n33023 );
xor ( n33025 , n32986 , n33024 );
not ( n33026 , n24921 );
nand ( n33027 , n33026 , n25034 );
nand ( n33028 , n33026 , n24987 );
nand ( n33029 , n25034 , n24987 );
nand ( n33030 , n33027 , n33028 , n33029 );
buf ( n33031 , n33030 );
and ( n33032 , n33025 , n33031 );
and ( n33033 , n32986 , n33024 );
or ( n33034 , n33032 , n33033 );
buf ( n33035 , n33034 );
buf ( n33036 , n33035 );
xor ( n33037 , n32999 , n33014 );
and ( n33038 , n33037 , n33021 );
and ( n33039 , n32999 , n33014 );
or ( n33040 , n33038 , n33039 );
buf ( n33041 , n33040 );
buf ( n33042 , n33041 );
buf ( n33043 , n32947 );
buf ( n33044 , n853 );
buf ( n33045 , n864 );
and ( n33046 , n33044 , n33045 );
buf ( n33047 , n33046 );
buf ( n33048 , n33047 );
buf ( n33049 , n25009 );
not ( n33050 , n33049 );
buf ( n33051 , n19614 );
not ( n33052 , n33051 );
or ( n33053 , n33050 , n33052 );
buf ( n33054 , n18860 );
buf ( n33055 , n32248 );
nand ( n33056 , n33054 , n33055 );
buf ( n33057 , n33056 );
buf ( n33058 , n33057 );
nand ( n33059 , n33053 , n33058 );
buf ( n33060 , n33059 );
buf ( n33061 , n33060 );
xor ( n33062 , n33048 , n33061 );
buf ( n33063 , n25029 );
not ( n33064 , n33063 );
buf ( n33065 , n25022 );
not ( n33066 , n33065 );
or ( n33067 , n33064 , n33066 );
buf ( n33068 , n25263 );
buf ( n33069 , n884 );
nand ( n33070 , n33068 , n33069 );
buf ( n33071 , n33070 );
buf ( n33072 , n33071 );
nand ( n33073 , n33067 , n33072 );
buf ( n33074 , n33073 );
buf ( n33075 , n33074 );
and ( n33076 , n33062 , n33075 );
and ( n33077 , n33048 , n33061 );
or ( n33078 , n33076 , n33077 );
buf ( n33079 , n33078 );
buf ( n33080 , n33079 );
xor ( n33081 , n33043 , n33080 );
buf ( n33082 , n24935 );
not ( n33083 , n33082 );
buf ( n33084 , n19122 );
not ( n33085 , n33084 );
or ( n33086 , n33083 , n33085 );
buf ( n33087 , n19131 );
buf ( n33088 , n32383 );
nand ( n33089 , n33087 , n33088 );
buf ( n33090 , n33089 );
buf ( n33091 , n33090 );
nand ( n33092 , n33086 , n33091 );
buf ( n33093 , n33092 );
buf ( n33094 , n33093 );
buf ( n33095 , n24978 );
not ( n33096 , n33095 );
buf ( n33097 , n19479 );
not ( n33098 , n33097 );
or ( n33099 , n33096 , n33098 );
buf ( n33100 , n19265 );
buf ( n33101 , n32428 );
nand ( n33102 , n33100 , n33101 );
buf ( n33103 , n33102 );
buf ( n33104 , n33103 );
nand ( n33105 , n33099 , n33104 );
buf ( n33106 , n33105 );
buf ( n33107 , n33106 );
xor ( n33108 , n33094 , n33107 );
buf ( n33109 , n24889 );
not ( n33110 , n33109 );
buf ( n33111 , n18887 );
not ( n33112 , n33111 );
or ( n33113 , n33110 , n33112 );
buf ( n33114 , n19461 );
buf ( n33115 , n32348 );
nand ( n33116 , n33114 , n33115 );
buf ( n33117 , n33116 );
buf ( n33118 , n33117 );
nand ( n33119 , n33113 , n33118 );
buf ( n33120 , n33119 );
buf ( n33121 , n33120 );
and ( n33122 , n33108 , n33121 );
and ( n33123 , n33094 , n33107 );
or ( n33124 , n33122 , n33123 );
buf ( n33125 , n33124 );
buf ( n33126 , n33125 );
xor ( n33127 , n33081 , n33126 );
buf ( n33128 , n33127 );
buf ( n33129 , n33128 );
xor ( n33130 , n33042 , n33129 );
xor ( n33131 , n33048 , n33061 );
xor ( n33132 , n33131 , n33075 );
buf ( n33133 , n33132 );
buf ( n33134 , n33133 );
xor ( n33135 , n24942 , n24963 );
and ( n33136 , n33135 , n24985 );
and ( n33137 , n24942 , n24963 );
or ( n33138 , n33136 , n33137 );
buf ( n33139 , n33138 );
buf ( n33140 , n33139 );
xor ( n33141 , n33134 , n33140 );
xor ( n33142 , n33094 , n33107 );
xor ( n33143 , n33142 , n33121 );
buf ( n33144 , n33143 );
buf ( n33145 , n33144 );
and ( n33146 , n33141 , n33145 );
and ( n33147 , n33134 , n33140 );
or ( n33148 , n33146 , n33147 );
buf ( n33149 , n33148 );
buf ( n33150 , n33149 );
xor ( n33151 , n33130 , n33150 );
buf ( n33152 , n33151 );
buf ( n33153 , n33152 );
xor ( n33154 , n33036 , n33153 );
xor ( n33155 , n33134 , n33140 );
xor ( n33156 , n33155 , n33145 );
buf ( n33157 , n33156 );
buf ( n33158 , n33157 );
xor ( n33159 , n32866 , n32879 );
xor ( n33160 , n33159 , n32894 );
buf ( n33161 , n33160 );
buf ( n33162 , n33161 );
xor ( n33163 , n32921 , n32934 );
xor ( n33164 , n33163 , n32951 );
buf ( n33165 , n33164 );
buf ( n33166 , n33165 );
xor ( n33167 , n33162 , n33166 );
xor ( n33168 , n26084 , n26090 );
and ( n33169 , n33168 , n26132 );
and ( n33170 , n26084 , n26090 );
or ( n33171 , n33169 , n33170 );
buf ( n33172 , n33171 );
buf ( n33173 , n33172 );
xor ( n33174 , n33167 , n33173 );
buf ( n33175 , n33174 );
buf ( n33176 , n33175 );
xor ( n33177 , n33158 , n33176 );
xor ( n33178 , n25086 , n25186 );
and ( n33179 , n33178 , n25350 );
and ( n33180 , n25086 , n25186 );
or ( n33181 , n33179 , n33180 );
buf ( n33182 , n33181 );
buf ( n33183 , n33182 );
and ( n33184 , n33177 , n33183 );
and ( n33185 , n33158 , n33176 );
or ( n33186 , n33184 , n33185 );
buf ( n33187 , n33186 );
buf ( n33188 , n33187 );
and ( n33189 , n33154 , n33188 );
and ( n33190 , n33036 , n33153 );
or ( n33191 , n33189 , n33190 );
buf ( n33192 , n33191 );
buf ( n33193 , n33192 );
xor ( n33194 , n32980 , n33193 );
xor ( n33195 , n33042 , n33129 );
and ( n33196 , n33195 , n33150 );
and ( n33197 , n33042 , n33129 );
or ( n33198 , n33196 , n33197 );
buf ( n33199 , n33198 );
buf ( n33200 , n33199 );
xor ( n33201 , n32208 , n32225 );
xor ( n33202 , n33201 , n32289 );
buf ( n33203 , n33202 );
buf ( n33204 , n33203 );
xor ( n33205 , n33043 , n33080 );
and ( n33206 , n33205 , n33126 );
and ( n33207 , n33043 , n33080 );
or ( n33208 , n33206 , n33207 );
buf ( n33209 , n33208 );
buf ( n33210 , n33209 );
xor ( n33211 , n33204 , n33210 );
xor ( n33212 , n32344 , n32401 );
xor ( n33213 , n33212 , n32446 );
buf ( n33214 , n33213 );
buf ( n33215 , n33214 );
xor ( n33216 , n33211 , n33215 );
buf ( n33217 , n33216 );
buf ( n33218 , n33217 );
xor ( n33219 , n33200 , n33218 );
xor ( n33220 , n32956 , n32960 );
xor ( n33221 , n33220 , n32965 );
buf ( n33222 , n33221 );
buf ( n33223 , n33222 );
not ( n33224 , n33223 );
buf ( n33225 , n33224 );
buf ( n33226 , n33225 );
not ( n33227 , n33226 );
xor ( n33228 , n32843 , n32898 );
xor ( n33229 , n33228 , n32850 );
buf ( n33230 , n33229 );
not ( n33231 , n33230 );
or ( n33232 , n33227 , n33231 );
xor ( n33233 , n33162 , n33166 );
and ( n33234 , n33233 , n33173 );
and ( n33235 , n33162 , n33166 );
or ( n33236 , n33234 , n33235 );
buf ( n33237 , n33236 );
buf ( n33238 , n33237 );
nand ( n33239 , n33232 , n33238 );
buf ( n33240 , n33239 );
buf ( n33241 , n33240 );
buf ( n33242 , n33222 );
buf ( n33243 , n33229 );
not ( n33244 , n33243 );
buf ( n33245 , n33244 );
buf ( n33246 , n33245 );
nand ( n33247 , n33242 , n33246 );
buf ( n33248 , n33247 );
buf ( n33249 , n33248 );
nand ( n33250 , n33241 , n33249 );
buf ( n33251 , n33250 );
buf ( n33252 , n33251 );
xor ( n33253 , n33219 , n33252 );
buf ( n33254 , n33253 );
buf ( n33255 , n33254 );
xor ( n33256 , n33194 , n33255 );
buf ( n33257 , n33256 );
not ( n33258 , n33257 );
buf ( n33259 , n33245 );
not ( n33260 , n33259 );
buf ( n33261 , n33225 );
not ( n33262 , n33261 );
or ( n33263 , n33260 , n33262 );
buf ( n33264 , n33222 );
buf ( n33265 , n33229 );
nand ( n33266 , n33264 , n33265 );
buf ( n33267 , n33266 );
buf ( n33268 , n33267 );
nand ( n33269 , n33263 , n33268 );
buf ( n33270 , n33269 );
buf ( n33271 , n33270 );
buf ( n33272 , n33237 );
and ( n33273 , n33271 , n33272 );
not ( n33274 , n33271 );
buf ( n33275 , n33237 );
not ( n33276 , n33275 );
buf ( n33277 , n33276 );
buf ( n33278 , n33277 );
and ( n33279 , n33274 , n33278 );
nor ( n33280 , n33273 , n33279 );
buf ( n33281 , n33280 );
buf ( n33282 , n33281 );
xor ( n33283 , n32986 , n33024 );
xor ( n33284 , n33283 , n33031 );
buf ( n33285 , n33284 );
buf ( n33286 , n33285 );
xor ( n33287 , n26032 , n26135 );
and ( n33288 , n33287 , n26157 );
and ( n33289 , n26032 , n26135 );
or ( n33290 , n33288 , n33289 );
buf ( n33291 , n33290 );
buf ( n33292 , n33291 );
xor ( n33293 , n33286 , n33292 );
nand ( n33294 , n25035 , n25352 );
nand ( n33295 , n25035 , n25585 );
nand ( n33296 , n25352 , n25585 );
nand ( n33297 , n33294 , n33295 , n33296 );
buf ( n33298 , n33297 );
and ( n33299 , n33293 , n33298 );
and ( n33300 , n33286 , n33292 );
or ( n33301 , n33299 , n33300 );
buf ( n33302 , n33301 );
buf ( n33303 , n33302 );
xor ( n33304 , n33282 , n33303 );
xor ( n33305 , n33036 , n33153 );
xor ( n33306 , n33305 , n33188 );
buf ( n33307 , n33306 );
buf ( n33308 , n33307 );
and ( n33309 , n33304 , n33308 );
and ( n33310 , n33282 , n33303 );
or ( n33311 , n33309 , n33310 );
buf ( n33312 , n33311 );
not ( n33313 , n33312 );
nand ( n33314 , n33258 , n33313 );
xor ( n33315 , n32908 , n32970 );
and ( n33316 , n33315 , n32977 );
and ( n33317 , n32908 , n32970 );
or ( n33318 , n33316 , n33317 );
buf ( n33319 , n33318 );
buf ( n33320 , n33319 );
xor ( n33321 , n33200 , n33218 );
and ( n33322 , n33321 , n33252 );
and ( n33323 , n33200 , n33218 );
or ( n33324 , n33322 , n33323 );
buf ( n33325 , n33324 );
buf ( n33326 , n33325 );
xor ( n33327 , n33320 , n33326 );
xor ( n33328 , n32294 , n32298 );
xor ( n33329 , n33328 , n32451 );
buf ( n33330 , n33329 );
buf ( n33331 , n33330 );
xor ( n33332 , n33204 , n33210 );
and ( n33333 , n33332 , n33215 );
and ( n33334 , n33204 , n33210 );
or ( n33335 , n33333 , n33334 );
buf ( n33336 , n33335 );
buf ( n33337 , n33336 );
xor ( n33338 , n33331 , n33337 );
xor ( n33339 , n32483 , n32487 );
xor ( n33340 , n33339 , n32491 );
buf ( n33341 , n33340 );
buf ( n33342 , n33341 );
xor ( n33343 , n33338 , n33342 );
buf ( n33344 , n33343 );
buf ( n33345 , n33344 );
xor ( n33346 , n33327 , n33345 );
buf ( n33347 , n33346 );
not ( n33348 , n33347 );
xor ( n33349 , n32980 , n33193 );
and ( n33350 , n33349 , n33255 );
and ( n33351 , n32980 , n33193 );
or ( n33352 , n33350 , n33351 );
buf ( n33353 , n33352 );
not ( n33354 , n33353 );
nand ( n33355 , n33348 , n33354 );
nand ( n33356 , n33314 , n33355 );
xor ( n33357 , n33320 , n33326 );
and ( n33358 , n33357 , n33345 );
and ( n33359 , n33320 , n33326 );
or ( n33360 , n33358 , n33359 );
buf ( n33361 , n33360 );
not ( n33362 , n33361 );
buf ( n33363 , n20073 );
not ( n33364 , n33363 );
buf ( n33365 , n20044 );
not ( n33366 , n33365 );
or ( n33367 , n33364 , n33366 );
buf ( n33368 , n20044 );
buf ( n33369 , n20073 );
or ( n33370 , n33368 , n33369 );
nand ( n33371 , n33367 , n33370 );
buf ( n33372 , n33371 );
xor ( n33373 , n20053 , n33372 );
xor ( n33374 , n32455 , n32458 );
xor ( n33375 , n33374 , n32495 );
xor ( n33376 , n33373 , n33375 );
xor ( n33377 , n33331 , n33337 );
and ( n33378 , n33377 , n33342 );
and ( n33379 , n33331 , n33337 );
or ( n33380 , n33378 , n33379 );
buf ( n33381 , n33380 );
xor ( n33382 , n33376 , n33381 );
not ( n33383 , n33382 );
nand ( n33384 , n33362 , n33383 );
xor ( n33385 , n32207 , n32498 );
xor ( n33386 , n33385 , n32502 );
not ( n33387 , n33386 );
xor ( n33388 , n33373 , n33375 );
and ( n33389 , n33388 , n33381 );
and ( n33390 , n33373 , n33375 );
or ( n33391 , n33389 , n33390 );
not ( n33392 , n33391 );
nand ( n33393 , n33387 , n33392 );
nand ( n33394 , n33384 , n33393 );
nor ( n33395 , n33356 , n33394 );
not ( n33396 , n33395 );
xor ( n33397 , n33282 , n33303 );
xor ( n33398 , n33397 , n33308 );
buf ( n33399 , n33398 );
not ( n33400 , n33399 );
xor ( n33401 , n33158 , n33176 );
xor ( n33402 , n33401 , n33183 );
buf ( n33403 , n33402 );
buf ( n33404 , n33403 );
xor ( n33405 , n26026 , n26160 );
and ( n33406 , n33405 , n26177 );
and ( n33407 , n26026 , n26160 );
or ( n33408 , n33406 , n33407 );
buf ( n33409 , n33408 );
buf ( n33410 , n33409 );
xor ( n33411 , n33404 , n33410 );
xor ( n33412 , n33286 , n33292 );
xor ( n33413 , n33412 , n33298 );
buf ( n33414 , n33413 );
buf ( n33415 , n33414 );
and ( n33416 , n33411 , n33415 );
and ( n33417 , n33404 , n33410 );
or ( n33418 , n33416 , n33417 );
buf ( n33419 , n33418 );
not ( n33420 , n33419 );
nand ( n33421 , n33400 , n33420 );
not ( n33422 , n26384 );
xor ( n33423 , n33404 , n33410 );
xor ( n33424 , n33423 , n33415 );
buf ( n33425 , n33424 );
not ( n33426 , n33425 );
nand ( n33427 , n33422 , n33426 );
nand ( n33428 , n33421 , n33427 );
not ( n33429 , n33428 );
not ( n33430 , n33429 );
xor ( n33431 , n26164 , n26167 );
xor ( n33432 , n33431 , n26173 );
buf ( n33433 , n33432 );
xor ( n33434 , n25837 , n25876 );
xor ( n33435 , n33434 , n26014 );
buf ( n33436 , n33435 );
buf ( n33437 , n33436 );
xor ( n33438 , n33433 , n33437 );
xor ( n33439 , n23836 , n23870 );
and ( n33440 , n33439 , n23931 );
and ( n33441 , n23836 , n23870 );
or ( n33442 , n33440 , n33441 );
buf ( n33443 , n33442 );
xor ( n33444 , n25847 , n25851 );
xor ( n33445 , n33444 , n25861 );
buf ( n33446 , n33445 );
buf ( n33447 , n33446 );
xor ( n33448 , n33443 , n33447 );
xor ( n33449 , n23940 , n23991 );
and ( n33450 , n33449 , n23998 );
and ( n33451 , n23940 , n23991 );
or ( n33452 , n33450 , n33451 );
buf ( n33453 , n33452 );
buf ( n33454 , n33453 );
and ( n33455 , n33448 , n33454 );
and ( n33456 , n33443 , n33447 );
or ( n33457 , n33455 , n33456 );
buf ( n33458 , n33457 );
buf ( n33459 , n33458 );
xor ( n33460 , n25841 , n25866 );
xor ( n33461 , n33460 , n25871 );
buf ( n33462 , n33461 );
buf ( n33463 , n33462 );
xor ( n33464 , n33459 , n33463 );
xor ( n33465 , n25938 , n25988 );
xor ( n33466 , n33465 , n26009 );
buf ( n33467 , n33466 );
buf ( n33468 , n33467 );
and ( n33469 , n33464 , n33468 );
and ( n33470 , n33459 , n33463 );
or ( n33471 , n33469 , n33470 );
buf ( n33472 , n33471 );
buf ( n33473 , n33472 );
xor ( n33474 , n33438 , n33473 );
buf ( n33475 , n33474 );
not ( n33476 , n33475 );
xor ( n33477 , n25893 , n25896 );
xor ( n33478 , n33477 , n25933 );
buf ( n33479 , n33478 );
buf ( n33480 , n33479 );
xor ( n33481 , n23482 , n23544 );
and ( n33482 , n33481 , n23682 );
and ( n33483 , n23482 , n23544 );
or ( n33484 , n33482 , n33483 );
buf ( n33485 , n33484 );
xor ( n33486 , n33480 , n33485 );
xor ( n33487 , n25944 , n25953 );
xor ( n33488 , n33487 , n25983 );
buf ( n33489 , n33488 );
buf ( n33490 , n33489 );
and ( n33491 , n33486 , n33490 );
and ( n33492 , n33480 , n33485 );
or ( n33493 , n33491 , n33492 );
buf ( n33494 , n33493 );
buf ( n33495 , n33494 );
xor ( n33496 , n23794 , n23933 );
and ( n33497 , n33496 , n24001 );
and ( n33498 , n23794 , n23933 );
or ( n33499 , n33497 , n33498 );
buf ( n33500 , n33499 );
buf ( n33501 , n33500 );
xor ( n33502 , n33443 , n33447 );
xor ( n33503 , n33502 , n33454 );
buf ( n33504 , n33503 );
buf ( n33505 , n33504 );
xor ( n33506 , n33501 , n33505 );
xor ( n33507 , n33480 , n33485 );
xor ( n33508 , n33507 , n33490 );
buf ( n33509 , n33508 );
buf ( n33510 , n33509 );
and ( n33511 , n33506 , n33510 );
and ( n33512 , n33501 , n33505 );
or ( n33513 , n33511 , n33512 );
buf ( n33514 , n33513 );
buf ( n33515 , n33514 );
xor ( n33516 , n33495 , n33515 );
xor ( n33517 , n33459 , n33463 );
xor ( n33518 , n33517 , n33468 );
buf ( n33519 , n33518 );
buf ( n33520 , n33519 );
and ( n33521 , n33516 , n33520 );
and ( n33522 , n33495 , n33515 );
or ( n33523 , n33521 , n33522 );
buf ( n33524 , n33523 );
not ( n33525 , n33524 );
nor ( n33526 , n33476 , n33525 );
not ( n33527 , n33526 );
not ( n33528 , n26182 );
xor ( n33529 , n33433 , n33437 );
and ( n33530 , n33529 , n33473 );
and ( n33531 , n33433 , n33437 );
or ( n33532 , n33530 , n33531 );
buf ( n33533 , n33532 );
not ( n33534 , n33533 );
nand ( n33535 , n33528 , n33534 );
not ( n33536 , n33535 );
or ( n33537 , n33527 , n33536 );
not ( n33538 , n33534 );
not ( n33539 , n33528 );
nand ( n33540 , n33538 , n33539 );
nand ( n33541 , n33537 , n33540 );
not ( n33542 , n33541 );
or ( n33543 , n33430 , n33542 );
nor ( n33544 , n33399 , n33419 );
not ( n33545 , n33544 );
nand ( n33546 , n26384 , n33425 );
not ( n33547 , n33546 );
and ( n33548 , n33545 , n33547 );
nand ( n33549 , n33399 , n33419 );
not ( n33550 , n33549 );
nor ( n33551 , n33548 , n33550 );
nand ( n33552 , n33543 , n33551 );
not ( n33553 , n33552 );
or ( n33554 , n33396 , n33553 );
not ( n33555 , n33394 );
not ( n33556 , n33355 );
not ( n33557 , n33313 );
buf ( n33558 , n33257 );
nand ( n33559 , n33557 , n33558 );
or ( n33560 , n33556 , n33559 );
not ( n33561 , n33354 );
nand ( n33562 , n33561 , n33347 );
nand ( n33563 , n33560 , n33562 );
and ( n33564 , n33555 , n33563 );
not ( n33565 , n33393 );
nand ( n33566 , n33361 , n33382 );
or ( n33567 , n33565 , n33566 );
or ( n33568 , n33387 , n33392 );
nand ( n33569 , n33567 , n33568 );
nor ( n33570 , n33564 , n33569 );
nand ( n33571 , n33554 , n33570 );
not ( n33572 , n33571 );
xor ( n33573 , n24008 , n24017 );
xor ( n33574 , n33573 , n24022 );
buf ( n33575 , n33574 );
buf ( n33576 , n33575 );
xor ( n33577 , n22129 , n22468 );
and ( n33578 , n33577 , n22511 );
and ( n33579 , n22129 , n22468 );
or ( n33580 , n33578 , n33579 );
buf ( n33581 , n33580 );
buf ( n33582 , n33581 );
xor ( n33583 , n33576 , n33582 );
not ( n33584 , n24039 );
not ( n33585 , n24044 );
or ( n33586 , n33584 , n33585 );
nand ( n33587 , n24042 , n24033 );
nand ( n33588 , n33586 , n33587 );
and ( n33589 , n33588 , n24068 );
not ( n33590 , n33588 );
not ( n33591 , n24068 );
and ( n33592 , n33590 , n33591 );
nor ( n33593 , n33589 , n33592 );
buf ( n33594 , n33593 );
and ( n33595 , n33583 , n33594 );
and ( n33596 , n33576 , n33582 );
or ( n33597 , n33595 , n33596 );
buf ( n33598 , n33597 );
not ( n33599 , n33598 );
not ( n33600 , n33599 );
not ( n33601 , n33600 );
xor ( n33602 , n23742 , n24070 );
xor ( n33603 , n33602 , n24027 );
buf ( n33604 , n33603 );
not ( n33605 , n33604 );
or ( n33606 , n33601 , n33605 );
not ( n33607 , n33603 );
not ( n33608 , n33607 );
not ( n33609 , n33599 );
or ( n33610 , n33608 , n33609 );
xor ( n33611 , n33576 , n33582 );
xor ( n33612 , n33611 , n33594 );
buf ( n33613 , n33612 );
and ( n33614 , n33613 , n22525 );
nand ( n33615 , n33610 , n33614 );
nand ( n33616 , n33606 , n33615 );
buf ( n33617 , n22101 );
buf ( n33618 , n33617 );
not ( n33619 , n33618 );
not ( n33620 , n22096 );
not ( n33621 , n21915 );
or ( n33622 , n33620 , n33621 );
or ( n33623 , n22096 , n21915 );
nand ( n33624 , n33622 , n33623 );
buf ( n33625 , n33624 );
not ( n33626 , n33625 );
or ( n33627 , n33619 , n33626 );
buf ( n33628 , n33617 );
buf ( n33629 , n33624 );
or ( n33630 , n33628 , n33629 );
nand ( n33631 , n33627 , n33630 );
buf ( n33632 , n33631 );
buf ( n33633 , n33632 );
xor ( n33634 , n24840 , n24844 );
and ( n33635 , n33634 , n24849 );
and ( n33636 , n24840 , n24844 );
or ( n33637 , n33635 , n33636 );
buf ( n33638 , n33637 );
buf ( n33639 , n33638 );
xor ( n33640 , n33633 , n33639 );
xor ( n33641 , n22745 , n22748 );
xor ( n33642 , n33641 , n23007 );
buf ( n33643 , n33642 );
buf ( n33644 , n33643 );
xor ( n33645 , n33640 , n33644 );
buf ( n33646 , n33645 );
not ( n33647 , n33646 );
not ( n33648 , n27513 );
nand ( n33649 , n33647 , n33648 );
xor ( n33650 , n24091 , n24308 );
xor ( n33651 , n33650 , n24444 );
buf ( n33652 , n33651 );
buf ( n33653 , n33652 );
xor ( n33654 , n24322 , n24435 );
xor ( n33655 , n33654 , n24439 );
buf ( n33656 , n33655 );
buf ( n33657 , n33656 );
xor ( n33658 , n24095 , n24267 );
xor ( n33659 , n33658 , n24303 );
buf ( n33660 , n33659 );
buf ( n33661 , n33660 );
xor ( n33662 , n33657 , n33661 );
xor ( n33663 , n24280 , n24290 );
xor ( n33664 , n33663 , n24299 );
buf ( n33665 , n33664 );
not ( n33666 , n24422 );
not ( n33667 , n33666 );
not ( n33668 , n24394 );
not ( n33669 , n20694 );
or ( n33670 , n33668 , n33669 );
nand ( n33671 , n33670 , n24403 );
xor ( n33672 , n33671 , n24388 );
not ( n33673 , n33672 );
or ( n33674 , n33667 , n33673 );
or ( n33675 , n33666 , n33672 );
nand ( n33676 , n33674 , n33675 );
buf ( n33677 , n849 );
buf ( n33678 , n882 );
xor ( n33679 , n33677 , n33678 );
buf ( n33680 , n33679 );
buf ( n33681 , n33680 );
not ( n33682 , n33681 );
buf ( n33683 , n19580 );
not ( n33684 , n33683 );
or ( n33685 , n33682 , n33684 );
buf ( n33686 , n26538 );
buf ( n33687 , n24326 );
nand ( n33688 , n33686 , n33687 );
buf ( n33689 , n33688 );
buf ( n33690 , n33689 );
nand ( n33691 , n33685 , n33690 );
buf ( n33692 , n33691 );
not ( n33693 , n33692 );
not ( n33694 , n24488 );
not ( n33695 , n24476 );
or ( n33696 , n33694 , n33695 );
or ( n33697 , n24476 , n24488 );
nand ( n33698 , n33696 , n33697 );
not ( n33699 , n33698 );
not ( n33700 , n33699 );
or ( n33701 , n33693 , n33700 );
buf ( n33702 , n33692 );
not ( n33703 , n33702 );
buf ( n33704 , n33703 );
buf ( n33705 , n33704 );
not ( n33706 , n33705 );
buf ( n33707 , n33698 );
not ( n33708 , n33707 );
or ( n33709 , n33706 , n33708 );
buf ( n33710 , n18892 );
buf ( n33711 , n863 );
and ( n33712 , n33710 , n33711 );
buf ( n33713 , n33712 );
buf ( n33714 , n33713 );
xor ( n33715 , n888 , n844 );
buf ( n33716 , n33715 );
not ( n33717 , n33716 );
buf ( n33718 , n23144 );
not ( n33719 , n33718 );
or ( n33720 , n33717 , n33719 );
buf ( n33721 , n20363 );
buf ( n33722 , n24509 );
nand ( n33723 , n33721 , n33722 );
buf ( n33724 , n33723 );
buf ( n33725 , n33724 );
nand ( n33726 , n33720 , n33725 );
buf ( n33727 , n33726 );
buf ( n33728 , n33727 );
xor ( n33729 , n33714 , n33728 );
xor ( n33730 , n892 , n840 );
buf ( n33731 , n33730 );
not ( n33732 , n33731 );
buf ( n33733 , n23175 );
not ( n33734 , n33733 );
or ( n33735 , n33732 , n33734 );
buf ( n33736 , n22818 );
buf ( n33737 , n24468 );
nand ( n33738 , n33736 , n33737 );
buf ( n33739 , n33738 );
buf ( n33740 , n33739 );
nand ( n33741 , n33735 , n33740 );
buf ( n33742 , n33741 );
buf ( n33743 , n33742 );
and ( n33744 , n33729 , n33743 );
and ( n33745 , n33714 , n33728 );
or ( n33746 , n33744 , n33745 );
buf ( n33747 , n33746 );
buf ( n33748 , n33747 );
nand ( n33749 , n33709 , n33748 );
buf ( n33750 , n33749 );
nand ( n33751 , n33701 , n33750 );
xor ( n33752 , n33676 , n33751 );
buf ( n33753 , n852 );
buf ( n33754 , n880 );
xor ( n33755 , n33753 , n33754 );
buf ( n33756 , n33755 );
buf ( n33757 , n33756 );
not ( n33758 , n33757 );
buf ( n33759 , n18850 );
not ( n33760 , n33759 );
or ( n33761 , n33758 , n33760 );
buf ( n33762 , n18860 );
buf ( n33763 , n24499 );
nand ( n33764 , n33762 , n33763 );
buf ( n33765 , n33764 );
buf ( n33766 , n33765 );
nand ( n33767 , n33761 , n33766 );
buf ( n33768 , n33767 );
buf ( n33769 , n846 );
buf ( n33770 , n886 );
xor ( n33771 , n33769 , n33770 );
buf ( n33772 , n33771 );
buf ( n33773 , n33772 );
not ( n33774 , n33773 );
buf ( n33775 , n20521 );
not ( n33776 , n33775 );
or ( n33777 , n33774 , n33776 );
buf ( n33778 , n20525 );
buf ( n33779 , n24553 );
nand ( n33780 , n33778 , n33779 );
buf ( n33781 , n33780 );
buf ( n33782 , n33781 );
nand ( n33783 , n33777 , n33782 );
buf ( n33784 , n33783 );
or ( n33785 , n33768 , n33784 );
buf ( n33786 , n854 );
buf ( n33787 , n878 );
xor ( n33788 , n33786 , n33787 );
buf ( n33789 , n33788 );
buf ( n33790 , n33789 );
not ( n33791 , n33790 );
buf ( n33792 , n19259 );
not ( n33793 , n33792 );
or ( n33794 , n33791 , n33793 );
buf ( n33795 , n19265 );
buf ( n33796 , n24530 );
nand ( n33797 , n33795 , n33796 );
buf ( n33798 , n33797 );
buf ( n33799 , n33798 );
nand ( n33800 , n33794 , n33799 );
buf ( n33801 , n33800 );
nand ( n33802 , n33785 , n33801 );
buf ( n33803 , n33784 );
buf ( n33804 , n33768 );
nand ( n33805 , n33803 , n33804 );
buf ( n33806 , n33805 );
nand ( n33807 , n33802 , n33806 );
not ( n33808 , n33807 );
xor ( n33809 , n872 , n860 );
buf ( n33810 , n33809 );
not ( n33811 , n33810 );
buf ( n33812 , n20211 );
not ( n33813 , n33812 );
or ( n33814 , n33811 , n33813 );
buf ( n33815 , n19234 );
buf ( n33816 , n24720 );
nand ( n33817 , n33815 , n33816 );
buf ( n33818 , n33817 );
buf ( n33819 , n33818 );
nand ( n33820 , n33814 , n33819 );
buf ( n33821 , n33820 );
buf ( n33822 , n33821 );
buf ( n33823 , n848 );
buf ( n33824 , n884 );
xor ( n33825 , n33823 , n33824 );
buf ( n33826 , n33825 );
buf ( n33827 , n33826 );
not ( n33828 , n33827 );
buf ( n33829 , n20694 );
not ( n33830 , n33829 );
or ( n33831 , n33828 , n33830 );
buf ( n33832 , n23233 );
buf ( n33833 , n24705 );
nand ( n33834 , n33832 , n33833 );
buf ( n33835 , n33834 );
buf ( n33836 , n33835 );
nand ( n33837 , n33831 , n33836 );
buf ( n33838 , n33837 );
buf ( n33839 , n33838 );
xor ( n33840 , n33822 , n33839 );
buf ( n33841 , n862 );
buf ( n33842 , n870 );
xor ( n33843 , n33841 , n33842 );
buf ( n33844 , n33843 );
buf ( n33845 , n33844 );
not ( n33846 , n33845 );
buf ( n33847 , n19122 );
not ( n33848 , n33847 );
or ( n33849 , n33846 , n33848 );
buf ( n33850 , n19134 );
buf ( n33851 , n24782 );
nand ( n33852 , n33850 , n33851 );
buf ( n33853 , n33852 );
buf ( n33854 , n33853 );
nand ( n33855 , n33849 , n33854 );
buf ( n33856 , n33855 );
buf ( n33857 , n33856 );
and ( n33858 , n33840 , n33857 );
and ( n33859 , n33822 , n33839 );
or ( n33860 , n33858 , n33859 );
buf ( n33861 , n33860 );
not ( n33862 , n33861 );
or ( n33863 , n33808 , n33862 );
nor ( n33864 , n33807 , n33861 );
buf ( n33865 , n838 );
buf ( n33866 , n894 );
xor ( n33867 , n33865 , n33866 );
buf ( n33868 , n33867 );
buf ( n33869 , n33868 );
not ( n33870 , n33869 );
buf ( n33871 , n21297 );
not ( n33872 , n33871 );
or ( n33873 , n33870 , n33872 );
buf ( n33874 , n24688 );
buf ( n33875 , n895 );
nand ( n33876 , n33874 , n33875 );
buf ( n33877 , n33876 );
buf ( n33878 , n33877 );
nand ( n33879 , n33873 , n33878 );
buf ( n33880 , n33879 );
buf ( n33881 , n33880 );
xor ( n33882 , n858 , n874 );
not ( n33883 , n33882 );
not ( n33884 , n18974 );
or ( n33885 , n33883 , n33884 );
nand ( n33886 , n24593 , n21513 );
nand ( n33887 , n33885 , n33886 );
buf ( n33888 , n33887 );
xor ( n33889 , n33881 , n33888 );
buf ( n33890 , n856 );
buf ( n33891 , n876 );
xor ( n33892 , n33890 , n33891 );
buf ( n33893 , n33892 );
not ( n33894 , n33893 );
not ( n33895 , n19153 );
or ( n33896 , n33894 , n33895 );
nand ( n33897 , n24570 , n19082 );
nand ( n33898 , n33896 , n33897 );
buf ( n33899 , n33898 );
and ( n33900 , n33889 , n33899 );
and ( n33901 , n33881 , n33888 );
or ( n33902 , n33900 , n33901 );
buf ( n33903 , n33902 );
buf ( n33904 , n33903 );
not ( n33905 , n33904 );
buf ( n33906 , n33905 );
or ( n33907 , n33864 , n33906 );
nand ( n33908 , n33863 , n33907 );
and ( n33909 , n33752 , n33908 );
and ( n33910 , n33676 , n33751 );
or ( n33911 , n33909 , n33910 );
buf ( n33912 , n33911 );
xor ( n33913 , n33665 , n33912 );
xor ( n33914 , n24491 , n24548 );
xor ( n33915 , n33914 , n24602 );
not ( n33916 , n33915 );
xor ( n33917 , n24738 , n24801 );
xor ( n33918 , n33917 , n24806 );
buf ( n33919 , n33918 );
not ( n33920 , n33919 );
or ( n33921 , n33916 , n33920 );
or ( n33922 , n33919 , n33915 );
buf ( n33923 , n24524 );
not ( n33924 , n33923 );
buf ( n33925 , n24501 );
not ( n33926 , n33925 );
or ( n33927 , n33924 , n33926 );
buf ( n33928 , n24504 );
buf ( n33929 , n24521 );
nand ( n33930 , n33928 , n33929 );
buf ( n33931 , n33930 );
buf ( n33932 , n33931 );
nand ( n33933 , n33927 , n33932 );
buf ( n33934 , n33933 );
not ( n33935 , n24542 );
and ( n33936 , n33934 , n33935 );
not ( n33937 , n33934 );
and ( n33938 , n33937 , n24542 );
nor ( n33939 , n33936 , n33938 );
not ( n33940 , n33939 );
not ( n33941 , n33940 );
xor ( n33942 , n24701 , n24718 );
xor ( n33943 , n33942 , n24733 );
buf ( n33944 , n33943 );
not ( n33945 , n33944 );
or ( n33946 , n33941 , n33945 );
not ( n33947 , n33939 );
buf ( n33948 , n33944 );
not ( n33949 , n33948 );
buf ( n33950 , n33949 );
not ( n33951 , n33950 );
or ( n33952 , n33947 , n33951 );
xor ( n33953 , n24772 , n24754 );
xor ( n33954 , n33953 , n24794 );
nand ( n33955 , n33952 , n33954 );
nand ( n33956 , n33946 , n33955 );
nand ( n33957 , n33922 , n33956 );
nand ( n33958 , n33921 , n33957 );
buf ( n33959 , n33958 );
and ( n33960 , n33913 , n33959 );
and ( n33961 , n33665 , n33912 );
or ( n33962 , n33960 , n33961 );
buf ( n33963 , n33962 );
buf ( n33964 , n33963 );
and ( n33965 , n33662 , n33964 );
and ( n33966 , n33657 , n33661 );
or ( n33967 , n33965 , n33966 );
buf ( n33968 , n33967 );
buf ( n33969 , n33968 );
xor ( n33970 , n33653 , n33969 );
xor ( n33971 , n24453 , n24457 );
xor ( n33972 , n33971 , n24831 );
buf ( n33973 , n33972 );
buf ( n33974 , n33973 );
and ( n33975 , n33970 , n33974 );
and ( n33976 , n33653 , n33969 );
or ( n33977 , n33975 , n33976 );
buf ( n33978 , n33977 );
and ( n33979 , n24854 , n33978 );
nand ( n33980 , n33649 , n33979 );
xor ( n33981 , n33633 , n33639 );
and ( n33982 , n33981 , n33644 );
and ( n33983 , n33633 , n33639 );
or ( n33984 , n33982 , n33983 );
buf ( n33985 , n33984 );
nand ( n33986 , n23014 , n33985 );
nand ( n33987 , n27513 , n33646 );
nand ( n33988 , n33986 , n33987 );
not ( n33989 , n33988 );
buf ( n33990 , n21187 );
buf ( n33991 , n22117 );
xor ( n33992 , n33990 , n33991 );
buf ( n33993 , n22513 );
xor ( n33994 , n33992 , n33993 );
buf ( n33995 , n33994 );
xor ( n33996 , n22544 , n22548 );
and ( n33997 , n33996 , n23012 );
and ( n33998 , n22544 , n22548 );
or ( n33999 , n33997 , n33998 );
buf ( n34000 , n33999 );
nand ( n34001 , n33995 , n34000 );
nand ( n34002 , n33980 , n33989 , n34001 );
nor ( n34003 , n33616 , n34002 );
xor ( n34004 , n23401 , n23683 );
and ( n34005 , n34004 , n23741 );
and ( n34006 , n23401 , n23683 );
or ( n34007 , n34005 , n34006 );
buf ( n34008 , n34007 );
xor ( n34009 , n23788 , n24003 );
and ( n34010 , n34009 , n24026 );
and ( n34011 , n23788 , n24003 );
or ( n34012 , n34010 , n34011 );
buf ( n34013 , n34012 );
xor ( n34014 , n34008 , n34013 );
xor ( n34015 , n33501 , n33505 );
xor ( n34016 , n34015 , n33510 );
buf ( n34017 , n34016 );
buf ( n34018 , n34017 );
and ( n34019 , n34014 , n34018 );
and ( n34020 , n34008 , n34013 );
or ( n34021 , n34019 , n34020 );
buf ( n34022 , n34021 );
not ( n34023 , n34022 );
not ( n34024 , n34023 );
xor ( n34025 , n33495 , n33515 );
xor ( n34026 , n34025 , n33520 );
buf ( n34027 , n34026 );
not ( n34028 , n34027 );
not ( n34029 , n34028 );
or ( n34030 , n34024 , n34029 );
xor ( n34031 , n34008 , n34013 );
xor ( n34032 , n34031 , n34018 );
buf ( n34033 , n34032 );
or ( n34034 , n34033 , n24074 );
nand ( n34035 , n34030 , n34034 );
not ( n34036 , n34035 );
not ( n34037 , n34036 );
or ( n34038 , n34003 , n34037 );
not ( n34039 , n34023 );
nor ( n34040 , n34039 , n34027 );
nand ( n34041 , n34033 , n24074 );
or ( n34042 , n34040 , n34041 );
not ( n34043 , n34023 );
buf ( n34044 , n34027 );
nand ( n34045 , n34043 , n34044 );
nand ( n34046 , n34042 , n34045 );
not ( n34047 , n34046 );
nand ( n34048 , n34038 , n34047 );
not ( n34049 , n33616 );
not ( n34050 , n33603 );
nand ( n34051 , n34050 , n33599 );
not ( n34052 , n33613 );
not ( n34053 , n22525 );
nand ( n34054 , n34052 , n34053 );
nand ( n34055 , n34051 , n34054 );
not ( n34056 , n34055 );
nor ( n34057 , n33995 , n34000 );
nor ( n34058 , n23014 , n33985 );
or ( n34059 , n34057 , n34058 );
nand ( n34060 , n34059 , n34001 );
nand ( n34061 , n34056 , n34060 );
nand ( n34062 , n34049 , n34061 , n34047 );
nand ( n34063 , n33476 , n33525 );
nand ( n34064 , n34063 , n33535 );
nor ( n34065 , n33428 , n34064 );
nand ( n34066 , n34065 , n33395 );
not ( n34067 , n34066 );
nand ( n34068 , n34048 , n34062 , n34067 );
nand ( n34069 , n33572 , n34068 );
not ( n34070 , n34069 );
or ( n34071 , n32840 , n34070 );
not ( n34072 , n33646 );
not ( n34073 , n27513 );
and ( n34074 , n34072 , n34073 );
nor ( n34075 , n24854 , n33978 );
nor ( n34076 , n34074 , n34075 );
not ( n34077 , n34076 );
not ( n34078 , n33995 );
not ( n34079 , n34000 );
nand ( n34080 , n34078 , n34079 );
not ( n34081 , n23014 );
not ( n34082 , n33985 );
nand ( n34083 , n34081 , n34082 );
nand ( n34084 , n34080 , n34083 );
nor ( n34085 , n34077 , n34084 );
not ( n34086 , n34053 );
not ( n34087 , n34052 );
or ( n34088 , n34086 , n34087 );
nand ( n34089 , n34088 , n34051 );
nor ( n34090 , n34035 , n34089 );
nand ( n34091 , n34085 , n34090 );
nor ( n34092 , n34091 , n34066 );
not ( n34093 , n34092 );
not ( n34094 , n34093 );
and ( n34095 , n34094 , n32839 );
buf ( n34096 , n842 );
buf ( n34097 , n890 );
xor ( n34098 , n34096 , n34097 );
buf ( n34099 , n34098 );
buf ( n34100 , n34099 );
not ( n34101 , n34100 );
buf ( n34102 , n21441 );
not ( n34103 , n34102 );
or ( n34104 , n34101 , n34103 );
buf ( n34105 , n20869 );
buf ( n34106 , n24742 );
nand ( n34107 , n34105 , n34106 );
buf ( n34108 , n34107 );
buf ( n34109 , n34108 );
nand ( n34110 , n34104 , n34109 );
buf ( n34111 , n34110 );
not ( n34112 , n34111 );
buf ( n34113 , n850 );
buf ( n34114 , n882 );
xor ( n34115 , n34113 , n34114 );
buf ( n34116 , n34115 );
buf ( n34117 , n34116 );
not ( n34118 , n34117 );
buf ( n34119 , n19580 );
not ( n34120 , n34119 );
or ( n34121 , n34118 , n34120 );
buf ( n34122 , n26538 );
buf ( n34123 , n33680 );
nand ( n34124 , n34122 , n34123 );
buf ( n34125 , n34124 );
buf ( n34126 , n34125 );
nand ( n34127 , n34121 , n34126 );
buf ( n34128 , n34127 );
not ( n34129 , n34128 );
nand ( n34130 , n34112 , n34129 );
not ( n34131 , n34130 );
buf ( n34132 , n863 );
buf ( n34133 , n871 );
or ( n34134 , n34132 , n34133 );
buf ( n34135 , n872 );
nand ( n34136 , n34134 , n34135 );
buf ( n34137 , n34136 );
buf ( n34138 , n34137 );
buf ( n34139 , n863 );
buf ( n34140 , n871 );
nand ( n34141 , n34139 , n34140 );
buf ( n34142 , n34141 );
buf ( n34143 , n34142 );
buf ( n34144 , n870 );
nand ( n34145 , n34138 , n34143 , n34144 );
buf ( n34146 , n34145 );
not ( n34147 , n34146 );
buf ( n34148 , n841 );
buf ( n34149 , n892 );
xor ( n34150 , n34148 , n34149 );
buf ( n34151 , n34150 );
buf ( n34152 , n34151 );
not ( n34153 , n34152 );
buf ( n34154 , n23175 );
not ( n34155 , n34154 );
or ( n34156 , n34153 , n34155 );
buf ( n34157 , n22818 );
buf ( n34158 , n33730 );
nand ( n34159 , n34157 , n34158 );
buf ( n34160 , n34159 );
buf ( n34161 , n34160 );
nand ( n34162 , n34156 , n34161 );
buf ( n34163 , n34162 );
nand ( n34164 , n34147 , n34163 );
not ( n34165 , n34164 );
not ( n34166 , n34165 );
or ( n34167 , n34131 , n34166 );
nand ( n34168 , n34128 , n34111 );
nand ( n34169 , n34167 , n34168 );
xor ( n34170 , n24565 , n24582 );
buf ( n34171 , n34170 );
buf ( n34172 , n24600 );
xnor ( n34173 , n34171 , n34172 );
buf ( n34174 , n34173 );
xor ( n34175 , n34169 , n34174 );
and ( n34176 , n33699 , n33692 );
not ( n34177 , n33699 );
and ( n34178 , n34177 , n33704 );
nor ( n34179 , n34176 , n34178 );
buf ( n34180 , n33747 );
and ( n34181 , n34179 , n34180 );
not ( n34182 , n34179 );
not ( n34183 , n34180 );
and ( n34184 , n34182 , n34183 );
nor ( n34185 , n34181 , n34184 );
xor ( n34186 , n34175 , n34185 );
buf ( n34187 , n34186 );
buf ( n34188 , n34187 );
not ( n34189 , n34188 );
xor ( n34190 , n33822 , n33839 );
xor ( n34191 , n34190 , n33857 );
buf ( n34192 , n34191 );
buf ( n34193 , n34192 );
xor ( n34194 , n33768 , n33784 );
and ( n34195 , n34194 , n33801 );
not ( n34196 , n34194 );
buf ( n34197 , n33801 );
not ( n34198 , n34197 );
buf ( n34199 , n34198 );
and ( n34200 , n34196 , n34199 );
nor ( n34201 , n34195 , n34200 );
buf ( n34202 , n34201 );
xor ( n34203 , n34193 , n34202 );
xor ( n34204 , n34111 , n34129 );
xor ( n34205 , n34204 , n34164 );
buf ( n34206 , n34205 );
and ( n34207 , n34203 , n34206 );
and ( n34208 , n34193 , n34202 );
or ( n34209 , n34207 , n34208 );
buf ( n34210 , n34209 );
buf ( n34211 , n34210 );
not ( n34212 , n34211 );
not ( n34213 , n33940 );
and ( n34214 , n33954 , n34213 );
not ( n34215 , n33954 );
and ( n34216 , n34215 , n33940 );
nor ( n34217 , n34214 , n34216 );
buf ( n34218 , n34217 );
buf ( n34219 , n33944 );
and ( n34220 , n34218 , n34219 );
not ( n34221 , n34218 );
buf ( n34222 , n33950 );
buf ( n34223 , n34222 );
and ( n34224 , n34221 , n34223 );
nor ( n34225 , n34220 , n34224 );
buf ( n34226 , n34225 );
buf ( n34227 , n34226 );
not ( n34228 , n34227 );
and ( n34229 , n34212 , n34228 );
buf ( n34230 , n34210 );
buf ( n34231 , n34226 );
and ( n34232 , n34230 , n34231 );
nor ( n34233 , n34229 , n34232 );
buf ( n34234 , n34233 );
buf ( n34235 , n34234 );
not ( n34236 , n34235 );
or ( n34237 , n34189 , n34236 );
buf ( n34238 , n34234 );
buf ( n34239 , n34187 );
or ( n34240 , n34238 , n34239 );
nand ( n34241 , n34237 , n34240 );
buf ( n34242 , n34241 );
buf ( n34243 , n34242 );
buf ( n34244 , n852 );
buf ( n34245 , n882 );
xor ( n34246 , n34244 , n34245 );
buf ( n34247 , n34246 );
buf ( n34248 , n34247 );
not ( n34249 , n34248 );
buf ( n34250 , n26534 );
not ( n34251 , n34250 );
or ( n34252 , n34249 , n34251 );
buf ( n34253 , n26538 );
buf ( n34254 , n851 );
buf ( n34255 , n882 );
xor ( n34256 , n34254 , n34255 );
buf ( n34257 , n34256 );
buf ( n34258 , n34257 );
nand ( n34259 , n34253 , n34258 );
buf ( n34260 , n34259 );
buf ( n34261 , n34260 );
nand ( n34262 , n34252 , n34261 );
buf ( n34263 , n34262 );
buf ( n34264 , n34263 );
buf ( n34265 , n29776 );
not ( n34266 , n34265 );
buf ( n34267 , n20599 );
not ( n34268 , n34267 );
or ( n34269 , n34266 , n34268 );
buf ( n34270 , n23181 );
buf ( n34271 , n842 );
buf ( n34272 , n892 );
xor ( n34273 , n34271 , n34272 );
buf ( n34274 , n34273 );
buf ( n34275 , n34274 );
nand ( n34276 , n34270 , n34275 );
buf ( n34277 , n34276 );
buf ( n34278 , n34277 );
nand ( n34279 , n34269 , n34278 );
buf ( n34280 , n34279 );
buf ( n34281 , n34280 );
not ( n34282 , n34281 );
buf ( n34283 , n863 );
buf ( n34284 , n873 );
or ( n34285 , n34283 , n34284 );
buf ( n34286 , n874 );
nand ( n34287 , n34285 , n34286 );
buf ( n34288 , n34287 );
buf ( n34289 , n34288 );
buf ( n34290 , n863 );
buf ( n34291 , n873 );
nand ( n34292 , n34290 , n34291 );
buf ( n34293 , n34292 );
buf ( n34294 , n34293 );
buf ( n34295 , n872 );
nand ( n34296 , n34289 , n34294 , n34295 );
buf ( n34297 , n34296 );
buf ( n34298 , n34297 );
nor ( n34299 , n34282 , n34298 );
buf ( n34300 , n34299 );
buf ( n34301 , n34300 );
xor ( n34302 , n34264 , n34301 );
buf ( n34303 , n29813 );
not ( n34304 , n34303 );
buf ( n34305 , n19077 );
not ( n34306 , n34305 );
or ( n34307 , n34304 , n34306 );
buf ( n34308 , n20246 );
buf ( n34309 , n858 );
buf ( n34310 , n876 );
xor ( n34311 , n34309 , n34310 );
buf ( n34312 , n34311 );
buf ( n34313 , n34312 );
nand ( n34314 , n34308 , n34313 );
buf ( n34315 , n34314 );
buf ( n34316 , n34315 );
nand ( n34317 , n34307 , n34316 );
buf ( n34318 , n34317 );
buf ( n34319 , n34318 );
buf ( n34320 , n29831 );
not ( n34321 , n34320 );
buf ( n34322 , n18974 );
not ( n34323 , n34322 );
or ( n34324 , n34321 , n34323 );
buf ( n34325 , n21513 );
buf ( n34326 , n860 );
buf ( n34327 , n874 );
xor ( n34328 , n34326 , n34327 );
buf ( n34329 , n34328 );
buf ( n34330 , n34329 );
nand ( n34331 , n34325 , n34330 );
buf ( n34332 , n34331 );
buf ( n34333 , n34332 );
nand ( n34334 , n34324 , n34333 );
buf ( n34335 , n34334 );
buf ( n34336 , n34335 );
xor ( n34337 , n34319 , n34336 );
not ( n34338 , n23320 );
buf ( n34339 , n848 );
buf ( n34340 , n886 );
xor ( n34341 , n34339 , n34340 );
buf ( n34342 , n34341 );
not ( n34343 , n34342 );
or ( n34344 , n34338 , n34343 );
buf ( n34345 , n29706 );
not ( n34346 , n34345 );
buf ( n34347 , n34346 );
or ( n34348 , n23024 , n34347 );
nand ( n34349 , n34344 , n34348 );
buf ( n34350 , n34349 );
and ( n34351 , n34337 , n34350 );
and ( n34352 , n34319 , n34336 );
or ( n34353 , n34351 , n34352 );
buf ( n34354 , n34353 );
buf ( n34355 , n34354 );
and ( n34356 , n34302 , n34355 );
and ( n34357 , n34264 , n34301 );
or ( n34358 , n34356 , n34357 );
buf ( n34359 , n34358 );
buf ( n34360 , n34359 );
buf ( n34361 , n19131 );
buf ( n34362 , n863 );
and ( n34363 , n34361 , n34362 );
buf ( n34364 , n34363 );
buf ( n34365 , n34364 );
not ( n34366 , n34365 );
buf ( n34367 , n846 );
buf ( n34368 , n888 );
xor ( n34369 , n34367 , n34368 );
buf ( n34370 , n34369 );
buf ( n34371 , n34370 );
not ( n34372 , n34371 );
buf ( n34373 , n22303 );
not ( n34374 , n34373 );
or ( n34375 , n34372 , n34374 );
buf ( n34376 , n20363 );
buf ( n34377 , n845 );
buf ( n34378 , n888 );
xor ( n34379 , n34377 , n34378 );
buf ( n34380 , n34379 );
buf ( n34381 , n34380 );
nand ( n34382 , n34376 , n34381 );
buf ( n34383 , n34382 );
buf ( n34384 , n34383 );
nand ( n34385 , n34375 , n34384 );
buf ( n34386 , n34385 );
buf ( n34387 , n34386 );
not ( n34388 , n34387 );
or ( n34389 , n34366 , n34388 );
buf ( n34390 , n34386 );
buf ( n34391 , n34364 );
or ( n34392 , n34390 , n34391 );
buf ( n34393 , n34274 );
not ( n34394 , n34393 );
buf ( n34395 , n23175 );
not ( n34396 , n34395 );
or ( n34397 , n34394 , n34396 );
buf ( n34398 , n22818 );
buf ( n34399 , n34151 );
nand ( n34400 , n34398 , n34399 );
buf ( n34401 , n34400 );
buf ( n34402 , n34401 );
nand ( n34403 , n34397 , n34402 );
buf ( n34404 , n34403 );
buf ( n34405 , n34404 );
nand ( n34406 , n34392 , n34405 );
buf ( n34407 , n34406 );
buf ( n34408 , n34407 );
nand ( n34409 , n34389 , n34408 );
buf ( n34410 , n34409 );
buf ( n34411 , n34410 );
buf ( n34412 , n862 );
buf ( n34413 , n872 );
xor ( n34414 , n34412 , n34413 );
buf ( n34415 , n34414 );
buf ( n34416 , n34415 );
not ( n34417 , n34416 );
buf ( n34418 , n25285 );
not ( n34419 , n34418 );
or ( n34420 , n34417 , n34419 );
buf ( n34421 , n19234 );
buf ( n34422 , n861 );
buf ( n34423 , n872 );
xor ( n34424 , n34422 , n34423 );
buf ( n34425 , n34424 );
buf ( n34426 , n34425 );
nand ( n34427 , n34421 , n34426 );
buf ( n34428 , n34427 );
buf ( n34429 , n34428 );
nand ( n34430 , n34420 , n34429 );
buf ( n34431 , n34430 );
buf ( n34432 , n34431 );
not ( n34433 , n34432 );
buf ( n34434 , n844 );
buf ( n34435 , n890 );
xor ( n34436 , n34434 , n34435 );
buf ( n34437 , n34436 );
buf ( n34438 , n34437 );
not ( n34439 , n34438 );
buf ( n34440 , n21441 );
not ( n34441 , n34440 );
or ( n34442 , n34439 , n34441 );
buf ( n34443 , n20869 );
buf ( n34444 , n843 );
buf ( n34445 , n890 );
xor ( n34446 , n34444 , n34445 );
buf ( n34447 , n34446 );
buf ( n34448 , n34447 );
nand ( n34449 , n34443 , n34448 );
buf ( n34450 , n34449 );
buf ( n34451 , n34450 );
nand ( n34452 , n34442 , n34451 );
buf ( n34453 , n34452 );
buf ( n34454 , n34453 );
not ( n34455 , n34454 );
or ( n34456 , n34433 , n34455 );
buf ( n34457 , n34453 );
buf ( n34458 , n34431 );
or ( n34459 , n34457 , n34458 );
buf ( n34460 , n850 );
buf ( n34461 , n884 );
xor ( n34462 , n34460 , n34461 );
buf ( n34463 , n34462 );
buf ( n34464 , n34463 );
not ( n34465 , n34464 );
buf ( n34466 , n20694 );
not ( n34467 , n34466 );
or ( n34468 , n34465 , n34467 );
buf ( n34469 , n25263 );
buf ( n34470 , n849 );
buf ( n34471 , n884 );
xor ( n34472 , n34470 , n34471 );
buf ( n34473 , n34472 );
buf ( n34474 , n34473 );
nand ( n34475 , n34469 , n34474 );
buf ( n34476 , n34475 );
buf ( n34477 , n34476 );
nand ( n34478 , n34468 , n34477 );
buf ( n34479 , n34478 );
buf ( n34480 , n34479 );
nand ( n34481 , n34459 , n34480 );
buf ( n34482 , n34481 );
buf ( n34483 , n34482 );
nand ( n34484 , n34456 , n34483 );
buf ( n34485 , n34484 );
buf ( n34486 , n34485 );
xor ( n34487 , n34411 , n34486 );
buf ( n34488 , n34257 );
not ( n34489 , n34488 );
buf ( n34490 , n19580 );
not ( n34491 , n34490 );
or ( n34492 , n34489 , n34491 );
buf ( n34493 , n19909 );
buf ( n34494 , n34116 );
nand ( n34495 , n34493 , n34494 );
buf ( n34496 , n34495 );
buf ( n34497 , n34496 );
nand ( n34498 , n34492 , n34497 );
buf ( n34499 , n34498 );
buf ( n34500 , n34499 );
buf ( n34501 , n863 );
buf ( n34502 , n870 );
xor ( n34503 , n34501 , n34502 );
buf ( n34504 , n34503 );
buf ( n34505 , n34504 );
not ( n34506 , n34505 );
buf ( n34507 , n19122 );
not ( n34508 , n34507 );
or ( n34509 , n34506 , n34508 );
buf ( n34510 , n19131 );
buf ( n34511 , n33844 );
nand ( n34512 , n34510 , n34511 );
buf ( n34513 , n34512 );
buf ( n34514 , n34513 );
nand ( n34515 , n34509 , n34514 );
buf ( n34516 , n34515 );
buf ( n34517 , n34516 );
xor ( n34518 , n34500 , n34517 );
buf ( n34519 , n34447 );
not ( n34520 , n34519 );
buf ( n34521 , n21441 );
not ( n34522 , n34521 );
or ( n34523 , n34520 , n34522 );
buf ( n34524 , n20869 );
buf ( n34525 , n34099 );
nand ( n34526 , n34524 , n34525 );
buf ( n34527 , n34526 );
buf ( n34528 , n34527 );
nand ( n34529 , n34523 , n34528 );
buf ( n34530 , n34529 );
buf ( n34531 , n34530 );
xor ( n34532 , n34518 , n34531 );
buf ( n34533 , n34532 );
buf ( n34534 , n34533 );
xor ( n34535 , n34487 , n34534 );
buf ( n34536 , n34535 );
buf ( n34537 , n34536 );
xor ( n34538 , n34360 , n34537 );
buf ( n34539 , n34404 );
buf ( n34540 , n21727 );
buf ( n34541 , n863 );
and ( n34542 , n34540 , n34541 );
buf ( n34543 , n34542 );
buf ( n34544 , n34543 );
and ( n34545 , n34539 , n34544 );
not ( n34546 , n34539 );
buf ( n34547 , n34543 );
not ( n34548 , n34547 );
buf ( n34549 , n34548 );
buf ( n34550 , n34549 );
and ( n34551 , n34546 , n34550 );
nor ( n34552 , n34545 , n34551 );
buf ( n34553 , n34552 );
buf ( n34554 , n34553 );
buf ( n34555 , n34386 );
and ( n34556 , n34554 , n34555 );
not ( n34557 , n34554 );
buf ( n34558 , n34386 );
not ( n34559 , n34558 );
buf ( n34560 , n34559 );
buf ( n34561 , n34560 );
and ( n34562 , n34557 , n34561 );
nor ( n34563 , n34556 , n34562 );
buf ( n34564 , n34563 );
buf ( n34565 , n34564 );
not ( n34566 , n34565 );
not ( n34567 , n34342 );
not ( n34568 , n20521 );
or ( n34569 , n34567 , n34568 );
buf ( n34570 , n20525 );
buf ( n34571 , n847 );
buf ( n34572 , n886 );
xor ( n34573 , n34571 , n34572 );
buf ( n34574 , n34573 );
buf ( n34575 , n34574 );
nand ( n34576 , n34570 , n34575 );
buf ( n34577 , n34576 );
nand ( n34578 , n34569 , n34577 );
buf ( n34579 , n854 );
buf ( n34580 , n880 );
xor ( n34581 , n34579 , n34580 );
buf ( n34582 , n34581 );
not ( n34583 , n34582 );
not ( n34584 , n18850 );
or ( n34585 , n34583 , n34584 );
buf ( n34586 , n20325 );
buf ( n34587 , n853 );
buf ( n34588 , n880 );
xor ( n34589 , n34587 , n34588 );
buf ( n34590 , n34589 );
buf ( n34591 , n34590 );
nand ( n34592 , n34586 , n34591 );
buf ( n34593 , n34592 );
nand ( n34594 , n34585 , n34593 );
xor ( n34595 , n34578 , n34594 );
buf ( n34596 , n856 );
buf ( n34597 , n878 );
xor ( n34598 , n34596 , n34597 );
buf ( n34599 , n34598 );
not ( n34600 , n34599 );
not ( n34601 , n19259 );
or ( n34602 , n34600 , n34601 );
buf ( n34603 , n19265 );
buf ( n34604 , n855 );
buf ( n34605 , n878 );
xor ( n34606 , n34604 , n34605 );
buf ( n34607 , n34606 );
buf ( n34608 , n34607 );
nand ( n34609 , n34603 , n34608 );
buf ( n34610 , n34609 );
nand ( n34611 , n34602 , n34610 );
xor ( n34612 , n34595 , n34611 );
buf ( n34613 , n34612 );
not ( n34614 , n34613 );
or ( n34615 , n34566 , n34614 );
buf ( n34616 , n34612 );
buf ( n34617 , n34564 );
or ( n34618 , n34616 , n34617 );
buf ( n34619 , n840 );
buf ( n34620 , n894 );
xor ( n34621 , n34619 , n34620 );
buf ( n34622 , n34621 );
buf ( n34623 , n34622 );
not ( n34624 , n34623 );
buf ( n34625 , n21297 );
not ( n34626 , n34625 );
or ( n34627 , n34624 , n34626 );
buf ( n34628 , n839 );
buf ( n34629 , n894 );
xor ( n34630 , n34628 , n34629 );
buf ( n34631 , n34630 );
buf ( n34632 , n34631 );
buf ( n34633 , n895 );
nand ( n34634 , n34632 , n34633 );
buf ( n34635 , n34634 );
buf ( n34636 , n34635 );
nand ( n34637 , n34627 , n34636 );
buf ( n34638 , n34637 );
buf ( n34639 , n34638 );
buf ( n34640 , n34312 );
not ( n34641 , n34640 );
buf ( n34642 , n19077 );
not ( n34643 , n34642 );
or ( n34644 , n34641 , n34643 );
buf ( n34645 , n19082 );
buf ( n34646 , n857 );
buf ( n34647 , n876 );
xor ( n34648 , n34646 , n34647 );
buf ( n34649 , n34648 );
buf ( n34650 , n34649 );
nand ( n34651 , n34645 , n34650 );
buf ( n34652 , n34651 );
buf ( n34653 , n34652 );
nand ( n34654 , n34644 , n34653 );
buf ( n34655 , n34654 );
buf ( n34656 , n34655 );
xor ( n34657 , n34639 , n34656 );
buf ( n34658 , n34329 );
not ( n34659 , n34658 );
buf ( n34660 , n18977 );
not ( n34661 , n34660 );
or ( n34662 , n34659 , n34661 );
buf ( n34663 , n18987 );
xor ( n34664 , n874 , n859 );
buf ( n34665 , n34664 );
nand ( n34666 , n34663 , n34665 );
buf ( n34667 , n34666 );
buf ( n34668 , n34667 );
nand ( n34669 , n34662 , n34668 );
buf ( n34670 , n34669 );
buf ( n34671 , n34670 );
xor ( n34672 , n34657 , n34671 );
buf ( n34673 , n34672 );
buf ( n34674 , n34673 );
nand ( n34675 , n34618 , n34674 );
buf ( n34676 , n34675 );
buf ( n34677 , n34676 );
nand ( n34678 , n34615 , n34677 );
buf ( n34679 , n34678 );
buf ( n34680 , n34679 );
and ( n34681 , n34538 , n34680 );
and ( n34682 , n34360 , n34537 );
or ( n34683 , n34681 , n34682 );
buf ( n34684 , n34683 );
buf ( n34685 , n34684 );
not ( n34686 , n23288 );
not ( n34687 , n29795 );
or ( n34688 , n34686 , n34687 );
buf ( n34689 , n34622 );
buf ( n34690 , n895 );
nand ( n34691 , n34689 , n34690 );
buf ( n34692 , n34691 );
nand ( n34693 , n34688 , n34692 );
not ( n34694 , n29650 );
not ( n34695 , n21441 );
or ( n34696 , n34694 , n34695 );
buf ( n34697 , n20869 );
buf ( n34698 , n34437 );
nand ( n34699 , n34697 , n34698 );
buf ( n34700 , n34699 );
nand ( n34701 , n34696 , n34700 );
xor ( n34702 , n34693 , n34701 );
not ( n34703 , n19235 );
not ( n34704 , n34415 );
or ( n34705 , n34703 , n34704 );
buf ( n34706 , n863 );
buf ( n34707 , n872 );
xor ( n34708 , n34706 , n34707 );
buf ( n34709 , n34708 );
nand ( n34710 , n19230 , n34709 );
nand ( n34711 , n34705 , n34710 );
and ( n34712 , n34702 , n34711 );
and ( n34713 , n34693 , n34701 );
or ( n34714 , n34712 , n34713 );
buf ( n34715 , n34714 );
xor ( n34716 , n34431 , n34453 );
xor ( n34717 , n34716 , n34479 );
buf ( n34718 , n34717 );
xor ( n34719 , n34715 , n34718 );
not ( n34720 , n29757 );
not ( n34721 , n23144 );
or ( n34722 , n34720 , n34721 );
buf ( n34723 , n20363 );
buf ( n34724 , n34370 );
nand ( n34725 , n34723 , n34724 );
buf ( n34726 , n34725 );
nand ( n34727 , n34722 , n34726 );
not ( n34728 , n34727 );
not ( n34729 , n34728 );
buf ( n34730 , n29735 );
not ( n34731 , n34730 );
buf ( n34732 , n19259 );
not ( n34733 , n34732 );
or ( n34734 , n34731 , n34733 );
buf ( n34735 , n19265 );
buf ( n34736 , n34599 );
nand ( n34737 , n34735 , n34736 );
buf ( n34738 , n34737 );
buf ( n34739 , n34738 );
nand ( n34740 , n34734 , n34739 );
buf ( n34741 , n34740 );
not ( n34742 , n34741 );
not ( n34743 , n34742 );
or ( n34744 , n34729 , n34743 );
buf ( n34745 , n29720 );
not ( n34746 , n34745 );
buf ( n34747 , n19614 );
not ( n34748 , n34747 );
or ( n34749 , n34746 , n34748 );
buf ( n34750 , n22271 );
buf ( n34751 , n34582 );
nand ( n34752 , n34750 , n34751 );
buf ( n34753 , n34752 );
buf ( n34754 , n34753 );
nand ( n34755 , n34749 , n34754 );
buf ( n34756 , n34755 );
nand ( n34757 , n34744 , n34756 );
nand ( n34758 , n34741 , n34727 );
nand ( n34759 , n34757 , n34758 );
buf ( n34760 , n34759 );
and ( n34761 , n34719 , n34760 );
and ( n34762 , n34715 , n34718 );
or ( n34763 , n34761 , n34762 );
buf ( n34764 , n34763 );
buf ( n34765 , n34764 );
not ( n34766 , n34765 );
or ( n34767 , n34594 , n34578 );
nand ( n34768 , n34767 , n34611 );
nand ( n34769 , n34594 , n34578 );
nand ( n34770 , n34768 , n34769 );
not ( n34771 , n34146 );
not ( n34772 , n34771 );
not ( n34773 , n34163 );
or ( n34774 , n34772 , n34773 );
or ( n34775 , n34163 , n34771 );
nand ( n34776 , n34774 , n34775 );
xor ( n34777 , n34770 , n34776 );
xor ( n34778 , n34639 , n34656 );
and ( n34779 , n34778 , n34671 );
and ( n34780 , n34639 , n34656 );
or ( n34781 , n34779 , n34780 );
buf ( n34782 , n34781 );
xor ( n34783 , n34777 , n34782 );
buf ( n34784 , n34783 );
not ( n34785 , n34784 );
buf ( n34786 , n34785 );
buf ( n34787 , n34786 );
not ( n34788 , n34787 );
or ( n34789 , n34766 , n34788 );
buf ( n34790 , n34783 );
not ( n34791 , n34790 );
buf ( n34792 , n34764 );
not ( n34793 , n34792 );
buf ( n34794 , n34793 );
buf ( n34795 , n34794 );
not ( n34796 , n34795 );
or ( n34797 , n34791 , n34796 );
buf ( n34798 , n34631 );
not ( n34799 , n34798 );
buf ( n34800 , n20132 );
not ( n34801 , n34800 );
or ( n34802 , n34799 , n34801 );
buf ( n34803 , n33868 );
buf ( n34804 , n895 );
nand ( n34805 , n34803 , n34804 );
buf ( n34806 , n34805 );
buf ( n34807 , n34806 );
nand ( n34808 , n34802 , n34807 );
buf ( n34809 , n34808 );
buf ( n34810 , n34809 );
buf ( n34811 , n34473 );
not ( n34812 , n34811 );
buf ( n34813 , n20694 );
not ( n34814 , n34813 );
or ( n34815 , n34812 , n34814 );
buf ( n34816 , n20700 );
buf ( n34817 , n33826 );
nand ( n34818 , n34816 , n34817 );
buf ( n34819 , n34818 );
buf ( n34820 , n34819 );
nand ( n34821 , n34815 , n34820 );
buf ( n34822 , n34821 );
buf ( n34823 , n34822 );
xor ( n34824 , n34810 , n34823 );
buf ( n34825 , n34425 );
not ( n34826 , n34825 );
buf ( n34827 , n25285 );
not ( n34828 , n34827 );
or ( n34829 , n34826 , n34828 );
buf ( n34830 , n19235 );
buf ( n34831 , n33809 );
nand ( n34832 , n34830 , n34831 );
buf ( n34833 , n34832 );
buf ( n34834 , n34833 );
nand ( n34835 , n34829 , n34834 );
buf ( n34836 , n34835 );
buf ( n34837 , n34836 );
xor ( n34838 , n34824 , n34837 );
buf ( n34839 , n34838 );
buf ( n34840 , n34839 );
buf ( n34841 , n34590 );
not ( n34842 , n34841 );
buf ( n34843 , n18850 );
not ( n34844 , n34843 );
or ( n34845 , n34842 , n34844 );
buf ( n34846 , n18860 );
buf ( n34847 , n33756 );
nand ( n34848 , n34846 , n34847 );
buf ( n34849 , n34848 );
buf ( n34850 , n34849 );
nand ( n34851 , n34845 , n34850 );
buf ( n34852 , n34851 );
buf ( n34853 , n34380 );
not ( n34854 , n34853 );
buf ( n34855 , n22303 );
not ( n34856 , n34855 );
or ( n34857 , n34854 , n34856 );
buf ( n34858 , n20363 );
buf ( n34859 , n33715 );
nand ( n34860 , n34858 , n34859 );
buf ( n34861 , n34860 );
buf ( n34862 , n34861 );
nand ( n34863 , n34857 , n34862 );
buf ( n34864 , n34863 );
xor ( n34865 , n34852 , n34864 );
buf ( n34866 , n34607 );
not ( n34867 , n34866 );
buf ( n34868 , n19259 );
not ( n34869 , n34868 );
or ( n34870 , n34867 , n34869 );
buf ( n34871 , n19265 );
buf ( n34872 , n33789 );
nand ( n34873 , n34871 , n34872 );
buf ( n34874 , n34873 );
buf ( n34875 , n34874 );
nand ( n34876 , n34870 , n34875 );
buf ( n34877 , n34876 );
xor ( n34878 , n34865 , n34877 );
buf ( n34879 , n34878 );
xor ( n34880 , n34840 , n34879 );
buf ( n34881 , n34649 );
not ( n34882 , n34881 );
buf ( n34883 , n19153 );
not ( n34884 , n34883 );
or ( n34885 , n34882 , n34884 );
buf ( n34886 , n19082 );
buf ( n34887 , n33893 );
nand ( n34888 , n34886 , n34887 );
buf ( n34889 , n34888 );
buf ( n34890 , n34889 );
nand ( n34891 , n34885 , n34890 );
buf ( n34892 , n34891 );
buf ( n34893 , n34574 );
not ( n34894 , n34893 );
buf ( n34895 , n21817 );
not ( n34896 , n34895 );
or ( n34897 , n34894 , n34896 );
buf ( n34898 , n20525 );
buf ( n34899 , n33772 );
nand ( n34900 , n34898 , n34899 );
buf ( n34901 , n34900 );
buf ( n34902 , n34901 );
nand ( n34903 , n34897 , n34902 );
buf ( n34904 , n34903 );
xor ( n34905 , n34892 , n34904 );
buf ( n34906 , n18977 );
buf ( n34907 , n34664 );
and ( n34908 , n34906 , n34907 );
buf ( n34909 , n20555 );
buf ( n34910 , n33882 );
and ( n34911 , n34909 , n34910 );
nor ( n34912 , n34908 , n34911 );
buf ( n34913 , n34912 );
xnor ( n34914 , n34905 , n34913 );
buf ( n34915 , n34914 );
xor ( n34916 , n34880 , n34915 );
buf ( n34917 , n34916 );
buf ( n34918 , n34917 );
nand ( n34919 , n34797 , n34918 );
buf ( n34920 , n34919 );
buf ( n34921 , n34920 );
nand ( n34922 , n34789 , n34921 );
buf ( n34923 , n34922 );
buf ( n34924 , n34923 );
xor ( n34925 , n34685 , n34924 );
buf ( n34926 , n34776 );
not ( n34927 , n34926 );
buf ( n34928 , n34770 );
not ( n34929 , n34928 );
buf ( n34930 , n34929 );
buf ( n34931 , n34930 );
not ( n34932 , n34931 );
or ( n34933 , n34927 , n34932 );
buf ( n34934 , n34782 );
nand ( n34935 , n34933 , n34934 );
buf ( n34936 , n34935 );
buf ( n34937 , n34936 );
not ( n34938 , n34769 );
not ( n34939 , n34768 );
or ( n34940 , n34938 , n34939 );
not ( n34941 , n34776 );
nand ( n34942 , n34940 , n34941 );
buf ( n34943 , n34942 );
nand ( n34944 , n34937 , n34943 );
buf ( n34945 , n34944 );
buf ( n34946 , n34945 );
xor ( n34947 , n34411 , n34486 );
and ( n34948 , n34947 , n34534 );
and ( n34949 , n34411 , n34486 );
or ( n34950 , n34948 , n34949 );
buf ( n34951 , n34950 );
buf ( n34952 , n34951 );
xor ( n34953 , n34946 , n34952 );
xor ( n34954 , n34840 , n34879 );
and ( n34955 , n34954 , n34915 );
and ( n34956 , n34840 , n34879 );
or ( n34957 , n34955 , n34956 );
buf ( n34958 , n34957 );
buf ( n34959 , n34958 );
xor ( n34960 , n34953 , n34959 );
buf ( n34961 , n34960 );
buf ( n34962 , n34961 );
and ( n34963 , n34925 , n34962 );
and ( n34964 , n34685 , n34924 );
or ( n34965 , n34963 , n34964 );
buf ( n34966 , n34965 );
buf ( n34967 , n34966 );
xor ( n34968 , n34243 , n34967 );
xor ( n34969 , n34946 , n34952 );
and ( n34970 , n34969 , n34959 );
and ( n34971 , n34946 , n34952 );
or ( n34972 , n34970 , n34971 );
buf ( n34973 , n34972 );
buf ( n34974 , n34973 );
buf ( n34975 , n34852 );
not ( n34976 , n34975 );
buf ( n34977 , n34864 );
not ( n34978 , n34977 );
or ( n34979 , n34976 , n34978 );
buf ( n34980 , n34864 );
buf ( n34981 , n34852 );
or ( n34982 , n34980 , n34981 );
buf ( n34983 , n34877 );
nand ( n34984 , n34982 , n34983 );
buf ( n34985 , n34984 );
buf ( n34986 , n34985 );
nand ( n34987 , n34979 , n34986 );
buf ( n34988 , n34987 );
not ( n34989 , n34988 );
xor ( n34990 , n34810 , n34823 );
and ( n34991 , n34990 , n34837 );
and ( n34992 , n34810 , n34823 );
or ( n34993 , n34991 , n34992 );
buf ( n34994 , n34993 );
buf ( n34995 , n34994 );
not ( n34996 , n34995 );
buf ( n34997 , n34996 );
nand ( n34998 , n34989 , n34997 );
not ( n34999 , n34998 );
not ( n35000 , n34904 );
not ( n35001 , n34892 );
or ( n35002 , n35000 , n35001 );
buf ( n35003 , n34904 );
buf ( n35004 , n34892 );
nor ( n35005 , n35003 , n35004 );
buf ( n35006 , n35005 );
or ( n35007 , n35006 , n34913 );
nand ( n35008 , n35002 , n35007 );
not ( n35009 , n35008 );
or ( n35010 , n34999 , n35009 );
buf ( n35011 , n34988 );
buf ( n35012 , n34994 );
nand ( n35013 , n35011 , n35012 );
buf ( n35014 , n35013 );
nand ( n35015 , n35010 , n35014 );
buf ( n35016 , n35015 );
xor ( n35017 , n33714 , n33728 );
xor ( n35018 , n35017 , n33743 );
buf ( n35019 , n35018 );
not ( n35020 , n35019 );
xor ( n35021 , n34500 , n34517 );
and ( n35022 , n35021 , n34531 );
and ( n35023 , n34500 , n34517 );
or ( n35024 , n35022 , n35023 );
buf ( n35025 , n35024 );
not ( n35026 , n35025 );
or ( n35027 , n35020 , n35026 );
or ( n35028 , n35019 , n35025 );
xor ( n35029 , n33881 , n33888 );
xor ( n35030 , n35029 , n33899 );
buf ( n35031 , n35030 );
nand ( n35032 , n35028 , n35031 );
nand ( n35033 , n35027 , n35032 );
buf ( n35034 , n35033 );
xor ( n35035 , n35016 , n35034 );
and ( n35036 , n33807 , n33906 );
not ( n35037 , n33807 );
and ( n35038 , n35037 , n33903 );
nor ( n35039 , n35036 , n35038 );
buf ( n35040 , n35039 );
buf ( n35041 , n33861 );
not ( n35042 , n35041 );
buf ( n35043 , n35042 );
buf ( n35044 , n35043 );
and ( n35045 , n35040 , n35044 );
not ( n35046 , n35040 );
buf ( n35047 , n33861 );
and ( n35048 , n35046 , n35047 );
nor ( n35049 , n35045 , n35048 );
buf ( n35050 , n35049 );
buf ( n35051 , n35050 );
xor ( n35052 , n35035 , n35051 );
buf ( n35053 , n35052 );
buf ( n35054 , n35053 );
xor ( n35055 , n34974 , n35054 );
xor ( n35056 , n34193 , n34202 );
xor ( n35057 , n35056 , n34206 );
buf ( n35058 , n35057 );
buf ( n35059 , n35058 );
buf ( n35060 , n34988 );
not ( n35061 , n35060 );
buf ( n35062 , n35008 );
not ( n35063 , n35062 );
buf ( n35064 , n35063 );
buf ( n35065 , n35064 );
not ( n35066 , n35065 );
or ( n35067 , n35061 , n35066 );
buf ( n35068 , n35064 );
buf ( n35069 , n34988 );
or ( n35070 , n35068 , n35069 );
nand ( n35071 , n35067 , n35070 );
buf ( n35072 , n35071 );
buf ( n35073 , n35072 );
buf ( n35074 , n34997 );
and ( n35075 , n35073 , n35074 );
not ( n35076 , n35073 );
buf ( n35077 , n34994 );
and ( n35078 , n35076 , n35077 );
nor ( n35079 , n35075 , n35078 );
buf ( n35080 , n35079 );
buf ( n35081 , n35080 );
not ( n35082 , n35081 );
buf ( n35083 , n35082 );
buf ( n35084 , n35083 );
or ( n35085 , n35059 , n35084 );
xor ( n35086 , n35025 , n35019 );
xor ( n35087 , n35086 , n35031 );
buf ( n35088 , n35087 );
nand ( n35089 , n35085 , n35088 );
buf ( n35090 , n35089 );
buf ( n35091 , n35090 );
buf ( n35092 , n35083 );
buf ( n35093 , n35058 );
nand ( n35094 , n35092 , n35093 );
buf ( n35095 , n35094 );
buf ( n35096 , n35095 );
nand ( n35097 , n35091 , n35096 );
buf ( n35098 , n35097 );
buf ( n35099 , n35098 );
xor ( n35100 , n35055 , n35099 );
buf ( n35101 , n35100 );
buf ( n35102 , n35101 );
and ( n35103 , n34968 , n35102 );
and ( n35104 , n34243 , n34967 );
or ( n35105 , n35103 , n35104 );
buf ( n35106 , n35105 );
not ( n35107 , n35106 );
xor ( n35108 , n34169 , n34174 );
and ( n35109 , n35108 , n34185 );
and ( n35110 , n34169 , n34174 );
or ( n35111 , n35109 , n35110 );
buf ( n35112 , n35111 );
buf ( n35113 , n24629 );
not ( n35114 , n35113 );
buf ( n35115 , n24638 );
not ( n35116 , n35115 );
or ( n35117 , n35114 , n35116 );
buf ( n35118 , n24629 );
buf ( n35119 , n24638 );
or ( n35120 , n35118 , n35119 );
nand ( n35121 , n35117 , n35120 );
buf ( n35122 , n35121 );
buf ( n35123 , n35122 );
buf ( n35124 , n24647 );
and ( n35125 , n35123 , n35124 );
not ( n35126 , n35123 );
buf ( n35127 , n24617 );
buf ( n35128 , n35127 );
and ( n35129 , n35126 , n35128 );
nor ( n35130 , n35125 , n35129 );
buf ( n35131 , n35130 );
buf ( n35132 , n35131 );
xor ( n35133 , n35112 , n35132 );
xor ( n35134 , n35016 , n35034 );
and ( n35135 , n35134 , n35051 );
and ( n35136 , n35016 , n35034 );
or ( n35137 , n35135 , n35136 );
buf ( n35138 , n35137 );
buf ( n35139 , n35138 );
xor ( n35140 , n35133 , n35139 );
buf ( n35141 , n35140 );
buf ( n35142 , n35141 );
xor ( n35143 , n34974 , n35054 );
and ( n35144 , n35143 , n35099 );
and ( n35145 , n34974 , n35054 );
or ( n35146 , n35144 , n35145 );
buf ( n35147 , n35146 );
buf ( n35148 , n35147 );
xor ( n35149 , n35142 , n35148 );
xor ( n35150 , n33676 , n33751 );
xor ( n35151 , n35150 , n33908 );
buf ( n35152 , n35151 );
buf ( n35153 , n33956 );
not ( n35154 , n35153 );
buf ( n35155 , n33915 );
not ( n35156 , n35155 );
buf ( n35157 , n35156 );
buf ( n35158 , n35157 );
not ( n35159 , n35158 );
or ( n35160 , n35154 , n35159 );
not ( n35161 , n33956 );
nand ( n35162 , n35161 , n33915 );
buf ( n35163 , n35162 );
nand ( n35164 , n35160 , n35163 );
buf ( n35165 , n35164 );
buf ( n35166 , n35165 );
buf ( n35167 , n33919 );
buf ( n35168 , n35167 );
buf ( n35169 , n35168 );
buf ( n35170 , n35169 );
xor ( n35171 , n35166 , n35170 );
buf ( n35172 , n35171 );
buf ( n35173 , n35172 );
xor ( n35174 , n35152 , n35173 );
not ( n35175 , n34210 );
not ( n35176 , n34186 );
or ( n35177 , n35175 , n35176 );
buf ( n35178 , n34186 );
buf ( n35179 , n34210 );
or ( n35180 , n35178 , n35179 );
buf ( n35181 , n34226 );
not ( n35182 , n35181 );
buf ( n35183 , n35182 );
buf ( n35184 , n35183 );
nand ( n35185 , n35180 , n35184 );
buf ( n35186 , n35185 );
nand ( n35187 , n35177 , n35186 );
buf ( n35188 , n35187 );
xor ( n35189 , n35174 , n35188 );
buf ( n35190 , n35189 );
buf ( n35191 , n35190 );
xor ( n35192 , n35149 , n35191 );
buf ( n35193 , n35192 );
not ( n35194 , n35193 );
nand ( n35195 , n35107 , n35194 );
xor ( n35196 , n35112 , n35132 );
and ( n35197 , n35196 , n35139 );
and ( n35198 , n35112 , n35132 );
or ( n35199 , n35197 , n35198 );
buf ( n35200 , n35199 );
buf ( n35201 , n35200 );
xor ( n35202 , n35152 , n35173 );
and ( n35203 , n35202 , n35188 );
and ( n35204 , n35152 , n35173 );
or ( n35205 , n35203 , n35204 );
buf ( n35206 , n35205 );
buf ( n35207 , n35206 );
xor ( n35208 , n35201 , n35207 );
xor ( n35209 , n24464 , n24606 );
xor ( n35210 , n35209 , n24654 );
buf ( n35211 , n35210 );
buf ( n35212 , n35211 );
buf ( n35213 , n24673 );
not ( n35214 , n35213 );
buf ( n35215 , n24810 );
not ( n35216 , n35215 );
and ( n35217 , n35214 , n35216 );
buf ( n35218 , n24673 );
buf ( n35219 , n24810 );
and ( n35220 , n35218 , n35219 );
nor ( n35221 , n35217 , n35220 );
buf ( n35222 , n35221 );
buf ( n35223 , n35222 );
buf ( n35224 , n24681 );
and ( n35225 , n35223 , n35224 );
not ( n35226 , n35223 );
buf ( n35227 , n24819 );
and ( n35228 , n35226 , n35227 );
nor ( n35229 , n35225 , n35228 );
buf ( n35230 , n35229 );
buf ( n35231 , n35230 );
xor ( n35232 , n35212 , n35231 );
xor ( n35233 , n33665 , n33912 );
xor ( n35234 , n35233 , n33959 );
buf ( n35235 , n35234 );
buf ( n35236 , n35235 );
xor ( n35237 , n35232 , n35236 );
buf ( n35238 , n35237 );
buf ( n35239 , n35238 );
xor ( n35240 , n35208 , n35239 );
buf ( n35241 , n35240 );
not ( n35242 , n35241 );
xor ( n35243 , n35142 , n35148 );
and ( n35244 , n35243 , n35191 );
and ( n35245 , n35142 , n35148 );
or ( n35246 , n35244 , n35245 );
buf ( n35247 , n35246 );
not ( n35248 , n35247 );
nand ( n35249 , n35242 , n35248 );
nand ( n35250 , n35195 , n35249 );
not ( n35251 , n35250 );
xor ( n35252 , n35201 , n35207 );
and ( n35253 , n35252 , n35239 );
and ( n35254 , n35201 , n35207 );
or ( n35255 , n35253 , n35254 );
buf ( n35256 , n35255 );
xor ( n35257 , n24461 , n24659 );
xor ( n35258 , n35257 , n24826 );
buf ( n35259 , n35258 );
buf ( n35260 , n35259 );
xor ( n35261 , n33657 , n33661 );
xor ( n35262 , n35261 , n33964 );
buf ( n35263 , n35262 );
buf ( n35264 , n35263 );
xor ( n35265 , n35260 , n35264 );
xor ( n35266 , n35212 , n35231 );
and ( n35267 , n35266 , n35236 );
and ( n35268 , n35212 , n35231 );
or ( n35269 , n35267 , n35268 );
buf ( n35270 , n35269 );
buf ( n35271 , n35270 );
xor ( n35272 , n35265 , n35271 );
buf ( n35273 , n35272 );
nor ( n35274 , n35256 , n35273 );
xor ( n35275 , n33653 , n33969 );
xor ( n35276 , n35275 , n33974 );
buf ( n35277 , n35276 );
xor ( n35278 , n35260 , n35264 );
and ( n35279 , n35278 , n35271 );
and ( n35280 , n35260 , n35264 );
or ( n35281 , n35279 , n35280 );
buf ( n35282 , n35281 );
nor ( n35283 , n35277 , n35282 );
nor ( n35284 , n35274 , n35283 );
nand ( n35285 , n35251 , n35284 );
not ( n35286 , n35285 );
xor ( n35287 , n34243 , n34967 );
xor ( n35288 , n35287 , n35102 );
buf ( n35289 , n35288 );
xor ( n35290 , n35080 , n35058 );
xnor ( n35291 , n35290 , n35087 );
buf ( n35292 , n35291 );
buf ( n35293 , n29667 );
not ( n35294 , n35293 );
buf ( n35295 , n25022 );
not ( n35296 , n35295 );
or ( n35297 , n35294 , n35296 );
buf ( n35298 , n25263 );
buf ( n35299 , n34463 );
nand ( n35300 , n35298 , n35299 );
buf ( n35301 , n35300 );
buf ( n35302 , n35301 );
nand ( n35303 , n35297 , n35302 );
buf ( n35304 , n35303 );
buf ( n35305 , n35304 );
buf ( n35306 , n29685 );
not ( n35307 , n35306 );
buf ( n35308 , n19580 );
not ( n35309 , n35308 );
or ( n35310 , n35307 , n35309 );
buf ( n35311 , n26538 );
buf ( n35312 , n34247 );
nand ( n35313 , n35311 , n35312 );
buf ( n35314 , n35313 );
buf ( n35315 , n35314 );
nand ( n35316 , n35310 , n35315 );
buf ( n35317 , n35316 );
buf ( n35318 , n35317 );
xor ( n35319 , n35305 , n35318 );
buf ( n35320 , n34280 );
not ( n35321 , n35320 );
buf ( n35322 , n34297 );
not ( n35323 , n35322 );
or ( n35324 , n35321 , n35323 );
buf ( n35325 , n34280 );
buf ( n35326 , n34297 );
or ( n35327 , n35325 , n35326 );
nand ( n35328 , n35324 , n35327 );
buf ( n35329 , n35328 );
buf ( n35330 , n35329 );
and ( n35331 , n35319 , n35330 );
and ( n35332 , n35305 , n35318 );
or ( n35333 , n35331 , n35332 );
buf ( n35334 , n35333 );
buf ( n35335 , n35334 );
xor ( n35336 , n34264 , n34301 );
xor ( n35337 , n35336 , n34355 );
buf ( n35338 , n35337 );
buf ( n35339 , n35338 );
xor ( n35340 , n35335 , n35339 );
xor ( n35341 , n29748 , n29765 );
and ( n35342 , n35341 , n29783 );
and ( n35343 , n29748 , n29765 );
or ( n35344 , n35342 , n35343 );
buf ( n35345 , n35344 );
buf ( n35346 , n35345 );
xor ( n35347 , n29803 , n29820 );
and ( n35348 , n35347 , n29838 );
and ( n35349 , n29803 , n29820 );
or ( n35350 , n35348 , n35349 );
buf ( n35351 , n35350 );
buf ( n35352 , n35351 );
xor ( n35353 , n35346 , n35352 );
xor ( n35354 , n29657 , n29674 );
and ( n35355 , n35354 , n29692 );
and ( n35356 , n29657 , n29674 );
or ( n35357 , n35355 , n35356 );
buf ( n35358 , n35357 );
buf ( n35359 , n35358 );
and ( n35360 , n35353 , n35359 );
and ( n35361 , n35346 , n35352 );
or ( n35362 , n35360 , n35361 );
buf ( n35363 , n35362 );
buf ( n35364 , n35363 );
and ( n35365 , n35340 , n35364 );
and ( n35366 , n35335 , n35339 );
or ( n35367 , n35365 , n35366 );
buf ( n35368 , n35367 );
buf ( n35369 , n35368 );
xor ( n35370 , n34360 , n34537 );
xor ( n35371 , n35370 , n34680 );
buf ( n35372 , n35371 );
buf ( n35373 , n35372 );
xor ( n35374 , n35369 , n35373 );
buf ( n35375 , n29724 );
buf ( n35376 , n29712 );
or ( n35377 , n35375 , n35376 );
buf ( n35378 , n29741 );
nand ( n35379 , n35377 , n35378 );
buf ( n35380 , n35379 );
buf ( n35381 , n35380 );
buf ( n35382 , n29724 );
buf ( n35383 , n29712 );
nand ( n35384 , n35382 , n35383 );
buf ( n35385 , n35384 );
buf ( n35386 , n35385 );
nand ( n35387 , n35381 , n35386 );
buf ( n35388 , n35387 );
buf ( n35389 , n35388 );
xor ( n35390 , n34693 , n34701 );
xor ( n35391 , n35390 , n34711 );
buf ( n35392 , n35391 );
xor ( n35393 , n35389 , n35392 );
xor ( n35394 , n34319 , n34336 );
xor ( n35395 , n35394 , n34350 );
buf ( n35396 , n35395 );
buf ( n35397 , n35396 );
and ( n35398 , n35393 , n35397 );
and ( n35399 , n35389 , n35392 );
or ( n35400 , n35398 , n35399 );
buf ( n35401 , n35400 );
buf ( n35402 , n35401 );
not ( n35403 , n35402 );
buf ( n35404 , n35403 );
buf ( n35405 , n35404 );
not ( n35406 , n35405 );
xor ( n35407 , n34715 , n34718 );
xor ( n35408 , n35407 , n34760 );
buf ( n35409 , n35408 );
buf ( n35410 , n35409 );
not ( n35411 , n35410 );
buf ( n35412 , n35411 );
buf ( n35413 , n35412 );
not ( n35414 , n35413 );
or ( n35415 , n35406 , n35414 );
xor ( n35416 , n34673 , n34564 );
xor ( n35417 , n35416 , n34612 );
buf ( n35418 , n35417 );
nand ( n35419 , n35415 , n35418 );
buf ( n35420 , n35419 );
buf ( n35421 , n35420 );
buf ( n35422 , n35409 );
buf ( n35423 , n35401 );
nand ( n35424 , n35422 , n35423 );
buf ( n35425 , n35424 );
buf ( n35426 , n35425 );
nand ( n35427 , n35421 , n35426 );
buf ( n35428 , n35427 );
buf ( n35429 , n35428 );
and ( n35430 , n35374 , n35429 );
and ( n35431 , n35369 , n35373 );
or ( n35432 , n35430 , n35431 );
buf ( n35433 , n35432 );
buf ( n35434 , n35433 );
xor ( n35435 , n35292 , n35434 );
xor ( n35436 , n34685 , n34924 );
xor ( n35437 , n35436 , n34962 );
buf ( n35438 , n35437 );
buf ( n35439 , n35438 );
and ( n35440 , n35435 , n35439 );
and ( n35441 , n35292 , n35434 );
or ( n35442 , n35440 , n35441 );
buf ( n35443 , n35442 );
nor ( n35444 , n35289 , n35443 );
xor ( n35445 , n35292 , n35434 );
xor ( n35446 , n35445 , n35439 );
buf ( n35447 , n35446 );
xor ( n35448 , n34794 , n34786 );
not ( n35449 , n34917 );
xor ( n35450 , n35448 , n35449 );
xor ( n35451 , n34727 , n34742 );
not ( n35452 , n34756 );
xor ( n35453 , n35451 , n35452 );
buf ( n35454 , n35453 );
xor ( n35455 , n35305 , n35318 );
xor ( n35456 , n35455 , n35330 );
buf ( n35457 , n35456 );
buf ( n35458 , n35457 );
xor ( n35459 , n35454 , n35458 );
xor ( n35460 , n29574 , n29594 );
and ( n35461 , n35460 , n29601 );
and ( n35462 , n29574 , n29594 );
or ( n35463 , n35461 , n35462 );
buf ( n35464 , n35463 );
buf ( n35465 , n35464 );
and ( n35466 , n35459 , n35465 );
and ( n35467 , n35454 , n35458 );
or ( n35468 , n35466 , n35467 );
buf ( n35469 , n35468 );
buf ( n35470 , n35469 );
xor ( n35471 , n35335 , n35339 );
xor ( n35472 , n35471 , n35364 );
buf ( n35473 , n35472 );
buf ( n35474 , n35473 );
xor ( n35475 , n35470 , n35474 );
xor ( n35476 , n35346 , n35352 );
xor ( n35477 , n35476 , n35359 );
buf ( n35478 , n35477 );
buf ( n35479 , n35478 );
xor ( n35480 , n29640 , n29695 );
and ( n35481 , n35480 , n29743 );
and ( n35482 , n29640 , n29695 );
or ( n35483 , n35481 , n35482 );
buf ( n35484 , n35483 );
buf ( n35485 , n35484 );
xor ( n35486 , n35479 , n35485 );
xor ( n35487 , n35389 , n35392 );
xor ( n35488 , n35487 , n35397 );
buf ( n35489 , n35488 );
buf ( n35490 , n35489 );
and ( n35491 , n35486 , n35490 );
and ( n35492 , n35479 , n35485 );
or ( n35493 , n35491 , n35492 );
buf ( n35494 , n35493 );
buf ( n35495 , n35494 );
and ( n35496 , n35475 , n35495 );
and ( n35497 , n35470 , n35474 );
or ( n35498 , n35496 , n35497 );
buf ( n35499 , n35498 );
xor ( n35500 , n35450 , n35499 );
xor ( n35501 , n35369 , n35373 );
xor ( n35502 , n35501 , n35429 );
buf ( n35503 , n35502 );
and ( n35504 , n35500 , n35503 );
and ( n35505 , n35450 , n35499 );
or ( n35506 , n35504 , n35505 );
nor ( n35507 , n35447 , n35506 );
nor ( n35508 , n35444 , n35507 );
xor ( n35509 , n35450 , n35499 );
xor ( n35510 , n35509 , n35503 );
xor ( n35511 , n35404 , n35409 );
xnor ( n35512 , n35511 , n35417 );
buf ( n35513 , n35512 );
xor ( n35514 , n29786 , n29841 );
and ( n35515 , n35514 , n29848 );
and ( n35516 , n29786 , n29841 );
or ( n35517 , n35515 , n35516 );
buf ( n35518 , n35517 );
xor ( n35519 , n35454 , n35458 );
xor ( n35520 , n35519 , n35465 );
buf ( n35521 , n35520 );
xor ( n35522 , n35518 , n35521 );
xor ( n35523 , n35479 , n35485 );
xor ( n35524 , n35523 , n35490 );
buf ( n35525 , n35524 );
and ( n35526 , n35522 , n35525 );
and ( n35527 , n35518 , n35521 );
or ( n35528 , n35526 , n35527 );
buf ( n35529 , n35528 );
xor ( n35530 , n35513 , n35529 );
xor ( n35531 , n35470 , n35474 );
xor ( n35532 , n35531 , n35495 );
buf ( n35533 , n35532 );
buf ( n35534 , n35533 );
and ( n35535 , n35530 , n35534 );
and ( n35536 , n35513 , n35529 );
or ( n35537 , n35535 , n35536 );
buf ( n35538 , n35537 );
nor ( n35539 , n35510 , n35538 );
xor ( n35540 , n35513 , n35529 );
xor ( n35541 , n35540 , n35534 );
buf ( n35542 , n35541 );
xor ( n35543 , n29604 , n29610 );
and ( n35544 , n35543 , n29617 );
and ( n35545 , n29604 , n29610 );
or ( n35546 , n35544 , n35545 );
buf ( n35547 , n35546 );
buf ( n35548 , n35547 );
not ( n35549 , n35548 );
not ( n35550 , n35549 );
xor ( n35551 , n29746 , n29851 );
and ( n35552 , n35551 , n29858 );
and ( n35553 , n29746 , n29851 );
or ( n35554 , n35552 , n35553 );
buf ( n35555 , n35554 );
not ( n35556 , n35555 );
not ( n35557 , n35556 );
or ( n35558 , n35550 , n35557 );
xor ( n35559 , n35518 , n35521 );
xor ( n35560 , n35559 , n35525 );
nand ( n35561 , n35558 , n35560 );
nand ( n35562 , n35555 , n35548 );
nand ( n35563 , n35561 , n35562 );
nor ( n35564 , n35542 , n35563 );
nor ( n35565 , n35539 , n35564 );
and ( n35566 , n35508 , n35565 );
nand ( n35567 , n35286 , n35566 );
xor ( n35568 , n28004 , n28281 );
xor ( n35569 , n35568 , n28563 );
buf ( n35570 , n35569 );
not ( n35571 , n35570 );
xor ( n35572 , n28705 , n28875 );
and ( n35573 , n35572 , n28897 );
and ( n35574 , n28705 , n28875 );
or ( n35575 , n35573 , n35574 );
buf ( n35576 , n35575 );
not ( n35577 , n35576 );
nand ( n35578 , n35571 , n35577 );
or ( n35579 , n28899 , n28988 );
nand ( n35580 , n35578 , n35579 );
not ( n35581 , n29872 );
not ( n35582 , n35581 );
xor ( n35583 , n35547 , n35555 );
xnor ( n35584 , n35583 , n35560 );
not ( n35585 , n35584 );
or ( n35586 , n35582 , n35585 );
xor ( n35587 , n29620 , n29861 );
xor ( n35588 , n35587 , n29868 );
buf ( n35589 , n35588 );
not ( n35590 , n35589 );
not ( n35591 , n28567 );
nand ( n35592 , n35590 , n35591 );
nand ( n35593 , n35586 , n35592 );
nor ( n35594 , n35580 , n35593 );
not ( n35595 , n35594 );
xor ( n35596 , n28955 , n28962 );
xnor ( n35597 , n35596 , n28950 );
buf ( n35598 , n35597 );
xor ( n35599 , n26882 , n26993 );
and ( n35600 , n35599 , n27048 );
and ( n35601 , n26882 , n26993 );
or ( n35602 , n35600 , n35601 );
buf ( n35603 , n35602 );
buf ( n35604 , n35603 );
xor ( n35605 , n35598 , n35604 );
xor ( n35606 , n26885 , n26933 );
and ( n35607 , n35606 , n26990 );
and ( n35608 , n26885 , n26933 );
or ( n35609 , n35607 , n35608 );
buf ( n35610 , n35609 );
buf ( n35611 , n35610 );
xor ( n35612 , n28911 , n28915 );
xor ( n35613 , n35612 , n28930 );
buf ( n35614 , n35613 );
xor ( n35615 , n35611 , n35614 );
not ( n35616 , n26554 );
not ( n35617 , n26440 );
or ( n35618 , n35616 , n35617 );
nand ( n35619 , n26486 , n26550 );
nand ( n35620 , n35618 , n35619 );
buf ( n35621 , n35620 );
xor ( n35622 , n35615 , n35621 );
buf ( n35623 , n35622 );
buf ( n35624 , n35623 );
and ( n35625 , n35605 , n35624 );
and ( n35626 , n35598 , n35604 );
or ( n35627 , n35625 , n35626 );
buf ( n35628 , n35627 );
xor ( n35629 , n28746 , n28750 );
xor ( n35630 , n35629 , n28766 );
buf ( n35631 , n35630 );
buf ( n35632 , n35631 );
xor ( n35633 , n35611 , n35614 );
and ( n35634 , n35633 , n35621 );
and ( n35635 , n35611 , n35614 );
or ( n35636 , n35634 , n35635 );
buf ( n35637 , n35636 );
buf ( n35638 , n35637 );
xor ( n35639 , n35632 , n35638 );
xor ( n35640 , n28934 , n28938 );
xor ( n35641 , n35640 , n28969 );
buf ( n35642 , n35641 );
buf ( n35643 , n35642 );
xor ( n35644 , n35639 , n35643 );
buf ( n35645 , n35644 );
nor ( n35646 , n35628 , n35645 );
xor ( n35647 , n28904 , n28974 );
xor ( n35648 , n35647 , n28984 );
buf ( n35649 , n35648 );
xor ( n35650 , n35632 , n35638 );
and ( n35651 , n35650 , n35643 );
and ( n35652 , n35632 , n35638 );
or ( n35653 , n35651 , n35652 );
buf ( n35654 , n35653 );
nor ( n35655 , n35649 , n35654 );
nor ( n35656 , n35646 , n35655 );
not ( n35657 , n35656 );
xor ( n35658 , n27058 , n27175 );
and ( n35659 , n35658 , n27180 );
and ( n35660 , n27058 , n27175 );
or ( n35661 , n35659 , n35660 );
buf ( n35662 , n35661 );
nand ( n35663 , n27053 , n35662 );
not ( n35664 , n35663 );
xor ( n35665 , n35598 , n35604 );
xor ( n35666 , n35665 , n35624 );
buf ( n35667 , n35666 );
xor ( n35668 , n26563 , n26875 );
and ( n35669 , n35668 , n27051 );
and ( n35670 , n26563 , n26875 );
or ( n35671 , n35669 , n35670 );
buf ( n35672 , n35671 );
nand ( n35673 , n35667 , n35672 );
not ( n35674 , n35673 );
or ( n35675 , n35664 , n35674 );
not ( n35676 , n35667 );
not ( n35677 , n35672 );
nand ( n35678 , n35676 , n35677 );
nand ( n35679 , n35675 , n35678 );
not ( n35680 , n35679 );
not ( n35681 , n35680 );
or ( n35682 , n35657 , n35681 );
not ( n35683 , n35655 );
nand ( n35684 , n35628 , n35645 );
not ( n35685 , n35684 );
and ( n35686 , n35683 , n35685 );
and ( n35687 , n35649 , n35654 );
nor ( n35688 , n35686 , n35687 );
nand ( n35689 , n35682 , n35688 );
not ( n35690 , n35689 );
or ( n35691 , n35595 , n35690 );
xor ( n35692 , n35547 , n35555 );
xor ( n35693 , n35692 , n35560 );
not ( n35694 , n35693 );
and ( n35695 , n35694 , n35581 );
nor ( n35696 , n35589 , n28567 );
nor ( n35697 , n35695 , n35696 );
not ( n35698 , n35697 );
not ( n35699 , n35578 );
and ( n35700 , n28899 , n28988 );
not ( n35701 , n35700 );
or ( n35702 , n35699 , n35701 );
not ( n35703 , n35571 );
not ( n35704 , n35577 );
nand ( n35705 , n35703 , n35704 );
nand ( n35706 , n35702 , n35705 );
not ( n35707 , n35706 );
or ( n35708 , n35698 , n35707 );
and ( n35709 , n35589 , n28567 );
nand ( n35710 , n35584 , n35581 );
and ( n35711 , n35709 , n35710 );
nand ( n35712 , n35693 , n29872 );
not ( n35713 , n35712 );
nor ( n35714 , n35711 , n35713 );
nand ( n35715 , n35708 , n35714 );
not ( n35716 , n35715 );
nand ( n35717 , n35691 , n35716 );
not ( n35718 , n35655 );
not ( n35719 , n35667 );
not ( n35720 , n35672 );
and ( n35721 , n35719 , n35720 );
nor ( n35722 , n27053 , n35662 );
nor ( n35723 , n35721 , n35722 );
not ( n35724 , n35646 );
and ( n35725 , n35718 , n35723 , n35724 );
not ( n35726 , n35580 );
xor ( n35727 , n26744 , n26812 );
xor ( n35728 , n35727 , n26865 );
buf ( n35729 , n35728 );
buf ( n35730 , n35729 );
xor ( n35731 , n27559 , n27563 );
and ( n35732 , n35731 , n27596 );
and ( n35733 , n27559 , n27563 );
or ( n35734 , n35732 , n35733 );
buf ( n35735 , n35734 );
buf ( n35736 , n35735 );
xor ( n35737 , n35730 , n35736 );
xor ( n35738 , n27062 , n27066 );
xor ( n35739 , n35738 , n27170 );
buf ( n35740 , n35739 );
buf ( n35741 , n35740 );
xor ( n35742 , n35737 , n35741 );
buf ( n35743 , n35742 );
not ( n35744 , n35743 );
xor ( n35745 , n27518 , n27545 );
and ( n35746 , n35745 , n27599 );
and ( n35747 , n27518 , n27545 );
or ( n35748 , n35746 , n35747 );
buf ( n35749 , n35748 );
not ( n35750 , n35749 );
and ( n35751 , n35744 , n35750 );
xor ( n35752 , n27578 , n27584 );
xor ( n35753 , n35752 , n27591 );
buf ( n35754 , n35753 );
buf ( n35755 , n35754 );
xor ( n35756 , n27258 , n27273 );
and ( n35757 , n35756 , n27317 );
and ( n35758 , n27258 , n27273 );
or ( n35759 , n35757 , n35758 );
buf ( n35760 , n35759 );
buf ( n35761 , n35760 );
xor ( n35762 , n35755 , n35761 );
xor ( n35763 , n27522 , n27526 );
xor ( n35764 , n35763 , n27540 );
buf ( n35765 , n35764 );
buf ( n35766 , n35765 );
and ( n35767 , n35762 , n35766 );
and ( n35768 , n35755 , n35761 );
or ( n35769 , n35767 , n35768 );
buf ( n35770 , n35769 );
not ( n35771 , n35770 );
not ( n35772 , n35771 );
not ( n35773 , n27601 );
not ( n35774 , n35773 );
or ( n35775 , n35772 , n35774 );
xor ( n35776 , n35755 , n35761 );
xor ( n35777 , n35776 , n35766 );
buf ( n35778 , n35777 );
xor ( n35779 , n27252 , n27320 );
and ( n35780 , n35779 , n27327 );
and ( n35781 , n27252 , n27320 );
or ( n35782 , n35780 , n35781 );
buf ( n35783 , n35782 );
or ( n35784 , n35778 , n35783 );
nand ( n35785 , n35775 , n35784 );
nor ( n35786 , n35751 , n35785 );
not ( n35787 , n27329 );
xor ( n35788 , n23084 , n23223 );
and ( n35789 , n35788 , n23336 );
and ( n35790 , n23084 , n23223 );
or ( n35791 , n35789 , n35790 );
buf ( n35792 , n35791 );
not ( n35793 , n35792 );
nand ( n35794 , n35787 , n35793 );
buf ( n35795 , n35794 );
buf ( n35796 , n20869 );
buf ( n35797 , n863 );
and ( n35798 , n35796 , n35797 );
buf ( n35799 , n35798 );
buf ( n35800 , n35799 );
buf ( n35801 , n27497 );
not ( n35802 , n35801 );
buf ( n35803 , n21297 );
not ( n35804 , n35803 );
or ( n35805 , n35802 , n35804 );
buf ( n35806 , n859 );
buf ( n35807 , n894 );
xor ( n35808 , n35806 , n35807 );
buf ( n35809 , n35808 );
buf ( n35810 , n35809 );
buf ( n35811 , n895 );
nand ( n35812 , n35810 , n35811 );
buf ( n35813 , n35812 );
buf ( n35814 , n35813 );
nand ( n35815 , n35805 , n35814 );
buf ( n35816 , n35815 );
buf ( n35817 , n35816 );
xor ( n35818 , n35800 , n35817 );
buf ( n35819 , n862 );
buf ( n35820 , n892 );
xor ( n35821 , n35819 , n35820 );
buf ( n35822 , n35821 );
buf ( n35823 , n35822 );
not ( n35824 , n35823 );
buf ( n35825 , n23175 );
not ( n35826 , n35825 );
or ( n35827 , n35824 , n35826 );
buf ( n35828 , n23181 );
buf ( n35829 , n861 );
buf ( n35830 , n892 );
xor ( n35831 , n35829 , n35830 );
buf ( n35832 , n35831 );
buf ( n35833 , n35832 );
nand ( n35834 , n35828 , n35833 );
buf ( n35835 , n35834 );
buf ( n35836 , n35835 );
nand ( n35837 , n35827 , n35836 );
buf ( n35838 , n35837 );
buf ( n35839 , n35838 );
xor ( n35840 , n35818 , n35839 );
buf ( n35841 , n35840 );
and ( n35842 , n27484 , n27505 );
buf ( n35843 , n35842 );
nand ( n35844 , n35841 , n35843 );
not ( n35845 , n35844 );
not ( n35846 , n35845 );
buf ( n35847 , n35832 );
not ( n35848 , n35847 );
buf ( n35849 , n23175 );
not ( n35850 , n35849 );
or ( n35851 , n35848 , n35850 );
buf ( n35852 , n23181 );
buf ( n35853 , n860 );
buf ( n35854 , n892 );
xor ( n35855 , n35853 , n35854 );
buf ( n35856 , n35855 );
buf ( n35857 , n35856 );
nand ( n35858 , n35852 , n35857 );
buf ( n35859 , n35858 );
buf ( n35860 , n35859 );
nand ( n35861 , n35851 , n35860 );
buf ( n35862 , n35861 );
buf ( n35863 , n35862 );
buf ( n35864 , n863 );
buf ( n35865 , n890 );
xor ( n35866 , n35864 , n35865 );
buf ( n35867 , n35866 );
buf ( n35868 , n35867 );
not ( n35869 , n35868 );
buf ( n35870 , n21441 );
not ( n35871 , n35870 );
or ( n35872 , n35869 , n35871 );
buf ( n35873 , n20869 );
buf ( n35874 , n862 );
buf ( n35875 , n890 );
xor ( n35876 , n35874 , n35875 );
buf ( n35877 , n35876 );
buf ( n35878 , n35877 );
nand ( n35879 , n35873 , n35878 );
buf ( n35880 , n35879 );
buf ( n35881 , n35880 );
nand ( n35882 , n35872 , n35881 );
buf ( n35883 , n35882 );
buf ( n35884 , n35883 );
xor ( n35885 , n35863 , n35884 );
not ( n35886 , n35809 );
not ( n35887 , n21297 );
or ( n35888 , n35886 , n35887 );
buf ( n35889 , n858 );
buf ( n35890 , n894 );
xor ( n35891 , n35889 , n35890 );
buf ( n35892 , n35891 );
buf ( n35893 , n35892 );
buf ( n35894 , n895 );
nand ( n35895 , n35893 , n35894 );
buf ( n35896 , n35895 );
nand ( n35897 , n35888 , n35896 );
buf ( n35898 , n863 );
buf ( n35899 , n891 );
or ( n35900 , n35898 , n35899 );
buf ( n35901 , n892 );
nand ( n35902 , n35900 , n35901 );
buf ( n35903 , n35902 );
buf ( n35904 , n863 );
buf ( n35905 , n891 );
nand ( n35906 , n35904 , n35905 );
buf ( n35907 , n35906 );
nand ( n35908 , n35903 , n35907 , n890 );
not ( n35909 , n35908 );
and ( n35910 , n35897 , n35909 );
not ( n35911 , n35897 );
and ( n35912 , n35911 , n35908 );
nor ( n35913 , n35910 , n35912 );
buf ( n35914 , n35913 );
xor ( n35915 , n35885 , n35914 );
buf ( n35916 , n35915 );
not ( n35917 , n35916 );
xor ( n35918 , n35800 , n35817 );
and ( n35919 , n35918 , n35839 );
and ( n35920 , n35800 , n35817 );
or ( n35921 , n35919 , n35920 );
buf ( n35922 , n35921 );
not ( n35923 , n35922 );
nand ( n35924 , n35917 , n35923 );
not ( n35925 , n35924 );
or ( n35926 , n35846 , n35925 );
nand ( n35927 , n35916 , n35922 );
nand ( n35928 , n35926 , n35927 );
not ( n35929 , n35916 );
nand ( n35930 , n35929 , n35923 );
buf ( n35931 , n863 );
buf ( n35932 , n892 );
xor ( n35933 , n35931 , n35932 );
buf ( n35934 , n35933 );
buf ( n35935 , n35934 );
not ( n35936 , n35935 );
buf ( n35937 , n20599 );
not ( n35938 , n35937 );
or ( n35939 , n35936 , n35938 );
buf ( n35940 , n23181 );
buf ( n35941 , n35822 );
nand ( n35942 , n35940 , n35941 );
buf ( n35943 , n35942 );
buf ( n35944 , n35943 );
nand ( n35945 , n35939 , n35944 );
buf ( n35946 , n35945 );
nand ( n35947 , n27507 , n35946 );
buf ( n35948 , n28998 );
not ( n35949 , n35948 );
buf ( n35950 , n22776 );
not ( n35951 , n35950 );
or ( n35952 , n35949 , n35951 );
buf ( n35953 , n27488 );
buf ( n35954 , n895 );
nand ( n35955 , n35953 , n35954 );
buf ( n35956 , n35955 );
buf ( n35957 , n35956 );
nand ( n35958 , n35952 , n35957 );
buf ( n35959 , n35958 );
buf ( n35960 , n23181 );
buf ( n35961 , n863 );
and ( n35962 , n35960 , n35961 );
buf ( n35963 , n35962 );
nor ( n35964 , n35959 , n35963 );
buf ( n35965 , n863 );
buf ( n35966 , n895 );
nand ( n35967 , n35965 , n35966 );
buf ( n35968 , n35967 );
buf ( n35969 , n35968 );
buf ( n35970 , n894 );
and ( n35971 , n35969 , n35970 );
buf ( n35972 , n35971 );
nand ( n35973 , n35972 , n29005 );
nor ( n35974 , n35964 , n35973 );
and ( n35975 , n35959 , n35963 );
or ( n35976 , n35974 , n35975 );
or ( n35977 , n35946 , n27507 );
nand ( n35978 , n35976 , n35977 );
nand ( n35979 , n35947 , n35978 );
or ( n35980 , n35841 , n35843 );
nand ( n35981 , n35930 , n35979 , n35980 );
not ( n35982 , n35981 );
or ( n35983 , n35928 , n35982 );
buf ( n35984 , n863 );
buf ( n35985 , n20363 );
nand ( n35986 , n35984 , n35985 );
buf ( n35987 , n35986 );
buf ( n35988 , n35987 );
not ( n35989 , n35988 );
buf ( n35990 , n35989 );
buf ( n35991 , n35990 );
not ( n35992 , n35991 );
buf ( n35993 , n35892 );
not ( n35994 , n35993 );
buf ( n35995 , n23288 );
not ( n35996 , n35995 );
or ( n35997 , n35994 , n35996 );
buf ( n35998 , n27424 );
buf ( n35999 , n895 );
nand ( n36000 , n35998 , n35999 );
buf ( n36001 , n36000 );
buf ( n36002 , n36001 );
nand ( n36003 , n35997 , n36002 );
buf ( n36004 , n36003 );
buf ( n36005 , n36004 );
not ( n36006 , n36005 );
or ( n36007 , n35992 , n36006 );
buf ( n36008 , n36004 );
not ( n36009 , n36008 );
buf ( n36010 , n36009 );
buf ( n36011 , n36010 );
not ( n36012 , n36011 );
buf ( n36013 , n35987 );
not ( n36014 , n36013 );
or ( n36015 , n36012 , n36014 );
buf ( n36016 , n35856 );
not ( n36017 , n36016 );
buf ( n36018 , n23175 );
not ( n36019 , n36018 );
or ( n36020 , n36017 , n36019 );
buf ( n36021 , n23181 );
buf ( n36022 , n27334 );
nand ( n36023 , n36021 , n36022 );
buf ( n36024 , n36023 );
buf ( n36025 , n36024 );
nand ( n36026 , n36020 , n36025 );
buf ( n36027 , n36026 );
buf ( n36028 , n36027 );
nand ( n36029 , n36015 , n36028 );
buf ( n36030 , n36029 );
buf ( n36031 , n36030 );
nand ( n36032 , n36007 , n36031 );
buf ( n36033 , n36032 );
buf ( n36034 , n36033 );
not ( n36035 , n36034 );
buf ( n36036 , n27436 );
buf ( n36037 , n27452 );
and ( n36038 , n36036 , n36037 );
not ( n36039 , n36036 );
buf ( n36040 , n27455 );
and ( n36041 , n36039 , n36040 );
nor ( n36042 , n36038 , n36041 );
buf ( n36043 , n36042 );
buf ( n36044 , n36043 );
not ( n36045 , n36044 );
and ( n36046 , n36035 , n36045 );
buf ( n36047 , n36033 );
buf ( n36048 , n36043 );
and ( n36049 , n36047 , n36048 );
nor ( n36050 , n36046 , n36049 );
buf ( n36051 , n36050 );
xor ( n36052 , n27346 , n27362 );
xor ( n36053 , n36052 , n27376 );
xnor ( n36054 , n36051 , n36053 );
not ( n36055 , n36054 );
buf ( n36056 , n35877 );
not ( n36057 , n36056 );
buf ( n36058 , n21441 );
not ( n36059 , n36058 );
or ( n36060 , n36057 , n36059 );
buf ( n36061 , n20869 );
buf ( n36062 , n27350 );
nand ( n36063 , n36061 , n36062 );
buf ( n36064 , n36063 );
buf ( n36065 , n36064 );
nand ( n36066 , n36060 , n36065 );
buf ( n36067 , n36066 );
buf ( n36068 , n36067 );
not ( n36069 , n36068 );
buf ( n36070 , n36069 );
nand ( n36071 , n35897 , n35909 );
nand ( n36072 , n36070 , n36071 );
buf ( n36073 , n36072 );
not ( n36074 , n36073 );
xor ( n36075 , n35990 , n36010 );
xor ( n36076 , n36075 , n36027 );
buf ( n36077 , n36076 );
not ( n36078 , n36077 );
buf ( n36079 , n36078 );
buf ( n36080 , n36079 );
not ( n36081 , n36080 );
or ( n36082 , n36074 , n36081 );
not ( n36083 , n36071 );
nand ( n36084 , n36083 , n36067 );
buf ( n36085 , n36084 );
nand ( n36086 , n36082 , n36085 );
buf ( n36087 , n36086 );
not ( n36088 , n36087 );
nand ( n36089 , n36055 , n36088 );
and ( n36090 , n36071 , n36070 );
not ( n36091 , n36071 );
and ( n36092 , n36091 , n36067 );
nor ( n36093 , n36090 , n36092 );
buf ( n36094 , n36093 );
not ( n36095 , n36094 );
buf ( n36096 , n36095 );
buf ( n36097 , n36096 );
not ( n36098 , n36097 );
buf ( n36099 , n36079 );
not ( n36100 , n36099 );
or ( n36101 , n36098 , n36100 );
buf ( n36102 , n36076 );
buf ( n36103 , n36093 );
nand ( n36104 , n36102 , n36103 );
buf ( n36105 , n36104 );
buf ( n36106 , n36105 );
nand ( n36107 , n36101 , n36106 );
buf ( n36108 , n36107 );
not ( n36109 , n36108 );
xor ( n36110 , n35863 , n35884 );
and ( n36111 , n36110 , n35914 );
and ( n36112 , n35863 , n35884 );
or ( n36113 , n36111 , n36112 );
buf ( n36114 , n36113 );
not ( n36115 , n36114 );
nand ( n36116 , n36109 , n36115 );
nand ( n36117 , n35983 , n36089 , n36116 );
nand ( n36118 , n36108 , n36114 );
not ( n36119 , n36118 );
or ( n36120 , n36054 , n36087 );
and ( n36121 , n36119 , n36120 );
nand ( n36122 , n36054 , n36087 );
not ( n36123 , n36122 );
nor ( n36124 , n36121 , n36123 );
nand ( n36125 , n36117 , n36124 );
buf ( n36126 , n27407 );
buf ( n36127 , n27461 );
or ( n36128 , n36126 , n36127 );
buf ( n36129 , n27419 );
nand ( n36130 , n36128 , n36129 );
buf ( n36131 , n36130 );
buf ( n36132 , n36131 );
buf ( n36133 , n27407 );
buf ( n36134 , n27461 );
nand ( n36135 , n36133 , n36134 );
buf ( n36136 , n36135 );
buf ( n36137 , n36136 );
nand ( n36138 , n36132 , n36137 );
buf ( n36139 , n36138 );
buf ( n36140 , n36139 );
xor ( n36141 , n23299 , n23312 );
xor ( n36142 , n36141 , n23328 );
buf ( n36143 , n36142 );
buf ( n36144 , n36143 );
xor ( n36145 , n36140 , n36144 );
xor ( n36146 , n23102 , n23165 );
xor ( n36147 , n36146 , n23218 );
buf ( n36148 , n36147 );
buf ( n36149 , n36148 );
and ( n36150 , n36145 , n36149 );
and ( n36151 , n36140 , n36144 );
or ( n36152 , n36150 , n36151 );
buf ( n36153 , n36152 );
not ( n36154 , n36153 );
not ( n36155 , n23338 );
nand ( n36156 , n36154 , n36155 );
xor ( n36157 , n36140 , n36144 );
xor ( n36158 , n36157 , n36149 );
buf ( n36159 , n36158 );
not ( n36160 , n27394 );
not ( n36161 , n27465 );
or ( n36162 , n36160 , n36161 );
nand ( n36163 , n36162 , n27379 );
or ( n36164 , n27465 , n27394 );
nand ( n36165 , n36163 , n36164 );
nor ( n36166 , n36159 , n36165 );
buf ( n36167 , n36033 );
not ( n36168 , n36167 );
buf ( n36169 , n36043 );
nand ( n36170 , n36168 , n36169 );
buf ( n36171 , n36170 );
buf ( n36172 , n36171 );
not ( n36173 , n36172 );
buf ( n36174 , n36053 );
not ( n36175 , n36174 );
or ( n36176 , n36173 , n36175 );
buf ( n36177 , n36043 );
not ( n36178 , n36177 );
buf ( n36179 , n36033 );
nand ( n36180 , n36178 , n36179 );
buf ( n36181 , n36180 );
buf ( n36182 , n36181 );
nand ( n36183 , n36176 , n36182 );
buf ( n36184 , n36183 );
nor ( n36185 , n27467 , n36184 );
nor ( n36186 , n36166 , n36185 );
and ( n36187 , n35795 , n36125 , n36156 , n36186 );
xor ( n36188 , n35730 , n35736 );
and ( n36189 , n36188 , n35741 );
and ( n36190 , n35730 , n35736 );
or ( n36191 , n36189 , n36190 );
buf ( n36192 , n36191 );
or ( n36193 , n27182 , n36192 );
nand ( n36194 , n35786 , n36187 , n36193 );
nor ( n36195 , n27182 , n36192 );
nor ( n36196 , n35743 , n35749 );
nor ( n36197 , n36195 , n36196 );
nand ( n36198 , n35778 , n35783 );
not ( n36199 , n36198 );
not ( n36200 , n36199 );
nand ( n36201 , n35773 , n35771 );
not ( n36202 , n36201 );
or ( n36203 , n36200 , n36202 );
nand ( n36204 , n27601 , n35770 );
nand ( n36205 , n36203 , n36204 );
and ( n36206 , n36197 , n36205 );
nand ( n36207 , n35743 , n35749 );
or ( n36208 , n36195 , n36207 );
nand ( n36209 , n27182 , n36192 );
nand ( n36210 , n36208 , n36209 );
nor ( n36211 , n36206 , n36210 );
nand ( n36212 , n27467 , n36184 );
nor ( n36213 , n36159 , n36165 );
or ( n36214 , n36212 , n36213 );
nand ( n36215 , n36159 , n36165 );
nand ( n36216 , n36214 , n36215 );
not ( n36217 , n36216 );
not ( n36218 , n36153 );
nand ( n36219 , n36218 , n36155 );
and ( n36220 , n35794 , n36219 );
not ( n36221 , n36220 );
or ( n36222 , n36217 , n36221 );
nand ( n36223 , n23338 , n36153 );
not ( n36224 , n36223 );
not ( n36225 , n36224 );
not ( n36226 , n35794 );
or ( n36227 , n36225 , n36226 );
not ( n36228 , n35787 );
nand ( n36229 , n36228 , n35792 );
nand ( n36230 , n36227 , n36229 );
not ( n36231 , n36230 );
nand ( n36232 , n36222 , n36231 );
not ( n36233 , n35785 );
nand ( n36234 , n36232 , n36197 , n36233 );
nand ( n36235 , n36194 , n36211 , n36234 );
and ( n36236 , n35725 , n35726 , n36235 , n35697 );
nor ( n36237 , n35717 , n36236 );
or ( n36238 , n35567 , n36237 );
nand ( n36239 , n35542 , n35563 );
nand ( n36240 , n35510 , n35538 );
nand ( n36241 , n36239 , n36240 );
not ( n36242 , n35506 );
not ( n36243 , n35447 );
nand ( n36244 , n36242 , n36243 );
nand ( n36245 , n36241 , n36244 );
not ( n36246 , n36245 );
not ( n36247 , n36246 );
nor ( n36248 , n35444 , n35539 );
not ( n36249 , n36248 );
or ( n36250 , n36247 , n36249 );
nand ( n36251 , n35447 , n35506 );
not ( n36252 , n36251 );
not ( n36253 , n36252 );
not ( n36254 , n35289 );
not ( n36255 , n35443 );
nand ( n36256 , n36254 , n36255 );
not ( n36257 , n36256 );
or ( n36258 , n36253 , n36257 );
nand ( n36259 , n35289 , n35443 );
nand ( n36260 , n36258 , n36259 );
not ( n36261 , n36260 );
nand ( n36262 , n36250 , n36261 );
and ( n36263 , n35286 , n36262 );
not ( n36264 , n35284 );
not ( n36265 , n35106 );
nor ( n36266 , n36265 , n35194 );
not ( n36267 , n36266 );
not ( n36268 , n35249 );
or ( n36269 , n36267 , n36268 );
not ( n36270 , n35248 );
buf ( n36271 , n35241 );
nand ( n36272 , n36270 , n36271 );
nand ( n36273 , n36269 , n36272 );
not ( n36274 , n36273 );
or ( n36275 , n36264 , n36274 );
and ( n36276 , n35273 , n35256 );
not ( n36277 , n35277 );
not ( n36278 , n35282 );
nand ( n36279 , n36277 , n36278 );
and ( n36280 , n36276 , n36279 );
and ( n36281 , n35277 , n35282 );
nor ( n36282 , n36280 , n36281 );
nand ( n36283 , n36275 , n36282 );
nor ( n36284 , n36263 , n36283 );
nand ( n36285 , n36238 , n36284 );
buf ( n36286 , n36285 );
buf ( n36287 , n36286 );
and ( n36288 , n34095 , n36287 );
not ( n36289 , n32838 );
not ( n36290 , n36289 );
not ( n36291 , n32773 );
not ( n36292 , n36291 );
nand ( n36293 , n32505 , n20095 );
nor ( n36294 , n32513 , n26378 );
or ( n36295 , n36293 , n36294 );
nand ( n36296 , n32513 , n26378 );
nand ( n36297 , n36295 , n36296 );
not ( n36298 , n36297 );
or ( n36299 , n36292 , n36298 );
and ( n36300 , n32522 , n32688 );
and ( n36301 , n32772 , n36300 );
not ( n36302 , n32764 );
nor ( n36303 , n36302 , n32771 );
nor ( n36304 , n36301 , n36303 );
nand ( n36305 , n36299 , n36304 );
not ( n36306 , n36305 );
not ( n36307 , n36306 );
not ( n36308 , n36307 );
or ( n36309 , n36290 , n36308 );
nand ( n36310 , n32831 , n32836 );
not ( n36311 , n36310 );
not ( n36312 , n36311 );
not ( n36313 , n32828 );
or ( n36314 , n36312 , n36313 );
nand ( n36315 , n32810 , n32827 );
nand ( n36316 , n36314 , n36315 );
not ( n36317 , n36316 );
nand ( n36318 , n36309 , n36317 );
nor ( n36319 , n36288 , n36318 );
nand ( n36320 , n34071 , n36319 );
not ( n36321 , n29570 );
xor ( n36322 , n32814 , n32818 );
and ( n36323 , n36322 , n32825 );
and ( n36324 , n32814 , n32818 );
or ( n36325 , n36323 , n36324 );
buf ( n36326 , n36325 );
not ( n36327 , n36326 );
nand ( n36328 , n36321 , n36327 );
not ( n36329 , n29570 );
nor ( n36330 , n36329 , n36327 );
not ( n36331 , n36330 );
nand ( n36332 , n36328 , n36331 );
not ( n36333 , n36332 );
and ( n36334 , n36320 , n36333 );
not ( n36335 , n36320 );
and ( n36336 , n36335 , n36332 );
nor ( n36337 , n36334 , n36336 );
not ( n36338 , n34093 );
not ( n36339 , n32775 );
and ( n36340 , n36338 , n36339 );
buf ( n36341 , n36286 );
and ( n36342 , n36340 , n36341 );
nor ( n36343 , n36342 , n36307 );
not ( n36344 , n32775 );
not ( n36345 , n33571 );
nand ( n36346 , n34048 , n34062 , n34067 );
nand ( n36347 , n36345 , n36346 );
nand ( n36348 , n36344 , n36347 );
nand ( n36349 , n36343 , n36348 );
not ( n36350 , n32837 );
or ( n36351 , n36311 , n36350 );
not ( n36352 , n36351 );
and ( n36353 , n36349 , n36352 );
not ( n36354 , n36349 );
and ( n36355 , n36354 , n36351 );
nor ( n36356 , n36353 , n36355 );
not ( n36357 , n34076 );
nor ( n36358 , n36357 , n34058 );
not ( n36359 , n36358 );
not ( n36360 , n36286 );
or ( n36361 , n36359 , n36360 );
buf ( n36362 , n34083 );
not ( n36363 , n36362 );
not ( n36364 , n33987 );
not ( n36365 , n36364 );
nand ( n36366 , n33980 , n36365 );
not ( n36367 , n36366 );
or ( n36368 , n36363 , n36367 );
buf ( n36369 , n33986 );
nand ( n36370 , n36368 , n36369 );
not ( n36371 , n36370 );
nand ( n36372 , n36361 , n36371 );
buf ( n36373 , n34001 );
nand ( n36374 , n34080 , n36373 );
nand ( n36375 , n36372 , n36374 );
nor ( n36376 , n32775 , n36350 );
not ( n36377 , n36376 );
not ( n36378 , n36347 );
or ( n36379 , n36377 , n36378 );
not ( n36380 , n36286 );
buf ( n36381 , n34092 );
nand ( n36382 , n36381 , n36376 );
nor ( n36383 , n36380 , n36382 );
not ( n36384 , n32837 );
not ( n36385 , n36305 );
or ( n36386 , n36384 , n36385 );
nand ( n36387 , n36386 , n36310 );
nor ( n36388 , n36383 , n36387 );
nand ( n36389 , n36379 , n36388 );
xor ( n36390 , n29190 , n29380 );
and ( n36391 , n36390 , n29568 );
and ( n36392 , n29190 , n29380 );
or ( n36393 , n36391 , n36392 );
buf ( n36394 , n36393 );
xor ( n36395 , n29073 , n29130 );
and ( n36396 , n36395 , n29187 );
and ( n36397 , n29073 , n29130 );
or ( n36398 , n36396 , n36397 );
buf ( n36399 , n36398 );
buf ( n36400 , n36399 );
xor ( n36401 , n29193 , n29210 );
and ( n36402 , n36401 , n29231 );
and ( n36403 , n29193 , n29210 );
or ( n36404 , n36402 , n36403 );
buf ( n36405 , n36404 );
buf ( n36406 , n36405 );
buf ( n36407 , n29147 );
not ( n36408 , n36407 );
buf ( n36409 , n29139 );
not ( n36410 , n36409 );
or ( n36411 , n36408 , n36410 );
buf ( n36412 , n18944 );
xor ( n36413 , n866 , n836 );
buf ( n36414 , n36413 );
nand ( n36415 , n36412 , n36414 );
buf ( n36416 , n36415 );
buf ( n36417 , n36416 );
nand ( n36418 , n36411 , n36417 );
buf ( n36419 , n36418 );
buf ( n36420 , n36419 );
not ( n36421 , n19229 );
buf ( n36422 , n19235 );
not ( n36423 , n36422 );
buf ( n36424 , n36423 );
not ( n36425 , n36424 );
or ( n36426 , n36421 , n36425 );
nand ( n36427 , n36426 , n872 );
buf ( n36428 , n36427 );
xor ( n36429 , n36420 , n36428 );
buf ( n36430 , n29221 );
not ( n36431 , n36430 );
buf ( n36432 , n19125 );
not ( n36433 , n36432 );
or ( n36434 , n36431 , n36433 );
buf ( n36435 , n19134 );
buf ( n36436 , n832 );
buf ( n36437 , n870 );
xor ( n36438 , n36436 , n36437 );
buf ( n36439 , n36438 );
buf ( n36440 , n36439 );
nand ( n36441 , n36435 , n36440 );
buf ( n36442 , n36441 );
buf ( n36443 , n36442 );
nand ( n36444 , n36434 , n36443 );
buf ( n36445 , n36444 );
buf ( n36446 , n36445 );
xor ( n36447 , n36429 , n36446 );
buf ( n36448 , n36447 );
buf ( n36449 , n36448 );
xor ( n36450 , n36406 , n36449 );
buf ( n36451 , n29227 );
buf ( n36452 , n29183 );
buf ( n36453 , n29153 );
or ( n36454 , n36452 , n36453 );
buf ( n36455 , n29165 );
nand ( n36456 , n36454 , n36455 );
buf ( n36457 , n36456 );
buf ( n36458 , n36457 );
buf ( n36459 , n29183 );
buf ( n36460 , n29153 );
nand ( n36461 , n36459 , n36460 );
buf ( n36462 , n36461 );
buf ( n36463 , n36462 );
nand ( n36464 , n36458 , n36463 );
buf ( n36465 , n36464 );
buf ( n36466 , n36465 );
xor ( n36467 , n36451 , n36466 );
and ( n36468 , n29058 , n29059 );
buf ( n36469 , n36468 );
buf ( n36470 , n36469 );
buf ( n36471 , n29177 );
not ( n36472 , n36471 );
buf ( n36473 , n19330 );
not ( n36474 , n36473 );
or ( n36475 , n36472 , n36474 );
buf ( n36476 , n19030 );
buf ( n36477 , n864 );
buf ( n36478 , n838 );
xor ( n36479 , n36477 , n36478 );
buf ( n36480 , n36479 );
buf ( n36481 , n36480 );
nand ( n36482 , n36476 , n36481 );
buf ( n36483 , n36482 );
buf ( n36484 , n36483 );
nand ( n36485 , n36475 , n36484 );
buf ( n36486 , n36485 );
buf ( n36487 , n36486 );
xor ( n36488 , n36470 , n36487 );
buf ( n36489 , n29203 );
not ( n36490 , n36489 );
buf ( n36491 , n18887 );
not ( n36492 , n36491 );
or ( n36493 , n36490 , n36492 );
buf ( n36494 , n18898 );
buf ( n36495 , n834 );
buf ( n36496 , n868 );
xor ( n36497 , n36495 , n36496 );
buf ( n36498 , n36497 );
buf ( n36499 , n36498 );
nand ( n36500 , n36494 , n36499 );
buf ( n36501 , n36500 );
buf ( n36502 , n36501 );
nand ( n36503 , n36493 , n36502 );
buf ( n36504 , n36503 );
buf ( n36505 , n36504 );
xor ( n36506 , n36488 , n36505 );
buf ( n36507 , n36506 );
buf ( n36508 , n36507 );
xor ( n36509 , n36467 , n36508 );
buf ( n36510 , n36509 );
buf ( n36511 , n36510 );
xor ( n36512 , n36450 , n36511 );
buf ( n36513 , n36512 );
buf ( n36514 , n36513 );
xor ( n36515 , n36400 , n36514 );
xor ( n36516 , n29234 , n29319 );
and ( n36517 , n36516 , n29377 );
and ( n36518 , n29234 , n29319 );
or ( n36519 , n36517 , n36518 );
buf ( n36520 , n36519 );
buf ( n36521 , n36520 );
xor ( n36522 , n36515 , n36521 );
buf ( n36523 , n36522 );
or ( n36524 , n36394 , n36523 );
nand ( n36525 , n36328 , n36524 );
nor ( n36526 , n32838 , n36525 );
and ( n36527 , n32774 , n36526 );
buf ( n36528 , n36527 );
not ( n36529 , n36528 );
not ( n36530 , n34069 );
or ( n36531 , n36529 , n36530 );
nand ( n36532 , n36381 , n36527 );
nor ( n36533 , n36532 , n36380 );
not ( n36534 , n36526 );
not ( n36535 , n36305 );
or ( n36536 , n36534 , n36535 );
not ( n36537 , n36525 );
not ( n36538 , n36537 );
not ( n36539 , n36316 );
or ( n36540 , n36538 , n36539 );
and ( n36541 , n36330 , n36524 );
and ( n36542 , n36394 , n36523 );
nor ( n36543 , n36541 , n36542 );
nand ( n36544 , n36540 , n36543 );
not ( n36545 , n36544 );
nand ( n36546 , n36536 , n36545 );
buf ( n36547 , n36546 );
nor ( n36548 , n36533 , n36547 );
nand ( n36549 , n36531 , n36548 );
buf ( n36550 , n34075 );
not ( n36551 , n36550 );
not ( n36552 , n36551 );
not ( n36553 , n36286 );
or ( n36554 , n36552 , n36553 );
not ( n36555 , n33979 );
nand ( n36556 , n36554 , n36555 );
and ( n36557 , n34065 , n33314 );
not ( n36558 , n36557 );
not ( n36559 , n34091 );
not ( n36560 , n36559 );
nor ( n36561 , n36558 , n36560 );
not ( n36562 , n36561 );
not ( n36563 , n36286 );
or ( n36564 , n36562 , n36563 );
not ( n36565 , n36557 );
buf ( n36566 , n34090 );
not ( n36567 , n36566 );
and ( n36568 , n34002 , n34060 );
not ( n36569 , n36568 );
or ( n36570 , n36567 , n36569 );
not ( n36571 , n33616 );
not ( n36572 , n34036 );
or ( n36573 , n36571 , n36572 );
nand ( n36574 , n36573 , n34047 );
not ( n36575 , n36574 );
nand ( n36576 , n36570 , n36575 );
not ( n36577 , n36576 );
or ( n36578 , n36565 , n36577 );
buf ( n36579 , n33552 );
not ( n36580 , n33257 );
buf ( n36581 , n33313 );
nand ( n36582 , n36580 , n36581 );
and ( n36583 , n36579 , n36582 );
buf ( n36584 , n33559 );
not ( n36585 , n36584 );
nor ( n36586 , n36583 , n36585 );
nand ( n36587 , n36578 , n36586 );
not ( n36588 , n36587 );
nand ( n36589 , n36564 , n36588 );
buf ( n36590 , n34064 );
nor ( n36591 , n36560 , n36590 );
not ( n36592 , n36591 );
not ( n36593 , n36341 );
or ( n36594 , n36592 , n36593 );
not ( n36595 , n36590 );
not ( n36596 , n36595 );
not ( n36597 , n36566 );
not ( n36598 , n36568 );
or ( n36599 , n36597 , n36598 );
nand ( n36600 , n36599 , n36575 );
not ( n36601 , n36600 );
or ( n36602 , n36596 , n36601 );
buf ( n36603 , n33541 );
not ( n36604 , n36603 );
nand ( n36605 , n36602 , n36604 );
not ( n36606 , n36605 );
nand ( n36607 , n36594 , n36606 );
not ( n36608 , n36372 );
not ( n36609 , n36248 );
not ( n36610 , n36246 );
or ( n36611 , n36609 , n36610 );
nand ( n36612 , n36611 , n36261 );
not ( n36613 , n36612 );
not ( n36614 , n35717 );
not ( n36615 , n36614 );
not ( n36616 , n35566 );
not ( n36617 , n36616 );
nand ( n36618 , n36615 , n36617 );
not ( n36619 , n35725 );
not ( n36620 , n36619 );
not ( n36621 , n35726 );
not ( n36622 , n36621 );
buf ( n36623 , n35697 );
nand ( n36624 , n36620 , n36622 , n36623 );
not ( n36625 , n36624 );
buf ( n36626 , n36235 );
buf ( n36627 , n36626 );
nand ( n36628 , n36625 , n36617 , n36627 );
nand ( n36629 , n36613 , n36618 , n36628 );
buf ( n36630 , n35195 );
not ( n36631 , n36266 );
nand ( n36632 , n36630 , n36631 );
not ( n36633 , n36632 );
and ( n36634 , n36629 , n36633 );
not ( n36635 , n36629 );
and ( n36636 , n36635 , n36632 );
nor ( n36637 , n36634 , n36636 );
buf ( n36638 , n33356 );
not ( n36639 , n36638 );
buf ( n36640 , n34065 );
nand ( n36641 , n36639 , n36640 );
nor ( n36642 , n36560 , n36641 );
not ( n36643 , n36642 );
not ( n36644 , n36341 );
or ( n36645 , n36643 , n36644 );
not ( n36646 , n36600 );
not ( n36647 , n36641 );
not ( n36648 , n36647 );
or ( n36649 , n36646 , n36648 );
and ( n36650 , n36639 , n36579 );
buf ( n36651 , n33563 );
nor ( n36652 , n36650 , n36651 );
nand ( n36653 , n36649 , n36652 );
not ( n36654 , n36653 );
nand ( n36655 , n36645 , n36654 );
buf ( n36656 , n33427 );
not ( n36657 , n36656 );
nor ( n36658 , n36657 , n36590 );
not ( n36659 , n36658 );
nor ( n36660 , n36659 , n36560 );
not ( n36661 , n36660 );
not ( n36662 , n36286 );
or ( n36663 , n36661 , n36662 );
not ( n36664 , n36658 );
not ( n36665 , n36576 );
or ( n36666 , n36664 , n36665 );
not ( n36667 , n36656 );
not ( n36668 , n36603 );
or ( n36669 , n36667 , n36668 );
buf ( n36670 , n33546 );
nand ( n36671 , n36669 , n36670 );
not ( n36672 , n36671 );
nand ( n36673 , n36666 , n36672 );
not ( n36674 , n36673 );
nand ( n36675 , n36663 , n36674 );
not ( n36676 , n36236 );
not ( n36677 , n36676 );
or ( n36678 , n36677 , n36615 );
buf ( n36679 , n35250 );
not ( n36680 , n36679 );
not ( n36681 , n35274 );
nand ( n36682 , n36680 , n36681 );
nor ( n36683 , n36682 , n36616 );
nand ( n36684 , n36678 , n36683 );
not ( n36685 , n36682 );
and ( n36686 , n36685 , n36612 );
not ( n36687 , n36681 );
buf ( n36688 , n36273 );
not ( n36689 , n36688 );
or ( n36690 , n36687 , n36689 );
buf ( n36691 , n36276 );
not ( n36692 , n36691 );
nand ( n36693 , n36690 , n36692 );
nor ( n36694 , n36686 , n36693 );
nand ( n36695 , n36684 , n36694 );
not ( n36696 , n36695 );
not ( n36697 , n36381 );
and ( n36698 , n32774 , n36526 );
buf ( n36699 , n36413 );
not ( n36700 , n36699 );
buf ( n36701 , n29139 );
not ( n36702 , n36701 );
or ( n36703 , n36700 , n36702 );
buf ( n36704 , n18944 );
buf ( n36705 , n835 );
buf ( n36706 , n866 );
xor ( n36707 , n36705 , n36706 );
buf ( n36708 , n36707 );
buf ( n36709 , n36708 );
nand ( n36710 , n36704 , n36709 );
buf ( n36711 , n36710 );
buf ( n36712 , n36711 );
nand ( n36713 , n36703 , n36712 );
buf ( n36714 , n36713 );
buf ( n36715 , n36714 );
buf ( n36716 , n36498 );
not ( n36717 , n36716 );
buf ( n36718 , n18887 );
not ( n36719 , n36718 );
or ( n36720 , n36717 , n36719 );
buf ( n36721 , n833 );
buf ( n36722 , n868 );
xnor ( n36723 , n36721 , n36722 );
buf ( n36724 , n36723 );
buf ( n36725 , n36724 );
not ( n36726 , n36725 );
buf ( n36727 , n18898 );
nand ( n36728 , n36726 , n36727 );
buf ( n36729 , n36728 );
buf ( n36730 , n36729 );
nand ( n36731 , n36720 , n36730 );
buf ( n36732 , n36731 );
buf ( n36733 , n36732 );
not ( n36734 , n36733 );
buf ( n36735 , n36734 );
buf ( n36736 , n36735 );
xor ( n36737 , n36715 , n36736 );
xor ( n36738 , n36470 , n36487 );
and ( n36739 , n36738 , n36505 );
and ( n36740 , n36470 , n36487 );
or ( n36741 , n36739 , n36740 );
buf ( n36742 , n36741 );
buf ( n36743 , n36742 );
and ( n36744 , n36737 , n36743 );
and ( n36745 , n36715 , n36736 );
or ( n36746 , n36744 , n36745 );
buf ( n36747 , n36746 );
buf ( n36748 , n36747 );
and ( n36749 , n29174 , n29175 );
buf ( n36750 , n36749 );
buf ( n36751 , n36750 );
buf ( n36752 , n36480 );
not ( n36753 , n36752 );
buf ( n36754 , n19330 );
not ( n36755 , n36754 );
or ( n36756 , n36753 , n36755 );
buf ( n36757 , n19030 );
buf ( n36758 , n864 );
buf ( n36759 , n837 );
xor ( n36760 , n36758 , n36759 );
buf ( n36761 , n36760 );
buf ( n36762 , n36761 );
nand ( n36763 , n36757 , n36762 );
buf ( n36764 , n36763 );
buf ( n36765 , n36764 );
nand ( n36766 , n36756 , n36765 );
buf ( n36767 , n36766 );
buf ( n36768 , n36767 );
xor ( n36769 , n36751 , n36768 );
buf ( n36770 , n36439 );
not ( n36771 , n36770 );
buf ( n36772 , n19125 );
not ( n36773 , n36772 );
or ( n36774 , n36771 , n36773 );
buf ( n36775 , n19134 );
buf ( n36776 , n870 );
nand ( n36777 , n36775 , n36776 );
buf ( n36778 , n36777 );
buf ( n36779 , n36778 );
nand ( n36780 , n36774 , n36779 );
buf ( n36781 , n36780 );
buf ( n36782 , n36781 );
xor ( n36783 , n36769 , n36782 );
buf ( n36784 , n36783 );
buf ( n36785 , n36784 );
xor ( n36786 , n36420 , n36428 );
and ( n36787 , n36786 , n36446 );
and ( n36788 , n36420 , n36428 );
or ( n36789 , n36787 , n36788 );
buf ( n36790 , n36789 );
buf ( n36791 , n36790 );
xor ( n36792 , n36785 , n36791 );
xor ( n36793 , n36715 , n36736 );
xor ( n36794 , n36793 , n36743 );
buf ( n36795 , n36794 );
buf ( n36796 , n36795 );
and ( n36797 , n36792 , n36796 );
and ( n36798 , n36785 , n36791 );
or ( n36799 , n36797 , n36798 );
buf ( n36800 , n36799 );
buf ( n36801 , n36800 );
xor ( n36802 , n36748 , n36801 );
xor ( n36803 , n36751 , n36768 );
and ( n36804 , n36803 , n36782 );
and ( n36805 , n36751 , n36768 );
or ( n36806 , n36804 , n36805 );
buf ( n36807 , n36806 );
buf ( n36808 , n36807 );
and ( n36809 , n36477 , n36478 );
buf ( n36810 , n36809 );
buf ( n36811 , n36810 );
buf ( n36812 , n36708 );
not ( n36813 , n36812 );
buf ( n36814 , n29139 );
not ( n36815 , n36814 );
or ( n36816 , n36813 , n36815 );
buf ( n36817 , n834 );
buf ( n36818 , n866 );
xnor ( n36819 , n36817 , n36818 );
buf ( n36820 , n36819 );
buf ( n36821 , n36820 );
not ( n36822 , n36821 );
buf ( n36823 , n18944 );
nand ( n36824 , n36822 , n36823 );
buf ( n36825 , n36824 );
buf ( n36826 , n36825 );
nand ( n36827 , n36816 , n36826 );
buf ( n36828 , n36827 );
buf ( n36829 , n36828 );
xor ( n36830 , n36811 , n36829 );
buf ( n36831 , n36732 );
xor ( n36832 , n36830 , n36831 );
buf ( n36833 , n36832 );
buf ( n36834 , n36833 );
xor ( n36835 , n36808 , n36834 );
buf ( n36836 , n36761 );
not ( n36837 , n36836 );
buf ( n36838 , n19330 );
not ( n36839 , n36838 );
or ( n36840 , n36837 , n36839 );
buf ( n36841 , n19030 );
buf ( n36842 , n864 );
buf ( n36843 , n836 );
xor ( n36844 , n36842 , n36843 );
buf ( n36845 , n36844 );
buf ( n36846 , n36845 );
nand ( n36847 , n36841 , n36846 );
buf ( n36848 , n36847 );
buf ( n36849 , n36848 );
nand ( n36850 , n36840 , n36849 );
buf ( n36851 , n36850 );
buf ( n36852 , n36851 );
buf ( n36853 , n19134 );
buf ( n36854 , n19125 );
or ( n36855 , n36853 , n36854 );
buf ( n36856 , n870 );
nand ( n36857 , n36855 , n36856 );
buf ( n36858 , n36857 );
buf ( n36859 , n36858 );
xor ( n36860 , n36852 , n36859 );
buf ( n36861 , n18887 );
not ( n36862 , n36861 );
buf ( n36863 , n36862 );
buf ( n36864 , n36863 );
buf ( n36865 , n36724 );
or ( n36866 , n36864 , n36865 );
buf ( n36867 , n18895 );
buf ( n36868 , n868 );
buf ( n36869 , n832 );
not ( n36870 , n36869 );
buf ( n36871 , n36870 );
buf ( n36872 , n36871 );
and ( n36873 , n36868 , n36872 );
not ( n36874 , n36868 );
buf ( n36875 , n832 );
and ( n36876 , n36874 , n36875 );
nor ( n36877 , n36873 , n36876 );
buf ( n36878 , n36877 );
buf ( n36879 , n36878 );
or ( n36880 , n36867 , n36879 );
nand ( n36881 , n36866 , n36880 );
buf ( n36882 , n36881 );
buf ( n36883 , n36882 );
xor ( n36884 , n36860 , n36883 );
buf ( n36885 , n36884 );
buf ( n36886 , n36885 );
xor ( n36887 , n36835 , n36886 );
buf ( n36888 , n36887 );
buf ( n36889 , n36888 );
xor ( n36890 , n36802 , n36889 );
buf ( n36891 , n36890 );
xor ( n36892 , n36451 , n36466 );
and ( n36893 , n36892 , n36508 );
and ( n36894 , n36451 , n36466 );
or ( n36895 , n36893 , n36894 );
buf ( n36896 , n36895 );
buf ( n36897 , n36896 );
xor ( n36898 , n36785 , n36791 );
xor ( n36899 , n36898 , n36796 );
buf ( n36900 , n36899 );
buf ( n36901 , n36900 );
xor ( n36902 , n36897 , n36901 );
xor ( n36903 , n36406 , n36449 );
and ( n36904 , n36903 , n36511 );
and ( n36905 , n36406 , n36449 );
or ( n36906 , n36904 , n36905 );
buf ( n36907 , n36906 );
buf ( n36908 , n36907 );
and ( n36909 , n36902 , n36908 );
and ( n36910 , n36897 , n36901 );
or ( n36911 , n36909 , n36910 );
buf ( n36912 , n36911 );
or ( n36913 , n36891 , n36912 );
xor ( n36914 , n36400 , n36514 );
and ( n36915 , n36914 , n36521 );
and ( n36916 , n36400 , n36514 );
or ( n36917 , n36915 , n36916 );
buf ( n36918 , n36917 );
xor ( n36919 , n36897 , n36901 );
xor ( n36920 , n36919 , n36908 );
buf ( n36921 , n36920 );
or ( n36922 , n36918 , n36921 );
nand ( n36923 , n36913 , n36922 );
not ( n36924 , n36923 );
nand ( n36925 , n36698 , n36924 );
nor ( n36926 , n36697 , n36925 );
nand ( n36927 , n36926 , n36341 );
not ( n36928 , n35723 );
not ( n36929 , n36626 );
or ( n36930 , n36928 , n36929 );
buf ( n36931 , n35679 );
nand ( n36932 , n36930 , n36931 );
nand ( n36933 , n35724 , n35684 );
not ( n36934 , n36933 );
and ( n36935 , n36932 , n36934 );
not ( n36936 , n36932 );
and ( n36937 , n36936 , n36933 );
nor ( n36938 , n36935 , n36937 );
nor ( n36939 , n36621 , n35696 );
nand ( n36940 , n36939 , n36626 , n36620 );
buf ( n36941 , n35689 );
nand ( n36942 , n36939 , n36941 );
not ( n36943 , n35592 );
buf ( n36944 , n35706 );
not ( n36945 , n36944 );
or ( n36946 , n36943 , n36945 );
not ( n36947 , n35709 );
nand ( n36948 , n36946 , n36947 );
not ( n36949 , n36948 );
nand ( n36950 , n36940 , n36942 , n36949 );
nand ( n36951 , n35710 , n35712 );
nand ( n36952 , n36950 , n36951 );
not ( n36953 , n36614 );
and ( n36954 , n35565 , n36244 );
nand ( n36955 , n36953 , n36954 );
nand ( n36956 , n36625 , n36954 , n36627 );
not ( n36957 , n35538 );
not ( n36958 , n35510 );
nand ( n36959 , n36957 , n36958 );
and ( n36960 , n36959 , n36241 );
not ( n36961 , n35507 );
and ( n36962 , n36960 , n36961 );
nor ( n36963 , n36962 , n36252 );
nand ( n36964 , n36955 , n36956 , n36963 );
nand ( n36965 , n36676 , n36614 );
buf ( n36966 , n36965 );
nor ( n36967 , n36616 , n36679 );
nand ( n36968 , n36677 , n36967 );
not ( n36969 , n36630 );
nor ( n36970 , n36969 , n36616 );
nand ( n36971 , n36970 , n36677 );
buf ( n36972 , n35579 );
not ( n36973 , n36972 );
nor ( n36974 , n36619 , n36973 );
not ( n36975 , n36974 );
not ( n36976 , n36626 );
or ( n36977 , n36975 , n36976 );
not ( n36978 , n36972 );
not ( n36979 , n35689 );
or ( n36980 , n36978 , n36979 );
not ( n36981 , n35700 );
nand ( n36982 , n36980 , n36981 );
not ( n36983 , n36982 );
nand ( n36984 , n36977 , n36983 );
not ( n36985 , n36950 );
not ( n36986 , n36626 );
buf ( n36987 , n35564 );
nor ( n36988 , n36986 , n36987 );
nand ( n36989 , n36625 , n36988 );
not ( n36990 , n36216 );
not ( n36991 , n36220 );
or ( n36992 , n36990 , n36991 );
nand ( n36993 , n36992 , n36231 );
nand ( n36994 , n36993 , n35784 );
and ( n36995 , n36220 , n36186 );
not ( n36996 , n36125 );
not ( n36997 , n36996 );
nand ( n36998 , n36995 , n36997 , n35784 );
buf ( n36999 , n36198 );
nand ( n37000 , n36994 , n36998 , n36999 );
and ( n37001 , n36201 , n36204 );
and ( n37002 , n37000 , n37001 );
not ( n37003 , n37000 );
not ( n37004 , n37001 );
and ( n37005 , n37003 , n37004 );
nor ( n37006 , n37002 , n37005 );
not ( n37007 , n35722 );
nand ( n37008 , n37007 , n35663 );
not ( n37009 , n37008 );
not ( n37010 , n36626 );
or ( n37011 , n37009 , n37010 );
or ( n37012 , n36626 , n37008 );
nand ( n37013 , n37011 , n37012 );
and ( n37014 , n35723 , n35724 );
not ( n37015 , n37014 );
not ( n37016 , n36626 );
or ( n37017 , n37015 , n37016 );
not ( n37018 , n36931 );
and ( n37019 , n37018 , n35724 );
not ( n37020 , n35684 );
nor ( n37021 , n37019 , n37020 );
nand ( n37022 , n37017 , n37021 );
not ( n37023 , n36620 );
not ( n37024 , n36626 );
or ( n37025 , n37023 , n37024 );
not ( n37026 , n36941 );
nand ( n37027 , n37025 , n37026 );
not ( n37028 , n36205 );
nand ( n37029 , n36995 , n36233 , n36997 );
nand ( n37030 , n36993 , n36233 );
nand ( n37031 , n37028 , n37029 , n37030 );
nand ( n37032 , n35744 , n35750 );
buf ( n37033 , n36207 );
nand ( n37034 , n37032 , n37033 );
not ( n37035 , n37034 );
and ( n37036 , n37031 , n37035 );
not ( n37037 , n37031 );
and ( n37038 , n37037 , n37034 );
nor ( n37039 , n37036 , n37038 );
not ( n37040 , n36186 );
not ( n37041 , n36125 );
or ( n37042 , n37040 , n37041 );
not ( n37043 , n36216 );
nand ( n37044 , n37042 , n37043 );
buf ( n37045 , n36223 );
nand ( n37046 , n36156 , n37045 );
not ( n37047 , n37046 );
and ( n37048 , n37044 , n37047 );
not ( n37049 , n37044 );
and ( n37050 , n37049 , n37046 );
nor ( n37051 , n37048 , n37050 );
not ( n37052 , n36185 );
not ( n37053 , n37052 );
not ( n37054 , n36125 );
or ( n37055 , n37053 , n37054 );
nand ( n37056 , n37055 , n36212 );
not ( n37057 , n36166 );
nand ( n37058 , n37057 , n36215 );
not ( n37059 , n37058 );
and ( n37060 , n37056 , n37059 );
not ( n37061 , n37056 );
and ( n37062 , n37061 , n37058 );
nor ( n37063 , n37060 , n37062 );
nand ( n37064 , n36922 , n36527 );
not ( n37065 , n37064 );
nand ( n37066 , n36347 , n37065 );
buf ( n37067 , n34069 );
xor ( n37068 , n36811 , n36829 );
and ( n37069 , n37068 , n36831 );
and ( n37070 , n36811 , n36829 );
or ( n37071 , n37069 , n37070 );
buf ( n37072 , n37071 );
buf ( n37073 , n37072 );
xor ( n37074 , n36808 , n36834 );
and ( n37075 , n37074 , n36886 );
and ( n37076 , n36808 , n36834 );
or ( n37077 , n37075 , n37076 );
buf ( n37078 , n37077 );
buf ( n37079 , n37078 );
xor ( n37080 , n37073 , n37079 );
buf ( n37081 , n36878 );
not ( n37082 , n37081 );
buf ( n37083 , n37082 );
buf ( n37084 , n37083 );
not ( n37085 , n37084 );
buf ( n37086 , n18887 );
not ( n37087 , n37086 );
or ( n37088 , n37085 , n37087 );
buf ( n37089 , n18898 );
buf ( n37090 , n868 );
nand ( n37091 , n37089 , n37090 );
buf ( n37092 , n37091 );
buf ( n37093 , n37092 );
nand ( n37094 , n37088 , n37093 );
buf ( n37095 , n37094 );
buf ( n37096 , n37095 );
not ( n37097 , n37096 );
buf ( n37098 , n37097 );
buf ( n37099 , n37098 );
xor ( n37100 , n36852 , n36859 );
and ( n37101 , n37100 , n36883 );
and ( n37102 , n36852 , n36859 );
or ( n37103 , n37101 , n37102 );
buf ( n37104 , n37103 );
buf ( n37105 , n37104 );
xor ( n37106 , n37099 , n37105 );
and ( n37107 , n36758 , n36759 );
buf ( n37108 , n37107 );
buf ( n37109 , n37108 );
buf ( n37110 , n36845 );
not ( n37111 , n37110 );
buf ( n37112 , n19330 );
not ( n37113 , n37112 );
or ( n37114 , n37111 , n37113 );
buf ( n37115 , n864 );
buf ( n37116 , n835 );
xnor ( n37117 , n37115 , n37116 );
buf ( n37118 , n37117 );
buf ( n37119 , n37118 );
not ( n37120 , n37119 );
buf ( n37121 , n19030 );
nand ( n37122 , n37120 , n37121 );
buf ( n37123 , n37122 );
buf ( n37124 , n37123 );
nand ( n37125 , n37114 , n37124 );
buf ( n37126 , n37125 );
buf ( n37127 , n37126 );
xor ( n37128 , n37109 , n37127 );
buf ( n37129 , n29136 );
buf ( n37130 , n36820 );
or ( n37131 , n37129 , n37130 );
buf ( n37132 , n18941 );
buf ( n37133 , n866 );
buf ( n37134 , n833 );
not ( n37135 , n37134 );
buf ( n37136 , n37135 );
buf ( n37137 , n37136 );
and ( n37138 , n37133 , n37137 );
not ( n37139 , n37133 );
buf ( n37140 , n833 );
and ( n37141 , n37139 , n37140 );
nor ( n37142 , n37138 , n37141 );
buf ( n37143 , n37142 );
buf ( n37144 , n37143 );
or ( n37145 , n37132 , n37144 );
nand ( n37146 , n37131 , n37145 );
buf ( n37147 , n37146 );
buf ( n37148 , n37147 );
xor ( n37149 , n37128 , n37148 );
buf ( n37150 , n37149 );
buf ( n37151 , n37150 );
xor ( n37152 , n37106 , n37151 );
buf ( n37153 , n37152 );
buf ( n37154 , n37153 );
and ( n37155 , n37080 , n37154 );
and ( n37156 , n37073 , n37079 );
or ( n37157 , n37155 , n37156 );
buf ( n37158 , n37157 );
and ( n37159 , n36842 , n36843 );
buf ( n37160 , n37159 );
buf ( n37161 , n37160 );
buf ( n37162 , n18895 );
not ( n37163 , n37162 );
buf ( n37164 , n36863 );
not ( n37165 , n37164 );
or ( n37166 , n37163 , n37165 );
buf ( n37167 , n868 );
nand ( n37168 , n37166 , n37167 );
buf ( n37169 , n37168 );
buf ( n37170 , n37169 );
xor ( n37171 , n37161 , n37170 );
buf ( n37172 , n29136 );
buf ( n37173 , n37143 );
or ( n37174 , n37172 , n37173 );
buf ( n37175 , n18941 );
buf ( n37176 , n832 );
buf ( n37177 , n866 );
xnor ( n37178 , n37176 , n37177 );
buf ( n37179 , n37178 );
buf ( n37180 , n37179 );
or ( n37181 , n37175 , n37180 );
nand ( n37182 , n37174 , n37181 );
buf ( n37183 , n37182 );
buf ( n37184 , n37183 );
xor ( n37185 , n37171 , n37184 );
buf ( n37186 , n37185 );
buf ( n37187 , n37186 );
buf ( n37188 , n37095 );
buf ( n37189 , n19016 );
buf ( n37190 , n37118 );
or ( n37191 , n37189 , n37190 );
buf ( n37192 , n19033 );
buf ( n37193 , n864 );
buf ( n37194 , n834 );
xnor ( n37195 , n37193 , n37194 );
buf ( n37196 , n37195 );
buf ( n37197 , n37196 );
or ( n37198 , n37192 , n37197 );
nand ( n37199 , n37191 , n37198 );
buf ( n37200 , n37199 );
buf ( n37201 , n37200 );
xor ( n37202 , n37188 , n37201 );
xor ( n37203 , n37109 , n37127 );
and ( n37204 , n37203 , n37148 );
and ( n37205 , n37109 , n37127 );
or ( n37206 , n37204 , n37205 );
buf ( n37207 , n37206 );
buf ( n37208 , n37207 );
xor ( n37209 , n37202 , n37208 );
buf ( n37210 , n37209 );
buf ( n37211 , n37210 );
xor ( n37212 , n37187 , n37211 );
xor ( n37213 , n37099 , n37105 );
and ( n37214 , n37213 , n37151 );
and ( n37215 , n37099 , n37105 );
or ( n37216 , n37214 , n37215 );
buf ( n37217 , n37216 );
buf ( n37218 , n37217 );
xor ( n37219 , n37212 , n37218 );
buf ( n37220 , n37219 );
nor ( n37221 , n37158 , n37220 );
not ( n37222 , n37221 );
xor ( n37223 , n36748 , n36801 );
and ( n37224 , n37223 , n36889 );
and ( n37225 , n36748 , n36801 );
or ( n37226 , n37224 , n37225 );
buf ( n37227 , n37226 );
xor ( n37228 , n37073 , n37079 );
xor ( n37229 , n37228 , n37154 );
buf ( n37230 , n37229 );
or ( n37231 , n37227 , n37230 );
nand ( n37232 , n37222 , n37231 );
nor ( n37233 , n36923 , n37232 );
xor ( n37234 , n37187 , n37211 );
and ( n37235 , n37234 , n37218 );
and ( n37236 , n37187 , n37211 );
or ( n37237 , n37235 , n37236 );
buf ( n37238 , n37237 );
xor ( n37239 , n37161 , n37170 );
and ( n37240 , n37239 , n37184 );
and ( n37241 , n37161 , n37170 );
or ( n37242 , n37240 , n37241 );
buf ( n37243 , n37242 );
buf ( n37244 , n37243 );
buf ( n37245 , n835 );
buf ( n37246 , n864 );
and ( n37247 , n37245 , n37246 );
buf ( n37248 , n37247 );
buf ( n37249 , n37248 );
buf ( n37250 , n37179 );
not ( n37251 , n37250 );
buf ( n37252 , n29139 );
nand ( n37253 , n37251 , n37252 );
buf ( n37254 , n37253 );
buf ( n37255 , n37254 );
buf ( n37256 , n18944 );
buf ( n37257 , n866 );
nand ( n37258 , n37256 , n37257 );
buf ( n37259 , n37258 );
buf ( n37260 , n37259 );
and ( n37261 , n37255 , n37260 );
buf ( n37262 , n37261 );
buf ( n37263 , n37262 );
xor ( n37264 , n37249 , n37263 );
buf ( n37265 , n19016 );
buf ( n37266 , n37196 );
or ( n37267 , n37265 , n37266 );
buf ( n37268 , n19033 );
buf ( n37269 , n864 );
buf ( n37270 , n37136 );
and ( n37271 , n37269 , n37270 );
not ( n37272 , n37269 );
buf ( n37273 , n833 );
and ( n37274 , n37272 , n37273 );
nor ( n37275 , n37271 , n37274 );
buf ( n37276 , n37275 );
buf ( n37277 , n37276 );
or ( n37278 , n37268 , n37277 );
nand ( n37279 , n37267 , n37278 );
buf ( n37280 , n37279 );
buf ( n37281 , n37280 );
xor ( n37282 , n37264 , n37281 );
buf ( n37283 , n37282 );
buf ( n37284 , n37283 );
xor ( n37285 , n37244 , n37284 );
xor ( n37286 , n37188 , n37201 );
and ( n37287 , n37286 , n37208 );
and ( n37288 , n37188 , n37201 );
or ( n37289 , n37287 , n37288 );
buf ( n37290 , n37289 );
buf ( n37291 , n37290 );
xor ( n37292 , n37285 , n37291 );
buf ( n37293 , n37292 );
nor ( n37294 , n37238 , n37293 );
xor ( n37295 , n37244 , n37284 );
and ( n37296 , n37295 , n37291 );
and ( n37297 , n37244 , n37284 );
or ( n37298 , n37296 , n37297 );
buf ( n37299 , n37298 );
buf ( n37300 , n37262 );
not ( n37301 , n37300 );
buf ( n37302 , n37301 );
buf ( n37303 , n37302 );
xor ( n37304 , n37249 , n37263 );
and ( n37305 , n37304 , n37281 );
and ( n37306 , n37249 , n37263 );
or ( n37307 , n37305 , n37306 );
buf ( n37308 , n37307 );
buf ( n37309 , n37308 );
xor ( n37310 , n37303 , n37309 );
buf ( n37311 , n29139 );
buf ( n37312 , n18944 );
or ( n37313 , n37311 , n37312 );
buf ( n37314 , n866 );
nand ( n37315 , n37313 , n37314 );
buf ( n37316 , n37315 );
buf ( n37317 , n37316 );
buf ( n37318 , n834 );
buf ( n37319 , n864 );
and ( n37320 , n37318 , n37319 );
buf ( n37321 , n37320 );
buf ( n37322 , n37321 );
xor ( n37323 , n37317 , n37322 );
buf ( n37324 , n19016 );
buf ( n37325 , n37276 );
or ( n37326 , n37324 , n37325 );
buf ( n37327 , n19033 );
buf ( n37328 , n864 );
buf ( n37329 , n36871 );
and ( n37330 , n37328 , n37329 );
not ( n37331 , n37328 );
buf ( n37332 , n832 );
and ( n37333 , n37331 , n37332 );
nor ( n37334 , n37330 , n37333 );
buf ( n37335 , n37334 );
buf ( n37336 , n37335 );
or ( n37337 , n37327 , n37336 );
nand ( n37338 , n37326 , n37337 );
buf ( n37339 , n37338 );
buf ( n37340 , n37339 );
xor ( n37341 , n37323 , n37340 );
buf ( n37342 , n37341 );
buf ( n37343 , n37342 );
xor ( n37344 , n37310 , n37343 );
buf ( n37345 , n37344 );
nor ( n37346 , n37299 , n37345 );
nor ( n37347 , n37294 , n37346 );
xor ( n37348 , n37303 , n37309 );
and ( n37349 , n37348 , n37343 );
and ( n37350 , n37303 , n37309 );
or ( n37351 , n37349 , n37350 );
buf ( n37352 , n37351 );
buf ( n37353 , n833 );
buf ( n37354 , n864 );
nand ( n37355 , n37353 , n37354 );
buf ( n37356 , n37355 );
buf ( n37357 , n37356 );
buf ( n37358 , n19016 );
buf ( n37359 , n37335 );
or ( n37360 , n37358 , n37359 );
buf ( n37361 , n19033 );
buf ( n37362 , n864 );
not ( n37363 , n37362 );
buf ( n37364 , n37363 );
buf ( n37365 , n37364 );
or ( n37366 , n37361 , n37365 );
nand ( n37367 , n37360 , n37366 );
buf ( n37368 , n37367 );
buf ( n37369 , n37368 );
xor ( n37370 , n37357 , n37369 );
xor ( n37371 , n37317 , n37322 );
and ( n37372 , n37371 , n37340 );
and ( n37373 , n37317 , n37322 );
or ( n37374 , n37372 , n37373 );
buf ( n37375 , n37374 );
buf ( n37376 , n37375 );
xor ( n37377 , n37370 , n37376 );
buf ( n37378 , n37377 );
or ( n37379 , n37352 , n37378 );
and ( n37380 , n37347 , n37379 );
and ( n37381 , n37233 , n37380 );
and ( n37382 , n36528 , n37381 );
nand ( n37383 , n37067 , n37382 );
and ( n37384 , n36219 , n36186 );
not ( n37385 , n37384 );
not ( n37386 , n36125 );
or ( n37387 , n37385 , n37386 );
not ( n37388 , n36156 );
not ( n37389 , n36216 );
or ( n37390 , n37388 , n37389 );
nand ( n37391 , n37390 , n37045 );
not ( n37392 , n37391 );
nand ( n37393 , n37387 , n37392 );
not ( n37394 , n36347 );
not ( n37395 , n36640 );
not ( n37396 , n36576 );
or ( n37397 , n37395 , n37396 );
not ( n37398 , n36579 );
nand ( n37399 , n37397 , n37398 );
not ( n37400 , n37399 );
not ( n37401 , n36924 );
not ( n37402 , n36546 );
or ( n37403 , n37401 , n37402 );
not ( n37404 , n36913 );
and ( n37405 , n36921 , n36918 );
not ( n37406 , n37405 );
or ( n37407 , n37404 , n37406 );
nand ( n37408 , n36891 , n36912 );
nand ( n37409 , n37407 , n37408 );
not ( n37410 , n37409 );
nand ( n37411 , n37403 , n37410 );
not ( n37412 , n37411 );
not ( n37413 , n36922 );
not ( n37414 , n36546 );
or ( n37415 , n37413 , n37414 );
not ( n37416 , n37405 );
nand ( n37417 , n37415 , n37416 );
not ( n37418 , n37417 );
buf ( n37419 , n34063 );
not ( n37420 , n37419 );
not ( n37421 , n36600 );
or ( n37422 , n37420 , n37421 );
not ( n37423 , n33526 );
nand ( n37424 , n37422 , n37423 );
not ( n37425 , n37424 );
buf ( n37426 , n33384 );
not ( n37427 , n37426 );
nor ( n37428 , n37427 , n36638 );
nand ( n37429 , n37428 , n36640 );
not ( n37430 , n37429 );
not ( n37431 , n37430 );
not ( n37432 , n36600 );
or ( n37433 , n37431 , n37432 );
not ( n37434 , n37428 );
not ( n37435 , n36579 );
or ( n37436 , n37434 , n37435 );
and ( n37437 , n36651 , n37426 );
not ( n37438 , n33566 );
nor ( n37439 , n37437 , n37438 );
nand ( n37440 , n37436 , n37439 );
not ( n37441 , n37440 );
nand ( n37442 , n37433 , n37441 );
not ( n37443 , n37442 );
not ( n37444 , n37231 );
nor ( n37445 , n37444 , n36923 );
not ( n37446 , n37445 );
not ( n37447 , n36546 );
or ( n37448 , n37446 , n37447 );
not ( n37449 , n37231 );
not ( n37450 , n37409 );
or ( n37451 , n37449 , n37450 );
nand ( n37452 , n37227 , n37230 );
nand ( n37453 , n37451 , n37452 );
not ( n37454 , n37453 );
nand ( n37455 , n37448 , n37454 );
nand ( n37456 , n36967 , n36615 );
not ( n37457 , n35564 );
nand ( n37458 , n36615 , n37457 );
nand ( n37459 , n36970 , n36615 );
not ( n37460 , n35979 );
not ( n37461 , n35980 );
or ( n37462 , n37460 , n37461 );
nand ( n37463 , n37462 , n35844 );
not ( n37464 , n36630 );
not ( n37465 , n36612 );
or ( n37466 , n37464 , n37465 );
nand ( n37467 , n37466 , n36631 );
nand ( n37468 , n35980 , n35844 );
buf ( n37469 , n35979 );
nand ( n37470 , n37468 , n37469 );
not ( n37471 , n36679 );
not ( n37472 , n37471 );
not ( n37473 , n36612 );
or ( n37474 , n37472 , n37473 );
not ( n37475 , n36688 );
nand ( n37476 , n37474 , n37475 );
not ( n37477 , n37347 );
not ( n37478 , n37232 );
not ( n37479 , n37478 );
not ( n37480 , n37409 );
or ( n37481 , n37479 , n37480 );
not ( n37482 , n37452 );
not ( n37483 , n37221 );
and ( n37484 , n37482 , n37483 );
and ( n37485 , n37158 , n37220 );
nor ( n37486 , n37484 , n37485 );
nand ( n37487 , n37481 , n37486 );
not ( n37488 , n37487 );
or ( n37489 , n37477 , n37488 );
nand ( n37490 , n37238 , n37293 );
or ( n37491 , n37490 , n37346 );
nand ( n37492 , n37299 , n37345 );
nand ( n37493 , n37491 , n37492 );
not ( n37494 , n37493 );
nand ( n37495 , n37489 , n37494 );
not ( n37496 , n37294 );
not ( n37497 , n37496 );
not ( n37498 , n37487 );
or ( n37499 , n37497 , n37498 );
nand ( n37500 , n37499 , n37490 );
not ( n37501 , n37500 );
not ( n37502 , n36576 );
not ( n37503 , n37380 );
not ( n37504 , n37487 );
or ( n37505 , n37503 , n37504 );
and ( n37506 , n37493 , n37379 );
and ( n37507 , n37352 , n37378 );
nor ( n37508 , n37506 , n37507 );
nand ( n37509 , n37505 , n37508 );
buf ( n37510 , n34033 );
or ( n37511 , n37510 , n24074 );
not ( n37512 , n34055 );
nand ( n37513 , n37511 , n37512 );
not ( n37514 , n37513 );
buf ( n37515 , n36568 );
and ( n37516 , n37514 , n37515 );
not ( n37517 , n37511 );
not ( n37518 , n34049 );
not ( n37519 , n37518 );
or ( n37520 , n37517 , n37519 );
nand ( n37521 , n37520 , n34041 );
nor ( n37522 , n37516 , n37521 );
not ( n37523 , n36381 );
nor ( n37524 , n37523 , n37064 );
not ( n37525 , n34094 );
and ( n37526 , n36289 , n36328 );
nand ( n37527 , n36339 , n37526 );
nor ( n37528 , n37525 , n37527 );
not ( n37529 , n32690 );
buf ( n37530 , n32517 );
nor ( n37531 , n37529 , n37530 );
and ( n37532 , n36338 , n37531 );
nand ( n37533 , n35977 , n35947 );
not ( n37534 , n35974 );
not ( n37535 , n35975 );
nand ( n37536 , n37534 , n37535 );
nand ( n37537 , n37533 , n37536 );
not ( n37538 , n37515 );
nor ( n37539 , n36560 , n37429 );
and ( n37540 , n37233 , n37347 );
nand ( n37541 , n36528 , n37540 );
nand ( n37542 , n36528 , n37233 );
and ( n37543 , n37233 , n37496 );
nand ( n37544 , n36528 , n37543 );
not ( n37545 , n32690 );
not ( n37546 , n36297 );
or ( n37547 , n37545 , n37546 );
not ( n37548 , n36300 );
nand ( n37549 , n37547 , n37548 );
buf ( n37550 , n34085 );
not ( n37551 , n37550 );
nor ( n37552 , n37551 , n34055 );
not ( n37553 , n36366 );
and ( n37554 , n35924 , n35845 );
not ( n37555 , n35927 );
nor ( n37556 , n37554 , n37555 );
nand ( n37557 , n33604 , n33600 );
and ( n37558 , n37557 , n34051 );
not ( n37559 , n37558 );
nand ( n37560 , n35678 , n35673 );
not ( n37561 , n37560 );
nand ( n37562 , n37426 , n33566 );
not ( n37563 , n37562 );
nand ( n37564 , n36656 , n36670 );
not ( n37565 , n37564 );
nand ( n37566 , n36681 , n36692 );
not ( n37567 , n37566 );
not ( n37568 , n36357 );
nand ( n37569 , n36922 , n37416 );
nand ( n37570 , n37231 , n37452 );
nand ( n37571 , n36972 , n36981 );
nand ( n37572 , n32828 , n36315 );
not ( n37573 , n35795 );
not ( n37574 , n37573 );
nand ( n37575 , n37574 , n36229 );
nand ( n37576 , n37419 , n37423 );
nand ( n37577 , n35924 , n35927 );
not ( n37578 , n36281 );
nand ( n37579 , n37578 , n36279 );
not ( n37580 , n37579 );
nand ( n37581 , n35784 , n36198 );
not ( n37582 , n37581 );
not ( n37583 , n36951 );
buf ( n37584 , n37221 );
nor ( n37585 , n37485 , n37584 );
not ( n37586 , n37585 );
not ( n37587 , n35718 );
nor ( n37588 , n37587 , n35687 );
not ( n37589 , n37588 );
not ( n37590 , n36374 );
not ( n37591 , n36055 );
not ( n37592 , n36088 );
or ( n37593 , n37591 , n37592 );
nand ( n37594 , n37593 , n36122 );
not ( n37595 , n37594 );
not ( n37596 , n37530 );
nand ( n37597 , n36551 , n36555 );
buf ( n37598 , n37356 );
not ( n37599 , n37598 );
buf ( n37600 , n832 );
buf ( n37601 , n864 );
nand ( n37602 , n37600 , n37601 );
buf ( n37603 , n37602 );
buf ( n37604 , n37603 );
not ( n37605 , n37604 );
buf ( n37606 , n19330 );
buf ( n37607 , n19030 );
or ( n37608 , n37606 , n37607 );
buf ( n37609 , n864 );
nand ( n37610 , n37608 , n37609 );
buf ( n37611 , n37610 );
buf ( n37612 , n37611 );
not ( n37613 , n37612 );
or ( n37614 , n37605 , n37613 );
buf ( n37615 , n37611 );
buf ( n37616 , n37603 );
or ( n37617 , n37615 , n37616 );
nand ( n37618 , n37614 , n37617 );
buf ( n37619 , n37618 );
buf ( n37620 , n37619 );
not ( n37621 , n37620 );
or ( n37622 , n37599 , n37621 );
buf ( n37623 , n37619 );
buf ( n37624 , n37356 );
or ( n37625 , n37623 , n37624 );
nand ( n37626 , n37622 , n37625 );
buf ( n37627 , n37626 );
not ( n37628 , n37627 );
xor ( n37629 , n37357 , n37369 );
and ( n37630 , n37629 , n37376 );
and ( n37631 , n37357 , n37369 );
or ( n37632 , n37630 , n37631 );
buf ( n37633 , n37632 );
not ( n37634 , n37633 );
or ( n37635 , n37628 , n37634 );
or ( n37636 , n37633 , n37627 );
nand ( n37637 , n37635 , n37636 );
not ( n37638 , n37346 );
nand ( n37639 , n37638 , n37492 );
nand ( n37640 , n36959 , n36240 );
nand ( n37641 , n37052 , n36212 );
not ( n37642 , n36108 );
nand ( n37643 , n37642 , n36115 );
and ( n37644 , n37233 , n36547 );
nor ( n37645 , n37644 , n37487 );
and ( n37646 , n37381 , n36547 );
nor ( n37647 , n37646 , n37509 );
and ( n37648 , n35726 , n36941 );
nor ( n37649 , n37648 , n36944 );
or ( n37650 , n35972 , n29005 );
and ( n37651 , n35973 , n37650 );
not ( n37652 , n37476 );
nand ( n37653 , n37652 , n37456 , n36968 );
nand ( n37654 , n36698 , n37445 );
not ( n37655 , n37654 );
nand ( n37656 , n37655 , n36347 );
not ( n37657 , n36925 );
nand ( n37658 , n37657 , n34069 );
not ( n37659 , n37542 );
nand ( n37660 , n37659 , n37067 );
not ( n37661 , n37527 );
nand ( n37662 , n37661 , n34069 );
not ( n37663 , n35964 );
nand ( n37664 , n37663 , n37535 );
xor ( n37665 , n37664 , n35973 );
not ( n37666 , n36233 );
nor ( n37667 , n37666 , n36196 );
not ( n37668 , n33556 );
nand ( n37669 , n37668 , n33562 );
not ( n37670 , n37419 );
nor ( n37671 , n37670 , n36560 );
not ( n37672 , n36252 );
nand ( n37673 , n37672 , n36244 );
and ( n37674 , n31796 , n30976 );
xor ( n37675 , n16684 , n16678 );
not ( n37676 , n37675 );
buf ( n37677 , n16216 );
buf ( n37678 , n15956 );
and ( n37679 , n37677 , n37678 );
buf ( n37680 , n37679 );
not ( n37681 , n37680 );
and ( n37682 , n37676 , n37681 );
and ( n37683 , n15949 , n15650 );
buf ( n37684 , n37683 );
xor ( n37685 , n15956 , n16216 );
buf ( n37686 , n37685 );
nor ( n37687 , n37684 , n37686 );
buf ( n37688 , n37687 );
nor ( n37689 , n37682 , n37688 );
nand ( n37690 , n37674 , n37689 );
buf ( n37691 , n37690 );
not ( n37692 , n37691 );
buf ( n37693 , n37692 );
not ( n37694 , n31759 );
and ( n37695 , n37693 , n37694 );
nor ( n37696 , n37680 , n37675 );
nor ( n37697 , n37696 , n37688 );
not ( n37698 , n37697 );
not ( n37699 , n31766 );
or ( n37700 , n31793 , n31795 );
not ( n37701 , n37700 );
or ( n37702 , n37699 , n37701 );
nand ( n37703 , n37702 , n31798 );
not ( n37704 , n37703 );
or ( n37705 , n37698 , n37704 );
not ( n37706 , n37696 );
buf ( n37707 , n37683 );
buf ( n37708 , n37685 );
nand ( n37709 , n37707 , n37708 );
buf ( n37710 , n37709 );
not ( n37711 , n37710 );
and ( n37712 , n37706 , n37711 );
nand ( n37713 , n37675 , n37680 );
not ( n37714 , n37713 );
nor ( n37715 , n37712 , n37714 );
nand ( n37716 , n37705 , n37715 );
nor ( n37717 , n37695 , n37716 );
buf ( n37718 , n37717 );
buf ( n37719 , n31748 );
buf ( n37720 , n37690 );
or ( n37721 , n37719 , n37720 );
buf ( n37722 , n37721 );
buf ( n37723 , n37722 );
not ( n37724 , n31032 );
nand ( n37725 , n37724 , n37693 );
buf ( n37726 , n37725 );
nand ( n37727 , n37718 , n37723 , n37726 );
buf ( n37728 , n37727 );
buf ( n37729 , n37728 );
buf ( n37730 , n31716 );
not ( n37731 , n37697 );
not ( n37732 , n37703 );
or ( n37733 , n37731 , n37732 );
nand ( n37734 , n37733 , n37715 );
buf ( n37735 , n37734 );
not ( n37736 , n37735 );
buf ( n37737 , n37736 );
buf ( n37738 , n37737 );
and ( n37739 , n37730 , n37738 );
buf ( n37740 , n37739 );
buf ( n37741 , n37740 );
buf ( n37742 , n31748 );
buf ( n37743 , n31693 );
buf ( n37744 , n31758 );
nor ( n37745 , n37743 , n37744 );
buf ( n37746 , n37745 );
buf ( n37747 , n37746 );
and ( n37748 , n37742 , n37747 );
buf ( n37749 , n37748 );
buf ( n37750 , n37749 );
buf ( n37751 , n31670 );
nand ( n37752 , n37741 , n37750 , n37751 );
buf ( n37753 , n37752 );
buf ( n37754 , n37753 );
nand ( n37755 , n37729 , n37754 );
buf ( n37756 , n37755 );
buf ( n37757 , n37756 );
buf ( n37758 , n37757 );
buf ( n37759 , n37758 );
buf ( n37760 , n37759 );
not ( n37761 , n37760 );
buf ( n37762 , n37761 );
not ( n37763 , n37762 );
buf ( n37764 , n17461 );
buf ( n37765 , n17590 );
xor ( n37766 , n37764 , n37765 );
buf ( n37767 , n37766 );
buf ( n37768 , n37767 );
buf ( n37769 , n17600 );
buf ( n37770 , n17636 );
and ( n37771 , n37769 , n37770 );
buf ( n37772 , n37771 );
buf ( n37773 , n37772 );
nor ( n37774 , n37768 , n37773 );
buf ( n37775 , n37774 );
buf ( n37776 , n37775 );
buf ( n37777 , n17672 );
xor ( n37778 , n37769 , n37770 );
buf ( n37779 , n37778 );
buf ( n37780 , n37779 );
nor ( n37781 , n37777 , n37780 );
buf ( n37782 , n37781 );
buf ( n37783 , n37782 );
nor ( n37784 , n37776 , n37783 );
buf ( n37785 , n37784 );
buf ( n37786 , n37785 );
buf ( n37787 , n16678 );
buf ( n37788 , n16684 );
and ( n37789 , n37787 , n37788 );
buf ( n37790 , n37789 );
buf ( n37791 , n37790 );
xor ( n37792 , n17691 , n17694 );
buf ( n37793 , n37792 );
nor ( n37794 , n37791 , n37793 );
buf ( n37795 , n37794 );
buf ( n37796 , n37795 );
buf ( n37797 , n17694 );
buf ( n37798 , n17691 );
and ( n37799 , n37797 , n37798 );
buf ( n37800 , n37799 );
buf ( n37801 , n37800 );
buf ( n37802 , n17723 );
nor ( n37803 , n37801 , n37802 );
buf ( n37804 , n37803 );
buf ( n37805 , n37804 );
nor ( n37806 , n37796 , n37805 );
buf ( n37807 , n37806 );
buf ( n37808 , n37807 );
nand ( n37809 , n37786 , n37808 );
buf ( n37810 , n37809 );
buf ( n37811 , n37810 );
and ( n37812 , n37764 , n37765 );
buf ( n37813 , n37812 );
buf ( n37814 , n37813 );
not ( n37815 , n37814 );
buf ( n37816 , n17921 );
buf ( n37817 , n17748 );
xor ( n37818 , n37816 , n37817 );
buf ( n37819 , n37818 );
buf ( n37820 , n37819 );
not ( n37821 , n37820 );
buf ( n37822 , n37821 );
buf ( n37823 , n37822 );
nand ( n37824 , n37815 , n37823 );
buf ( n37825 , n37824 );
buf ( n37826 , n37825 );
xor ( n37827 , n18089 , n18083 );
buf ( n37828 , n37827 );
and ( n37829 , n37816 , n37817 );
buf ( n37830 , n37829 );
buf ( n37831 , n37830 );
or ( n37832 , n37828 , n37831 );
buf ( n37833 , n37832 );
buf ( n37834 , n37833 );
and ( n37835 , n37826 , n37834 );
buf ( n37836 , n37835 );
buf ( n37837 , n37836 );
and ( n37838 , n18089 , n18083 );
buf ( n37839 , n37838 );
buf ( n37840 , n18351 );
buf ( n37841 , n18357 );
xor ( n37842 , n37840 , n37841 );
buf ( n37843 , n37842 );
buf ( n37844 , n37843 );
nor ( n37845 , n37839 , n37844 );
buf ( n37846 , n37845 );
buf ( n37847 , n37846 );
and ( n37848 , n37840 , n37841 );
buf ( n37849 , n37848 );
buf ( n37850 , n37849 );
xor ( n37851 , n18228 , n18234 );
and ( n37852 , n37851 , n18282 );
and ( n37853 , n18228 , n18234 );
or ( n37854 , n37852 , n37853 );
buf ( n37855 , n37854 );
buf ( n37856 , n37855 );
xor ( n37857 , n18288 , n18305 );
and ( n37858 , n37857 , n18323 );
and ( n37859 , n18288 , n18305 );
or ( n37860 , n37858 , n37859 );
buf ( n37861 , n37860 );
buf ( n37862 , n37861 );
or ( n37863 , n2709 , n2713 );
nand ( n37864 , n37863 , n808 );
buf ( n37865 , n37864 );
buf ( n37866 , n18313 );
not ( n37867 , n37866 );
buf ( n37868 , n14278 );
not ( n37869 , n37868 );
or ( n37870 , n37867 , n37869 );
buf ( n37871 , n14284 );
buf ( n37872 , n806 );
buf ( n37873 , n768 );
and ( n37874 , n37872 , n37873 );
not ( n37875 , n37872 );
buf ( n37876 , n768 );
not ( n37877 , n37876 );
buf ( n37878 , n37877 );
buf ( n37879 , n37878 );
and ( n37880 , n37875 , n37879 );
nor ( n37881 , n37874 , n37880 );
buf ( n37882 , n37881 );
buf ( n37883 , n37882 );
nand ( n37884 , n37871 , n37883 );
buf ( n37885 , n37884 );
buf ( n37886 , n37885 );
nand ( n37887 , n37870 , n37886 );
buf ( n37888 , n37887 );
buf ( n37889 , n37888 );
xor ( n37890 , n37865 , n37889 );
buf ( n37891 , n18274 );
not ( n37892 , n37891 );
buf ( n37893 , n3109 );
not ( n37894 , n37893 );
or ( n37895 , n37892 , n37894 );
buf ( n37896 , n1560 );
buf ( n37897 , n772 );
buf ( n37898 , n802 );
xor ( n37899 , n37897 , n37898 );
buf ( n37900 , n37899 );
buf ( n37901 , n37900 );
nand ( n37902 , n37896 , n37901 );
buf ( n37903 , n37902 );
buf ( n37904 , n37903 );
nand ( n37905 , n37895 , n37904 );
buf ( n37906 , n37905 );
buf ( n37907 , n37906 );
xor ( n37908 , n37890 , n37907 );
buf ( n37909 , n37908 );
buf ( n37910 , n37909 );
xor ( n37911 , n37862 , n37910 );
buf ( n37912 , n18319 );
xor ( n37913 , n18251 , n18263 );
and ( n37914 , n37913 , n18280 );
and ( n37915 , n18251 , n18263 );
or ( n37916 , n37914 , n37915 );
buf ( n37917 , n37916 );
xor ( n37918 , n37912 , n37917 );
and ( n37919 , n17993 , n17994 );
buf ( n37920 , n37919 );
buf ( n37921 , n37920 );
buf ( n37922 , n18245 );
not ( n37923 , n37922 );
buf ( n37924 , n10509 );
not ( n37925 , n37924 );
or ( n37926 , n37923 , n37925 );
buf ( n37927 , n3662 );
buf ( n37928 , n774 );
buf ( n37929 , n800 );
xor ( n37930 , n37928 , n37929 );
buf ( n37931 , n37930 );
buf ( n37932 , n37931 );
nand ( n37933 , n37927 , n37932 );
buf ( n37934 , n37933 );
buf ( n37935 , n37934 );
nand ( n37936 , n37926 , n37935 );
buf ( n37937 , n37936 );
buf ( n37938 , n37937 );
xor ( n37939 , n37921 , n37938 );
buf ( n37940 , n18298 );
not ( n37941 , n37940 );
buf ( n37942 , n15873 );
not ( n37943 , n37942 );
or ( n37944 , n37941 , n37943 );
buf ( n37945 , n11137 );
buf ( n37946 , n770 );
buf ( n37947 , n804 );
xor ( n37948 , n37946 , n37947 );
buf ( n37949 , n37948 );
buf ( n37950 , n37949 );
nand ( n37951 , n37945 , n37950 );
buf ( n37952 , n37951 );
buf ( n37953 , n37952 );
nand ( n37954 , n37944 , n37953 );
buf ( n37955 , n37954 );
buf ( n37956 , n37955 );
xor ( n37957 , n37939 , n37956 );
buf ( n37958 , n37957 );
buf ( n37959 , n37958 );
xor ( n37960 , n37918 , n37959 );
buf ( n37961 , n37960 );
buf ( n37962 , n37961 );
xor ( n37963 , n37911 , n37962 );
buf ( n37964 , n37963 );
buf ( n37965 , n37964 );
xor ( n37966 , n37856 , n37965 );
xor ( n37967 , n18326 , n18332 );
and ( n37968 , n37967 , n18339 );
and ( n37969 , n18326 , n18332 );
or ( n37970 , n37968 , n37969 );
buf ( n37971 , n37970 );
buf ( n37972 , n37971 );
xor ( n37973 , n37966 , n37972 );
buf ( n37974 , n37973 );
buf ( n37975 , n37974 );
xor ( n37976 , n18285 , n18342 );
and ( n37977 , n37976 , n18349 );
and ( n37978 , n18285 , n18342 );
or ( n37979 , n37977 , n37978 );
buf ( n37980 , n37979 );
buf ( n37981 , n37980 );
xor ( n37982 , n37975 , n37981 );
buf ( n37983 , n37982 );
buf ( n37984 , n37983 );
nor ( n37985 , n37850 , n37984 );
buf ( n37986 , n37985 );
buf ( n37987 , n37986 );
nor ( n37988 , n37847 , n37987 );
buf ( n37989 , n37988 );
buf ( n37990 , n37989 );
nand ( n37991 , n37837 , n37990 );
buf ( n37992 , n37991 );
buf ( n37993 , n37992 );
nor ( n37994 , n37811 , n37993 );
buf ( n37995 , n37994 );
buf ( n37996 , n37995 );
and ( n37997 , n37975 , n37981 );
buf ( n37998 , n37997 );
buf ( n37999 , n37998 );
xor ( n38000 , n37912 , n37917 );
and ( n38001 , n38000 , n37959 );
and ( n38002 , n37912 , n37917 );
or ( n38003 , n38001 , n38002 );
buf ( n38004 , n38003 );
buf ( n38005 , n38004 );
and ( n38006 , n18242 , n18243 );
buf ( n38007 , n38006 );
buf ( n38008 , n38007 );
buf ( n38009 , n37931 );
not ( n38010 , n38009 );
buf ( n38011 , n10509 );
not ( n38012 , n38011 );
or ( n38013 , n38010 , n38012 );
buf ( n38014 , n800 );
buf ( n38015 , n773 );
xnor ( n38016 , n38014 , n38015 );
buf ( n38017 , n38016 );
buf ( n38018 , n38017 );
not ( n38019 , n38018 );
buf ( n38020 , n3662 );
nand ( n38021 , n38019 , n38020 );
buf ( n38022 , n38021 );
buf ( n38023 , n38022 );
nand ( n38024 , n38013 , n38023 );
buf ( n38025 , n38024 );
buf ( n38026 , n38025 );
xor ( n38027 , n38008 , n38026 );
buf ( n38028 , n37882 );
not ( n38029 , n38028 );
buf ( n38030 , n14278 );
not ( n38031 , n38030 );
or ( n38032 , n38029 , n38031 );
buf ( n38033 , n14284 );
buf ( n38034 , n806 );
nand ( n38035 , n38033 , n38034 );
buf ( n38036 , n38035 );
buf ( n38037 , n38036 );
nand ( n38038 , n38032 , n38037 );
buf ( n38039 , n38038 );
buf ( n38040 , n38039 );
xor ( n38041 , n38027 , n38040 );
buf ( n38042 , n38041 );
buf ( n38043 , n38042 );
xor ( n38044 , n37865 , n37889 );
and ( n38045 , n38044 , n37907 );
and ( n38046 , n37865 , n37889 );
or ( n38047 , n38045 , n38046 );
buf ( n38048 , n38047 );
buf ( n38049 , n38048 );
xor ( n38050 , n38043 , n38049 );
buf ( n38051 , n37949 );
not ( n38052 , n38051 );
buf ( n38053 , n15873 );
not ( n38054 , n38053 );
or ( n38055 , n38052 , n38054 );
buf ( n38056 , n11137 );
buf ( n38057 , n769 );
buf ( n38058 , n804 );
xor ( n38059 , n38057 , n38058 );
buf ( n38060 , n38059 );
buf ( n38061 , n38060 );
nand ( n38062 , n38056 , n38061 );
buf ( n38063 , n38062 );
buf ( n38064 , n38063 );
nand ( n38065 , n38055 , n38064 );
buf ( n38066 , n38065 );
buf ( n38067 , n38066 );
not ( n38068 , n38067 );
buf ( n38069 , n38068 );
buf ( n38070 , n38069 );
buf ( n38071 , n37900 );
not ( n38072 , n38071 );
buf ( n38073 , n3109 );
not ( n38074 , n38073 );
or ( n38075 , n38072 , n38074 );
buf ( n38076 , n1560 );
buf ( n38077 , n771 );
buf ( n38078 , n802 );
xor ( n38079 , n38077 , n38078 );
buf ( n38080 , n38079 );
buf ( n38081 , n38080 );
nand ( n38082 , n38076 , n38081 );
buf ( n38083 , n38082 );
buf ( n38084 , n38083 );
nand ( n38085 , n38075 , n38084 );
buf ( n38086 , n38085 );
buf ( n38087 , n38086 );
xor ( n38088 , n38070 , n38087 );
xor ( n38089 , n37921 , n37938 );
and ( n38090 , n38089 , n37956 );
and ( n38091 , n37921 , n37938 );
or ( n38092 , n38090 , n38091 );
buf ( n38093 , n38092 );
buf ( n38094 , n38093 );
xor ( n38095 , n38088 , n38094 );
buf ( n38096 , n38095 );
buf ( n38097 , n38096 );
xor ( n38098 , n38050 , n38097 );
buf ( n38099 , n38098 );
buf ( n38100 , n38099 );
xor ( n38101 , n38005 , n38100 );
xor ( n38102 , n37862 , n37910 );
and ( n38103 , n38102 , n37962 );
and ( n38104 , n37862 , n37910 );
or ( n38105 , n38103 , n38104 );
buf ( n38106 , n38105 );
buf ( n38107 , n38106 );
xor ( n38108 , n38101 , n38107 );
buf ( n38109 , n38108 );
buf ( n38110 , n38109 );
xor ( n38111 , n37856 , n37965 );
and ( n38112 , n38111 , n37972 );
and ( n38113 , n37856 , n37965 );
or ( n38114 , n38112 , n38113 );
buf ( n38115 , n38114 );
buf ( n38116 , n38115 );
xor ( n38117 , n38110 , n38116 );
buf ( n38118 , n38117 );
buf ( n38119 , n38118 );
nor ( n38120 , n37999 , n38119 );
buf ( n38121 , n38120 );
buf ( n38122 , n38121 );
not ( n38123 , n38122 );
buf ( n38124 , n38123 );
buf ( n38125 , n38124 );
and ( n38126 , n37996 , n38125 );
buf ( n38127 , n38126 );
not ( n38128 , n38127 );
or ( n38129 , n37763 , n38128 );
not ( n38130 , n31032 );
and ( n38131 , n31715 , n31113 );
and ( n38132 , n32140 , n37674 , n37689 );
not ( n38133 , n31167 );
and ( n38134 , n31080 , n38133 );
nand ( n38135 , n38130 , n38131 , n38132 , n38134 );
not ( n38136 , n38135 );
buf ( n38137 , n38136 );
buf ( n38138 , n38127 );
and ( n38139 , n38137 , n38138 );
buf ( n38140 , n38139 );
and ( n38141 , n31968 , n38140 );
buf ( n38142 , n38124 );
not ( n38143 , n38142 );
buf ( n38144 , n37992 );
not ( n38145 , n38144 );
buf ( n38146 , n38145 );
buf ( n38147 , n38146 );
not ( n38148 , n38147 );
buf ( n38149 , n37785 );
not ( n38150 , n38149 );
not ( n38151 , n37800 );
not ( n38152 , n17723 );
or ( n38153 , n38151 , n38152 );
not ( n38154 , n37804 );
nand ( n38155 , n38154 , n37792 , n37790 );
nand ( n38156 , n38153 , n38155 );
buf ( n38157 , n38156 );
not ( n38158 , n38157 );
or ( n38159 , n38150 , n38158 );
buf ( n38160 , n37775 );
not ( n38161 , n38160 );
buf ( n38162 , n38161 );
buf ( n38163 , n38162 );
buf ( n38164 , n17672 );
buf ( n38165 , n37779 );
and ( n38166 , n38164 , n38165 );
buf ( n38167 , n38166 );
buf ( n38168 , n38167 );
and ( n38169 , n38163 , n38168 );
buf ( n38170 , n37767 );
buf ( n38171 , n37772 );
and ( n38172 , n38170 , n38171 );
buf ( n38173 , n38172 );
buf ( n38174 , n38173 );
nor ( n38175 , n38169 , n38174 );
buf ( n38176 , n38175 );
buf ( n38177 , n38176 );
nand ( n38178 , n38159 , n38177 );
buf ( n38179 , n38178 );
buf ( n38180 , n38179 );
not ( n38181 , n38180 );
or ( n38182 , n38148 , n38181 );
buf ( n38183 , n37989 );
not ( n38184 , n38183 );
buf ( n38185 , n37833 );
not ( n38186 , n38185 );
buf ( n38187 , n37822 );
not ( n38188 , n38187 );
buf ( n38189 , n37813 );
nand ( n38190 , n38188 , n38189 );
buf ( n38191 , n38190 );
buf ( n38192 , n38191 );
not ( n38193 , n38192 );
buf ( n38194 , n38193 );
buf ( n38195 , n38194 );
not ( n38196 , n38195 );
or ( n38197 , n38186 , n38196 );
nand ( n38198 , n37830 , n37827 );
buf ( n38199 , n38198 );
nand ( n38200 , n38197 , n38199 );
buf ( n38201 , n38200 );
buf ( n38202 , n38201 );
not ( n38203 , n38202 );
or ( n38204 , n38184 , n38203 );
buf ( n38205 , n37838 );
buf ( n38206 , n37843 );
and ( n38207 , n38205 , n38206 );
buf ( n38208 , n38207 );
buf ( n38209 , n38208 );
buf ( n38210 , n37986 );
not ( n38211 , n38210 );
buf ( n38212 , n38211 );
buf ( n38213 , n38212 );
and ( n38214 , n38209 , n38213 );
buf ( n38215 , n37849 );
buf ( n38216 , n37983 );
and ( n38217 , n38215 , n38216 );
buf ( n38218 , n38217 );
buf ( n38219 , n38218 );
nor ( n38220 , n38214 , n38219 );
buf ( n38221 , n38220 );
buf ( n38222 , n38221 );
nand ( n38223 , n38204 , n38222 );
buf ( n38224 , n38223 );
buf ( n38225 , n38224 );
not ( n38226 , n38225 );
buf ( n38227 , n38226 );
buf ( n38228 , n38227 );
nand ( n38229 , n38182 , n38228 );
buf ( n38230 , n38229 );
buf ( n38231 , n38230 );
not ( n38232 , n38231 );
or ( n38233 , n38143 , n38232 );
buf ( n38234 , n37998 );
buf ( n38235 , n38118 );
and ( n38236 , n38234 , n38235 );
buf ( n38237 , n38236 );
buf ( n38238 , n38237 );
not ( n38239 , n38238 );
buf ( n38240 , n38239 );
buf ( n38241 , n38240 );
nand ( n38242 , n38233 , n38241 );
buf ( n38243 , n38242 );
nor ( n38244 , n38141 , n38243 );
nand ( n38245 , n38129 , n38244 );
not ( n38246 , n38245 );
and ( n38247 , n38110 , n38116 );
buf ( n38248 , n38247 );
buf ( n38249 , n38248 );
xor ( n38250 , n38005 , n38100 );
and ( n38251 , n38250 , n38107 );
and ( n38252 , n38005 , n38100 );
or ( n38253 , n38251 , n38252 );
buf ( n38254 , n38253 );
buf ( n38255 , n38254 );
xor ( n38256 , n38070 , n38087 );
and ( n38257 , n38256 , n38094 );
and ( n38258 , n38070 , n38087 );
or ( n38259 , n38257 , n38258 );
buf ( n38260 , n38259 );
buf ( n38261 , n38260 );
xor ( n38262 , n38043 , n38049 );
and ( n38263 , n38262 , n38097 );
and ( n38264 , n38043 , n38049 );
or ( n38265 , n38263 , n38264 );
buf ( n38266 , n38265 );
buf ( n38267 , n38266 );
xor ( n38268 , n38261 , n38267 );
xor ( n38269 , n38008 , n38026 );
and ( n38270 , n38269 , n38040 );
and ( n38271 , n38008 , n38026 );
or ( n38272 , n38270 , n38271 );
buf ( n38273 , n38272 );
buf ( n38274 , n38273 );
and ( n38275 , n37928 , n37929 );
buf ( n38276 , n38275 );
buf ( n38277 , n38276 );
buf ( n38278 , n38066 );
xor ( n38279 , n38277 , n38278 );
buf ( n38280 , n802 );
buf ( n38281 , n770 );
and ( n38282 , n38280 , n38281 );
not ( n38283 , n38280 );
buf ( n38284 , n770 );
not ( n38285 , n38284 );
buf ( n38286 , n38285 );
buf ( n38287 , n38286 );
and ( n38288 , n38283 , n38287 );
nor ( n38289 , n38282 , n38288 );
buf ( n38290 , n38289 );
buf ( n38291 , n38290 );
not ( n38292 , n38291 );
buf ( n38293 , n1560 );
not ( n38294 , n38293 );
or ( n38295 , n38292 , n38294 );
buf ( n38296 , n3109 );
buf ( n38297 , n38080 );
nand ( n38298 , n38296 , n38297 );
buf ( n38299 , n38298 );
buf ( n38300 , n38299 );
nand ( n38301 , n38295 , n38300 );
buf ( n38302 , n38301 );
buf ( n38303 , n38302 );
xor ( n38304 , n38279 , n38303 );
buf ( n38305 , n38304 );
buf ( n38306 , n38305 );
xor ( n38307 , n38274 , n38306 );
buf ( n38308 , n38060 );
not ( n38309 , n38308 );
buf ( n38310 , n15873 );
not ( n38311 , n38310 );
or ( n38312 , n38309 , n38311 );
buf ( n38313 , n804 );
buf ( n38314 , n768 );
xnor ( n38315 , n38313 , n38314 );
buf ( n38316 , n38315 );
buf ( n38317 , n38316 );
not ( n38318 , n38317 );
buf ( n38319 , n11137 );
nand ( n38320 , n38318 , n38319 );
buf ( n38321 , n38320 );
buf ( n38322 , n38321 );
nand ( n38323 , n38312 , n38322 );
buf ( n38324 , n38323 );
buf ( n38325 , n38324 );
buf ( n38326 , n14284 );
buf ( n38327 , n14278 );
or ( n38328 , n38326 , n38327 );
buf ( n38329 , n806 );
nand ( n38330 , n38328 , n38329 );
buf ( n38331 , n38330 );
buf ( n38332 , n38331 );
xor ( n38333 , n38325 , n38332 );
buf ( n38334 , n10509 );
not ( n38335 , n38334 );
buf ( n38336 , n38335 );
buf ( n38337 , n38336 );
buf ( n38338 , n38017 );
or ( n38339 , n38337 , n38338 );
buf ( n38340 , n3662 );
not ( n38341 , n38340 );
buf ( n38342 , n38341 );
buf ( n38343 , n38342 );
buf ( n38344 , n800 );
buf ( n38345 , n772 );
xor ( n38346 , n38344 , n38345 );
buf ( n38347 , n38346 );
buf ( n38348 , n38347 );
not ( n38349 , n38348 );
buf ( n38350 , n38349 );
buf ( n38351 , n38350 );
or ( n38352 , n38343 , n38351 );
nand ( n38353 , n38339 , n38352 );
buf ( n38354 , n38353 );
buf ( n38355 , n38354 );
xor ( n38356 , n38333 , n38355 );
buf ( n38357 , n38356 );
buf ( n38358 , n38357 );
xor ( n38359 , n38307 , n38358 );
buf ( n38360 , n38359 );
buf ( n38361 , n38360 );
xor ( n38362 , n38268 , n38361 );
buf ( n38363 , n38362 );
buf ( n38364 , n38363 );
xor ( n38365 , n38255 , n38364 );
buf ( n38366 , n38365 );
buf ( n38367 , n38366 );
nor ( n38368 , n38249 , n38367 );
buf ( n38369 , n38368 );
buf ( n38370 , n38369 );
not ( n38371 , n38370 );
buf ( n38372 , n38371 );
buf ( n38373 , n38372 );
buf ( n38374 , n38248 );
buf ( n38375 , n38366 );
nand ( n38376 , n38374 , n38375 );
buf ( n38377 , n38376 );
buf ( n38378 , n38377 );
nand ( n38379 , n38373 , n38378 );
buf ( n38380 , n38379 );
not ( n38381 , n38380 );
nor ( n38382 , n38381 , n831 );
nand ( n38383 , n38246 , n38382 );
buf ( n38384 , n37974 );
buf ( n38385 , n37980 );
and ( n38386 , n38384 , n38385 );
buf ( n38387 , n38386 );
buf ( n38388 , n38387 );
buf ( n38389 , n38109 );
buf ( n38390 , n38115 );
xor ( n38391 , n38389 , n38390 );
buf ( n38392 , n38391 );
buf ( n38393 , n38392 );
nor ( n38394 , n38388 , n38393 );
buf ( n38395 , n38394 );
buf ( n38396 , n38395 );
not ( n38397 , n38396 );
buf ( n38398 , n38397 );
not ( n38399 , n38398 );
buf ( n38400 , n18096 );
buf ( n38401 , n18363 );
xor ( n38402 , n37980 , n37974 );
buf ( n38403 , n38402 );
and ( n38404 , n18352 , n18358 );
buf ( n38405 , n38404 );
buf ( n38406 , n38405 );
nor ( n38407 , n38403 , n38406 );
buf ( n38408 , n38407 );
buf ( n38409 , n38408 );
nor ( n38410 , n38401 , n38409 );
buf ( n38411 , n38410 );
buf ( n38412 , n38411 );
nand ( n38413 , n38400 , n38412 );
buf ( n38414 , n38413 );
buf ( n38415 , n38414 );
not ( n38416 , n38415 );
buf ( n38417 , n38416 );
not ( n38418 , n38417 );
not ( n38419 , n18181 );
or ( n38420 , n38418 , n38419 );
buf ( n38421 , n38411 );
not ( n38422 , n38421 );
buf ( n38423 , n18209 );
not ( n38424 , n38423 );
or ( n38425 , n38422 , n38424 );
buf ( n38426 , n18370 );
buf ( n38427 , n38408 );
nor ( n38428 , n38426 , n38427 );
buf ( n38429 , n38428 );
buf ( n38430 , n38429 );
buf ( n38431 , n38405 );
buf ( n38432 , n38402 );
and ( n38433 , n38431 , n38432 );
buf ( n38434 , n38433 );
buf ( n38435 , n38434 );
nor ( n38436 , n38430 , n38435 );
buf ( n38437 , n38436 );
buf ( n38438 , n38437 );
nand ( n38439 , n38425 , n38438 );
buf ( n38440 , n38439 );
buf ( n38441 , n38440 );
not ( n38442 , n38441 );
buf ( n38443 , n38442 );
nand ( n38444 , n38420 , n38443 );
not ( n38445 , n38444 );
or ( n38446 , n38399 , n38445 );
buf ( n38447 , n38387 );
buf ( n38448 , n38392 );
nand ( n38449 , n38447 , n38448 );
buf ( n38450 , n38449 );
nand ( n38451 , n38446 , n38450 );
not ( n38452 , n38451 );
buf ( n38453 , n16833 );
buf ( n38454 , n17732 );
buf ( n38455 , n38414 );
nor ( n38456 , n38454 , n38455 );
buf ( n38457 , n38456 );
buf ( n38458 , n38457 );
buf ( n38459 , n38398 );
and ( n38460 , n38458 , n38459 );
buf ( n38461 , n38460 );
buf ( n38462 , n38461 );
nand ( n38463 , n38453 , n38462 );
buf ( n38464 , n38463 );
nand ( n38465 , n10417 , n18571 , n38461 );
nand ( n38466 , n38452 , n38464 , n38465 );
not ( n38467 , n38466 );
and ( n38468 , n38389 , n38390 );
buf ( n38469 , n38468 );
buf ( n38470 , n38469 );
buf ( n38471 , n38254 );
buf ( n38472 , n38363 );
xor ( n38473 , n38471 , n38472 );
buf ( n38474 , n38473 );
buf ( n38475 , n38474 );
nor ( n38476 , n38470 , n38475 );
buf ( n38477 , n38476 );
buf ( n38478 , n38477 );
not ( n38479 , n38478 );
buf ( n38480 , n38479 );
buf ( n38481 , n38480 );
buf ( n38482 , n38469 );
buf ( n38483 , n38474 );
nand ( n38484 , n38482 , n38483 );
buf ( n38485 , n38484 );
buf ( n38486 , n38485 );
nand ( n38487 , n38481 , n38486 );
buf ( n38488 , n38487 );
and ( n38489 , n38488 , n831 );
nand ( n38490 , n38467 , n38489 );
buf ( n38491 , n38488 );
not ( n38492 , n38491 );
buf ( n38493 , n38492 );
nand ( n38494 , n38466 , n38493 , n831 );
nor ( n38495 , n38380 , n831 );
nand ( n38496 , n38245 , n38495 );
nand ( n38497 , n38383 , n38490 , n38494 , n38496 );
not ( n38498 , n38497 );
buf ( n38499 , n38498 );
buf ( n38500 , n38499 );
buf ( n38501 , n3109 );
not ( n38502 , n38501 );
buf ( n38503 , n38502 );
buf ( n38504 , n38503 );
buf ( n38505 , n768 );
buf ( n38506 , n802 );
xnor ( n38507 , n38505 , n38506 );
buf ( n38508 , n38507 );
buf ( n38509 , n38508 );
or ( n38510 , n38504 , n38509 );
buf ( n38511 , n1560 );
not ( n38512 , n38511 );
buf ( n38513 , n38512 );
buf ( n38514 , n38513 );
buf ( n38515 , n802 );
not ( n38516 , n38515 );
buf ( n38517 , n38516 );
buf ( n38518 , n38517 );
or ( n38519 , n38514 , n38518 );
nand ( n38520 , n38510 , n38519 );
buf ( n38521 , n38520 );
buf ( n38522 , n38521 );
buf ( n38523 , n770 );
buf ( n38524 , n800 );
and ( n38525 , n38523 , n38524 );
buf ( n38526 , n38525 );
buf ( n38527 , n38526 );
buf ( n38528 , n38336 );
buf ( n38529 , n800 );
not ( n38530 , n38529 );
buf ( n38531 , n38530 );
buf ( n38532 , n38531 );
buf ( n38533 , n769 );
and ( n38534 , n38532 , n38533 );
buf ( n38535 , n11192 );
buf ( n38536 , n800 );
and ( n38537 , n38535 , n38536 );
nor ( n38538 , n38534 , n38537 );
buf ( n38539 , n38538 );
buf ( n38540 , n38539 );
or ( n38541 , n38528 , n38540 );
buf ( n38542 , n38342 );
buf ( n38543 , n38531 );
buf ( n38544 , n768 );
and ( n38545 , n38543 , n38544 );
buf ( n38546 , n37878 );
buf ( n38547 , n800 );
and ( n38548 , n38546 , n38547 );
nor ( n38549 , n38545 , n38548 );
buf ( n38550 , n38549 );
buf ( n38551 , n38550 );
or ( n38552 , n38542 , n38551 );
nand ( n38553 , n38541 , n38552 );
buf ( n38554 , n38553 );
buf ( n38555 , n38554 );
xor ( n38556 , n38527 , n38555 );
buf ( n38557 , n3109 );
buf ( n38558 , n1560 );
or ( n38559 , n38557 , n38558 );
buf ( n38560 , n802 );
nand ( n38561 , n38559 , n38560 );
buf ( n38562 , n38561 );
buf ( n38563 , n38562 );
xor ( n38564 , n38556 , n38563 );
buf ( n38565 , n38564 );
buf ( n38566 , n38565 );
xor ( n38567 , n38522 , n38566 );
buf ( n38568 , n771 );
buf ( n38569 , n800 );
and ( n38570 , n38568 , n38569 );
buf ( n38571 , n38570 );
buf ( n38572 , n38571 );
buf ( n38573 , n38336 );
buf ( n38574 , n38531 );
buf ( n38575 , n770 );
and ( n38576 , n38574 , n38575 );
buf ( n38577 , n38286 );
buf ( n38578 , n800 );
and ( n38579 , n38577 , n38578 );
nor ( n38580 , n38576 , n38579 );
buf ( n38581 , n38580 );
buf ( n38582 , n38581 );
or ( n38583 , n38573 , n38582 );
buf ( n38584 , n38342 );
buf ( n38585 , n38539 );
or ( n38586 , n38584 , n38585 );
nand ( n38587 , n38583 , n38586 );
buf ( n38588 , n38587 );
buf ( n38589 , n38588 );
xor ( n38590 , n38572 , n38589 );
buf ( n38591 , n38521 );
not ( n38592 , n38591 );
buf ( n38593 , n38592 );
buf ( n38594 , n38593 );
and ( n38595 , n38590 , n38594 );
and ( n38596 , n38572 , n38589 );
or ( n38597 , n38595 , n38596 );
buf ( n38598 , n38597 );
buf ( n38599 , n38598 );
xor ( n38600 , n38567 , n38599 );
buf ( n38601 , n38600 );
buf ( n38602 , n38601 );
and ( n38603 , n38344 , n38345 );
buf ( n38604 , n38603 );
buf ( n38605 , n38604 );
buf ( n38606 , n11137 );
not ( n38607 , n38606 );
buf ( n38608 , n38607 );
buf ( n38609 , n38608 );
not ( n38610 , n38609 );
buf ( n38611 , n15873 );
not ( n38612 , n38611 );
buf ( n38613 , n38612 );
buf ( n38614 , n38613 );
not ( n38615 , n38614 );
or ( n38616 , n38610 , n38615 );
buf ( n38617 , n804 );
nand ( n38618 , n38616 , n38617 );
buf ( n38619 , n38618 );
buf ( n38620 , n38619 );
xor ( n38621 , n38605 , n38620 );
buf ( n38622 , n38503 );
buf ( n38623 , n769 );
buf ( n38624 , n802 );
xnor ( n38625 , n38623 , n38624 );
buf ( n38626 , n38625 );
buf ( n38627 , n38626 );
or ( n38628 , n38622 , n38627 );
buf ( n38629 , n38513 );
buf ( n38630 , n38508 );
or ( n38631 , n38629 , n38630 );
nand ( n38632 , n38628 , n38631 );
buf ( n38633 , n38632 );
buf ( n38634 , n38633 );
and ( n38635 , n38621 , n38634 );
and ( n38636 , n38605 , n38620 );
or ( n38637 , n38635 , n38636 );
buf ( n38638 , n38637 );
buf ( n38639 , n38638 );
xor ( n38640 , n38572 , n38589 );
xor ( n38641 , n38640 , n38594 );
buf ( n38642 , n38641 );
buf ( n38643 , n38642 );
xor ( n38644 , n38639 , n38643 );
buf ( n38645 , n38613 );
buf ( n38646 , n38316 );
or ( n38647 , n38645 , n38646 );
buf ( n38648 , n38608 );
buf ( n38649 , n804 );
not ( n38650 , n38649 );
buf ( n38651 , n38650 );
buf ( n38652 , n38651 );
or ( n38653 , n38648 , n38652 );
nand ( n38654 , n38647 , n38653 );
buf ( n38655 , n38654 );
buf ( n38656 , n38655 );
buf ( n38657 , n38336 );
buf ( n38658 , n800 );
buf ( n38659 , n771 );
xnor ( n38660 , n38658 , n38659 );
buf ( n38661 , n38660 );
buf ( n38662 , n38661 );
or ( n38663 , n38657 , n38662 );
buf ( n38664 , n38342 );
buf ( n38665 , n38581 );
or ( n38666 , n38664 , n38665 );
nand ( n38667 , n38663 , n38666 );
buf ( n38668 , n38667 );
buf ( n38669 , n38668 );
xor ( n38670 , n38656 , n38669 );
buf ( n38671 , n773 );
buf ( n38672 , n800 );
and ( n38673 , n38671 , n38672 );
buf ( n38674 , n38673 );
buf ( n38675 , n38674 );
buf ( n38676 , n38347 );
not ( n38677 , n38676 );
buf ( n38678 , n10509 );
not ( n38679 , n38678 );
or ( n38680 , n38677 , n38679 );
buf ( n38681 , n38661 );
not ( n38682 , n38681 );
buf ( n38683 , n3662 );
nand ( n38684 , n38682 , n38683 );
buf ( n38685 , n38684 );
buf ( n38686 , n38685 );
nand ( n38687 , n38680 , n38686 );
buf ( n38688 , n38687 );
buf ( n38689 , n38688 );
xor ( n38690 , n38675 , n38689 );
buf ( n38691 , n38290 );
not ( n38692 , n38691 );
buf ( n38693 , n3109 );
not ( n38694 , n38693 );
or ( n38695 , n38692 , n38694 );
buf ( n38696 , n38626 );
not ( n38697 , n38696 );
buf ( n38698 , n1560 );
nand ( n38699 , n38697 , n38698 );
buf ( n38700 , n38699 );
buf ( n38701 , n38700 );
nand ( n38702 , n38695 , n38701 );
buf ( n38703 , n38702 );
buf ( n38704 , n38703 );
and ( n38705 , n38690 , n38704 );
and ( n38706 , n38675 , n38689 );
or ( n38707 , n38705 , n38706 );
buf ( n38708 , n38707 );
buf ( n38709 , n38708 );
and ( n38710 , n38670 , n38709 );
and ( n38711 , n38656 , n38669 );
or ( n38712 , n38710 , n38711 );
buf ( n38713 , n38712 );
buf ( n38714 , n38713 );
and ( n38715 , n38644 , n38714 );
and ( n38716 , n38639 , n38643 );
or ( n38717 , n38715 , n38716 );
buf ( n38718 , n38717 );
buf ( n38719 , n38718 );
and ( n38720 , n38602 , n38719 );
buf ( n38721 , n38720 );
buf ( n38722 , n38721 );
buf ( n38723 , n769 );
buf ( n38724 , n800 );
nand ( n38725 , n38723 , n38724 );
buf ( n38726 , n38725 );
buf ( n38727 , n38726 );
buf ( n38728 , n38336 );
buf ( n38729 , n38550 );
or ( n38730 , n38728 , n38729 );
buf ( n38731 , n38342 );
buf ( n38732 , n38531 );
or ( n38733 , n38731 , n38732 );
nand ( n38734 , n38730 , n38733 );
buf ( n38735 , n38734 );
buf ( n38736 , n38735 );
xor ( n38737 , n38727 , n38736 );
xor ( n38738 , n38527 , n38555 );
and ( n38739 , n38738 , n38563 );
and ( n38740 , n38527 , n38555 );
or ( n38741 , n38739 , n38740 );
buf ( n38742 , n38741 );
buf ( n38743 , n38742 );
xor ( n38744 , n38737 , n38743 );
buf ( n38745 , n38744 );
buf ( n38746 , n38745 );
xor ( n38747 , n38522 , n38566 );
and ( n38748 , n38747 , n38599 );
and ( n38749 , n38522 , n38566 );
or ( n38750 , n38748 , n38749 );
buf ( n38751 , n38750 );
buf ( n38752 , n38751 );
xor ( n38753 , n38746 , n38752 );
buf ( n38754 , n38753 );
buf ( n38755 , n38754 );
and ( n38756 , n38722 , n38755 );
buf ( n38757 , n38756 );
buf ( n38758 , n38757 );
not ( n38759 , n38758 );
buf ( n38760 , n38721 );
buf ( n38761 , n38754 );
or ( n38762 , n38760 , n38761 );
buf ( n38763 , n38762 );
buf ( n38764 , n38763 );
nand ( n38765 , n38759 , n38764 );
buf ( n38766 , n38765 );
not ( n38767 , n38766 );
buf ( n38768 , n10417 );
buf ( n38769 , n38768 );
buf ( n38770 , n38769 );
buf ( n38771 , n38770 );
buf ( n38772 , n18136 );
buf ( n38773 , n38457 );
buf ( n38774 , n38773 );
buf ( n38775 , n38774 );
buf ( n38776 , n38775 );
xor ( n38777 , n38605 , n38620 );
xor ( n38778 , n38777 , n38634 );
buf ( n38779 , n38778 );
buf ( n38780 , n38779 );
xor ( n38781 , n38656 , n38669 );
xor ( n38782 , n38781 , n38709 );
buf ( n38783 , n38782 );
buf ( n38784 , n38783 );
xor ( n38785 , n38780 , n38784 );
buf ( n38786 , n38655 );
not ( n38787 , n38786 );
buf ( n38788 , n38787 );
buf ( n38789 , n38788 );
xor ( n38790 , n38675 , n38689 );
xor ( n38791 , n38790 , n38704 );
buf ( n38792 , n38791 );
buf ( n38793 , n38792 );
xor ( n38794 , n38789 , n38793 );
xor ( n38795 , n38325 , n38332 );
and ( n38796 , n38795 , n38355 );
and ( n38797 , n38325 , n38332 );
or ( n38798 , n38796 , n38797 );
buf ( n38799 , n38798 );
buf ( n38800 , n38799 );
and ( n38801 , n38794 , n38800 );
and ( n38802 , n38789 , n38793 );
or ( n38803 , n38801 , n38802 );
buf ( n38804 , n38803 );
buf ( n38805 , n38804 );
xor ( n38806 , n38785 , n38805 );
buf ( n38807 , n38806 );
buf ( n38808 , n38807 );
xor ( n38809 , n38277 , n38278 );
and ( n38810 , n38809 , n38303 );
and ( n38811 , n38277 , n38278 );
or ( n38812 , n38810 , n38811 );
buf ( n38813 , n38812 );
buf ( n38814 , n38813 );
xor ( n38815 , n38789 , n38793 );
xor ( n38816 , n38815 , n38800 );
buf ( n38817 , n38816 );
buf ( n38818 , n38817 );
xor ( n38819 , n38814 , n38818 );
xor ( n38820 , n38274 , n38306 );
and ( n38821 , n38820 , n38358 );
and ( n38822 , n38274 , n38306 );
or ( n38823 , n38821 , n38822 );
buf ( n38824 , n38823 );
buf ( n38825 , n38824 );
and ( n38826 , n38819 , n38825 );
and ( n38827 , n38814 , n38818 );
or ( n38828 , n38826 , n38827 );
buf ( n38829 , n38828 );
buf ( n38830 , n38829 );
and ( n38831 , n38808 , n38830 );
buf ( n38832 , n38831 );
buf ( n38833 , n38832 );
xor ( n38834 , n38639 , n38643 );
xor ( n38835 , n38834 , n38714 );
buf ( n38836 , n38835 );
buf ( n38837 , n38836 );
xor ( n38838 , n38780 , n38784 );
and ( n38839 , n38838 , n38805 );
and ( n38840 , n38780 , n38784 );
or ( n38841 , n38839 , n38840 );
buf ( n38842 , n38841 );
buf ( n38843 , n38842 );
xor ( n38844 , n38837 , n38843 );
buf ( n38845 , n38844 );
buf ( n38846 , n38845 );
nor ( n38847 , n38833 , n38846 );
buf ( n38848 , n38847 );
buf ( n38849 , n38848 );
and ( n38850 , n38837 , n38843 );
buf ( n38851 , n38850 );
buf ( n38852 , n38851 );
xor ( n38853 , n38602 , n38719 );
buf ( n38854 , n38853 );
buf ( n38855 , n38854 );
nor ( n38856 , n38852 , n38855 );
buf ( n38857 , n38856 );
buf ( n38858 , n38857 );
nor ( n38859 , n38849 , n38858 );
buf ( n38860 , n38859 );
buf ( n38861 , n38860 );
not ( n38862 , n38861 );
xor ( n38863 , n38814 , n38818 );
xor ( n38864 , n38863 , n38825 );
buf ( n38865 , n38864 );
buf ( n38866 , n38865 );
xor ( n38867 , n38261 , n38267 );
and ( n38868 , n38867 , n38361 );
and ( n38869 , n38261 , n38267 );
or ( n38870 , n38868 , n38869 );
buf ( n38871 , n38870 );
buf ( n38872 , n38871 );
xor ( n38873 , n38866 , n38872 );
buf ( n38874 , n38873 );
buf ( n38875 , n38874 );
and ( n38876 , n38471 , n38472 );
buf ( n38877 , n38876 );
buf ( n38878 , n38877 );
nor ( n38879 , n38875 , n38878 );
buf ( n38880 , n38879 );
buf ( n38881 , n38880 );
and ( n38882 , n38866 , n38872 );
buf ( n38883 , n38882 );
buf ( n38884 , n38883 );
xor ( n38885 , n38808 , n38830 );
buf ( n38886 , n38885 );
buf ( n38887 , n38886 );
nor ( n38888 , n38884 , n38887 );
buf ( n38889 , n38888 );
buf ( n38890 , n38889 );
nor ( n38891 , n38881 , n38890 );
buf ( n38892 , n38891 );
buf ( n38893 , n38477 );
buf ( n38894 , n38395 );
nor ( n38895 , n38893 , n38894 );
buf ( n38896 , n38895 );
nand ( n38897 , n38892 , n38896 );
buf ( n38898 , n38897 );
nor ( n38899 , n38862 , n38898 );
buf ( n38900 , n38899 );
buf ( n38901 , n38900 );
nand ( n38902 , n38776 , n38901 );
buf ( n38903 , n38902 );
buf ( n38904 , n38903 );
nor ( n38905 , n38772 , n38904 );
buf ( n38906 , n38905 );
buf ( n38907 , n38906 );
nand ( n38908 , n38771 , n38907 );
buf ( n38909 , n38908 );
not ( n38910 , n38903 );
nand ( n38911 , n38910 , n18585 );
buf ( n38912 , n38900 );
not ( n38913 , n38912 );
buf ( n38914 , n38444 );
not ( n38915 , n38914 );
or ( n38916 , n38913 , n38915 );
not ( n38917 , n38892 );
buf ( n38918 , n38480 );
not ( n38919 , n38918 );
buf ( n38920 , n38450 );
not ( n38921 , n38920 );
buf ( n38922 , n38921 );
buf ( n38923 , n38922 );
not ( n38924 , n38923 );
or ( n38925 , n38919 , n38924 );
buf ( n38926 , n38485 );
nand ( n38927 , n38925 , n38926 );
buf ( n38928 , n38927 );
not ( n38929 , n38928 );
or ( n38930 , n38917 , n38929 );
buf ( n38931 , n38874 );
buf ( n38932 , n38877 );
and ( n38933 , n38931 , n38932 );
buf ( n38934 , n38933 );
buf ( n38935 , n38934 );
buf ( n38936 , n38889 );
not ( n38937 , n38936 );
buf ( n38938 , n38937 );
buf ( n38939 , n38938 );
and ( n38940 , n38935 , n38939 );
buf ( n38941 , n38883 );
buf ( n38942 , n38886 );
nand ( n38943 , n38941 , n38942 );
buf ( n38944 , n38943 );
buf ( n38945 , n38944 );
not ( n38946 , n38945 );
buf ( n38947 , n38946 );
buf ( n38948 , n38947 );
nor ( n38949 , n38940 , n38948 );
buf ( n38950 , n38949 );
nand ( n38951 , n38930 , n38950 );
and ( n38952 , n38860 , n38951 );
buf ( n38953 , n38832 );
buf ( n38954 , n38845 );
nand ( n38955 , n38953 , n38954 );
buf ( n38956 , n38955 );
buf ( n38957 , n38956 );
buf ( n38958 , n38857 );
or ( n38959 , n38957 , n38958 );
buf ( n38960 , n38851 );
buf ( n38961 , n38854 );
nand ( n38962 , n38960 , n38961 );
buf ( n38963 , n38962 );
buf ( n38964 , n38963 );
nand ( n38965 , n38959 , n38964 );
buf ( n38966 , n38965 );
nor ( n38967 , n38952 , n38966 );
buf ( n38968 , n38967 );
nand ( n38969 , n38916 , n38968 );
buf ( n38970 , n38969 );
buf ( n38971 , n38970 );
not ( n38972 , n38971 );
buf ( n38973 , n38972 );
nand ( n38974 , n38909 , n38911 , n38973 );
not ( n38975 , n38974 );
or ( n38976 , n38767 , n38975 );
not ( n38977 , n38766 );
and ( n38978 , n38973 , n38977 );
nand ( n38979 , n38978 , n38909 , n38911 );
nand ( n38980 , n38976 , n38979 );
nor ( n38981 , n38500 , n38980 );
buf ( n38982 , n38444 );
buf ( n38983 , n38982 );
buf ( n38984 , n38983 );
not ( n38985 , n38984 );
buf ( n38986 , n18571 );
buf ( n38987 , n38775 );
and ( n38988 , n38986 , n38987 );
buf ( n38989 , n38988 );
nand ( n38990 , n10430 , n38989 );
buf ( n38991 , n18585 );
buf ( n38992 , n38775 );
nand ( n38993 , n38991 , n38992 );
buf ( n38994 , n38993 );
nand ( n38995 , n38985 , n38990 , n38994 );
buf ( n38996 , n38398 );
buf ( n38997 , n38450 );
nand ( n38998 , n38996 , n38997 );
buf ( n38999 , n38998 );
buf ( n39000 , n38999 );
not ( n39001 , n39000 );
buf ( n39002 , n39001 );
and ( n39003 , n39002 , n831 );
and ( n39004 , n38995 , n39003 );
not ( n39005 , n38995 );
and ( n39006 , n38999 , n831 );
and ( n39007 , n39005 , n39006 );
nor ( n39008 , n39004 , n39007 );
buf ( n39009 , n37759 );
not ( n39010 , n39009 );
buf ( n39011 , n39010 );
buf ( n39012 , n39011 );
buf ( n39013 , n37995 );
buf ( n39014 , n39013 );
buf ( n39015 , n39014 );
buf ( n39016 , n39015 );
nand ( n39017 , n39012 , n39016 );
buf ( n39018 , n39017 );
not ( n39019 , n39018 );
buf ( n39020 , n38124 );
buf ( n39021 , n38240 );
nand ( n39022 , n39020 , n39021 );
buf ( n39023 , n39022 );
nand ( n39024 , n39019 , n39023 );
buf ( n39025 , n31968 );
buf ( n39026 , n38136 );
buf ( n39027 , n39015 );
and ( n39028 , n39026 , n39027 );
buf ( n39029 , n39028 );
buf ( n39030 , n39029 );
nand ( n39031 , n39025 , n39030 );
buf ( n39032 , n39031 );
not ( n39033 , n39032 );
nand ( n39034 , n39033 , n39023 );
buf ( n39035 , n38146 );
not ( n39036 , n39035 );
buf ( n39037 , n38179 );
not ( n39038 , n39037 );
or ( n39039 , n39036 , n39038 );
buf ( n39040 , n38227 );
nand ( n39041 , n39039 , n39040 );
buf ( n39042 , n39041 );
buf ( n39043 , n39042 );
not ( n39044 , n39043 );
buf ( n39045 , n39044 );
buf ( n39046 , n39023 );
not ( n39047 , n39046 );
buf ( n39048 , n39047 );
and ( n39049 , n39045 , n39048 );
nand ( n39050 , n39018 , n39032 , n39049 );
or ( n39051 , n39045 , n39048 );
and ( n39052 , n39051 , n2206 );
nand ( n39053 , n39024 , n39034 , n39050 , n39052 );
nand ( n39054 , n39008 , n39053 );
not ( n39055 , n39054 );
buf ( n39056 , n39055 );
buf ( n39057 , n18136 );
buf ( n39058 , n38775 );
buf ( n39059 , n38897 );
buf ( n39060 , n38848 );
nor ( n39061 , n39059 , n39060 );
buf ( n39062 , n39061 );
buf ( n39063 , n39062 );
nand ( n39064 , n39058 , n39063 );
buf ( n39065 , n39064 );
buf ( n39066 , n39065 );
nor ( n39067 , n39057 , n39066 );
buf ( n39068 , n39067 );
nand ( n39069 , n39068 , n38770 );
buf ( n39070 , n39065 );
not ( n39071 , n39070 );
buf ( n39072 , n18585 );
nand ( n39073 , n39071 , n39072 );
buf ( n39074 , n39073 );
buf ( n39075 , n39062 );
buf ( n39076 , n38444 );
and ( n39077 , n39075 , n39076 );
buf ( n39078 , n38848 );
not ( n39079 , n39078 );
buf ( n39080 , n39079 );
buf ( n39081 , n39080 );
not ( n39082 , n39081 );
buf ( n39083 , n38951 );
not ( n39084 , n39083 );
or ( n39085 , n39082 , n39084 );
buf ( n39086 , n38956 );
nand ( n39087 , n39085 , n39086 );
buf ( n39088 , n39087 );
buf ( n39089 , n39088 );
nor ( n39090 , n39077 , n39089 );
buf ( n39091 , n39090 );
nand ( n39092 , n39069 , n39074 , n39091 );
not ( n39093 , n38857 );
nand ( n39094 , n39093 , n38963 );
not ( n39095 , n39094 );
and ( n39096 , n39092 , n39095 );
not ( n39097 , n39092 );
and ( n39098 , n39097 , n39094 );
nor ( n39099 , n39096 , n39098 );
nor ( n39100 , n39056 , n39099 );
nor ( n39101 , n38981 , n39100 );
not ( n39102 , n39101 );
not ( n39103 , n831 );
buf ( n39104 , n38457 );
buf ( n39105 , n38896 );
not ( n39106 , n39105 );
buf ( n39107 , n39106 );
buf ( n39108 , n39107 );
buf ( n39109 , n38880 );
nor ( n39110 , n39108 , n39109 );
buf ( n39111 , n39110 );
buf ( n39112 , n39111 );
and ( n39113 , n39104 , n39112 );
buf ( n39114 , n39113 );
nand ( n39115 , n10417 , n18571 , n39114 );
buf ( n39116 , n39115 );
buf ( n39117 , n18585 );
buf ( n39118 , n39114 );
nand ( n39119 , n39117 , n39118 );
buf ( n39120 , n39119 );
buf ( n39121 , n39120 );
buf ( n39122 , n39111 );
not ( n39123 , n39122 );
buf ( n39124 , n38444 );
not ( n39125 , n39124 );
or ( n39126 , n39123 , n39125 );
buf ( n39127 , n38928 );
buf ( n39128 , n38880 );
not ( n39129 , n39128 );
buf ( n39130 , n39129 );
buf ( n39131 , n39130 );
and ( n39132 , n39127 , n39131 );
buf ( n39133 , n38934 );
nor ( n39134 , n39132 , n39133 );
buf ( n39135 , n39134 );
buf ( n39136 , n39135 );
nand ( n39137 , n39126 , n39136 );
buf ( n39138 , n39137 );
buf ( n39139 , n39138 );
not ( n39140 , n39139 );
buf ( n39141 , n39140 );
buf ( n39142 , n39141 );
nand ( n39143 , n39116 , n39121 , n39142 );
buf ( n39144 , n39143 );
buf ( n39145 , n38938 );
buf ( n39146 , n38944 );
nand ( n39147 , n39145 , n39146 );
buf ( n39148 , n39147 );
buf ( n39149 , n39148 );
not ( n39150 , n39149 );
buf ( n39151 , n39150 );
and ( n39152 , n39144 , n39151 );
not ( n39153 , n39144 );
and ( n39154 , n39153 , n39148 );
nor ( n39155 , n39152 , n39154 );
not ( n39156 , n39155 );
or ( n39157 , n39103 , n39156 );
buf ( n39158 , n38865 );
buf ( n39159 , n38871 );
and ( n39160 , n39158 , n39159 );
buf ( n39161 , n39160 );
buf ( n39162 , n39161 );
buf ( n39163 , n38807 );
buf ( n39164 , n38829 );
xor ( n39165 , n39163 , n39164 );
buf ( n39166 , n39165 );
buf ( n39167 , n39166 );
nor ( n39168 , n39162 , n39167 );
buf ( n39169 , n39168 );
buf ( n39170 , n39169 );
not ( n39171 , n39170 );
buf ( n39172 , n39171 );
buf ( n39173 , n39172 );
buf ( n39174 , n39161 );
buf ( n39175 , n39166 );
nand ( n39176 , n39174 , n39175 );
buf ( n39177 , n39176 );
buf ( n39178 , n39177 );
nand ( n39179 , n39173 , n39178 );
buf ( n39180 , n39179 );
not ( n39181 , n39180 );
buf ( n39182 , n38369 );
buf ( n39183 , n38121 );
nor ( n39184 , n39182 , n39183 );
buf ( n39185 , n39184 );
buf ( n39186 , n39185 );
not ( n39187 , n39186 );
buf ( n39188 , n39187 );
buf ( n39189 , n39188 );
xor ( n39190 , n39158 , n39159 );
buf ( n39191 , n39190 );
buf ( n39192 , n39191 );
and ( n39193 , n38255 , n38364 );
buf ( n39194 , n39193 );
buf ( n39195 , n39194 );
nor ( n39196 , n39192 , n39195 );
buf ( n39197 , n39196 );
buf ( n39198 , n39197 );
nor ( n39199 , n39189 , n39198 );
buf ( n39200 , n39199 );
buf ( n39201 , n39200 );
not ( n39202 , n39201 );
buf ( n39203 , n38230 );
not ( n39204 , n39203 );
or ( n39205 , n39202 , n39204 );
buf ( n39206 , n38372 );
not ( n39207 , n39206 );
buf ( n39208 , n38237 );
not ( n39209 , n39208 );
or ( n39210 , n39207 , n39209 );
buf ( n39211 , n38377 );
nand ( n39212 , n39210 , n39211 );
buf ( n39213 , n39212 );
buf ( n39214 , n39213 );
buf ( n39215 , n39197 );
not ( n39216 , n39215 );
buf ( n39217 , n39216 );
buf ( n39218 , n39217 );
and ( n39219 , n39214 , n39218 );
buf ( n39220 , n39191 );
buf ( n39221 , n39194 );
and ( n39222 , n39220 , n39221 );
buf ( n39223 , n39222 );
buf ( n39224 , n39223 );
nor ( n39225 , n39219 , n39224 );
buf ( n39226 , n39225 );
buf ( n39227 , n39226 );
nand ( n39228 , n39205 , n39227 );
buf ( n39229 , n39228 );
not ( n39230 , n39229 );
buf ( n39231 , n37759 );
not ( n39232 , n39231 );
buf ( n39233 , n39232 );
buf ( n39234 , n39233 );
buf ( n39235 , n37995 );
buf ( n39236 , n39200 );
and ( n39237 , n39235 , n39236 );
buf ( n39238 , n39237 );
buf ( n39239 , n39238 );
nand ( n39240 , n39234 , n39239 );
buf ( n39241 , n39240 );
not ( n39242 , n38135 );
nand ( n39243 , n31968 , n39242 , n39238 );
nand ( n39244 , n39230 , n39241 , n39243 );
not ( n39245 , n39244 );
or ( n39246 , n39181 , n39245 );
not ( n39247 , n39229 );
not ( n39248 , n39180 );
nand ( n39249 , n39241 , n39247 , n39243 , n39248 );
nand ( n39250 , n39246 , n39249 );
nand ( n39251 , n39250 , n1152 );
nand ( n39252 , n39157 , n39251 );
buf ( n39253 , n39252 );
not ( n39254 , n39253 );
not ( n39255 , n39254 );
buf ( n39256 , n16833 );
buf ( n39257 , n39107 );
not ( n39258 , n39257 );
buf ( n39259 , n38775 );
nand ( n39260 , n39258 , n39259 );
buf ( n39261 , n39260 );
buf ( n39262 , n39261 );
not ( n39263 , n39262 );
buf ( n39264 , n39263 );
buf ( n39265 , n39264 );
nand ( n39266 , n39256 , n39265 );
buf ( n39267 , n39266 );
buf ( n39268 , n10417 );
buf ( n39269 , n18136 );
buf ( n39270 , n39261 );
nor ( n39271 , n39269 , n39270 );
buf ( n39272 , n39271 );
buf ( n39273 , n39272 );
nand ( n39274 , n39268 , n39273 );
buf ( n39275 , n39274 );
and ( n39276 , n38896 , n38444 );
nor ( n39277 , n39276 , n38928 );
nand ( n39278 , n39267 , n39275 , n39277 );
buf ( n39279 , n38934 );
buf ( n39280 , n38880 );
nor ( n39281 , n39279 , n39280 );
buf ( n39282 , n39281 );
xor ( n39283 , n39278 , n39282 );
not ( n39284 , n831 );
or ( n39285 , n39283 , n39284 );
buf ( n39286 , n39185 );
not ( n39287 , n39286 );
buf ( n39288 , n39042 );
not ( n39289 , n39288 );
or ( n39290 , n39287 , n39289 );
buf ( n39291 , n39213 );
not ( n39292 , n39291 );
buf ( n39293 , n39292 );
buf ( n39294 , n39293 );
nand ( n39295 , n39290 , n39294 );
buf ( n39296 , n39295 );
buf ( n39297 , n39296 );
not ( n39298 , n39297 );
buf ( n39299 , n39298 );
nor ( n39300 , n39223 , n39197 );
not ( n39301 , n39300 );
nand ( n39302 , n39301 , n39284 );
and ( n39303 , n39299 , n39302 );
buf ( n39304 , n39188 );
not ( n39305 , n39304 );
buf ( n39306 , n39015 );
nand ( n39307 , n39305 , n39306 );
buf ( n39308 , n39307 );
not ( n39309 , n39308 );
nand ( n39310 , n39309 , n39011 );
buf ( n39311 , n31968 );
buf ( n39312 , n39242 );
not ( n39313 , n39312 );
buf ( n39314 , n39308 );
nor ( n39315 , n39313 , n39314 );
buf ( n39316 , n39315 );
buf ( n39317 , n39316 );
nand ( n39318 , n39311 , n39317 );
buf ( n39319 , n39318 );
nand ( n39320 , n39303 , n39310 , n39319 );
not ( n39321 , n39310 );
nand ( n39322 , n39300 , n39284 );
nand ( n39323 , n39321 , n39322 );
not ( n39324 , n39299 );
not ( n39325 , n39319 );
or ( n39326 , n39324 , n39325 );
nand ( n39327 , n39326 , n39322 );
nand ( n39328 , n39320 , n39323 , n39327 );
nand ( n39329 , n39285 , n39328 );
not ( n39330 , n39329 );
not ( n39331 , n39330 );
not ( n39332 , n39331 );
not ( n39333 , n39332 );
buf ( n39334 , n39333 );
not ( n39335 , n39334 );
and ( n39336 , n38746 , n38752 );
buf ( n39337 , n39336 );
buf ( n39338 , n39337 );
not ( n39339 , n39338 );
xor ( n39340 , n38727 , n38736 );
and ( n39341 , n39340 , n38743 );
and ( n39342 , n38727 , n38736 );
or ( n39343 , n39341 , n39342 );
buf ( n39344 , n39343 );
buf ( n39345 , n39344 );
buf ( n39346 , n38726 );
not ( n39347 , n39346 );
buf ( n39348 , n768 );
buf ( n39349 , n800 );
nand ( n39350 , n39348 , n39349 );
buf ( n39351 , n39350 );
buf ( n39352 , n39351 );
not ( n39353 , n39352 );
buf ( n39354 , n10509 );
buf ( n39355 , n3662 );
or ( n39356 , n39354 , n39355 );
buf ( n39357 , n800 );
nand ( n39358 , n39356 , n39357 );
buf ( n39359 , n39358 );
buf ( n39360 , n39359 );
not ( n39361 , n39360 );
or ( n39362 , n39353 , n39361 );
buf ( n39363 , n39359 );
buf ( n39364 , n39351 );
or ( n39365 , n39363 , n39364 );
nand ( n39366 , n39362 , n39365 );
buf ( n39367 , n39366 );
buf ( n39368 , n39367 );
not ( n39369 , n39368 );
or ( n39370 , n39347 , n39369 );
buf ( n39371 , n39367 );
buf ( n39372 , n38726 );
or ( n39373 , n39371 , n39372 );
nand ( n39374 , n39370 , n39373 );
buf ( n39375 , n39374 );
buf ( n39376 , n39375 );
xor ( n39377 , n39345 , n39376 );
buf ( n39378 , n39377 );
buf ( n39379 , n39378 );
not ( n39380 , n39379 );
and ( n39381 , n39339 , n39380 );
buf ( n39382 , n39337 );
buf ( n39383 , n39378 );
and ( n39384 , n39382 , n39383 );
nor ( n39385 , n39381 , n39384 );
buf ( n39386 , n39385 );
not ( n39387 , n39386 );
not ( n39388 , n39387 );
buf ( n39389 , n38770 );
buf ( n39390 , n18136 );
buf ( n39391 , n38775 );
buf ( n39392 , n38897 );
buf ( n39393 , n38860 );
buf ( n39394 , n38763 );
nand ( n39395 , n39393 , n39394 );
buf ( n39396 , n39395 );
buf ( n39397 , n39396 );
nor ( n39398 , n39392 , n39397 );
buf ( n39399 , n39398 );
buf ( n39400 , n39399 );
nand ( n39401 , n39391 , n39400 );
buf ( n39402 , n39401 );
buf ( n39403 , n39402 );
nor ( n39404 , n39390 , n39403 );
buf ( n39405 , n39404 );
buf ( n39406 , n39405 );
nand ( n39407 , n39389 , n39406 );
buf ( n39408 , n39407 );
buf ( n39409 , n39399 );
not ( n39410 , n39409 );
buf ( n39411 , n38984 );
not ( n39412 , n39411 );
or ( n39413 , n39410 , n39412 );
buf ( n39414 , n39396 );
not ( n39415 , n39414 );
buf ( n39416 , n39415 );
and ( n39417 , n39416 , n38951 );
and ( n39418 , n38966 , n38763 );
nor ( n39419 , n39417 , n39418 , n38757 );
buf ( n39420 , n39419 );
nand ( n39421 , n39413 , n39420 );
buf ( n39422 , n39421 );
buf ( n39423 , n39422 );
not ( n39424 , n39423 );
buf ( n39425 , n39424 );
not ( n39426 , n39402 );
nand ( n39427 , n39426 , n16833 );
nand ( n39428 , n39408 , n39425 , n39427 );
not ( n39429 , n39428 );
or ( n39430 , n39388 , n39429 );
nand ( n39431 , n39408 , n39425 , n39427 , n39386 );
nand ( n39432 , n39430 , n39431 );
buf ( n39433 , n39432 );
or ( n39434 , n39335 , n39433 );
nand ( n39435 , n39255 , n39434 );
nor ( n39436 , n39102 , n39435 );
not ( n39437 , n39436 );
buf ( n39438 , n38136 );
not ( n39439 , n39438 );
buf ( n39440 , n39439 );
buf ( n39441 , n39440 );
buf ( n39442 , n37810 );
buf ( n39443 , n39442 );
buf ( n39444 , n39443 );
buf ( n39445 , n39444 );
not ( n39446 , n39445 );
buf ( n39447 , n39446 );
buf ( n39448 , n39447 );
buf ( n39449 , n37836 );
not ( n39450 , n39449 );
buf ( n39451 , n37846 );
nor ( n39452 , n39450 , n39451 );
buf ( n39453 , n39452 );
buf ( n39454 , n39453 );
nand ( n39455 , n39448 , n39454 );
buf ( n39456 , n39455 );
buf ( n39457 , n39456 );
nor ( n39458 , n39441 , n39457 );
buf ( n39459 , n39458 );
buf ( n39460 , n39459 );
not ( n39461 , n39460 );
buf ( n39462 , n31968 );
not ( n39463 , n39462 );
or ( n39464 , n39461 , n39463 );
buf ( n39465 , n39453 );
not ( n39466 , n39465 );
buf ( n39467 , n38179 );
buf ( n39468 , n39467 );
buf ( n39469 , n39468 );
buf ( n39470 , n39469 );
not ( n39471 , n39470 );
or ( n39472 , n39466 , n39471 );
buf ( n39473 , n38201 );
buf ( n39474 , n37846 );
not ( n39475 , n39474 );
buf ( n39476 , n39475 );
buf ( n39477 , n39476 );
and ( n39478 , n39473 , n39477 );
buf ( n39479 , n38208 );
nor ( n39480 , n39478 , n39479 );
buf ( n39481 , n39480 );
buf ( n39482 , n39481 );
nand ( n39483 , n39472 , n39482 );
buf ( n39484 , n39483 );
buf ( n39485 , n39484 );
not ( n39486 , n39485 );
buf ( n39487 , n39486 );
buf ( n39488 , n39487 );
nand ( n39489 , n39464 , n39488 );
buf ( n39490 , n39489 );
not ( n39491 , n39490 );
buf ( n39492 , n38218 );
not ( n39493 , n39492 );
buf ( n39494 , n38212 );
nand ( n39495 , n39493 , n39494 );
buf ( n39496 , n39495 );
buf ( n39497 , n1152 );
and ( n39498 , n39496 , n39497 );
nor ( n39499 , n37759 , n39456 );
nor ( n39500 , n39498 , n39499 );
nand ( n39501 , n39491 , n39500 );
not ( n39502 , n39501 );
or ( n39503 , n39490 , n39499 );
not ( n39504 , n39496 );
nand ( n39505 , n39504 , n39497 );
nand ( n39506 , n39503 , n39505 );
not ( n39507 , n39506 );
or ( n39508 , n39502 , n39507 );
buf ( n39509 , n17735 );
buf ( n39510 , n18096 );
buf ( n39511 , n18366 );
nand ( n39512 , n39510 , n39511 );
buf ( n39513 , n39512 );
buf ( n39514 , n39513 );
nor ( n39515 , n39509 , n39514 );
buf ( n39516 , n39515 );
buf ( n39517 , n39516 );
not ( n39518 , n39517 );
buf ( n39519 , n18585 );
not ( n39520 , n39519 );
or ( n39521 , n39518 , n39520 );
buf ( n39522 , n10417 );
buf ( n39523 , n18571 );
buf ( n39524 , n39516 );
and ( n39525 , n39523 , n39524 );
buf ( n39526 , n39525 );
buf ( n39527 , n39526 );
and ( n39528 , n39522 , n39527 );
buf ( n39529 , n39513 );
not ( n39530 , n39529 );
buf ( n39531 , n39530 );
buf ( n39532 , n39531 );
not ( n39533 , n39532 );
buf ( n39534 , n18184 );
not ( n39535 , n39534 );
or ( n39536 , n39533 , n39535 );
buf ( n39537 , n18366 );
not ( n39538 , n39537 );
buf ( n39539 , n18209 );
not ( n39540 , n39539 );
or ( n39541 , n39538 , n39540 );
buf ( n39542 , n18370 );
nand ( n39543 , n39541 , n39542 );
buf ( n39544 , n39543 );
buf ( n39545 , n39544 );
not ( n39546 , n39545 );
buf ( n39547 , n39546 );
buf ( n39548 , n39547 );
nand ( n39549 , n39536 , n39548 );
buf ( n39550 , n39549 );
buf ( n39551 , n39550 );
nor ( n39552 , n39528 , n39551 );
buf ( n39553 , n39552 );
buf ( n39554 , n39553 );
nand ( n39555 , n39521 , n39554 );
buf ( n39556 , n39555 );
buf ( n39557 , n38434 );
buf ( n39558 , n38408 );
nor ( n39559 , n39557 , n39558 );
buf ( n39560 , n39559 );
not ( n39561 , n39560 );
nor ( n39562 , n39561 , n39497 );
and ( n39563 , n39556 , n39562 );
not ( n39564 , n39556 );
buf ( n39565 , n39560 );
not ( n39566 , n39565 );
buf ( n39567 , n39566 );
not ( n39568 , n39567 );
nor ( n39569 , n39568 , n39497 );
and ( n39570 , n39564 , n39569 );
nor ( n39571 , n39563 , n39570 );
nand ( n39572 , n39508 , n39571 );
not ( n39573 , n39572 );
buf ( n39574 , n39573 );
buf ( n39575 , n39574 );
buf ( n39576 , n10430 );
buf ( n39577 , n18571 );
buf ( n39578 , n38457 );
not ( n39579 , n38897 );
buf ( n39580 , n39579 );
and ( n39581 , n39578 , n39580 );
buf ( n39582 , n39581 );
buf ( n39583 , n39582 );
and ( n39584 , n39577 , n39583 );
buf ( n39585 , n39584 );
buf ( n39586 , n39585 );
nand ( n39587 , n39576 , n39586 );
buf ( n39588 , n39587 );
and ( n39589 , n39579 , n38444 );
nor ( n39590 , n39589 , n38951 );
buf ( n39591 , n18585 );
buf ( n39592 , n39582 );
nand ( n39593 , n39591 , n39592 );
buf ( n39594 , n39593 );
nand ( n39595 , n39588 , n39590 , n39594 );
buf ( n39596 , n39080 );
buf ( n39597 , n38956 );
nand ( n39598 , n39596 , n39597 );
buf ( n39599 , n39598 );
xnor ( n39600 , n39595 , n39599 );
or ( n39601 , n39575 , n39600 );
buf ( n39602 , n39283 );
buf ( n39603 , n39602 );
not ( n39604 , n1152 );
buf ( n39605 , n37825 );
not ( n39606 , n39605 );
buf ( n39607 , n39469 );
not ( n39608 , n39607 );
or ( n39609 , n39606 , n39608 );
buf ( n39610 , n38191 );
nand ( n39611 , n39609 , n39610 );
buf ( n39612 , n39611 );
not ( n39613 , n39612 );
buf ( n39614 , n37762 );
not ( n39615 , n37825 );
nor ( n39616 , n39615 , n39444 );
buf ( n39617 , n39616 );
nand ( n39618 , n39614 , n39617 );
buf ( n39619 , n39618 );
nand ( n39620 , n31968 , n38136 , n39616 );
nand ( n39621 , n39613 , n39619 , n39620 );
buf ( n39622 , n39621 );
buf ( n39623 , n37833 );
buf ( n39624 , n38198 );
nand ( n39625 , n39623 , n39624 );
buf ( n39626 , n39625 );
buf ( n39627 , n39626 );
not ( n39628 , n39627 );
buf ( n39629 , n39628 );
buf ( n39630 , n39629 );
and ( n39631 , n39622 , n39630 );
not ( n39632 , n39622 );
buf ( n39633 , n39626 );
and ( n39634 , n39632 , n39633 );
nor ( n39635 , n39631 , n39634 );
buf ( n39636 , n39635 );
not ( n39637 , n39636 );
or ( n39638 , n39604 , n39637 );
buf ( n39639 , n17930 );
not ( n39640 , n39639 );
buf ( n39641 , n18184 );
not ( n39642 , n39641 );
or ( n39643 , n39640 , n39642 );
buf ( n39644 , n18196 );
nand ( n39645 , n39643 , n39644 );
buf ( n39646 , n39645 );
not ( n39647 , n39646 );
buf ( n39648 , n18133 );
buf ( n39649 , n17930 );
not ( n39650 , n39649 );
buf ( n39651 , n17735 );
nor ( n39652 , n39650 , n39651 );
buf ( n39653 , n39652 );
buf ( n39654 , n39653 );
and ( n39655 , n39648 , n39654 );
buf ( n39656 , n39655 );
buf ( n39657 , n39656 );
buf ( n39658 , n10417 );
nand ( n39659 , n39657 , n39658 );
buf ( n39660 , n39659 );
buf ( n39661 , n16833 );
buf ( n39662 , n39653 );
nand ( n39663 , n39661 , n39662 );
buf ( n39664 , n39663 );
nand ( n39665 , n39647 , n39660 , n39664 );
buf ( n39666 , n18093 );
buf ( n39667 , n18206 );
nand ( n39668 , n39666 , n39667 );
buf ( n39669 , n39668 );
buf ( n39670 , n39669 );
not ( n39671 , n39670 );
buf ( n39672 , n39671 );
and ( n39673 , n39665 , n39672 );
not ( n39674 , n39665 );
and ( n39675 , n39674 , n39669 );
nor ( n39676 , n39673 , n39675 );
nand ( n39677 , n39676 , n831 );
nand ( n39678 , n39638 , n39677 );
not ( n39679 , n39678 );
not ( n39680 , n39679 );
buf ( n39681 , n39680 );
or ( n39682 , n39603 , n39681 );
and ( n39683 , n831 , n18376 );
not ( n39684 , n831 );
buf ( n39685 , n39476 );
buf ( n39686 , n38208 );
not ( n39687 , n39686 );
and ( n39688 , n39685 , n39687 );
buf ( n39689 , n39688 );
not ( n39690 , n39689 );
not ( n39691 , n39690 );
buf ( n39692 , n39440 );
buf ( n39693 , n37836 );
buf ( n39694 , n39447 );
nand ( n39695 , n39693 , n39694 );
buf ( n39696 , n39695 );
buf ( n39697 , n39696 );
nor ( n39698 , n39692 , n39697 );
buf ( n39699 , n39698 );
nand ( n39700 , n39699 , n31968 );
not ( n39701 , n37759 );
not ( n39702 , n39696 );
nand ( n39703 , n39701 , n39702 );
and ( n39704 , n37836 , n39469 );
nor ( n39705 , n39704 , n38201 );
nand ( n39706 , n39700 , n39703 , n39705 );
not ( n39707 , n39706 );
or ( n39708 , n39691 , n39707 );
nand ( n39709 , n39700 , n39703 , n39705 , n39689 );
nand ( n39710 , n39708 , n39709 );
and ( n39711 , n39684 , n39710 );
nor ( n39712 , n39683 , n39711 );
not ( n39713 , n39712 );
buf ( n39714 , n39713 );
not ( n39715 , n39714 );
not ( n39716 , n39715 );
buf ( n39717 , n39155 );
or ( n39718 , n39716 , n39717 );
not ( n39719 , n831 );
buf ( n39720 , n18184 );
not ( n39721 , n39720 );
buf ( n39722 , n10430 );
buf ( n39723 , n18571 );
buf ( n39724 , n17738 );
and ( n39725 , n39723 , n39724 );
buf ( n39726 , n39725 );
buf ( n39727 , n39726 );
nand ( n39728 , n39722 , n39727 );
buf ( n39729 , n39728 );
buf ( n39730 , n39729 );
buf ( n39731 , n16833 );
buf ( n39732 , n17738 );
nand ( n39733 , n39731 , n39732 );
buf ( n39734 , n39733 );
buf ( n39735 , n39734 );
nand ( n39736 , n39721 , n39730 , n39735 );
buf ( n39737 , n39736 );
buf ( n39738 , n39737 );
buf ( n39739 , n17930 );
buf ( n39740 , n18196 );
nand ( n39741 , n39739 , n39740 );
buf ( n39742 , n39741 );
buf ( n39743 , n39742 );
not ( n39744 , n39743 );
buf ( n39745 , n39744 );
buf ( n39746 , n39745 );
and ( n39747 , n39738 , n39746 );
not ( n39748 , n39738 );
buf ( n39749 , n39742 );
and ( n39750 , n39748 , n39749 );
nor ( n39751 , n39747 , n39750 );
buf ( n39752 , n39751 );
not ( n39753 , n39752 );
or ( n39754 , n39719 , n39753 );
not ( n39755 , n39469 );
buf ( n39756 , n39233 );
buf ( n39757 , n39447 );
nand ( n39758 , n39756 , n39757 );
buf ( n39759 , n39758 );
nand ( n39760 , n31968 , n39242 , n39447 );
nand ( n39761 , n39755 , n39759 , n39760 );
buf ( n39762 , n39761 );
buf ( n39763 , n37825 );
buf ( n39764 , n38191 );
nand ( n39765 , n39763 , n39764 );
buf ( n39766 , n39765 );
buf ( n39767 , n39766 );
not ( n39768 , n39767 );
buf ( n39769 , n39768 );
buf ( n39770 , n39769 );
and ( n39771 , n39762 , n39770 );
not ( n39772 , n39762 );
buf ( n39773 , n39766 );
and ( n39774 , n39772 , n39773 );
nor ( n39775 , n39771 , n39774 );
buf ( n39776 , n39775 );
nand ( n39777 , n39776 , n1152 );
nand ( n39778 , n39754 , n39777 );
buf ( n39779 , n39778 );
buf ( n39780 , n38466 );
and ( n39781 , n39780 , n38493 );
not ( n39782 , n39780 );
and ( n39783 , n39782 , n38488 );
nor ( n39784 , n39781 , n39783 );
or ( n39785 , n39779 , n39784 );
and ( n39786 , n39601 , n39682 , n39718 , n39785 );
not ( n39787 , n39786 );
buf ( n39788 , n39233 );
buf ( n39789 , n37807 );
nand ( n39790 , n39788 , n39789 );
buf ( n39791 , n39790 );
buf ( n39792 , n39791 );
nand ( n39793 , n31968 , n39242 , n37807 );
buf ( n39794 , n39793 );
buf ( n39795 , n38156 );
buf ( n39796 , n39795 );
buf ( n39797 , n39796 );
buf ( n39798 , n39797 );
not ( n39799 , n39798 );
buf ( n39800 , n39799 );
buf ( n39801 , n39800 );
nand ( n39802 , n39792 , n39794 , n39801 );
buf ( n39803 , n39802 );
not ( n39804 , n39803 );
buf ( n39805 , n38167 );
buf ( n39806 , n37782 );
buf ( n39807 , n39806 );
buf ( n39808 , n39807 );
buf ( n39809 , n39808 );
nor ( n39810 , n39805 , n39809 );
buf ( n39811 , n39810 );
nor ( n39812 , n39811 , n831 );
nand ( n39813 , n39804 , n39812 );
not ( n39814 , n18158 );
buf ( n39815 , n10430 );
buf ( n39816 , n18571 );
buf ( n39817 , n17729 );
and ( n39818 , n39816 , n39817 );
buf ( n39819 , n39818 );
buf ( n39820 , n39819 );
nand ( n39821 , n39815 , n39820 );
buf ( n39822 , n39821 );
buf ( n39823 , n16833 );
buf ( n39824 , n17729 );
nand ( n39825 , n39823 , n39824 );
buf ( n39826 , n39825 );
nand ( n39827 , n39814 , n39822 , n39826 );
not ( n39828 , n39827 );
buf ( n39829 , n18558 );
buf ( n39830 , n18166 );
nand ( n39831 , n39829 , n39830 );
buf ( n39832 , n39831 );
and ( n39833 , n39832 , n831 );
nand ( n39834 , n39828 , n39833 );
not ( n39835 , n39811 );
nor ( n39836 , n39835 , n831 );
nand ( n39837 , n39803 , n39836 );
buf ( n39838 , n39832 );
not ( n39839 , n39838 );
buf ( n39840 , n39839 );
and ( n39841 , n39840 , n831 );
nand ( n39842 , n39827 , n39841 );
nand ( n39843 , n39813 , n39834 , n39837 , n39842 );
buf ( n39844 , n39843 );
not ( n39845 , n39844 );
not ( n39846 , n39845 );
not ( n39847 , n39846 );
buf ( n39848 , n39556 );
and ( n39849 , n39848 , n39560 );
not ( n39850 , n39848 );
and ( n39851 , n39850 , n39567 );
nor ( n39852 , n39849 , n39851 );
or ( n39853 , n39847 , n39852 );
buf ( n39854 , n1152 );
buf ( n39855 , n39233 );
not ( n39856 , n37807 );
nor ( n39857 , n39856 , n39808 );
buf ( n39858 , n39857 );
nand ( n39859 , n39855 , n39858 );
buf ( n39860 , n39859 );
buf ( n39861 , n39860 );
buf ( n39862 , n39242 );
buf ( n39863 , n39857 );
and ( n39864 , n39862 , n39863 );
buf ( n39865 , n39864 );
buf ( n39866 , n39865 );
buf ( n39867 , n31968 );
nand ( n39868 , n39866 , n39867 );
buf ( n39869 , n39868 );
buf ( n39870 , n39869 );
buf ( n39871 , n39797 );
buf ( n39872 , n39808 );
not ( n39873 , n39872 );
buf ( n39874 , n39873 );
buf ( n39875 , n39874 );
and ( n39876 , n39871 , n39875 );
buf ( n39877 , n38167 );
nor ( n39878 , n39876 , n39877 );
buf ( n39879 , n39878 );
buf ( n39880 , n39879 );
nand ( n39881 , n39861 , n39870 , n39880 );
buf ( n39882 , n39881 );
buf ( n39883 , n38162 );
not ( n39884 , n39883 );
buf ( n39885 , n38173 );
nor ( n39886 , n39884 , n39885 );
buf ( n39887 , n39886 );
xor ( n39888 , n39882 , n39887 );
and ( n39889 , n39854 , n39888 );
not ( n39890 , n39854 );
and ( n39891 , n39890 , n18606 );
nor ( n39892 , n39889 , n39891 );
buf ( n39893 , n39892 );
buf ( n39894 , n39893 );
buf ( n39895 , n39894 );
not ( n39896 , n39895 );
and ( n39897 , n38995 , n39002 );
not ( n39898 , n38995 );
and ( n39899 , n39898 , n38999 );
nor ( n39900 , n39897 , n39899 );
or ( n39901 , n39896 , n39900 );
nand ( n39902 , n39853 , n39901 );
buf ( n39903 , n37725 );
buf ( n39904 , n37795 );
nor ( n39905 , n39903 , n39904 );
buf ( n39906 , n39905 );
buf ( n39907 , n39906 );
not ( n39908 , n39907 );
buf ( n39909 , n32124 );
not ( n39910 , n39909 );
or ( n39911 , n39908 , n39910 );
buf ( n39912 , n37795 );
not ( n39913 , n39912 );
buf ( n39914 , n39913 );
buf ( n39915 , n39914 );
not ( n39916 , n39915 );
buf ( n39917 , n37693 );
not ( n39918 , n39917 );
buf ( n39919 , n31762 );
not ( n39920 , n39919 );
or ( n39921 , n39918 , n39920 );
buf ( n39922 , n37737 );
nand ( n39923 , n39921 , n39922 );
buf ( n39924 , n39923 );
buf ( n39925 , n39924 );
not ( n39926 , n39925 );
or ( n39927 , n39916 , n39926 );
buf ( n39928 , n37792 );
buf ( n39929 , n37790 );
nand ( n39930 , n39928 , n39929 );
buf ( n39931 , n39930 );
buf ( n39932 , n39931 );
nand ( n39933 , n39927 , n39932 );
buf ( n39934 , n39933 );
buf ( n39935 , n39934 );
not ( n39936 , n39935 );
buf ( n39937 , n39936 );
buf ( n39938 , n39937 );
nand ( n39939 , n39911 , n39938 );
buf ( n39940 , n39939 );
buf ( n39941 , n37804 );
not ( n39942 , n39941 );
buf ( n39943 , n37800 );
buf ( n39944 , n17723 );
buf ( n39945 , n39944 );
nand ( n39946 , n39943 , n39945 );
buf ( n39947 , n39946 );
buf ( n39948 , n39947 );
nand ( n39949 , n39942 , n39948 );
buf ( n39950 , n39949 );
buf ( n39951 , n39950 );
not ( n39952 , n39951 );
buf ( n39953 , n39952 );
and ( n39954 , n39940 , n39953 );
not ( n39955 , n39940 );
and ( n39956 , n39955 , n39950 );
nor ( n39957 , n39954 , n39956 );
not ( n39958 , n39957 );
not ( n39959 , n1152 );
or ( n39960 , n39958 , n39959 );
nand ( n39961 , n39960 , n32036 );
buf ( n39962 , n39961 );
not ( n39963 , n39962 );
not ( n39964 , n39963 );
nor ( n39965 , n39964 , n18377 );
not ( n39966 , n39965 );
buf ( n39967 , n39242 );
not ( n39968 , n39967 );
buf ( n39969 , n31632 );
not ( n39970 , n39969 );
or ( n39971 , n39968 , n39970 );
buf ( n39972 , n37759 );
nand ( n39973 , n39971 , n39972 );
buf ( n39974 , n39973 );
not ( n39975 , n39974 );
buf ( n39976 , n39914 );
buf ( n39977 , n39931 );
nand ( n39978 , n39976 , n39977 );
buf ( n39979 , n39978 );
not ( n39980 , n39979 );
nor ( n39981 , n39980 , n831 );
nand ( n39982 , n39975 , n39981 );
buf ( n39983 , n18133 );
not ( n39984 , n39983 );
buf ( n39985 , n10427 );
not ( n39986 , n39985 );
or ( n39987 , n39984 , n39986 );
buf ( n39988 , n16784 );
not ( n39989 , n39988 );
buf ( n39990 , n16811 );
not ( n39991 , n39990 );
or ( n39992 , n39989 , n39991 );
buf ( n39993 , n16829 );
nand ( n39994 , n39992 , n39993 );
buf ( n39995 , n39994 );
buf ( n39996 , n39995 );
nand ( n39997 , n39987 , n39996 );
buf ( n39998 , n39997 );
not ( n39999 , n39998 );
buf ( n40000 , n18787 );
buf ( n40001 , n18151 );
nand ( n40002 , n40000 , n40001 );
buf ( n40003 , n40002 );
nand ( n40004 , n39999 , n40003 , n831 );
not ( n40005 , n831 );
nor ( n40006 , n40003 , n40005 );
nand ( n40007 , n39998 , n40006 );
not ( n40008 , n39979 );
nand ( n40009 , n40008 , n39974 , n40005 );
nand ( n40010 , n39982 , n40004 , n40007 , n40009 );
not ( n40011 , n40010 );
buf ( n40012 , n40011 );
buf ( n40013 , n39665 );
and ( n40014 , n40013 , n39672 );
not ( n40015 , n40013 );
and ( n40016 , n40015 , n39669 );
nor ( n40017 , n40014 , n40016 );
or ( n40018 , n40012 , n40017 );
nand ( n40019 , n39966 , n40018 );
nor ( n40020 , n39902 , n40019 );
not ( n40021 , n40020 );
buf ( n40022 , n16713 );
buf ( n40023 , n14550 );
buf ( n40024 , n40023 );
buf ( n40025 , n40024 );
buf ( n40026 , n40025 );
buf ( n40027 , n15319 );
not ( n40028 , n40027 );
buf ( n40029 , n40028 );
buf ( n40030 , n40029 );
nand ( n40031 , n40026 , n40030 );
buf ( n40032 , n40031 );
buf ( n40033 , n40032 );
nor ( n40034 , n40022 , n40033 );
buf ( n40035 , n40034 );
buf ( n40036 , n40035 );
not ( n40037 , n40036 );
buf ( n40038 , n10417 );
not ( n40039 , n40038 );
or ( n40040 , n40037 , n40039 );
buf ( n40041 , n40032 );
not ( n40042 , n40041 );
buf ( n40043 , n40042 );
buf ( n40044 , n40043 );
not ( n40045 , n40044 );
buf ( n40046 , n16736 );
not ( n40047 , n40046 );
or ( n40048 , n40045 , n40047 );
buf ( n40049 , n40029 );
not ( n40050 , n40049 );
buf ( n40051 , n16333 );
buf ( n40052 , n40051 );
not ( n40053 , n40052 );
or ( n40054 , n40050 , n40053 );
buf ( n40055 , n16352 );
not ( n40056 , n40055 );
buf ( n40057 , n40056 );
buf ( n40058 , n40057 );
nand ( n40059 , n40054 , n40058 );
buf ( n40060 , n40059 );
buf ( n40061 , n40060 );
not ( n40062 , n40061 );
buf ( n40063 , n40062 );
buf ( n40064 , n40063 );
nand ( n40065 , n40048 , n40064 );
buf ( n40066 , n40065 );
buf ( n40067 , n40066 );
not ( n40068 , n40067 );
buf ( n40069 , n40068 );
buf ( n40070 , n40069 );
nand ( n40071 , n40040 , n40070 );
buf ( n40072 , n40071 );
buf ( n40073 , n15296 );
buf ( n40074 , n16359 );
and ( n40075 , n40073 , n40074 );
buf ( n40076 , n40075 );
and ( n40077 , n40072 , n40076 );
not ( n40078 , n40072 );
buf ( n40079 , n40076 );
not ( n40080 , n40079 );
buf ( n40081 , n40080 );
and ( n40082 , n40078 , n40081 );
nor ( n40083 , n40077 , n40082 );
and ( n40084 , n831 , n40083 );
not ( n40085 , n831 );
buf ( n40086 , n31182 );
not ( n40087 , n40086 );
buf ( n40088 , n40087 );
buf ( n40089 , n40088 );
buf ( n40090 , n31010 );
buf ( n40091 , n40090 );
buf ( n40092 , n40091 );
buf ( n40093 , n40092 );
buf ( n40094 , n31020 );
buf ( n40095 , n40094 );
buf ( n40096 , n40095 );
buf ( n40097 , n40096 );
nand ( n40098 , n40093 , n40097 );
buf ( n40099 , n40098 );
buf ( n40100 , n40099 );
nor ( n40101 , n40089 , n40100 );
buf ( n40102 , n40101 );
not ( n40103 , n40102 );
not ( n40104 , n31632 );
or ( n40105 , n40103 , n40104 );
buf ( n40106 , n40099 );
not ( n40107 , n40106 );
buf ( n40108 , n40107 );
buf ( n40109 , n40108 );
not ( n40110 , n40109 );
buf ( n40111 , n31721 );
not ( n40112 , n40111 );
or ( n40113 , n40110 , n40112 );
buf ( n40114 , n40096 );
not ( n40115 , n40114 );
buf ( n40116 , n31744 );
buf ( n40117 , n40116 );
buf ( n40118 , n40117 );
buf ( n40119 , n40118 );
not ( n40120 , n40119 );
or ( n40121 , n40115 , n40120 );
buf ( n40122 , n31754 );
not ( n40123 , n40122 );
buf ( n40124 , n40123 );
buf ( n40125 , n40124 );
nand ( n40126 , n40121 , n40125 );
buf ( n40127 , n40126 );
buf ( n40128 , n40127 );
not ( n40129 , n40128 );
buf ( n40130 , n40129 );
buf ( n40131 , n40130 );
nand ( n40132 , n40113 , n40131 );
buf ( n40133 , n40132 );
buf ( n40134 , n40133 );
not ( n40135 , n40134 );
buf ( n40136 , n40135 );
nand ( n40137 , n40105 , n40136 );
buf ( n40138 , n31757 );
nand ( n40139 , n40138 , n31029 );
not ( n40140 , n40139 );
and ( n40141 , n40137 , n40140 );
not ( n40142 , n40137 );
and ( n40143 , n40142 , n40139 );
nor ( n40144 , n40141 , n40143 );
and ( n40145 , n40085 , n40144 );
nor ( n40146 , n40084 , n40145 );
not ( n40147 , n40146 );
not ( n40148 , n40147 );
not ( n40149 , n40148 );
xnor ( n40150 , n39998 , n40003 );
or ( n40151 , n40149 , n40150 );
buf ( n40152 , n40088 );
buf ( n40153 , n31009 );
nor ( n40154 , n40152 , n40153 );
buf ( n40155 , n40154 );
buf ( n40156 , n40155 );
not ( n40157 , n40156 );
buf ( n40158 , n31968 );
not ( n40159 , n40158 );
or ( n40160 , n40157 , n40159 );
buf ( n40161 , n32128 );
not ( n40162 , n40161 );
buf ( n40163 , n31721 );
not ( n40164 , n40163 );
or ( n40165 , n40162 , n40164 );
buf ( n40166 , n32132 );
nand ( n40167 , n40165 , n40166 );
buf ( n40168 , n40167 );
buf ( n40169 , n40168 );
not ( n40170 , n40169 );
buf ( n40171 , n40170 );
buf ( n40172 , n40171 );
nand ( n40173 , n40160 , n40172 );
buf ( n40174 , n40173 );
not ( n40175 , n40174 );
buf ( n40176 , n31728 );
buf ( n40177 , n31741 );
and ( n40178 , n40176 , n40177 );
buf ( n40179 , n40178 );
nor ( n40180 , n40179 , n831 );
nand ( n40181 , n40175 , n40180 );
buf ( n40182 , n16713 );
buf ( n40183 , n14549 );
buf ( n40184 , n40183 );
nor ( n40185 , n40182 , n40184 );
buf ( n40186 , n40185 );
buf ( n40187 , n40186 );
not ( n40188 , n40187 );
buf ( n40189 , n10417 );
not ( n40190 , n40189 );
or ( n40191 , n40188 , n40190 );
buf ( n40192 , n40183 );
not ( n40193 , n40192 );
buf ( n40194 , n40193 );
buf ( n40195 , n40194 );
not ( n40196 , n40195 );
buf ( n40197 , n16736 );
not ( n40198 , n40197 );
or ( n40199 , n40196 , n40198 );
buf ( n40200 , n16328 );
buf ( n40201 , n40200 );
nand ( n40202 , n40199 , n40201 );
buf ( n40203 , n40202 );
buf ( n40204 , n40203 );
not ( n40205 , n40204 );
buf ( n40206 , n40205 );
buf ( n40207 , n40206 );
nand ( n40208 , n40191 , n40207 );
buf ( n40209 , n40208 );
not ( n40210 , n40209 );
buf ( n40211 , n16326 );
buf ( n40212 , n16332 );
and ( n40213 , n40211 , n40212 );
buf ( n40214 , n40213 );
buf ( n40215 , n40214 );
not ( n40216 , n40215 );
buf ( n40217 , n40216 );
and ( n40218 , n40217 , n831 );
nand ( n40219 , n40210 , n40218 );
nand ( n40220 , n40209 , n40214 , n831 );
not ( n40221 , n40179 );
nor ( n40222 , n40221 , n831 );
nand ( n40223 , n40174 , n40222 );
nand ( n40224 , n40181 , n40219 , n40220 , n40223 );
buf ( n40225 , n40224 );
not ( n40226 , n40225 );
buf ( n40227 , n10427 );
not ( n40228 , n40227 );
buf ( n40229 , n13771 );
buf ( n40230 , n15325 );
not ( n40231 , n40230 );
buf ( n40232 , n15945 );
nand ( n40233 , n40231 , n40232 );
buf ( n40234 , n40233 );
buf ( n40235 , n40234 );
nor ( n40236 , n40229 , n40235 );
buf ( n40237 , n40236 );
buf ( n40238 , n40237 );
not ( n40239 , n40238 );
or ( n40240 , n40228 , n40239 );
buf ( n40241 , n40234 );
not ( n40242 , n40241 );
buf ( n40243 , n40242 );
buf ( n40244 , n40243 );
not ( n40245 , n40244 );
buf ( n40246 , n16736 );
not ( n40247 , n40246 );
or ( n40248 , n40245 , n40247 );
buf ( n40249 , n15945 );
not ( n40250 , n40249 );
buf ( n40251 , n16368 );
not ( n40252 , n40251 );
or ( n40253 , n40250 , n40252 );
buf ( n40254 , n16394 );
not ( n40255 , n40254 );
buf ( n40256 , n40255 );
buf ( n40257 , n40256 );
nand ( n40258 , n40253 , n40257 );
buf ( n40259 , n40258 );
buf ( n40260 , n40259 );
not ( n40261 , n40260 );
buf ( n40262 , n40261 );
buf ( n40263 , n40262 );
nand ( n40264 , n40248 , n40263 );
buf ( n40265 , n40264 );
buf ( n40266 , n40265 );
not ( n40267 , n40266 );
buf ( n40268 , n40267 );
buf ( n40269 , n40268 );
nand ( n40270 , n40240 , n40269 );
buf ( n40271 , n40270 );
buf ( n40272 , n16223 );
buf ( n40273 , n16401 );
nand ( n40274 , n40272 , n40273 );
buf ( n40275 , n40274 );
buf ( n40276 , n40275 );
not ( n40277 , n40276 );
buf ( n40278 , n40277 );
and ( n40279 , n40271 , n40278 );
not ( n40280 , n40271 );
and ( n40281 , n40280 , n40275 );
nor ( n40282 , n40279 , n40281 );
or ( n40283 , n40226 , n40282 );
not ( n40284 , n831 );
buf ( n40285 , n13771 );
buf ( n40286 , n40025 );
not ( n40287 , n40286 );
buf ( n40288 , n40287 );
buf ( n40289 , n40288 );
nor ( n40290 , n40285 , n40289 );
buf ( n40291 , n40290 );
buf ( n40292 , n40291 );
not ( n40293 , n40292 );
buf ( n40294 , n10417 );
not ( n40295 , n40294 );
or ( n40296 , n40293 , n40295 );
buf ( n40297 , n40025 );
buf ( n40298 , n16313 );
and ( n40299 , n40297 , n40298 );
buf ( n40300 , n40051 );
nor ( n40301 , n40299 , n40300 );
buf ( n40302 , n40301 );
buf ( n40303 , n40302 );
nand ( n40304 , n40296 , n40303 );
buf ( n40305 , n40304 );
buf ( n40306 , n40029 );
buf ( n40307 , n40057 );
nand ( n40308 , n40306 , n40307 );
buf ( n40309 , n40308 );
buf ( n40310 , n40309 );
not ( n40311 , n40310 );
buf ( n40312 , n40311 );
and ( n40313 , n40305 , n40312 );
not ( n40314 , n40305 );
and ( n40315 , n40314 , n40309 );
nor ( n40316 , n40313 , n40315 );
not ( n40317 , n40316 );
or ( n40318 , n40284 , n40317 );
buf ( n40319 , n40092 );
not ( n40320 , n40319 );
buf ( n40321 , n40088 );
nor ( n40322 , n40320 , n40321 );
buf ( n40323 , n40322 );
buf ( n40324 , n40323 );
not ( n40325 , n40324 );
buf ( n40326 , n31968 );
not ( n40327 , n40326 );
or ( n40328 , n40325 , n40327 );
buf ( n40329 , n40092 );
not ( n40330 , n40329 );
buf ( n40331 , n31721 );
not ( n40332 , n40331 );
or ( n40333 , n40330 , n40332 );
buf ( n40334 , n40118 );
not ( n40335 , n40334 );
buf ( n40336 , n40335 );
buf ( n40337 , n40336 );
nand ( n40338 , n40333 , n40337 );
buf ( n40339 , n40338 );
buf ( n40340 , n40339 );
not ( n40341 , n40340 );
buf ( n40342 , n40341 );
buf ( n40343 , n40342 );
nand ( n40344 , n40328 , n40343 );
buf ( n40345 , n40344 );
buf ( n40346 , n40345 );
buf ( n40347 , n40096 );
buf ( n40348 , n40124 );
nand ( n40349 , n40347 , n40348 );
buf ( n40350 , n40349 );
buf ( n40351 , n40350 );
not ( n40352 , n40351 );
buf ( n40353 , n40352 );
buf ( n40354 , n40353 );
and ( n40355 , n40346 , n40354 );
not ( n40356 , n40346 );
buf ( n40357 , n40350 );
and ( n40358 , n40356 , n40357 );
nor ( n40359 , n40355 , n40358 );
buf ( n40360 , n40359 );
nand ( n40361 , n40360 , n1152 );
nand ( n40362 , n40318 , n40361 );
buf ( n40363 , n40362 );
buf ( n40364 , n40363 );
or ( n40365 , n40364 , n16710 );
nand ( n40366 , n40194 , n40200 );
not ( n40367 , n40366 );
and ( n40368 , n18773 , n40367 );
not ( n40369 , n18773 );
and ( n40370 , n40369 , n40366 );
nor ( n40371 , n40368 , n40370 );
not ( n40372 , n40371 );
not ( n40373 , n831 );
or ( n40374 , n40372 , n40373 );
nand ( n40375 , n40374 , n32139 );
buf ( n40376 , n40375 );
buf ( n40377 , n40376 );
or ( n40378 , n16777 , n40377 );
and ( n40379 , n40151 , n40283 , n40365 , n40378 );
not ( n40380 , n31815 );
buf ( n40381 , n40380 );
buf ( n40382 , n40381 );
and ( n40383 , n39827 , n39840 );
not ( n40384 , n39827 );
and ( n40385 , n40384 , n39832 );
nor ( n40386 , n40383 , n40385 );
or ( n40387 , n40382 , n40386 );
buf ( n40388 , n31847 );
buf ( n40389 , n40388 );
or ( n40390 , n40389 , n18802 );
nand ( n40391 , n40387 , n40390 );
and ( n40392 , n40271 , n40278 );
nor ( n40393 , n40392 , n40005 );
not ( n40394 , n40393 );
not ( n40395 , n40271 );
nand ( n40396 , n40395 , n40275 );
not ( n40397 , n40396 );
or ( n40398 , n40394 , n40397 );
buf ( n40399 , n31036 );
buf ( n40400 , n37674 );
not ( n40401 , n40400 );
buf ( n40402 , n40401 );
buf ( n40403 , n40402 );
nor ( n40404 , n40399 , n40403 );
buf ( n40405 , n40404 );
buf ( n40406 , n40405 );
buf ( n40407 , n31182 );
nand ( n40408 , n40406 , n40407 );
buf ( n40409 , n40408 );
buf ( n40410 , n40409 );
not ( n40411 , n40410 );
buf ( n40412 , n31631 );
not ( n40413 , n40412 );
and ( n40414 , n40411 , n40413 );
not ( n40415 , n40405 );
nand ( n40416 , n31720 , n31670 );
not ( n40417 , n40416 );
or ( n40418 , n40415 , n40417 );
buf ( n40419 , n31827 );
not ( n40420 , n40419 );
buf ( n40421 , n40402 );
not ( n40422 , n40421 );
and ( n40423 , n40420 , n40422 );
buf ( n40424 , n37703 );
nor ( n40425 , n40423 , n40424 );
buf ( n40426 , n40425 );
nand ( n40427 , n40418 , n40426 );
buf ( n40428 , n40427 );
nor ( n40429 , n40414 , n40428 );
buf ( n40430 , n40429 );
buf ( n40431 , n40430 );
buf ( n40432 , n37688 );
not ( n40433 , n40432 );
buf ( n40434 , n40433 );
buf ( n40435 , n40434 );
buf ( n40436 , n37710 );
nand ( n40437 , n40435 , n40436 );
buf ( n40438 , n40437 );
buf ( n40439 , n40438 );
and ( n40440 , n40431 , n40439 );
not ( n40441 , n40431 );
buf ( n40442 , n40438 );
not ( n40443 , n40442 );
buf ( n40444 , n40443 );
buf ( n40445 , n40444 );
and ( n40446 , n40441 , n40445 );
nor ( n40447 , n40440 , n40446 );
buf ( n40448 , n40447 );
nand ( n40449 , n40448 , n1152 );
nand ( n40450 , n40398 , n40449 );
buf ( n40451 , n40450 );
buf ( n40452 , n40451 );
or ( n40453 , n40452 , n18607 );
not ( n40454 , n31817 );
buf ( n40455 , n31036 );
buf ( n40456 , n37674 );
buf ( n40457 , n40434 );
nand ( n40458 , n40456 , n40457 );
buf ( n40459 , n40458 );
buf ( n40460 , n40459 );
nor ( n40461 , n40455 , n40460 );
buf ( n40462 , n40461 );
buf ( n40463 , n40462 );
buf ( n40464 , n31182 );
nand ( n40465 , n40463 , n40464 );
buf ( n40466 , n40465 );
nor ( n40467 , n40454 , n40466 );
not ( n40468 , n40467 );
not ( n40469 , n40468 );
buf ( n40470 , n37713 );
not ( n40471 , n40470 );
nor ( n40472 , n37680 , n37675 );
buf ( n40473 , n40472 );
nor ( n40474 , n40471 , n40473 );
buf ( n40475 , n40474 );
not ( n40476 , n40475 );
buf ( n40477 , n40462 );
not ( n40478 , n40477 );
buf ( n40479 , n31721 );
not ( n40480 , n40479 );
or ( n40481 , n40478 , n40480 );
buf ( n40482 , n31827 );
not ( n40483 , n40482 );
buf ( n40484 , n40459 );
not ( n40485 , n40484 );
and ( n40486 , n40483 , n40485 );
buf ( n40487 , n40434 );
not ( n40488 , n40487 );
buf ( n40489 , n37703 );
not ( n40490 , n40489 );
or ( n40491 , n40488 , n40490 );
buf ( n40492 , n37710 );
nand ( n40493 , n40491 , n40492 );
buf ( n40494 , n40493 );
buf ( n40495 , n40494 );
nor ( n40496 , n40486 , n40495 );
buf ( n40497 , n40496 );
buf ( n40498 , n40497 );
nand ( n40499 , n40481 , n40498 );
buf ( n40500 , n40499 );
nor ( n40501 , n40476 , n40500 );
not ( n40502 , n40501 );
or ( n40503 , n40469 , n40502 );
or ( n40504 , n40467 , n40500 );
not ( n40505 , n40475 );
nand ( n40506 , n40504 , n40505 );
nand ( n40507 , n40503 , n40506 );
not ( n40508 , n40507 );
not ( n40509 , n1152 );
or ( n40510 , n40508 , n40509 );
nand ( n40511 , n40510 , n32056 );
buf ( n40512 , n40511 );
not ( n40513 , n40512 );
not ( n40514 , n40513 );
buf ( n40515 , n40514 );
buf ( n40516 , n39752 );
or ( n40517 , n40515 , n40516 );
nand ( n40518 , n40453 , n40517 );
nor ( n40519 , n40391 , n40518 );
and ( n40520 , n40379 , n40519 );
not ( n40521 , n40520 );
not ( n40522 , n18669 );
not ( n40523 , n831 );
or ( n40524 , n40522 , n40523 );
nand ( n40525 , n40524 , n32007 );
buf ( n40526 , n40525 );
not ( n40527 , n40526 );
buf ( n40528 , n40527 );
not ( n40529 , n40528 );
and ( n40530 , n40209 , n40214 );
not ( n40531 , n40209 );
and ( n40532 , n40531 , n40217 );
nor ( n40533 , n40530 , n40532 );
or ( n40534 , n40529 , n40533 );
buf ( n40535 , n1152 );
nor ( n40536 , n31114 , n31990 );
buf ( n40537 , n40536 );
not ( n40538 , n40537 );
buf ( n40539 , n31968 );
not ( n40540 , n40539 );
or ( n40541 , n40538 , n40540 );
not ( n40542 , n31990 );
not ( n40543 , n40542 );
not ( n40544 , n31982 );
or ( n40545 , n40543 , n40544 );
nand ( n40546 , n40545 , n31995 );
buf ( n40547 , n40546 );
not ( n40548 , n40547 );
buf ( n40549 , n40548 );
buf ( n40550 , n40549 );
nand ( n40551 , n40541 , n40550 );
buf ( n40552 , n40551 );
buf ( n40553 , n40552 );
nand ( n40554 , n32140 , n31708 );
buf ( n40555 , n40554 );
not ( n40556 , n40555 );
buf ( n40557 , n40556 );
buf ( n40558 , n40557 );
and ( n40559 , n40553 , n40558 );
not ( n40560 , n40553 );
buf ( n40561 , n40554 );
and ( n40562 , n40560 , n40561 );
nor ( n40563 , n40559 , n40562 );
buf ( n40564 , n40563 );
and ( n40565 , n40535 , n40564 );
not ( n40566 , n40535 );
buf ( n40567 , n18484 );
buf ( n40568 , n12808 );
nor ( n40569 , n40567 , n40568 );
buf ( n40570 , n40569 );
not ( n40571 , n40570 );
not ( n40572 , n10417 );
or ( n40573 , n40571 , n40572 );
not ( n40574 , n18655 );
not ( n40575 , n18504 );
or ( n40576 , n40574 , n40575 );
nand ( n40577 , n40576 , n16258 );
buf ( n40578 , n40577 );
not ( n40579 , n40578 );
buf ( n40580 , n40579 );
nand ( n40581 , n40573 , n40580 );
nand ( n40582 , n18119 , n16278 );
not ( n40583 , n40582 );
and ( n40584 , n40581 , n40583 );
not ( n40585 , n40581 );
and ( n40586 , n40585 , n40582 );
nor ( n40587 , n40584 , n40586 );
and ( n40588 , n40566 , n40587 );
nor ( n40589 , n40565 , n40588 );
not ( n40590 , n40589 );
buf ( n40591 , n40590 );
buf ( n40592 , n40591 );
buf ( n40593 , n40316 );
or ( n40594 , n40592 , n40593 );
nand ( n40595 , n40534 , n40594 );
not ( n40596 , n1152 );
buf ( n40597 , n32142 );
not ( n40598 , n40597 );
buf ( n40599 , n31114 );
nor ( n40600 , n40598 , n40599 );
buf ( n40601 , n40600 );
buf ( n40602 , n40601 );
not ( n40603 , n40602 );
buf ( n40604 , n31817 );
not ( n40605 , n40604 );
or ( n40606 , n40603 , n40605 );
and ( n40607 , n31982 , n32142 );
nor ( n40608 , n40607 , n32169 );
buf ( n40609 , n40608 );
nand ( n40610 , n40606 , n40609 );
buf ( n40611 , n40610 );
buf ( n40612 , n32146 );
buf ( n40613 , n31678 );
nand ( n40614 , n40612 , n40613 );
buf ( n40615 , n40614 );
buf ( n40616 , n40615 );
not ( n40617 , n40616 );
buf ( n40618 , n40617 );
and ( n40619 , n40611 , n40618 );
not ( n40620 , n40611 );
and ( n40621 , n40620 , n40615 );
nor ( n40622 , n40619 , n40621 );
not ( n40623 , n40622 );
or ( n40624 , n40596 , n40623 );
nand ( n40625 , n40624 , n32057 );
buf ( n40626 , n40625 );
not ( n40627 , n40626 );
not ( n40628 , n40627 );
buf ( n40629 , n40083 );
or ( n40630 , n40628 , n40629 );
not ( n40631 , n831 );
not ( n40632 , n18539 );
or ( n40633 , n40631 , n40632 );
nand ( n40634 , n40633 , n32204 );
buf ( n40635 , n40634 );
buf ( n40636 , n40635 );
or ( n40637 , n40636 , n18422 );
nand ( n40638 , n40630 , n40637 );
nor ( n40639 , n40595 , n40638 );
not ( n40640 , n40639 );
not ( n40641 , n1152 );
buf ( n40642 , n31063 );
not ( n40643 , n40642 );
buf ( n40644 , n40643 );
buf ( n40645 , n40644 );
not ( n40646 , n40645 );
buf ( n40647 , n31968 );
not ( n40648 , n40647 );
or ( n40649 , n40646 , n40648 );
nand ( n40650 , n31047 , n31060 );
buf ( n40651 , n40650 );
buf ( n40652 , n40651 );
buf ( n40653 , n40652 );
buf ( n40654 , n40653 );
nand ( n40655 , n40649 , n40654 );
buf ( n40656 , n40655 );
buf ( n40657 , n40656 );
buf ( n40658 , n31079 );
not ( n40659 , n40658 );
buf ( n40660 , n31652 );
nand ( n40661 , n40659 , n40660 );
buf ( n40662 , n40661 );
buf ( n40663 , n40662 );
not ( n40664 , n40663 );
buf ( n40665 , n40664 );
buf ( n40666 , n40665 );
and ( n40667 , n40657 , n40666 );
not ( n40668 , n40657 );
buf ( n40669 , n40662 );
and ( n40670 , n40668 , n40669 );
nor ( n40671 , n40667 , n40670 );
buf ( n40672 , n40671 );
not ( n40673 , n40672 );
or ( n40674 , n40641 , n40673 );
nand ( n40675 , n18477 , n831 );
nand ( n40676 , n40674 , n40675 );
buf ( n40677 , n40676 );
or ( n40678 , n40677 , n18642 );
not ( n40679 , n40678 );
not ( n40680 , n831 );
not ( n40681 , n10435 );
or ( n40682 , n40680 , n40681 );
buf ( n40683 , n40644 );
buf ( n40684 , n40653 );
nand ( n40685 , n40683 , n40684 );
buf ( n40686 , n40685 );
not ( n40687 , n31968 );
xor ( n40688 , n40686 , n40687 );
nand ( n40689 , n40688 , n10103 );
nand ( n40690 , n40682 , n40689 );
buf ( n40691 , n40690 );
buf ( n40692 , n40691 );
buf ( n40693 , n40587 );
and ( n40694 , n40692 , n40693 );
not ( n40695 , n40694 );
or ( n40696 , n40679 , n40695 );
nand ( n40697 , n40677 , n18642 );
nand ( n40698 , n40696 , n40697 );
not ( n40699 , n31080 );
not ( n40700 , n31817 );
or ( n40701 , n40699 , n40700 );
buf ( n40702 , n31654 );
not ( n40703 , n40702 );
buf ( n40704 , n40703 );
nand ( n40705 , n40701 , n40704 );
nand ( n40706 , n31646 , n31655 );
buf ( n40707 , n40706 );
not ( n40708 , n40707 );
buf ( n40709 , n40708 );
and ( n40710 , n40705 , n40709 );
not ( n40711 , n40705 );
and ( n40712 , n40711 , n40706 );
nor ( n40713 , n40710 , n40712 );
not ( n40714 , n40713 );
not ( n40715 , n1152 );
or ( n40716 , n40714 , n40715 );
not ( n40717 , n18683 );
not ( n40718 , n18673 );
nand ( n40719 , n40718 , n10417 );
nand ( n40720 , n40717 , n40719 );
not ( n40721 , n18677 );
nand ( n40722 , n40721 , n18689 );
buf ( n40723 , n40722 );
not ( n40724 , n40723 );
buf ( n40725 , n40724 );
and ( n40726 , n40720 , n40725 );
not ( n40727 , n40720 );
and ( n40728 , n40727 , n40722 );
nor ( n40729 , n40726 , n40728 );
nand ( n40730 , n40729 , n831 );
nand ( n40731 , n40716 , n40730 );
not ( n40732 , n40731 );
buf ( n40733 , n40732 );
not ( n40734 , n40733 );
not ( n40735 , n40734 );
not ( n40736 , n40735 );
or ( n40737 , n40736 , n18540 );
and ( n40738 , n40698 , n40737 );
and ( n40739 , n40736 , n18540 );
nor ( n40740 , n40738 , n40739 );
not ( n40741 , n831 );
not ( n40742 , n18701 );
or ( n40743 , n40741 , n40742 );
and ( n40744 , n31080 , n31655 );
buf ( n40745 , n40744 );
not ( n40746 , n40745 );
buf ( n40747 , n31817 );
not ( n40748 , n40747 );
or ( n40749 , n40746 , n40748 );
and ( n40750 , n31656 , n31646 );
buf ( n40751 , n40750 );
nand ( n40752 , n40749 , n40751 );
buf ( n40753 , n40752 );
buf ( n40754 , n40753 );
or ( n40755 , n31664 , n31980 );
buf ( n40756 , n40755 );
not ( n40757 , n40756 );
buf ( n40758 , n40757 );
buf ( n40759 , n40758 );
and ( n40760 , n40754 , n40759 );
not ( n40761 , n40754 );
buf ( n40762 , n40755 );
and ( n40763 , n40761 , n40762 );
nor ( n40764 , n40760 , n40763 );
buf ( n40765 , n40764 );
nand ( n40766 , n40765 , n1152 );
nand ( n40767 , n40743 , n40766 );
buf ( n40768 , n40767 );
buf ( n40769 , n40768 );
buf ( n40770 , n40371 );
or ( n40771 , n40769 , n40770 );
not ( n40772 , n40771 );
or ( n40773 , n40740 , n40772 );
nand ( n40774 , n40769 , n40770 );
nand ( n40775 , n40773 , n40774 );
not ( n40776 , n40775 );
or ( n40777 , n40640 , n40776 );
not ( n40778 , n831 );
not ( n40779 , n40778 );
buf ( n40780 , n32091 );
not ( n40781 , n40780 );
buf ( n40782 , n40781 );
buf ( n40783 , n31396 );
not ( n40784 , n40783 );
buf ( n40785 , n31548 );
not ( n40786 , n40785 );
or ( n40787 , n40784 , n40786 );
buf ( n40788 , n32109 );
nand ( n40789 , n40787 , n40788 );
buf ( n40790 , n40789 );
buf ( n40791 , n40790 );
buf ( n40792 , n32101 );
nand ( n40793 , n40791 , n40792 );
buf ( n40794 , n40793 );
buf ( n40795 , n32101 );
buf ( n40796 , n31393 );
not ( n40797 , n40796 );
buf ( n40798 , n40797 );
buf ( n40799 , n40798 );
buf ( n40800 , n31282 );
and ( n40801 , n40799 , n40800 );
buf ( n40802 , n40801 );
buf ( n40803 , n40802 );
buf ( n40804 , n31320 );
nand ( n40805 , n40795 , n40803 , n40804 );
buf ( n40806 , n40805 );
nand ( n40807 , n40782 , n40794 , n40806 );
buf ( n40808 , n31578 );
not ( n40809 , n40808 );
buf ( n40810 , n40809 );
buf ( n40811 , n31597 );
buf ( n40812 , n40811 );
buf ( n40813 , n40812 );
nand ( n40814 , n40810 , n40813 );
and ( n40815 , n40807 , n40814 );
not ( n40816 , n40807 );
not ( n40817 , n40814 );
and ( n40818 , n40816 , n40817 );
nor ( n40819 , n40815 , n40818 );
not ( n40820 , n40819 );
or ( n40821 , n40779 , n40820 );
buf ( n40822 , n18753 );
not ( n40823 , n40822 );
buf ( n40824 , n18715 );
buf ( n40825 , n18724 );
nand ( n40826 , n40824 , n40825 );
buf ( n40827 , n40826 );
buf ( n40828 , n40827 );
buf ( n40829 , n18715 );
buf ( n40830 , n18729 );
not ( n40831 , n40830 );
buf ( n40832 , n40831 );
buf ( n40833 , n40832 );
buf ( n40834 , n30951 );
nand ( n40835 , n40829 , n40833 , n40834 );
buf ( n40836 , n40835 );
buf ( n40837 , n40836 );
nand ( n40838 , n40823 , n40828 , n40837 );
buf ( n40839 , n40838 );
not ( n40840 , n40839 );
buf ( n40841 , n5878 );
buf ( n40842 , n10369 );
not ( n40843 , n40842 );
buf ( n40844 , n40843 );
buf ( n40845 , n40844 );
nand ( n40846 , n40841 , n40845 );
buf ( n40847 , n40846 );
not ( n40848 , n40847 );
nand ( n40849 , n40840 , n40848 );
nand ( n40850 , n40839 , n40847 );
nand ( n40851 , n40849 , n40850 , n831 );
nand ( n40852 , n40821 , n40851 );
not ( n40853 , n40852 );
buf ( n40854 , n40853 );
not ( n40855 , n40854 );
not ( n40856 , n40855 );
nor ( n40857 , n18478 , n40856 );
not ( n40858 , n831 );
buf ( n40859 , n18712 );
buf ( n40860 , n5878 );
and ( n40861 , n40859 , n40860 );
buf ( n40862 , n40861 );
buf ( n40863 , n40862 );
buf ( n40864 , n18721 );
buf ( n40865 , n8799 );
nand ( n40866 , n40864 , n40865 );
buf ( n40867 , n40866 );
buf ( n40868 , n40867 );
nand ( n40869 , n40863 , n40868 );
buf ( n40870 , n40869 );
buf ( n40871 , n40870 );
buf ( n40872 , n40862 );
buf ( n40873 , n18732 );
nand ( n40874 , n40872 , n40873 );
buf ( n40875 , n40874 );
buf ( n40876 , n40875 );
buf ( n40877 , n5878 );
not ( n40878 , n40877 );
buf ( n40879 , n18750 );
not ( n40880 , n40879 );
or ( n40881 , n40878 , n40880 );
buf ( n40882 , n40844 );
nand ( n40883 , n40881 , n40882 );
buf ( n40884 , n40883 );
buf ( n40885 , n40884 );
not ( n40886 , n40885 );
buf ( n40887 , n40886 );
buf ( n40888 , n40887 );
nand ( n40889 , n40871 , n40876 , n40888 );
buf ( n40890 , n40889 );
buf ( n40891 , n5503 );
buf ( n40892 , n10378 );
nand ( n40893 , n40891 , n40892 );
buf ( n40894 , n40893 );
and ( n40895 , n40890 , n40894 );
not ( n40896 , n40890 );
not ( n40897 , n40894 );
and ( n40898 , n40896 , n40897 );
nor ( n40899 , n40895 , n40898 );
not ( n40900 , n40899 );
or ( n40901 , n40858 , n40900 );
buf ( n40902 , n32098 );
buf ( n40903 , n40810 );
and ( n40904 , n40902 , n40903 );
buf ( n40905 , n40904 );
buf ( n40906 , n40905 );
buf ( n40907 , n40790 );
nand ( n40908 , n40906 , n40907 );
buf ( n40909 , n40908 );
buf ( n40910 , n40909 );
buf ( n40911 , n40905 );
buf ( n40912 , n31393 );
buf ( n40913 , n31279 );
nor ( n40914 , n40912 , n40913 );
buf ( n40915 , n40914 );
buf ( n40916 , n40915 );
buf ( n40917 , n30836 );
and ( n40918 , n40916 , n40917 );
buf ( n40919 , n40918 );
buf ( n40920 , n40919 );
nand ( n40921 , n40911 , n40920 );
buf ( n40922 , n40921 );
buf ( n40923 , n40922 );
buf ( n40924 , n40810 );
not ( n40925 , n40924 );
buf ( n40926 , n32088 );
not ( n40927 , n40926 );
or ( n40928 , n40925 , n40927 );
buf ( n40929 , n40813 );
nand ( n40930 , n40928 , n40929 );
buf ( n40931 , n40930 );
buf ( n40932 , n40931 );
not ( n40933 , n40932 );
buf ( n40934 , n40933 );
buf ( n40935 , n40934 );
nand ( n40936 , n40910 , n40923 , n40935 );
buf ( n40937 , n40936 );
buf ( n40938 , n31574 );
not ( n40939 , n40938 );
buf ( n40940 , n31610 );
nand ( n40941 , n40939 , n40940 );
buf ( n40942 , n40941 );
nor ( n40943 , n40937 , n40942 );
not ( n40944 , n40943 );
nand ( n40945 , n40937 , n40942 );
not ( n40946 , n831 );
nand ( n40947 , n40944 , n40945 , n40946 );
nand ( n40948 , n40901 , n40947 );
not ( n40949 , n40948 );
buf ( n40950 , n40949 );
buf ( n40951 , n40950 );
buf ( n40952 , n40720 );
and ( n40953 , n40952 , n40725 );
not ( n40954 , n40952 );
and ( n40955 , n40954 , n40722 );
nor ( n40956 , n40953 , n40955 );
nor ( n40957 , n40951 , n40956 );
nor ( n40958 , n40857 , n40957 );
not ( n40959 , n31273 );
not ( n40960 , n32088 );
or ( n40961 , n40959 , n40960 );
buf ( n40962 , n31613 );
not ( n40963 , n40962 );
buf ( n40964 , n40963 );
nand ( n40965 , n40961 , n40964 );
not ( n40966 , n40965 );
buf ( n40967 , n31273 );
buf ( n40968 , n32098 );
and ( n40969 , n40967 , n40968 );
buf ( n40970 , n40969 );
buf ( n40971 , n40970 );
buf ( n40972 , n40919 );
nand ( n40973 , n40971 , n40972 );
buf ( n40974 , n40973 );
buf ( n40975 , n40970 );
buf ( n40976 , n40790 );
nand ( n40977 , n40975 , n40976 );
buf ( n40978 , n40977 );
nand ( n40979 , n40966 , n40974 , n40978 );
not ( n40980 , n40979 );
not ( n40981 , n2206 );
not ( n40982 , n31421 );
and ( n40983 , n40982 , n31619 );
nor ( n40984 , n40981 , n40983 );
nand ( n40985 , n40980 , n40984 );
buf ( n40986 , n5884 );
not ( n40987 , n40986 );
buf ( n40988 , n18750 );
not ( n40989 , n40988 );
or ( n40990 , n40987 , n40989 );
buf ( n40991 , n10381 );
not ( n40992 , n40991 );
buf ( n40993 , n40992 );
buf ( n40994 , n40993 );
nand ( n40995 , n40990 , n40994 );
buf ( n40996 , n40995 );
not ( n40997 , n40996 );
buf ( n40998 , n18712 );
buf ( n40999 , n5884 );
and ( n41000 , n40998 , n40999 );
buf ( n41001 , n41000 );
buf ( n41002 , n41001 );
buf ( n41003 , n18732 );
nand ( n41004 , n41002 , n41003 );
buf ( n41005 , n41004 );
buf ( n41006 , n41001 );
buf ( n41007 , n40867 );
nand ( n41008 , n41006 , n41007 );
buf ( n41009 , n41008 );
nand ( n41010 , n40997 , n41005 , n41009 );
not ( n41011 , n41010 );
buf ( n41012 , n4852 );
buf ( n41013 , n5173 );
nor ( n41014 , n41012 , n41013 );
buf ( n41015 , n41014 );
buf ( n41016 , n41015 );
not ( n41017 , n41016 );
buf ( n41018 , n41017 );
buf ( n41019 , n41018 );
buf ( n41020 , n10393 );
buf ( n41021 , n41020 );
buf ( n41022 , n41021 );
buf ( n41023 , n41022 );
nand ( n41024 , n41019 , n41023 );
buf ( n41025 , n41024 );
and ( n41026 , n41025 , n831 );
nand ( n41027 , n41011 , n41026 );
buf ( n41028 , n41025 );
not ( n41029 , n41028 );
buf ( n41030 , n41029 );
nand ( n41031 , n41010 , n41030 , n831 );
and ( n41032 , n40983 , n2206 );
nand ( n41033 , n40979 , n41032 );
nand ( n41034 , n40985 , n41027 , n41031 , n41033 );
not ( n41035 , n41034 );
buf ( n41036 , n41035 );
not ( n41037 , n41036 );
not ( n41038 , n41037 );
nor ( n41039 , n18702 , n41038 );
nand ( n41040 , n10389 , n10401 );
not ( n41041 , n41040 );
buf ( n41042 , n5881 );
buf ( n41043 , n41015 );
nor ( n41044 , n41042 , n41043 );
buf ( n41045 , n41044 );
buf ( n41046 , n41045 );
not ( n41047 , n41046 );
buf ( n41048 , n18753 );
not ( n41049 , n41048 );
or ( n41050 , n41047 , n41049 );
buf ( n41051 , n41018 );
not ( n41052 , n41051 );
buf ( n41053 , n10381 );
not ( n41054 , n41053 );
or ( n41055 , n41052 , n41054 );
buf ( n41056 , n41022 );
nand ( n41057 , n41055 , n41056 );
buf ( n41058 , n41057 );
buf ( n41059 , n41058 );
not ( n41060 , n41059 );
buf ( n41061 , n41060 );
buf ( n41062 , n41061 );
nand ( n41063 , n41050 , n41062 );
buf ( n41064 , n41063 );
buf ( n41065 , n41064 );
not ( n41066 , n41065 );
buf ( n41067 , n41066 );
buf ( n41068 , n18715 );
buf ( n41069 , n41045 );
and ( n41070 , n41068 , n41069 );
buf ( n41071 , n41070 );
buf ( n41072 , n41071 );
buf ( n41073 , n18732 );
buf ( n41074 , n41073 );
nand ( n41075 , n41072 , n41074 );
buf ( n41076 , n41075 );
buf ( n41077 , n41071 );
not ( n41078 , n18724 );
not ( n41079 , n41078 );
buf ( n41080 , n41079 );
nand ( n41081 , n41077 , n41080 );
buf ( n41082 , n41081 );
nand ( n41083 , n41067 , n41076 , n41082 );
not ( n41084 , n41083 );
or ( n41085 , n41041 , n41084 );
not ( n41086 , n41040 );
nand ( n41087 , n41067 , n41076 , n41082 , n41086 );
nand ( n41088 , n41085 , n41087 );
and ( n41089 , n831 , n41088 );
not ( n41090 , n831 );
buf ( n41091 , n31551 );
buf ( n41092 , n32109 );
nand ( n41093 , n41091 , n41092 );
buf ( n41094 , n41093 );
not ( n41095 , n41094 );
buf ( n41096 , n40919 );
not ( n41097 , n41096 );
buf ( n41098 , n41097 );
nand ( n41099 , n41095 , n41098 );
not ( n41100 , n41099 );
buf ( n41101 , n32101 );
and ( n41102 , n31273 , n40982 );
buf ( n41103 , n41102 );
and ( n41104 , n41101 , n41103 );
buf ( n41105 , n41104 );
not ( n41106 , n41105 );
or ( n41107 , n41100 , n41106 );
and ( n41108 , n41102 , n32091 );
not ( n41109 , n31436 );
not ( n41110 , n31613 );
or ( n41111 , n41109 , n41110 );
nand ( n41112 , n41111 , n31619 );
nor ( n41113 , n41108 , n41112 );
nand ( n41114 , n41107 , n41113 );
buf ( n41115 , n41114 );
not ( n41116 , n31429 );
and ( n41117 , n31625 , n31405 );
nor ( n41118 , n41116 , n41117 );
buf ( n41119 , n41118 );
and ( n41120 , n41115 , n41119 );
not ( n41121 , n41115 );
buf ( n41122 , n41118 );
not ( n41123 , n41122 );
buf ( n41124 , n41123 );
buf ( n41125 , n41124 );
and ( n41126 , n41121 , n41125 );
nor ( n41127 , n41120 , n41126 );
buf ( n41128 , n41127 );
and ( n41129 , n41090 , n41128 );
nor ( n41130 , n41089 , n41129 );
not ( n41131 , n41130 );
buf ( n41132 , n41131 );
nor ( n41133 , n18670 , n41132 );
nor ( n41134 , n41039 , n41133 );
and ( n41135 , n40958 , n41134 );
not ( n41136 , n41135 );
buf ( n41137 , n31311 );
not ( n41138 , n41137 );
buf ( n41139 , n41138 );
buf ( n41140 , n41139 );
not ( n41141 , n41140 );
buf ( n41142 , n31533 );
not ( n41143 , n41142 );
or ( n41144 , n41141 , n41143 );
buf ( n41145 , n31443 );
nand ( n41146 , n41144 , n41145 );
buf ( n41147 , n41146 );
not ( n41148 , n41147 );
buf ( n41149 , n31228 );
buf ( n41150 , n41139 );
and ( n41151 , n41149 , n41150 );
buf ( n41152 , n41151 );
nand ( n41153 , n41094 , n41152 );
buf ( n41154 , n41152 );
buf ( n41155 , n40802 );
buf ( n41156 , n31879 );
nand ( n41157 , n41154 , n41155 , n41156 );
buf ( n41158 , n41157 );
nand ( n41159 , n41148 , n41153 , n41158 );
buf ( n41160 , n41159 );
buf ( n41161 , n31435 );
buf ( n41162 , n31566 );
nand ( n41163 , n41161 , n41162 );
buf ( n41164 , n41163 );
buf ( n41165 , n41164 );
not ( n41166 , n41165 );
buf ( n41167 , n41166 );
buf ( n41168 , n41167 );
and ( n41169 , n41160 , n41168 );
not ( n41170 , n41160 );
buf ( n41171 , n41164 );
and ( n41172 , n41170 , n41171 );
nor ( n41173 , n41169 , n41172 );
buf ( n41174 , n41173 );
and ( n41175 , n1152 , n41174 );
not ( n41176 , n1152 );
buf ( n41177 , n6860 );
buf ( n41178 , n8861 );
not ( n41179 , n41178 );
buf ( n41180 , n41179 );
buf ( n41181 , n41180 );
and ( n41182 , n41177 , n41181 );
buf ( n41183 , n41182 );
not ( n41184 , n41183 );
not ( n41185 , n40832 );
not ( n41186 , n30945 );
or ( n41187 , n41185 , n41186 );
nand ( n41188 , n41187 , n41078 );
not ( n41189 , n41188 );
or ( n41190 , n41184 , n41189 );
and ( n41191 , n6340 , n6352 );
not ( n41192 , n41191 );
not ( n41193 , n41180 );
buf ( n41194 , n6884 );
not ( n41195 , n41194 );
or ( n41196 , n41193 , n41195 );
buf ( n41197 , n6326 );
buf ( n41198 , n41197 );
buf ( n41199 , n41198 );
nand ( n41200 , n41196 , n41199 );
nor ( n41201 , n41192 , n41200 );
nand ( n41202 , n41190 , n41201 );
and ( n41203 , n41194 , n41180 );
not ( n41204 , n41199 );
nor ( n41205 , n41203 , n41204 );
not ( n41206 , n41205 );
not ( n41207 , n41191 );
and ( n41208 , n41206 , n41207 );
not ( n41209 , n41183 );
nor ( n41210 , n41209 , n41191 );
and ( n41211 , n41188 , n41210 );
nor ( n41212 , n41208 , n41211 );
nand ( n41213 , n41202 , n41212 );
and ( n41214 , n41176 , n41213 );
nor ( n41215 , n41175 , n41214 );
buf ( n41216 , n41215 );
not ( n41217 , n41216 );
nor ( n41218 , n10436 , n41217 );
buf ( n41219 , n31228 );
not ( n41220 , n41219 );
buf ( n41221 , n41094 );
not ( n41222 , n41221 );
or ( n41223 , n41220 , n41222 );
not ( n41224 , n31228 );
buf ( n41225 , n30833 );
buf ( n41226 , n30780 );
buf ( n41227 , n30226 );
nand ( n41228 , n41226 , n41227 );
buf ( n41229 , n41228 );
buf ( n41230 , n41229 );
and ( n41231 , n41225 , n41230 );
buf ( n41232 , n41231 );
nor ( n41233 , n41224 , n41232 );
buf ( n41234 , n41233 );
buf ( n41235 , n40802 );
and ( n41236 , n41234 , n41235 );
buf ( n41237 , n31533 );
buf ( n41238 , n41237 );
buf ( n41239 , n41238 );
buf ( n41240 , n41239 );
nor ( n41241 , n41236 , n41240 );
buf ( n41242 , n41241 );
buf ( n41243 , n41242 );
nand ( n41244 , n41223 , n41243 );
buf ( n41245 , n41244 );
not ( n41246 , n41245 );
buf ( n41247 , n31443 );
buf ( n41248 , n41139 );
nand ( n41249 , n41247 , n41248 );
buf ( n41250 , n41249 );
not ( n41251 , n831 );
and ( n41252 , n41250 , n41251 );
nand ( n41253 , n41246 , n41252 );
not ( n41254 , n6860 );
not ( n41255 , n40867 );
or ( n41256 , n41254 , n41255 );
buf ( n41257 , n40832 );
buf ( n41258 , n6863 );
buf ( n41259 , n30942 );
nor ( n41260 , n41258 , n41259 );
buf ( n41261 , n41260 );
buf ( n41262 , n41261 );
and ( n41263 , n41257 , n41262 );
buf ( n41264 , n41194 );
nor ( n41265 , n41263 , n41264 );
buf ( n41266 , n41265 );
nand ( n41267 , n41256 , n41266 );
not ( n41268 , n41267 );
buf ( n41269 , n41180 );
buf ( n41270 , n41199 );
nand ( n41271 , n41269 , n41270 );
buf ( n41272 , n41271 );
and ( n41273 , n41272 , n831 );
nand ( n41274 , n41268 , n41273 );
buf ( n41275 , n41272 );
not ( n41276 , n41275 );
buf ( n41277 , n41276 );
not ( n41278 , n41277 );
nor ( n41279 , n41278 , n41251 );
nand ( n41280 , n41267 , n41279 );
nor ( n41281 , n41250 , n831 );
nand ( n41282 , n41245 , n41281 );
nand ( n41283 , n41253 , n41274 , n41280 , n41282 );
buf ( n41284 , n41283 );
buf ( n41285 , n41284 );
not ( n41286 , n41285 );
not ( n41287 , n41286 );
not ( n41288 , n41287 );
buf ( n41289 , n41088 );
buf ( n41290 , n41289 );
or ( n41291 , n41288 , n41290 );
buf ( n41292 , n40915 );
buf ( n41293 , n30836 );
buf ( n41294 , n31219 );
not ( n41295 , n41294 );
buf ( n41296 , n41295 );
buf ( n41297 , n41296 );
nand ( n41298 , n41292 , n41293 , n41297 );
buf ( n41299 , n41298 );
buf ( n41300 , n41299 );
buf ( n41301 , n31512 );
nand ( n41302 , n41300 , n41301 );
buf ( n41303 , n41302 );
buf ( n41304 , n41303 );
not ( n41305 , n41304 );
buf ( n41306 , n40790 );
buf ( n41307 , n41296 );
nand ( n41308 , n41306 , n41307 );
buf ( n41309 , n41308 );
buf ( n41310 , n41309 );
nand ( n41311 , n41305 , n41310 );
buf ( n41312 , n41311 );
buf ( n41313 , n31530 );
buf ( n41314 , n31520 );
nand ( n41315 , n41313 , n41314 );
buf ( n41316 , n41315 );
buf ( n41317 , n41316 );
not ( n41318 , n41317 );
buf ( n41319 , n41318 );
and ( n41320 , n41312 , n41319 );
not ( n41321 , n41312 );
and ( n41322 , n41321 , n41316 );
nor ( n41323 , n41320 , n41322 );
not ( n41324 , n41323 );
not ( n41325 , n1152 );
or ( n41326 , n41324 , n41325 );
buf ( n41327 , n40867 );
buf ( n41328 , n6854 );
not ( n41329 , n41328 );
buf ( n41330 , n41329 );
buf ( n41331 , n41330 );
nand ( n41332 , n41327 , n41331 );
buf ( n41333 , n41332 );
buf ( n41334 , n41333 );
buf ( n41335 , n40832 );
buf ( n41336 , n30951 );
buf ( n41337 , n41330 );
nand ( n41338 , n41335 , n41336 , n41337 );
buf ( n41339 , n41338 );
buf ( n41340 , n41339 );
buf ( n41341 , n6867 );
nand ( n41342 , n41334 , n41340 , n41341 );
buf ( n41343 , n41342 );
buf ( n41344 , n41343 );
buf ( n41345 , n6874 );
buf ( n41346 , n41345 );
buf ( n41347 , n6883 );
buf ( n41348 , n41347 );
and ( n41349 , n41346 , n41348 );
buf ( n41350 , n41349 );
buf ( n41351 , n41350 );
and ( n41352 , n41344 , n41351 );
not ( n41353 , n41344 );
buf ( n41354 , n41350 );
not ( n41355 , n41354 );
buf ( n41356 , n41355 );
buf ( n41357 , n41356 );
and ( n41358 , n41353 , n41357 );
nor ( n41359 , n41352 , n41358 );
buf ( n41360 , n41359 );
nand ( n41361 , n41360 , n831 );
nand ( n41362 , n41326 , n41361 );
buf ( n41363 , n41362 );
buf ( n41364 , n41363 );
and ( n41365 , n41010 , n41030 );
not ( n41366 , n41010 );
and ( n41367 , n41366 , n41025 );
nor ( n41368 , n41365 , n41367 );
or ( n41369 , n41364 , n41368 );
not ( n41370 , n1152 );
buf ( n41371 , n41094 );
not ( n41372 , n41371 );
buf ( n41373 , n41098 );
nand ( n41374 , n41372 , n41373 );
buf ( n41375 , n41374 );
buf ( n41376 , n41375 );
buf ( n41377 , n41296 );
buf ( n41378 , n31512 );
nand ( n41379 , n41377 , n41378 );
buf ( n41380 , n41379 );
buf ( n41381 , n41380 );
not ( n41382 , n41381 );
buf ( n41383 , n41382 );
buf ( n41384 , n41383 );
and ( n41385 , n41376 , n41384 );
not ( n41386 , n41376 );
buf ( n41387 , n41380 );
and ( n41388 , n41386 , n41387 );
nor ( n41389 , n41385 , n41388 );
buf ( n41390 , n41389 );
not ( n41391 , n41390 );
or ( n41392 , n41370 , n41391 );
not ( n41393 , n18738 );
buf ( n41394 , n41330 );
buf ( n41395 , n6867 );
nand ( n41396 , n41394 , n41395 );
buf ( n41397 , n41396 );
nor ( n41398 , n41397 , n41251 );
and ( n41399 , n41393 , n41398 );
buf ( n41400 , n41397 );
not ( n41401 , n41400 );
buf ( n41402 , n41401 );
nor ( n41403 , n41402 , n41251 );
and ( n41404 , n18738 , n41403 );
nor ( n41405 , n41399 , n41404 );
nand ( n41406 , n41392 , n41405 );
buf ( n41407 , n41406 );
not ( n41408 , n41407 );
buf ( n41409 , n40899 );
nand ( n41410 , n41408 , n41409 );
nand ( n41411 , n41291 , n41369 , n41410 );
nor ( n41412 , n41218 , n41411 );
not ( n41413 , n41412 );
buf ( n41414 , n41360 );
buf ( n41415 , n31911 );
not ( n41416 , n41415 );
not ( n41417 , n41416 );
nor ( n41418 , n41414 , n41417 );
buf ( n41419 , n41232 );
not ( n41420 , n41419 );
buf ( n41421 , n31389 );
buf ( n41422 , n31351 );
buf ( n41423 , n41422 );
buf ( n41424 , n41423 );
buf ( n41425 , n41424 );
nor ( n41426 , n41421 , n41425 );
buf ( n41427 , n41426 );
buf ( n41428 , n41427 );
buf ( n41429 , n31282 );
nand ( n41430 , n41428 , n41429 );
buf ( n41431 , n41430 );
buf ( n41432 , n41431 );
not ( n41433 , n41432 );
and ( n41434 , n41420 , n41433 );
buf ( n41435 , n41427 );
not ( n41436 , n41435 );
buf ( n41437 , n31548 );
not ( n41438 , n41437 );
or ( n41439 , n41436 , n41438 );
buf ( n41440 , n41424 );
not ( n41441 , n41440 );
buf ( n41442 , n41441 );
buf ( n41443 , n41442 );
not ( n41444 , n41443 );
buf ( n41445 , n31481 );
not ( n41446 , n41445 );
or ( n41447 , n41444 , n41446 );
buf ( n41448 , n31492 );
not ( n41449 , n41448 );
buf ( n41450 , n41449 );
buf ( n41451 , n41450 );
nand ( n41452 , n41447 , n41451 );
buf ( n41453 , n41452 );
buf ( n41454 , n41453 );
not ( n41455 , n41454 );
buf ( n41456 , n41455 );
buf ( n41457 , n41456 );
nand ( n41458 , n41439 , n41457 );
buf ( n41459 , n41458 );
buf ( n41460 , n41459 );
nor ( n41461 , n41434 , n41460 );
buf ( n41462 , n41461 );
not ( n41463 , n41462 );
buf ( n41464 , n31487 );
buf ( n41465 , n31498 );
nand ( n41466 , n41464 , n41465 );
buf ( n41467 , n41466 );
nor ( n41468 , n41467 , n831 );
nand ( n41469 , n41463 , n41468 );
buf ( n41470 , n8848 );
not ( n41471 , n41470 );
buf ( n41472 , n8834 );
nand ( n41473 , n41471 , n41472 );
buf ( n41474 , n41473 );
buf ( n41475 , n41474 );
not ( n41476 , n41475 );
buf ( n41477 , n41476 );
nor ( n41478 , n7724 , n18425 );
buf ( n41479 , n8806 );
not ( n41480 , n41479 );
buf ( n41481 , n41480 );
nand ( n41482 , n41478 , n41481 );
buf ( n41483 , n41482 );
buf ( n41484 , n8891 );
nor ( n41485 , n41483 , n41484 );
buf ( n41486 , n41485 );
buf ( n41487 , n41486 );
not ( n41488 , n41487 );
buf ( n41489 , n30945 );
not ( n41490 , n41489 );
or ( n41491 , n41488 , n41490 );
buf ( n41492 , n41482 );
not ( n41493 , n41492 );
buf ( n41494 , n41493 );
buf ( n41495 , n41494 );
buf ( n41496 , n31856 );
and ( n41497 , n41495 , n41496 );
buf ( n41498 , n41481 );
not ( n41499 , n41498 );
buf ( n41500 , n8813 );
not ( n41501 , n41500 );
buf ( n41502 , n8820 );
not ( n41503 , n41502 );
or ( n41504 , n41501 , n41503 );
buf ( n41505 , n8825 );
nand ( n41506 , n41504 , n41505 );
buf ( n41507 , n41506 );
buf ( n41508 , n41507 );
not ( n41509 , n41508 );
or ( n41510 , n41499 , n41509 );
buf ( n41511 , n8842 );
not ( n41512 , n41511 );
buf ( n41513 , n41512 );
buf ( n41514 , n41513 );
nand ( n41515 , n41510 , n41514 );
buf ( n41516 , n41515 );
buf ( n41517 , n41516 );
nor ( n41518 , n41497 , n41517 );
buf ( n41519 , n41518 );
buf ( n41520 , n41519 );
nand ( n41521 , n41491 , n41520 );
buf ( n41522 , n41521 );
nand ( n41523 , n41477 , n41522 , n831 );
not ( n41524 , n41522 );
not ( n41525 , n831 );
nor ( n41526 , n41477 , n41525 );
nand ( n41527 , n41524 , n41526 );
nand ( n41528 , n41462 , n41467 , n41525 );
nand ( n41529 , n41469 , n41523 , n41527 , n41528 );
buf ( n41530 , n41529 );
not ( n41531 , n41530 );
buf ( n41532 , n41531 );
buf ( n41533 , n40849 );
nand ( n41534 , n41533 , n40850 );
nor ( n41535 , n41532 , n41534 );
nor ( n41536 , n41418 , n41535 );
buf ( n41537 , n31892 );
not ( n41538 , n41537 );
buf ( n41539 , n31548 );
not ( n41540 , n41539 );
or ( n41541 , n41538 , n41540 );
buf ( n41542 , n31896 );
nand ( n41543 , n41541 , n41542 );
buf ( n41544 , n41543 );
buf ( n41545 , n41544 );
buf ( n41546 , n31282 );
buf ( n41547 , n31892 );
nand ( n41548 , n41546 , n41547 );
buf ( n41549 , n41548 );
buf ( n41550 , n41549 );
buf ( n41551 , n41232 );
nor ( n41552 , n41550 , n41551 );
buf ( n41553 , n41552 );
buf ( n41554 , n41553 );
nor ( n41555 , n41545 , n41554 );
buf ( n41556 , n41555 );
buf ( n41557 , n41556 );
buf ( n41558 , n31470 );
buf ( n41559 , n31478 );
and ( n41560 , n41558 , n41559 );
buf ( n41561 , n41560 );
buf ( n41562 , n41561 );
not ( n41563 , n41562 );
buf ( n41564 , n41563 );
buf ( n41565 , n41564 );
and ( n41566 , n41557 , n41565 );
not ( n41567 , n41557 );
buf ( n41568 , n41561 );
and ( n41569 , n41567 , n41568 );
nor ( n41570 , n41566 , n41569 );
buf ( n41571 , n41570 );
nand ( n41572 , n41571 , n1152 );
nand ( n41573 , n18456 , n831 );
nand ( n41574 , n41572 , n41573 );
buf ( n41575 , n41574 );
buf ( n41576 , n41575 );
and ( n41577 , n41268 , n41272 );
not ( n41578 , n41268 );
and ( n41579 , n41578 , n41277 );
nor ( n41580 , n41577 , n41579 );
nor ( n41581 , n41576 , n41580 );
buf ( n41582 , n41213 );
not ( n41583 , n831 );
buf ( n41584 , n10359 );
not ( n41585 , n41584 );
not ( n41586 , n41478 );
nor ( n41587 , n41586 , n8891 );
buf ( n41588 , n41587 );
not ( n41589 , n41588 );
or ( n41590 , n41585 , n41589 );
not ( n41591 , n41478 );
not ( n41592 , n8798 );
or ( n41593 , n41591 , n41592 );
buf ( n41594 , n41507 );
not ( n41595 , n41594 );
buf ( n41596 , n41595 );
nand ( n41597 , n41593 , n41596 );
buf ( n41598 , n41597 );
not ( n41599 , n41598 );
buf ( n41600 , n41599 );
buf ( n41601 , n41600 );
nand ( n41602 , n41590 , n41601 );
buf ( n41603 , n41602 );
buf ( n41604 , n41603 );
buf ( n41605 , n41481 );
buf ( n41606 , n41513 );
nand ( n41607 , n41605 , n41606 );
buf ( n41608 , n41607 );
buf ( n41609 , n41608 );
not ( n41610 , n41609 );
buf ( n41611 , n41610 );
buf ( n41612 , n41611 );
and ( n41613 , n41604 , n41612 );
not ( n41614 , n41604 );
buf ( n41615 , n41608 );
and ( n41616 , n41614 , n41615 );
nor ( n41617 , n41613 , n41616 );
buf ( n41618 , n41617 );
not ( n41619 , n41618 );
or ( n41620 , n41583 , n41619 );
buf ( n41621 , n31282 );
buf ( n41622 , n31389 );
not ( n41623 , n41622 );
buf ( n41624 , n41623 );
buf ( n41625 , n41624 );
nand ( n41626 , n41621 , n41625 );
buf ( n41627 , n41626 );
buf ( n41628 , n41627 );
not ( n41629 , n41628 );
buf ( n41630 , n41232 );
not ( n41631 , n41630 );
and ( n41632 , n41629 , n41631 );
buf ( n41633 , n41624 );
not ( n41634 , n41633 );
buf ( n41635 , n31548 );
not ( n41636 , n41635 );
or ( n41637 , n41634 , n41636 );
buf ( n41638 , n31481 );
not ( n41639 , n41638 );
buf ( n41640 , n41639 );
buf ( n41641 , n41640 );
nand ( n41642 , n41637 , n41641 );
buf ( n41643 , n41642 );
buf ( n41644 , n41643 );
nor ( n41645 , n41632 , n41644 );
buf ( n41646 , n41645 );
buf ( n41647 , n41646 );
buf ( n41648 , n41442 );
buf ( n41649 , n41648 );
buf ( n41650 , n41649 );
buf ( n41651 , n41650 );
buf ( n41652 , n41450 );
nand ( n41653 , n41651 , n41652 );
buf ( n41654 , n41653 );
buf ( n41655 , n41654 );
and ( n41656 , n41647 , n41655 );
not ( n41657 , n41647 );
buf ( n41658 , n41654 );
not ( n41659 , n41658 );
buf ( n41660 , n41659 );
buf ( n41661 , n41660 );
and ( n41662 , n41657 , n41661 );
nor ( n41663 , n41656 , n41662 );
buf ( n41664 , n41663 );
nand ( n41665 , n41664 , n1152 );
nand ( n41666 , n41620 , n41665 );
buf ( n41667 , n41666 );
buf ( n41668 , n41667 );
nor ( n41669 , n41582 , n41668 );
nor ( n41670 , n41581 , n41669 );
and ( n41671 , n41536 , n41670 );
not ( n41672 , n41671 );
and ( n41673 , n18738 , n41402 );
not ( n41674 , n18738 );
and ( n41675 , n41674 , n41397 );
nor ( n41676 , n41673 , n41675 );
or ( n41677 , n30929 , n41676 );
not ( n41678 , n41677 );
not ( n41679 , n831 );
not ( n41680 , n18833 );
or ( n41681 , n41679 , n41680 );
nand ( n41682 , n41681 , n32079 );
buf ( n41683 , n41682 );
and ( n41684 , n41522 , n41477 );
not ( n41685 , n41522 );
and ( n41686 , n41685 , n41474 );
nor ( n41687 , n41684 , n41686 );
or ( n41688 , n41683 , n41687 );
not ( n41689 , n41688 );
and ( n41690 , n30964 , n18457 );
not ( n41691 , n41690 );
buf ( n41692 , n31958 );
buf ( n41693 , n41618 );
or ( n41694 , n41692 , n41693 );
not ( n41695 , n41694 );
or ( n41696 , n41691 , n41695 );
nand ( n41697 , n41692 , n41693 );
nand ( n41698 , n41696 , n41697 );
not ( n41699 , n41698 );
or ( n41700 , n41689 , n41699 );
nand ( n41701 , n41683 , n41687 );
nand ( n41702 , n41700 , n41701 );
not ( n41703 , n41702 );
or ( n41704 , n41678 , n41703 );
nand ( n41705 , n30929 , n41676 );
nand ( n41706 , n41704 , n41705 );
not ( n41707 , n41706 );
or ( n41708 , n41672 , n41707 );
buf ( n41709 , n31868 );
buf ( n41710 , n9368 );
buf ( n41711 , n9136 );
not ( n41712 , n41711 );
buf ( n41713 , n41712 );
buf ( n41714 , n41713 );
and ( n41715 , n41710 , n41714 );
buf ( n41716 , n41715 );
buf ( n41717 , n41716 );
buf ( n41718 , n9844 );
buf ( n41719 , n10255 );
nand ( n41720 , n41717 , n41718 , n41719 );
buf ( n41721 , n41720 );
buf ( n41722 , n41721 );
buf ( n41723 , n41716 );
buf ( n41724 , n10303 );
nand ( n41725 , n41723 , n41724 );
buf ( n41726 , n41725 );
buf ( n41727 , n41726 );
buf ( n41728 , n41713 );
not ( n41729 , n41728 );
buf ( n41730 , n10328 );
not ( n41731 , n41730 );
or ( n41732 , n41729 , n41731 );
buf ( n41733 , n10335 );
not ( n41734 , n41733 );
buf ( n41735 , n41734 );
buf ( n41736 , n41735 );
nand ( n41737 , n41732 , n41736 );
buf ( n41738 , n41737 );
buf ( n41739 , n41738 );
not ( n41740 , n41739 );
buf ( n41741 , n41740 );
buf ( n41742 , n41741 );
nand ( n41743 , n41722 , n41727 , n41742 );
buf ( n41744 , n41743 );
buf ( n41745 , n10351 );
not ( n41746 , n41745 );
buf ( n41747 , n10344 );
nand ( n41748 , n41746 , n41747 );
buf ( n41749 , n41748 );
buf ( n41750 , n41749 );
not ( n41751 , n41750 );
buf ( n41752 , n41751 );
and ( n41753 , n41744 , n41752 );
not ( n41754 , n41744 );
and ( n41755 , n41754 , n41749 );
nor ( n41756 , n41753 , n41755 );
and ( n41757 , n831 , n41756 );
not ( n41758 , n831 );
buf ( n41759 , n30799 );
not ( n41760 , n41759 );
buf ( n41761 , n30777 );
not ( n41762 , n41761 );
or ( n41763 , n41760 , n41762 );
buf ( n41764 , n30817 );
not ( n41765 , n41764 );
buf ( n41766 , n41765 );
buf ( n41767 , n41766 );
nand ( n41768 , n41763 , n41767 );
buf ( n41769 , n41768 );
buf ( n41770 , n41769 );
not ( n41771 , n41770 );
buf ( n41772 , n30761 );
buf ( n41773 , n30777 );
and ( n41774 , n41772 , n41773 );
buf ( n41775 , n41774 );
buf ( n41776 , n41775 );
buf ( n41777 , n30171 );
buf ( n41778 , n30101 );
nand ( n41779 , n41776 , n41777 , n41778 );
buf ( n41780 , n41779 );
buf ( n41781 , n41780 );
buf ( n41782 , n41775 );
buf ( n41783 , n30223 );
not ( n41784 , n41783 );
buf ( n41785 , n41784 );
buf ( n41786 , n41785 );
nand ( n41787 , n41782 , n41786 );
buf ( n41788 , n41787 );
buf ( n41789 , n41788 );
nand ( n41790 , n41771 , n41781 , n41789 );
buf ( n41791 , n41790 );
buf ( n41792 , n30824 );
not ( n41793 , n41792 );
buf ( n41794 , n30741 );
nand ( n41795 , n41793 , n41794 );
buf ( n41796 , n41795 );
xnor ( n41797 , n41791 , n41796 );
and ( n41798 , n41758 , n41797 );
nor ( n41799 , n41757 , n41798 );
not ( n41800 , n41799 );
buf ( n41801 , n41800 );
buf ( n41802 , n41801 );
or ( n41803 , n41709 , n41802 );
not ( n41804 , n41803 );
buf ( n41805 , n30669 );
not ( n41806 , n831 );
buf ( n41807 , n10328 );
not ( n41808 , n41807 );
buf ( n41809 , n10303 );
buf ( n41810 , n9368 );
nand ( n41811 , n41809 , n41810 );
buf ( n41812 , n41811 );
buf ( n41813 , n41812 );
buf ( n41814 , n9844 );
buf ( n41815 , n9368 );
buf ( n41816 , n10255 );
nand ( n41817 , n41814 , n41815 , n41816 );
buf ( n41818 , n41817 );
buf ( n41819 , n41818 );
nand ( n41820 , n41808 , n41813 , n41819 );
buf ( n41821 , n41820 );
buf ( n41822 , n41821 );
buf ( n41823 , n41713 );
buf ( n41824 , n41735 );
nand ( n41825 , n41823 , n41824 );
buf ( n41826 , n41825 );
buf ( n41827 , n41826 );
not ( n41828 , n41827 );
buf ( n41829 , n41828 );
buf ( n41830 , n41829 );
and ( n41831 , n41822 , n41830 );
not ( n41832 , n41822 );
buf ( n41833 , n41826 );
and ( n41834 , n41832 , n41833 );
nor ( n41835 , n41831 , n41834 );
buf ( n41836 , n41835 );
not ( n41837 , n41836 );
or ( n41838 , n41806 , n41837 );
buf ( n41839 , n41785 );
buf ( n41840 , n30761 );
buf ( n41841 , n41840 );
buf ( n41842 , n41841 );
buf ( n41843 , n41842 );
nand ( n41844 , n41839 , n41843 );
buf ( n41845 , n41844 );
buf ( n41846 , n30171 );
buf ( n41847 , n41842 );
buf ( n41848 , n30101 );
nand ( n41849 , n41846 , n41847 , n41848 );
buf ( n41850 , n41849 );
not ( n41851 , n30799 );
nand ( n41852 , n41845 , n41850 , n41851 );
nand ( n41853 , n41766 , n30777 );
not ( n41854 , n41853 );
and ( n41855 , n41852 , n41854 );
not ( n41856 , n41852 );
and ( n41857 , n41856 , n41853 );
nor ( n41858 , n41855 , n41857 );
nand ( n41859 , n41858 , n1152 );
nand ( n41860 , n41838 , n41859 );
buf ( n41861 , n41860 );
nor ( n41862 , n41805 , n41861 );
not ( n41863 , n41862 );
not ( n41864 , n41863 );
nand ( n41865 , n31956 , n30259 );
not ( n41866 , n41865 );
not ( n41867 , n41866 );
buf ( n41868 , n10303 );
buf ( n41869 , n18544 );
nand ( n41870 , n41868 , n41869 );
buf ( n41871 , n41870 );
buf ( n41872 , n41871 );
buf ( n41873 , n9844 );
buf ( n41874 , n10255 );
buf ( n41875 , n18544 );
nand ( n41876 , n41873 , n41874 , n41875 );
buf ( n41877 , n41876 );
buf ( n41878 , n41877 );
buf ( n41879 , n10319 );
nand ( n41880 , n41872 , n41878 , n41879 );
buf ( n41881 , n41880 );
buf ( n41882 , n41881 );
buf ( n41883 , n10314 );
not ( n41884 , n41883 );
buf ( n41885 , n10325 );
nand ( n41886 , n41884 , n41885 );
buf ( n41887 , n41886 );
buf ( n41888 , n41887 );
not ( n41889 , n41888 );
buf ( n41890 , n41889 );
buf ( n41891 , n41890 );
and ( n41892 , n41882 , n41891 );
not ( n41893 , n41882 );
buf ( n41894 , n41887 );
and ( n41895 , n41893 , n41894 );
nor ( n41896 , n41892 , n41895 );
buf ( n41897 , n41896 );
and ( n41898 , n831 , n41897 );
not ( n41899 , n831 );
buf ( n41900 , n30223 );
not ( n41901 , n41900 );
buf ( n41902 , n30244 );
nand ( n41903 , n41901 , n41902 );
buf ( n41904 , n41903 );
buf ( n41905 , n41904 );
buf ( n41906 , n30171 );
buf ( n41907 , n30101 );
buf ( n41908 , n30244 );
nand ( n41909 , n41906 , n41907 , n41908 );
buf ( n41910 , n41909 );
buf ( n41911 , n41910 );
buf ( n41912 , n30252 );
nand ( n41913 , n41905 , n41911 , n41912 );
buf ( n41914 , n41913 );
buf ( n41915 , n41914 );
buf ( n41916 , n30789 );
not ( n41917 , n41916 );
buf ( n41918 , n30796 );
nand ( n41919 , n41917 , n41918 );
buf ( n41920 , n41919 );
buf ( n41921 , n41920 );
not ( n41922 , n41921 );
buf ( n41923 , n41922 );
buf ( n41924 , n41923 );
and ( n41925 , n41915 , n41924 );
not ( n41926 , n41915 );
buf ( n41927 , n41920 );
and ( n41928 , n41926 , n41927 );
nor ( n41929 , n41925 , n41928 );
buf ( n41930 , n41929 );
and ( n41931 , n41899 , n41930 );
nor ( n41932 , n41898 , n41931 );
not ( n41933 , n41932 );
nor ( n41934 , n18834 , n41933 );
not ( n41935 , n41934 );
not ( n41936 , n41935 );
or ( n41937 , n41867 , n41936 );
not ( n41938 , n41933 );
not ( n41939 , n41938 );
nand ( n41940 , n18834 , n41939 );
nand ( n41941 , n41937 , n41940 );
not ( n41942 , n41941 );
nor ( n41943 , n30956 , n30351 );
buf ( n41944 , n41756 );
not ( n41945 , n30525 );
buf ( n41946 , n41945 );
or ( n41947 , n41944 , n41946 );
buf ( n41948 , n30577 );
nor ( n41949 , n41836 , n41948 );
not ( n41950 , n41949 );
nand ( n41951 , n41947 , n41950 );
nor ( n41952 , n41943 , n41951 );
not ( n41953 , n41952 );
buf ( n41954 , n30465 );
xor ( n41955 , n41954 , n18554 );
buf ( n41956 , n30022 );
buf ( n41957 , n30071 );
not ( n41958 , n41957 );
buf ( n41959 , n41958 );
buf ( n41960 , n41959 );
nand ( n41961 , n41956 , n41960 );
buf ( n41962 , n41961 );
buf ( n41963 , n41962 );
buf ( n41964 , n30082 );
buf ( n41965 , n30448 );
nand ( n41966 , n41964 , n41965 );
buf ( n41967 , n41966 );
buf ( n41968 , n41967 );
not ( n41969 , n41968 );
buf ( n41970 , n41969 );
buf ( n41971 , n41970 );
and ( n41972 , n41963 , n41971 );
not ( n41973 , n41963 );
buf ( n41974 , n41967 );
and ( n41975 , n41973 , n41974 );
nor ( n41976 , n41972 , n41975 );
buf ( n41977 , n41976 );
and ( n41978 , n1152 , n41977 );
not ( n41979 , n1152 );
buf ( n41980 , n10242 );
not ( n41981 , n41980 );
buf ( n41982 , n41981 );
buf ( n41983 , n41982 );
buf ( n41984 , n10135 );
not ( n41985 , n41984 );
buf ( n41986 , n41985 );
buf ( n41987 , n41986 );
nand ( n41988 , n41983 , n41987 );
buf ( n41989 , n41988 );
buf ( n41990 , n41989 );
buf ( n41991 , n10143 );
buf ( n41992 , n9997 );
nand ( n41993 , n41991 , n41992 );
buf ( n41994 , n41993 );
buf ( n41995 , n41994 );
not ( n41996 , n41995 );
buf ( n41997 , n41996 );
buf ( n41998 , n41997 );
and ( n41999 , n41990 , n41998 );
not ( n42000 , n41990 );
buf ( n42001 , n41994 );
and ( n42002 , n42000 , n42001 );
nor ( n42003 , n41999 , n42002 );
buf ( n42004 , n42003 );
and ( n42005 , n41979 , n42004 );
or ( n42006 , n41978 , n42005 );
buf ( n42007 , n42006 );
or ( n42008 , n30348 , n42007 );
not ( n42009 , n42008 );
not ( n42010 , n1152 );
buf ( n42011 , n32040 );
not ( n42012 , n42011 );
buf ( n42013 , n30021 );
not ( n42014 , n42013 );
or ( n42015 , n42012 , n42014 );
buf ( n42016 , n30062 );
nand ( n42017 , n42015 , n42016 );
buf ( n42018 , n42017 );
buf ( n42019 , n42018 );
buf ( n42020 , n30057 );
not ( n42021 , n42020 );
buf ( n42022 , n30068 );
nand ( n42023 , n42021 , n42022 );
buf ( n42024 , n42023 );
buf ( n42025 , n42024 );
not ( n42026 , n42025 );
buf ( n42027 , n42026 );
buf ( n42028 , n42027 );
and ( n42029 , n42019 , n42028 );
not ( n42030 , n42019 );
buf ( n42031 , n42024 );
and ( n42032 , n42030 , n42031 );
nor ( n42033 , n42029 , n42032 );
buf ( n42034 , n42033 );
not ( n42035 , n42034 );
or ( n42036 , n42010 , n42035 );
nand ( n42037 , n42036 , n32035 );
buf ( n42038 , n42037 );
or ( n42039 , n30523 , n42038 );
not ( n42040 , n42039 );
not ( n42041 , n831 );
buf ( n42042 , n32008 );
buf ( n42043 , n10123 );
nand ( n42044 , n42042 , n42043 );
buf ( n42045 , n42044 );
xor ( n42046 , n30391 , n42045 );
not ( n42047 , n42046 );
or ( n42048 , n42041 , n42047 );
nand ( n42049 , n42048 , n32055 );
buf ( n42050 , n42049 );
or ( n42051 , n30575 , n42050 );
not ( n42052 , n42051 );
or ( n42053 , n30366 , n30610 );
not ( n42054 , n42053 );
not ( n42055 , n30418 );
not ( n42056 , n30633 );
nand ( n42057 , n42055 , n42056 );
not ( n42058 , n42057 );
nor ( n42059 , n42004 , n1213 );
not ( n42060 , n831 );
xor ( n42061 , n1183 , n863 );
not ( n42062 , n42061 );
or ( n42063 , n42060 , n42062 );
nand ( n42064 , n895 , n1152 );
nand ( n42065 , n42063 , n42064 );
nand ( n42066 , n32034 , n42065 );
or ( n42067 , n42059 , n42066 );
nand ( n42068 , n42004 , n1213 );
nand ( n42069 , n42067 , n42068 );
not ( n42070 , n42069 );
or ( n42071 , n42058 , n42070 );
nand ( n42072 , n30633 , n30418 );
nand ( n42073 , n42071 , n42072 );
not ( n42074 , n42073 );
or ( n42075 , n42054 , n42074 );
nand ( n42076 , n30366 , n30610 );
nand ( n42077 , n42075 , n42076 );
not ( n42078 , n42077 );
or ( n42079 , n42052 , n42078 );
nand ( n42080 , n30575 , n42050 );
nand ( n42081 , n42079 , n42080 );
not ( n42082 , n42081 );
or ( n42083 , n42040 , n42082 );
nand ( n42084 , n30523 , n42038 );
nand ( n42085 , n42083 , n42084 );
not ( n42086 , n42085 );
or ( n42087 , n42009 , n42086 );
nand ( n42088 , n30348 , n42007 );
nand ( n42089 , n42087 , n42088 );
and ( n42090 , n41955 , n42089 );
and ( n42091 , n41954 , n18554 );
or ( n42092 , n42090 , n42091 );
or ( n42093 , n41897 , n30379 );
and ( n42094 , n42092 , n42093 );
not ( n42095 , n42094 );
or ( n42096 , n41953 , n42095 );
not ( n42097 , n41943 );
nand ( n42098 , n41897 , n30379 );
or ( n42099 , n41949 , n42098 );
nand ( n42100 , n41836 , n41948 );
nand ( n42101 , n42099 , n42100 );
not ( n42102 , n42101 );
not ( n42103 , n41947 );
or ( n42104 , n42102 , n42103 );
nand ( n42105 , n41944 , n41946 );
nand ( n42106 , n42104 , n42105 );
and ( n42107 , n42097 , n42106 );
and ( n42108 , n30956 , n30351 );
nor ( n42109 , n42107 , n42108 );
nand ( n42110 , n42096 , n42109 );
nor ( n42111 , n31956 , n30259 );
nor ( n42112 , n41934 , n42111 );
nand ( n42113 , n42110 , n42112 );
nand ( n42114 , n41942 , n42113 );
not ( n42115 , n42114 );
or ( n42116 , n41864 , n42115 );
nand ( n42117 , n41805 , n41861 );
nand ( n42118 , n42116 , n42117 );
not ( n42119 , n42118 );
or ( n42120 , n41804 , n42119 );
nand ( n42121 , n41709 , n41802 );
nand ( n42122 , n42120 , n42121 );
or ( n42123 , n30964 , n18457 );
and ( n42124 , n41677 , n41688 , n41694 , n42123 );
and ( n42125 , n42122 , n42124 );
and ( n42126 , n42125 , n41671 );
not ( n42127 , n41416 );
nand ( n42128 , n41414 , n42127 );
or ( n42129 , n41581 , n42128 );
nand ( n42130 , n41576 , n41580 );
nand ( n42131 , n42129 , n42130 );
not ( n42132 , n41669 );
and ( n42133 , n42131 , n42132 );
nand ( n42134 , n41582 , n41668 );
not ( n42135 , n42134 );
nor ( n42136 , n42133 , n42135 );
or ( n42137 , n42136 , n41535 );
nand ( n42138 , n41534 , n41532 );
nand ( n42139 , n42137 , n42138 );
nor ( n42140 , n42126 , n42139 );
nand ( n42141 , n41708 , n42140 );
not ( n42142 , n42141 );
or ( n42143 , n41413 , n42142 );
not ( n42144 , n41291 );
not ( n42145 , n41407 );
nor ( n42146 , n42145 , n41409 );
not ( n42147 , n42146 );
not ( n42148 , n41369 );
or ( n42149 , n42147 , n42148 );
buf ( n42150 , n41364 );
nand ( n42151 , n42150 , n41368 );
nand ( n42152 , n42149 , n42151 );
not ( n42153 , n42152 );
or ( n42154 , n42144 , n42153 );
nand ( n42155 , n41288 , n41290 );
nand ( n42156 , n42154 , n42155 );
not ( n42157 , n41218 );
and ( n42158 , n42156 , n42157 );
and ( n42159 , n10436 , n41217 );
nor ( n42160 , n42158 , n42159 );
nand ( n42161 , n42143 , n42160 );
not ( n42162 , n42161 );
or ( n42163 , n41136 , n42162 );
nand ( n42164 , n18478 , n40856 );
or ( n42165 , n42164 , n40957 );
nand ( n42166 , n40951 , n40956 );
nand ( n42167 , n42165 , n42166 );
not ( n42168 , n42167 );
not ( n42169 , n41039 );
not ( n42170 , n42169 );
or ( n42171 , n42168 , n42170 );
nand ( n42172 , n18702 , n41038 );
nand ( n42173 , n42171 , n42172 );
not ( n42174 , n41133 );
and ( n42175 , n42173 , n42174 );
and ( n42176 , n18670 , n41132 );
nor ( n42177 , n42175 , n42176 );
nand ( n42178 , n42163 , n42177 );
or ( n42179 , n40692 , n40693 );
and ( n42180 , n40771 , n40678 , n40737 , n42179 );
and ( n42181 , n42178 , n42180 , n40639 );
not ( n42182 , n40630 );
and ( n42183 , n40529 , n40533 );
not ( n42184 , n42183 );
not ( n42185 , n40594 );
or ( n42186 , n42184 , n42185 );
nand ( n42187 , n40592 , n40593 );
nand ( n42188 , n42186 , n42187 );
not ( n42189 , n42188 );
or ( n42190 , n42182 , n42189 );
nand ( n42191 , n40628 , n40629 );
nand ( n42192 , n42190 , n42191 );
and ( n42193 , n42192 , n40637 );
and ( n42194 , n40636 , n18422 );
nor ( n42195 , n42193 , n42194 );
not ( n42196 , n42195 );
nor ( n42197 , n42181 , n42196 );
nand ( n42198 , n40777 , n42197 );
not ( n42199 , n42198 );
or ( n42200 , n40521 , n42199 );
not ( n42201 , n40151 );
not ( n42202 , n40365 );
nand ( n42203 , n16777 , n40377 );
not ( n42204 , n42203 );
not ( n42205 , n42204 );
not ( n42206 , n40283 );
or ( n42207 , n42205 , n42206 );
nand ( n42208 , n40226 , n40282 );
nand ( n42209 , n42207 , n42208 );
not ( n42210 , n42209 );
or ( n42211 , n42202 , n42210 );
nand ( n42212 , n40364 , n16710 );
nand ( n42213 , n42211 , n42212 );
not ( n42214 , n42213 );
or ( n42215 , n42201 , n42214 );
nand ( n42216 , n40149 , n40150 );
nand ( n42217 , n42215 , n42216 );
and ( n42218 , n42217 , n40519 );
not ( n42219 , n40387 );
and ( n42220 , n40389 , n18802 );
not ( n42221 , n42220 );
or ( n42222 , n42219 , n42221 );
nand ( n42223 , n40382 , n40386 );
nand ( n42224 , n42222 , n42223 );
and ( n42225 , n42224 , n40453 );
and ( n42226 , n40452 , n18607 );
nor ( n42227 , n42225 , n42226 );
not ( n42228 , n40517 );
or ( n42229 , n42227 , n42228 );
nand ( n42230 , n40515 , n40516 );
nand ( n42231 , n42229 , n42230 );
nor ( n42232 , n42218 , n42231 );
nand ( n42233 , n42200 , n42232 );
not ( n42234 , n42233 );
or ( n42235 , n40021 , n42234 );
not ( n42236 , n39853 );
nand ( n42237 , n40012 , n40017 );
or ( n42238 , n42237 , n39965 );
nand ( n42239 , n39964 , n18377 );
nand ( n42240 , n42238 , n42239 );
not ( n42241 , n42240 );
or ( n42242 , n42236 , n42241 );
nand ( n42243 , n39847 , n39852 );
nand ( n42244 , n42242 , n42243 );
and ( n42245 , n42244 , n39901 );
and ( n42246 , n39896 , n39900 );
nor ( n42247 , n42245 , n42246 );
nand ( n42248 , n42235 , n42247 );
not ( n42249 , n42248 );
or ( n42250 , n39787 , n42249 );
not ( n42251 , n39718 );
not ( n42252 , n39682 );
nand ( n42253 , n39784 , n39779 );
not ( n42254 , n42253 );
not ( n42255 , n42254 );
or ( n42256 , n42252 , n42255 );
nand ( n42257 , n39681 , n39603 );
nand ( n42258 , n42256 , n42257 );
not ( n42259 , n42258 );
or ( n42260 , n42251 , n42259 );
nand ( n42261 , n39716 , n39717 );
nand ( n42262 , n42260 , n42261 );
and ( n42263 , n42262 , n39601 );
and ( n42264 , n39575 , n39600 );
nor ( n42265 , n42263 , n42264 );
nand ( n42266 , n42250 , n42265 );
not ( n42267 , n42266 );
or ( n42268 , n39437 , n42267 );
not ( n42269 , n39254 );
nand ( n42270 , n39335 , n39433 );
not ( n42271 , n42270 );
and ( n42272 , n42269 , n42271 );
not ( n42273 , n38981 );
nand ( n42274 , n39056 , n39099 );
not ( n42275 , n42274 );
and ( n42276 , n42273 , n42275 );
and ( n42277 , n38500 , n38980 );
nor ( n42278 , n42276 , n42277 );
nor ( n42279 , n42278 , n39435 );
nor ( n42280 , n42272 , n42279 );
nand ( n42281 , n42268 , n42280 );
not ( n42282 , n1152 );
not ( n42283 , n31968 );
buf ( n42284 , n39242 );
not ( n42285 , n42284 );
buf ( n42286 , n42285 );
buf ( n42287 , n42286 );
buf ( n42288 , n39015 );
buf ( n42289 , n39185 );
buf ( n42290 , n39197 );
buf ( n42291 , n39169 );
nor ( n42292 , n42290 , n42291 );
buf ( n42293 , n42292 );
buf ( n42294 , n42293 );
and ( n42295 , n42289 , n42294 );
buf ( n42296 , n42295 );
buf ( n42297 , n42296 );
not ( n42298 , n42297 );
buf ( n42299 , n42298 );
buf ( n42300 , n42299 );
and ( n42301 , n39163 , n39164 );
buf ( n42302 , n42301 );
buf ( n42303 , n42302 );
buf ( n42304 , n38836 );
buf ( n42305 , n38842 );
xor ( n42306 , n42304 , n42305 );
buf ( n42307 , n42306 );
buf ( n42308 , n42307 );
nor ( n42309 , n42303 , n42308 );
buf ( n42310 , n42309 );
buf ( n42311 , n42310 );
nor ( n42312 , n42300 , n42311 );
buf ( n42313 , n42312 );
buf ( n42314 , n42313 );
nand ( n42315 , n42288 , n42314 );
buf ( n42316 , n42315 );
buf ( n42317 , n42316 );
nor ( n42318 , n42287 , n42317 );
buf ( n42319 , n42318 );
not ( n42320 , n42319 );
or ( n42321 , n42283 , n42320 );
buf ( n42322 , n42313 );
buf ( n42323 , n38230 );
and ( n42324 , n42322 , n42323 );
buf ( n42325 , n42310 );
not ( n42326 , n42325 );
buf ( n42327 , n42326 );
buf ( n42328 , n42327 );
not ( n42329 , n42328 );
buf ( n42330 , n42293 );
not ( n42331 , n42330 );
buf ( n42332 , n39213 );
not ( n42333 , n42332 );
or ( n42334 , n42331 , n42333 );
buf ( n42335 , n39223 );
buf ( n42336 , n39172 );
and ( n42337 , n42335 , n42336 );
buf ( n42338 , n39177 );
not ( n42339 , n42338 );
buf ( n42340 , n42339 );
buf ( n42341 , n42340 );
nor ( n42342 , n42337 , n42341 );
buf ( n42343 , n42342 );
buf ( n42344 , n42343 );
nand ( n42345 , n42334 , n42344 );
buf ( n42346 , n42345 );
buf ( n42347 , n42346 );
not ( n42348 , n42347 );
or ( n42349 , n42329 , n42348 );
buf ( n42350 , n42302 );
buf ( n42351 , n42307 );
nand ( n42352 , n42350 , n42351 );
buf ( n42353 , n42352 );
buf ( n42354 , n42353 );
nand ( n42355 , n42349 , n42354 );
buf ( n42356 , n42355 );
buf ( n42357 , n42356 );
nor ( n42358 , n42324 , n42357 );
buf ( n42359 , n42358 );
nand ( n42360 , n42321 , n42359 );
and ( n42361 , n42304 , n42305 );
buf ( n42362 , n42361 );
buf ( n42363 , n42362 );
buf ( n42364 , n38601 );
buf ( n42365 , n38718 );
xor ( n42366 , n42364 , n42365 );
buf ( n42367 , n42366 );
buf ( n42368 , n42367 );
nor ( n42369 , n42363 , n42368 );
buf ( n42370 , n42369 );
buf ( n42371 , n42370 );
not ( n42372 , n42371 );
buf ( n42373 , n42362 );
buf ( n42374 , n42367 );
nand ( n42375 , n42373 , n42374 );
buf ( n42376 , n42375 );
buf ( n42377 , n42376 );
nand ( n42378 , n42372 , n42377 );
buf ( n42379 , n42378 );
nor ( n42380 , n42360 , n42379 );
not ( n42381 , n42380 );
buf ( n42382 , n39011 );
not ( n42383 , n42382 );
buf ( n42384 , n42383 );
nor ( n42385 , n42316 , n42384 );
not ( n42386 , n42385 );
not ( n42387 , n42386 );
or ( n42388 , n42381 , n42387 );
or ( n42389 , n42385 , n42360 );
nand ( n42390 , n42389 , n42379 );
nand ( n42391 , n42388 , n42390 );
not ( n42392 , n42391 );
or ( n42393 , n42282 , n42392 );
nand ( n42394 , n39069 , n39074 , n39091 , n39094 );
nand ( n42395 , n39092 , n39095 );
nand ( n42396 , n42394 , n42395 , n831 );
nand ( n42397 , n42393 , n42396 );
not ( n42398 , n42397 );
buf ( n42399 , n42398 );
not ( n42400 , n42399 );
buf ( n42401 , n42400 );
not ( n42402 , n42401 );
buf ( n42403 , n42327 );
buf ( n42404 , n42353 );
nand ( n42405 , n42403 , n42404 );
buf ( n42406 , n42405 );
and ( n42407 , n1152 , n42406 );
not ( n42408 , n42407 );
not ( n42409 , n42408 );
buf ( n42410 , n37762 );
buf ( n42411 , n37995 );
buf ( n42412 , n39185 );
buf ( n42413 , n42293 );
and ( n42414 , n42412 , n42413 );
buf ( n42415 , n42414 );
buf ( n42416 , n42415 );
and ( n42417 , n42411 , n42416 );
buf ( n42418 , n42417 );
buf ( n42419 , n42418 );
nand ( n42420 , n42410 , n42419 );
buf ( n42421 , n42420 );
buf ( n42422 , n42415 );
not ( n42423 , n42422 );
buf ( n42424 , n38230 );
not ( n42425 , n42424 );
or ( n42426 , n42423 , n42425 );
buf ( n42427 , n42346 );
not ( n42428 , n42427 );
buf ( n42429 , n42428 );
buf ( n42430 , n42429 );
nand ( n42431 , n42426 , n42430 );
buf ( n42432 , n42431 );
buf ( n42433 , n42432 );
not ( n42434 , n42433 );
buf ( n42435 , n42434 );
buf ( n42436 , n38136 );
buf ( n42437 , n42418 );
and ( n42438 , n42436 , n42437 );
buf ( n42439 , n42438 );
buf ( n42440 , n42439 );
buf ( n42441 , n31968 );
nand ( n42442 , n42440 , n42441 );
buf ( n42443 , n42442 );
nand ( n42444 , n42421 , n42435 , n42443 );
not ( n42445 , n42444 );
or ( n42446 , n42409 , n42445 );
not ( n42447 , n1152 );
nor ( n42448 , n42447 , n42406 );
not ( n42449 , n42448 );
nand ( n42450 , n42449 , n42421 , n42435 , n42443 );
nand ( n42451 , n42446 , n42450 );
or ( n42452 , n39590 , n39599 );
nand ( n42453 , n42452 , n831 );
not ( n42454 , n42453 );
nand ( n42455 , n39590 , n39588 , n39594 , n39599 );
or ( n42456 , n39588 , n39599 );
or ( n42457 , n39594 , n39599 );
nand ( n42458 , n42454 , n42455 , n42456 , n42457 );
nand ( n42459 , n42451 , n42458 );
buf ( n42460 , n42459 );
not ( n42461 , n42460 );
nor ( n42462 , n42402 , n42461 );
nand ( n42463 , n42281 , n42462 );
and ( n42464 , n831 , n38980 );
not ( n42465 , n831 );
buf ( n42466 , n42384 );
not ( n42467 , n42466 );
buf ( n42468 , n39015 );
buf ( n42469 , n42310 );
buf ( n42470 , n42370 );
nor ( n42471 , n42469 , n42470 );
buf ( n42472 , n42471 );
buf ( n42473 , n42472 );
not ( n42474 , n42473 );
buf ( n42475 , n42299 );
nor ( n42476 , n42474 , n42475 );
buf ( n42477 , n42476 );
buf ( n42478 , n42477 );
nand ( n42479 , n42468 , n42478 );
buf ( n42480 , n42479 );
buf ( n42481 , n42480 );
not ( n42482 , n42481 );
and ( n42483 , n42467 , n42482 );
buf ( n42484 , n42286 );
buf ( n42485 , n42480 );
nor ( n42486 , n42484 , n42485 );
buf ( n42487 , n42486 );
buf ( n42488 , n42487 );
not ( n42489 , n42488 );
buf ( n42490 , n31968 );
not ( n42491 , n42490 );
or ( n42492 , n42489 , n42491 );
buf ( n42493 , n42477 );
buf ( n42494 , n39042 );
and ( n42495 , n42493 , n42494 );
buf ( n42496 , n42472 );
not ( n42497 , n42496 );
buf ( n42498 , n42346 );
not ( n42499 , n42498 );
or ( n42500 , n42497 , n42499 );
buf ( n42501 , n42353 );
buf ( n42502 , n42370 );
or ( n42503 , n42501 , n42502 );
buf ( n42504 , n42376 );
nand ( n42505 , n42503 , n42504 );
buf ( n42506 , n42505 );
buf ( n42507 , n42506 );
not ( n42508 , n42507 );
buf ( n42509 , n42508 );
buf ( n42510 , n42509 );
nand ( n42511 , n42500 , n42510 );
buf ( n42512 , n42511 );
buf ( n42513 , n42512 );
nor ( n42514 , n42495 , n42513 );
buf ( n42515 , n42514 );
buf ( n42516 , n42515 );
nand ( n42517 , n42492 , n42516 );
buf ( n42518 , n42517 );
buf ( n42519 , n42518 );
nor ( n42520 , n42483 , n42519 );
buf ( n42521 , n42520 );
buf ( n42522 , n42521 );
and ( n42523 , n42364 , n42365 );
buf ( n42524 , n42523 );
buf ( n42525 , n42524 );
buf ( n42526 , n38745 );
buf ( n42527 , n38751 );
xor ( n42528 , n42526 , n42527 );
buf ( n42529 , n42528 );
buf ( n42530 , n42529 );
and ( n42531 , n42525 , n42530 );
buf ( n42532 , n42531 );
buf ( n42533 , n42532 );
not ( n42534 , n42533 );
buf ( n42535 , n42524 );
buf ( n42536 , n42529 );
or ( n42537 , n42535 , n42536 );
buf ( n42538 , n42537 );
buf ( n42539 , n42538 );
nand ( n42540 , n42534 , n42539 );
buf ( n42541 , n42540 );
buf ( n42542 , n42541 );
and ( n42543 , n42522 , n42542 );
not ( n42544 , n42522 );
buf ( n42545 , n42541 );
not ( n42546 , n42545 );
buf ( n42547 , n42546 );
buf ( n42548 , n42547 );
and ( n42549 , n42544 , n42548 );
nor ( n42550 , n42543 , n42549 );
buf ( n42551 , n42550 );
and ( n42552 , n42465 , n42551 );
nor ( n42553 , n42464 , n42552 );
not ( n42554 , n42553 );
buf ( n42555 , n42554 );
buf ( n42556 , n42555 );
buf ( n42557 , n42556 );
not ( n42558 , n42557 );
nor ( n42559 , n42463 , n42558 );
not ( n42560 , n831 );
not ( n42561 , n39432 );
or ( n42562 , n42560 , n42561 );
not ( n42563 , n831 );
buf ( n42564 , n42384 );
not ( n42565 , n42564 );
buf ( n42566 , n39015 );
buf ( n42567 , n42299 );
buf ( n42568 , n42472 );
buf ( n42569 , n42538 );
nand ( n42570 , n42568 , n42569 );
buf ( n42571 , n42570 );
buf ( n42572 , n42571 );
nor ( n42573 , n42567 , n42572 );
buf ( n42574 , n42573 );
buf ( n42575 , n42574 );
nand ( n42576 , n42566 , n42575 );
buf ( n42577 , n42576 );
buf ( n42578 , n42577 );
not ( n42579 , n42578 );
and ( n42580 , n42565 , n42579 );
buf ( n42581 , n42286 );
buf ( n42582 , n42577 );
nor ( n42583 , n42581 , n42582 );
buf ( n42584 , n42583 );
buf ( n42585 , n42584 );
not ( n42586 , n42585 );
buf ( n42587 , n31968 );
not ( n42588 , n42587 );
or ( n42589 , n42586 , n42588 );
buf ( n42590 , n42574 );
not ( n42591 , n42590 );
buf ( n42592 , n39042 );
not ( n42593 , n42592 );
or ( n42594 , n42591 , n42593 );
buf ( n42595 , n42571 );
not ( n42596 , n42595 );
buf ( n42597 , n42596 );
buf ( n42598 , n42597 );
not ( n42599 , n42598 );
buf ( n42600 , n42346 );
not ( n42601 , n42600 );
or ( n42602 , n42599 , n42601 );
buf ( n42603 , n42506 );
buf ( n42604 , n42538 );
and ( n42605 , n42603 , n42604 );
buf ( n42606 , n42532 );
nor ( n42607 , n42605 , n42606 );
buf ( n42608 , n42607 );
buf ( n42609 , n42608 );
nand ( n42610 , n42602 , n42609 );
buf ( n42611 , n42610 );
buf ( n42612 , n42611 );
not ( n42613 , n42612 );
buf ( n42614 , n42613 );
buf ( n42615 , n42614 );
nand ( n42616 , n42594 , n42615 );
buf ( n42617 , n42616 );
buf ( n42618 , n42617 );
not ( n42619 , n42618 );
buf ( n42620 , n42619 );
buf ( n42621 , n42620 );
nand ( n42622 , n42589 , n42621 );
buf ( n42623 , n42622 );
buf ( n42624 , n42623 );
nor ( n42625 , n42580 , n42624 );
buf ( n42626 , n42625 );
buf ( n42627 , n42626 );
buf ( n42628 , n39378 );
not ( n42629 , n42628 );
and ( n42630 , n42526 , n42527 );
buf ( n42631 , n42630 );
buf ( n42632 , n42631 );
not ( n42633 , n42632 );
or ( n42634 , n42629 , n42633 );
buf ( n42635 , n42631 );
buf ( n42636 , n39378 );
or ( n42637 , n42635 , n42636 );
nand ( n42638 , n42634 , n42637 );
buf ( n42639 , n42638 );
buf ( n42640 , n42639 );
and ( n42641 , n42627 , n42640 );
not ( n42642 , n42627 );
buf ( n42643 , n42639 );
not ( n42644 , n42643 );
buf ( n42645 , n42644 );
buf ( n42646 , n42645 );
and ( n42647 , n42642 , n42646 );
nor ( n42648 , n42641 , n42647 );
buf ( n42649 , n42648 );
nand ( n42650 , n42563 , n42649 );
nand ( n42651 , n42562 , n42650 );
buf ( n42652 , n42651 );
not ( n42653 , n42652 );
not ( n42654 , n42653 );
not ( n42655 , n42654 );
not ( n42656 , n42655 );
buf ( n42657 , n42656 );
not ( n42658 , n42657 );
buf ( n42659 , n42658 );
buf ( n42660 , n42659 );
buf ( n42661 , n42660 );
buf ( n42662 , n42661 );
buf ( n42663 , n42662 );
buf ( n42664 , n42663 );
not ( n42665 , n42664 );
and ( n42666 , n42559 , n42665 );
not ( n42667 , n42559 );
and ( n42668 , n42667 , n42664 );
nor ( n42669 , n42666 , n42668 );
and ( n42670 , n42463 , n42558 );
not ( n42671 , n42463 );
and ( n42672 , n42671 , n42557 );
nor ( n42673 , n42670 , n42672 );
and ( n42674 , n42281 , n42460 );
not ( n42675 , n42281 );
and ( n42676 , n42675 , n42461 );
nor ( n42677 , n42674 , n42676 );
not ( n42678 , n39434 );
not ( n42679 , n39101 );
not ( n42680 , n42266 );
or ( n42681 , n42679 , n42680 );
nand ( n42682 , n42681 , n42278 );
not ( n42683 , n42682 );
or ( n42684 , n42678 , n42683 );
nand ( n42685 , n42684 , n42270 );
and ( n42686 , n42685 , n39255 );
not ( n42687 , n42685 );
and ( n42688 , n42687 , n39254 );
nor ( n42689 , n42686 , n42688 );
nand ( n42690 , n39434 , n42270 );
not ( n42691 , n42690 );
and ( n42692 , n42682 , n42691 );
not ( n42693 , n42682 );
and ( n42694 , n42693 , n42690 );
nor ( n42695 , n42692 , n42694 );
not ( n42696 , n39718 );
not ( n42697 , n42258 );
and ( n42698 , n39682 , n39785 );
nand ( n42699 , n42248 , n42698 );
nand ( n42700 , n42697 , n42699 );
not ( n42701 , n42700 );
or ( n42702 , n42696 , n42701 );
nand ( n42703 , n42702 , n42261 );
not ( n42704 , n42264 );
nand ( n42705 , n42704 , n39601 );
not ( n42706 , n42705 );
and ( n42707 , n42703 , n42706 );
not ( n42708 , n42703 );
and ( n42709 , n42708 , n42705 );
nor ( n42710 , n42707 , n42709 );
not ( n42711 , n39100 );
not ( n42712 , n42711 );
not ( n42713 , n42266 );
or ( n42714 , n42712 , n42713 );
nand ( n42715 , n42714 , n42274 );
not ( n42716 , n42266 );
nand ( n42717 , n42711 , n42274 );
and ( n42718 , n42716 , n42717 );
not ( n42719 , n42716 );
not ( n42720 , n42717 );
and ( n42721 , n42719 , n42720 );
nor ( n42722 , n42718 , n42721 );
nand ( n42723 , n42248 , n39785 );
nand ( n42724 , n42723 , n42253 );
not ( n42725 , n39853 );
not ( n42726 , n40019 );
not ( n42727 , n42726 );
not ( n42728 , n42233 );
or ( n42729 , n42727 , n42728 );
not ( n42730 , n42240 );
nand ( n42731 , n42729 , n42730 );
not ( n42732 , n42731 );
or ( n42733 , n42725 , n42732 );
nand ( n42734 , n42733 , n42243 );
not ( n42735 , n40453 );
not ( n42736 , n40391 );
not ( n42737 , n42736 );
not ( n42738 , n40379 );
not ( n42739 , n42198 );
or ( n42740 , n42738 , n42739 );
not ( n42741 , n42217 );
nand ( n42742 , n42740 , n42741 );
not ( n42743 , n42742 );
or ( n42744 , n42737 , n42743 );
not ( n42745 , n42224 );
nand ( n42746 , n42744 , n42745 );
not ( n42747 , n42746 );
or ( n42748 , n42735 , n42747 );
not ( n42749 , n42226 );
nand ( n42750 , n42748 , n42749 );
not ( n42751 , n40365 );
nand ( n42752 , n40378 , n42198 );
not ( n42753 , n40283 );
or ( n42754 , n42752 , n42753 );
not ( n42755 , n42209 );
nand ( n42756 , n42754 , n42755 );
not ( n42757 , n42756 );
or ( n42758 , n42751 , n42757 );
nand ( n42759 , n42758 , n42212 );
not ( n42760 , n40018 );
not ( n42761 , n42233 );
or ( n42762 , n42760 , n42761 );
nand ( n42763 , n42762 , n42237 );
not ( n42764 , n40630 );
not ( n42765 , n40595 );
not ( n42766 , n42765 );
not ( n42767 , n42180 );
not ( n42768 , n42178 );
or ( n42769 , n42767 , n42768 );
not ( n42770 , n40775 );
nand ( n42771 , n42769 , n42770 );
not ( n42772 , n42771 );
or ( n42773 , n42766 , n42772 );
not ( n42774 , n42188 );
nand ( n42775 , n42773 , n42774 );
not ( n42776 , n42775 );
or ( n42777 , n42764 , n42776 );
nand ( n42778 , n42777 , n42191 );
not ( n42779 , n40390 );
not ( n42780 , n42742 );
or ( n42781 , n42779 , n42780 );
not ( n42782 , n42220 );
nand ( n42783 , n42781 , n42782 );
not ( n42784 , n40534 );
not ( n42785 , n42771 );
or ( n42786 , n42784 , n42785 );
not ( n42787 , n42183 );
nand ( n42788 , n42786 , n42787 );
not ( n42789 , n42788 );
nand ( n42790 , n40594 , n42187 );
not ( n42791 , n42790 );
or ( n42792 , n42789 , n42791 );
or ( n42793 , n42790 , n42788 );
nand ( n42794 , n42792 , n42793 );
nand ( n42795 , n40630 , n42191 );
not ( n42796 , n42795 );
not ( n42797 , n42775 );
or ( n42798 , n42796 , n42797 );
or ( n42799 , n42795 , n42775 );
nand ( n42800 , n42798 , n42799 );
nand ( n42801 , n40018 , n42237 );
not ( n42802 , n42801 );
not ( n42803 , n42233 );
or ( n42804 , n42802 , n42803 );
or ( n42805 , n42801 , n42233 );
nand ( n42806 , n42804 , n42805 );
nand ( n42807 , n40390 , n42782 );
not ( n42808 , n42807 );
not ( n42809 , n42742 );
or ( n42810 , n42808 , n42809 );
or ( n42811 , n42807 , n42742 );
nand ( n42812 , n42810 , n42811 );
and ( n42813 , n42178 , n42179 );
and ( n42814 , n42813 , n40678 );
nor ( n42815 , n42814 , n40698 );
not ( n42816 , n40737 );
or ( n42817 , n42815 , n42816 );
not ( n42818 , n40739 );
nand ( n42819 , n42817 , n42818 );
not ( n42820 , n42815 );
nor ( n42821 , n42816 , n40739 );
not ( n42822 , n42821 );
or ( n42823 , n42820 , n42822 );
or ( n42824 , n42821 , n42815 );
nand ( n42825 , n42823 , n42824 );
not ( n42826 , n42198 );
nand ( n42827 , n40378 , n42203 );
not ( n42828 , n42827 );
or ( n42829 , n42826 , n42828 );
or ( n42830 , n42827 , n42198 );
nand ( n42831 , n42829 , n42830 );
not ( n42832 , n42771 );
nand ( n42833 , n40534 , n42787 );
not ( n42834 , n42833 );
or ( n42835 , n42832 , n42834 );
or ( n42836 , n42833 , n42771 );
nand ( n42837 , n42835 , n42836 );
nand ( n42838 , n40678 , n40697 );
not ( n42839 , n42838 );
not ( n42840 , n42813 );
not ( n42841 , n40694 );
nand ( n42842 , n42840 , n42841 );
not ( n42843 , n42842 );
or ( n42844 , n42839 , n42843 );
or ( n42845 , n42838 , n42842 );
nand ( n42846 , n42844 , n42845 );
and ( n42847 , n42161 , n40958 );
nor ( n42848 , n42847 , n42167 );
or ( n42849 , n42848 , n41039 );
nand ( n42850 , n42849 , n42172 );
not ( n42851 , n42850 );
not ( n42852 , n42176 );
nand ( n42853 , n42852 , n42174 );
not ( n42854 , n42853 );
or ( n42855 , n42851 , n42854 );
or ( n42856 , n42853 , n42850 );
nand ( n42857 , n42855 , n42856 );
nand ( n42858 , n42179 , n42841 );
not ( n42859 , n42858 );
not ( n42860 , n42178 );
or ( n42861 , n42859 , n42860 );
or ( n42862 , n42858 , n42178 );
nand ( n42863 , n42861 , n42862 );
not ( n42864 , n40857 );
not ( n42865 , n42864 );
not ( n42866 , n42161 );
or ( n42867 , n42865 , n42866 );
nand ( n42868 , n42867 , n42164 );
not ( n42869 , n42868 );
not ( n42870 , n40957 );
nand ( n42871 , n42870 , n42166 );
not ( n42872 , n42871 );
or ( n42873 , n42869 , n42872 );
or ( n42874 , n42871 , n42868 );
nand ( n42875 , n42873 , n42874 );
not ( n42876 , n41369 );
not ( n42877 , n42141 );
not ( n42878 , n41410 );
nor ( n42879 , n42877 , n42878 );
not ( n42880 , n42879 );
or ( n42881 , n42876 , n42880 );
not ( n42882 , n42152 );
nand ( n42883 , n42881 , n42882 );
nand ( n42884 , n41291 , n42883 );
nand ( n42885 , n42884 , n42155 );
not ( n42886 , n42161 );
nand ( n42887 , n42864 , n42164 );
not ( n42888 , n42887 );
or ( n42889 , n42886 , n42888 );
or ( n42890 , n42887 , n42161 );
nand ( n42891 , n42889 , n42890 );
or ( n42892 , n42879 , n42146 );
not ( n42893 , n42892 );
nand ( n42894 , n41369 , n42151 );
not ( n42895 , n42894 );
or ( n42896 , n42893 , n42895 );
or ( n42897 , n42894 , n42892 );
nand ( n42898 , n42896 , n42897 );
and ( n42899 , n42122 , n42123 );
and ( n42900 , n42899 , n41694 );
nor ( n42901 , n42900 , n41698 );
not ( n42902 , n41688 );
or ( n42903 , n42901 , n42902 );
nand ( n42904 , n42903 , n41701 );
not ( n42905 , n42904 );
nand ( n42906 , n41677 , n41705 );
not ( n42907 , n42906 );
or ( n42908 , n42905 , n42907 );
or ( n42909 , n42906 , n42904 );
nand ( n42910 , n42908 , n42909 );
not ( n42911 , n41581 );
nand ( n42912 , n42911 , n42130 );
not ( n42913 , n42912 );
or ( n42914 , n42125 , n41706 );
not ( n42915 , n42914 );
not ( n42916 , n41418 );
not ( n42917 , n42916 );
or ( n42918 , n42915 , n42917 );
nand ( n42919 , n42918 , n42128 );
not ( n42920 , n42919 );
or ( n42921 , n42913 , n42920 );
or ( n42922 , n42912 , n42919 );
nand ( n42923 , n42921 , n42922 );
nor ( n42924 , n42878 , n42146 );
not ( n42925 , n42924 );
not ( n42926 , n42877 );
or ( n42927 , n42925 , n42926 );
or ( n42928 , n42924 , n42877 );
nand ( n42929 , n42927 , n42928 );
not ( n42930 , n42901 );
and ( n42931 , n41688 , n41701 );
not ( n42932 , n42931 );
or ( n42933 , n42930 , n42932 );
or ( n42934 , n42931 , n42901 );
nand ( n42935 , n42933 , n42934 );
nand ( n42936 , n41694 , n41697 );
not ( n42937 , n42936 );
not ( n42938 , n42899 );
not ( n42939 , n41690 );
nand ( n42940 , n42938 , n42939 );
not ( n42941 , n42940 );
or ( n42942 , n42937 , n42941 );
or ( n42943 , n42936 , n42940 );
nand ( n42944 , n42942 , n42943 );
nand ( n42945 , n42123 , n42939 );
not ( n42946 , n42945 );
not ( n42947 , n42122 );
or ( n42948 , n42946 , n42947 );
or ( n42949 , n42945 , n42122 );
nand ( n42950 , n42948 , n42949 );
nand ( n42951 , n41803 , n42121 );
not ( n42952 , n42951 );
not ( n42953 , n42111 );
and ( n42954 , n42110 , n42953 );
and ( n42955 , n42954 , n41935 );
nor ( n42956 , n42955 , n41941 );
or ( n42957 , n42956 , n41862 );
nand ( n42958 , n42957 , n42117 );
not ( n42959 , n42958 );
or ( n42960 , n42952 , n42959 );
or ( n42961 , n42951 , n42958 );
nand ( n42962 , n42960 , n42961 );
not ( n42963 , n42956 );
and ( n42964 , n41863 , n42117 );
not ( n42965 , n42964 );
or ( n42966 , n42963 , n42965 );
or ( n42967 , n42964 , n42956 );
nand ( n42968 , n42966 , n42967 );
nand ( n42969 , n41935 , n41940 );
not ( n42970 , n42969 );
not ( n42971 , n42954 );
nand ( n42972 , n42971 , n41865 );
not ( n42973 , n42972 );
or ( n42974 , n42970 , n42973 );
or ( n42975 , n42969 , n42972 );
nand ( n42976 , n42974 , n42975 );
not ( n42977 , n42108 );
nand ( n42978 , n42977 , n42097 );
not ( n42979 , n42978 );
and ( n42980 , n42094 , n41950 );
nor ( n42981 , n42980 , n42101 );
not ( n42982 , n41947 );
or ( n42983 , n42981 , n42982 );
nand ( n42984 , n42983 , n42105 );
not ( n42985 , n42984 );
or ( n42986 , n42979 , n42985 );
or ( n42987 , n42978 , n42984 );
nand ( n42988 , n42986 , n42987 );
nand ( n42989 , n42953 , n41865 );
not ( n42990 , n42989 );
not ( n42991 , n42110 );
or ( n42992 , n42990 , n42991 );
or ( n42993 , n42989 , n42110 );
nand ( n42994 , n42992 , n42993 );
not ( n42995 , n42981 );
and ( n42996 , n41947 , n42105 );
not ( n42997 , n42996 );
or ( n42998 , n42995 , n42997 );
or ( n42999 , n42996 , n42981 );
nand ( n43000 , n42998 , n42999 );
nand ( n43001 , n41950 , n42100 );
not ( n43002 , n43001 );
not ( n43003 , n42094 );
nand ( n43004 , n43003 , n42098 );
not ( n43005 , n43004 );
or ( n43006 , n43002 , n43005 );
or ( n43007 , n43001 , n43004 );
nand ( n43008 , n43006 , n43007 );
nand ( n43009 , n42093 , n42098 );
not ( n43010 , n43009 );
not ( n43011 , n42092 );
or ( n43012 , n43010 , n43011 );
or ( n43013 , n43009 , n42092 );
nand ( n43014 , n43012 , n43013 );
xor ( n43015 , n41954 , n18554 );
xor ( n43016 , n43015 , n42089 );
nand ( n43017 , n42008 , n42088 );
not ( n43018 , n43017 );
not ( n43019 , n42085 );
or ( n43020 , n43018 , n43019 );
or ( n43021 , n43017 , n42085 );
nand ( n43022 , n43020 , n43021 );
nand ( n43023 , n42039 , n42084 );
not ( n43024 , n43023 );
not ( n43025 , n42081 );
or ( n43026 , n43024 , n43025 );
or ( n43027 , n43023 , n42081 );
nand ( n43028 , n43026 , n43027 );
nand ( n43029 , n42051 , n42080 );
not ( n43030 , n43029 );
not ( n43031 , n42077 );
or ( n43032 , n43030 , n43031 );
or ( n43033 , n43029 , n42077 );
nand ( n43034 , n43032 , n43033 );
not ( n43035 , n42069 );
nand ( n43036 , n42057 , n42072 );
not ( n43037 , n43036 );
or ( n43038 , n43035 , n43037 );
or ( n43039 , n42069 , n43036 );
nand ( n43040 , n43038 , n43039 );
not ( n43041 , n42068 );
nor ( n43042 , n43041 , n42059 );
not ( n43043 , n43042 );
not ( n43044 , n42066 );
or ( n43045 , n43043 , n43044 );
or ( n43046 , n42066 , n43042 );
nand ( n43047 , n43045 , n43046 );
nand ( n43048 , n40771 , n40774 );
and ( n43049 , n41291 , n42155 );
not ( n43050 , n42194 );
nand ( n43051 , n43050 , n40637 );
nand ( n43052 , n39853 , n42243 );
not ( n43053 , n39965 );
nand ( n43054 , n43053 , n42239 );
nand ( n43055 , n39718 , n42261 );
nand ( n43056 , n39682 , n42257 );
nand ( n43057 , n39785 , n42253 );
not ( n43058 , n42246 );
nand ( n43059 , n43058 , n39901 );
not ( n43060 , n42228 );
nand ( n43061 , n43060 , n42230 );
nand ( n43062 , n40453 , n42749 );
nand ( n43063 , n40387 , n42223 );
nor ( n43064 , n42135 , n41669 );
nor ( n43065 , n41218 , n42159 );
nand ( n43066 , n40151 , n42216 );
nand ( n43067 , n40365 , n42212 );
nor ( n43068 , n38981 , n42277 );
xnor ( n43069 , n42700 , n43055 );
xnor ( n43070 , n42819 , n43048 );
xnor ( n43071 , n42778 , n43051 );
xnor ( n43072 , n42731 , n43052 );
xnor ( n43073 , n42763 , n43054 );
xnor ( n43074 , n42724 , n43056 );
xnor ( n43075 , n42248 , n43057 );
xnor ( n43076 , n42734 , n43059 );
xnor ( n43077 , n42750 , n43061 );
xnor ( n43078 , n42746 , n43062 );
xnor ( n43079 , n42783 , n43063 );
xor ( n43080 , n42885 , n43065 );
xnor ( n43081 , n42759 , n43066 );
xnor ( n43082 , n42756 , n43067 );
xor ( n43083 , n42715 , n43068 );
buf ( n43084 , n36912 );
buf ( n43085 , n36891 );
buf ( n43086 , n42557 );
xor ( n43087 , n43084 , n43085 );
xor ( n43088 , n43087 , n43086 );
buf ( n43089 , n43088 );
xor ( n43090 , n43084 , n43085 );
and ( n43091 , n43090 , n43086 );
and ( n43092 , n43084 , n43085 );
or ( n43093 , n43091 , n43092 );
buf ( n43094 , n43093 );
buf ( n43095 , n36921 );
buf ( n43096 , n36918 );
buf ( n43097 , n42401 );
xor ( n43098 , n43095 , n43096 );
xor ( n43099 , n43098 , n43097 );
buf ( n43100 , n43099 );
xor ( n43101 , n43095 , n43096 );
and ( n43102 , n43101 , n43097 );
and ( n43103 , n43095 , n43096 );
or ( n43104 , n43102 , n43103 );
buf ( n43105 , n43104 );
buf ( n43106 , n36326 );
buf ( n43107 , n29571 );
buf ( n43108 , n39255 );
xor ( n43109 , n43106 , n43107 );
xor ( n43110 , n43109 , n43108 );
buf ( n43111 , n43110 );
xor ( n43112 , n43106 , n43107 );
and ( n43113 , n43112 , n43108 );
and ( n43114 , n43106 , n43107 );
or ( n43115 , n43113 , n43114 );
buf ( n43116 , n43115 );
buf ( n43117 , n37227 );
buf ( n43118 , n37230 );
not ( n43119 , n42662 );
buf ( n43120 , n43119 );
xor ( n43121 , n43117 , n43118 );
xor ( n43122 , n43121 , n43120 );
buf ( n43123 , n43122 );
xor ( n43124 , n43117 , n43118 );
and ( n43125 , n43124 , n43120 );
and ( n43126 , n43117 , n43118 );
or ( n43127 , n43125 , n43126 );
buf ( n43128 , n43127 );
buf ( n43129 , n35946 );
buf ( n43130 , n27508 );
buf ( n43131 , n30379 );
xor ( n43132 , n43129 , n43130 );
xor ( n43133 , n43132 , n43131 );
buf ( n43134 , n43133 );
xor ( n43135 , n43129 , n43130 );
and ( n43136 , n43135 , n43131 );
and ( n43137 , n43129 , n43130 );
or ( n43138 , n43136 , n43137 );
buf ( n43139 , n43138 );
buf ( n43140 , n35843 );
buf ( n43141 , n35841 );
buf ( n43142 , n41948 );
xor ( n43143 , n43140 , n43141 );
xor ( n43144 , n43143 , n43142 );
buf ( n43145 , n43144 );
xor ( n43146 , n43140 , n43141 );
and ( n43147 , n43146 , n43142 );
and ( n43148 , n43140 , n43141 );
or ( n43149 , n43147 , n43148 );
buf ( n43150 , n43149 );
buf ( n43151 , n36114 );
buf ( n43152 , n36108 );
buf ( n43153 , n30351 );
xor ( n43154 , n43151 , n43152 );
xor ( n43155 , n43154 , n43153 );
buf ( n43156 , n43155 );
xor ( n43157 , n43151 , n43152 );
and ( n43158 , n43157 , n43153 );
and ( n43159 , n43151 , n43152 );
or ( n43160 , n43158 , n43159 );
buf ( n43161 , n43160 );
buf ( n43162 , n36054 );
buf ( n43163 , n36087 );
buf ( n43164 , n30259 );
xor ( n43165 , n43162 , n43163 );
xor ( n43166 , n43165 , n43164 );
buf ( n43167 , n43166 );
xor ( n43168 , n43162 , n43163 );
and ( n43169 , n43168 , n43164 );
and ( n43170 , n43162 , n43163 );
or ( n43171 , n43169 , n43170 );
buf ( n43172 , n43171 );
buf ( n43173 , n23339 );
buf ( n43174 , n36153 );
buf ( n43175 , n41801 );
xor ( n43176 , n43173 , n43174 );
xor ( n43177 , n43176 , n43175 );
buf ( n43178 , n43177 );
xor ( n43179 , n43173 , n43174 );
and ( n43180 , n43179 , n43175 );
and ( n43181 , n43173 , n43174 );
or ( n43182 , n43180 , n43181 );
buf ( n43183 , n43182 );
buf ( n43184 , n35792 );
buf ( n43185 , n27330 );
buf ( n43186 , n30964 );
xor ( n43187 , n43184 , n43185 );
xor ( n43188 , n43187 , n43186 );
buf ( n43189 , n43188 );
xor ( n43190 , n43184 , n43185 );
and ( n43191 , n43190 , n43186 );
and ( n43192 , n43184 , n43185 );
or ( n43193 , n43191 , n43192 );
buf ( n43194 , n43193 );
buf ( n43195 , n35783 );
buf ( n43196 , n35778 );
buf ( n43197 , n41692 );
xor ( n43198 , n43195 , n43196 );
xor ( n43199 , n43198 , n43197 );
buf ( n43200 , n43199 );
xor ( n43201 , n43195 , n43196 );
and ( n43202 , n43201 , n43197 );
and ( n43203 , n43195 , n43196 );
or ( n43204 , n43202 , n43203 );
buf ( n43205 , n43204 );
buf ( n43206 , n35770 );
buf ( n43207 , n27602 );
buf ( n43208 , n41683 );
xor ( n43209 , n43206 , n43207 );
xor ( n43210 , n43209 , n43208 );
buf ( n43211 , n43210 );
xor ( n43212 , n43206 , n43207 );
and ( n43213 , n43212 , n43208 );
and ( n43214 , n43206 , n43207 );
or ( n43215 , n43213 , n43214 );
buf ( n43216 , n43215 );
buf ( n43217 , n35749 );
buf ( n43218 , n35743 );
buf ( n43219 , n30929 );
xor ( n43220 , n43217 , n43218 );
xor ( n43221 , n43220 , n43219 );
buf ( n43222 , n43221 );
xor ( n43223 , n43217 , n43218 );
and ( n43224 , n43223 , n43219 );
and ( n43225 , n43217 , n43218 );
or ( n43226 , n43224 , n43225 );
buf ( n43227 , n43226 );
buf ( n43228 , n35654 );
buf ( n43229 , n35649 );
buf ( n43230 , n41407 );
xor ( n43231 , n43228 , n43229 );
xor ( n43232 , n43231 , n43230 );
buf ( n43233 , n43232 );
xor ( n43234 , n43228 , n43229 );
and ( n43235 , n43234 , n43230 );
and ( n43236 , n43228 , n43229 );
or ( n43237 , n43235 , n43236 );
buf ( n43238 , n43237 );
buf ( n43239 , n28568 );
buf ( n43240 , n35589 );
buf ( n43241 , n41217 );
xor ( n43242 , n43239 , n43240 );
xor ( n43243 , n43242 , n43241 );
buf ( n43244 , n43243 );
xor ( n43245 , n43239 , n43240 );
and ( n43246 , n43245 , n43241 );
and ( n43247 , n43239 , n43240 );
or ( n43248 , n43246 , n43247 );
buf ( n43249 , n43248 );
buf ( n43250 , n35538 );
not ( n43251 , n36958 );
buf ( n43252 , n43251 );
buf ( n43253 , n41038 );
xor ( n43254 , n43250 , n43252 );
xor ( n43255 , n43254 , n43253 );
buf ( n43256 , n43255 );
xor ( n43257 , n43250 , n43252 );
and ( n43258 , n43257 , n43253 );
and ( n43259 , n43250 , n43252 );
or ( n43260 , n43258 , n43259 );
buf ( n43261 , n43260 );
buf ( n43262 , n35563 );
buf ( n43263 , n35542 );
buf ( n43264 , n40951 );
xor ( n43265 , n43262 , n43263 );
xor ( n43266 , n43265 , n43264 );
buf ( n43267 , n43266 );
xor ( n43268 , n43262 , n43263 );
and ( n43269 , n43268 , n43264 );
and ( n43270 , n43262 , n43263 );
or ( n43271 , n43269 , n43270 );
buf ( n43272 , n43271 );
buf ( n43273 , n35443 );
not ( n43274 , n36254 );
buf ( n43275 , n43274 );
buf ( n43276 , n40692 );
xor ( n43277 , n43273 , n43275 );
xor ( n43278 , n43277 , n43276 );
buf ( n43279 , n43278 );
xor ( n43280 , n43273 , n43275 );
and ( n43281 , n43280 , n43276 );
and ( n43282 , n43273 , n43275 );
or ( n43283 , n43281 , n43282 );
buf ( n43284 , n43283 );
buf ( n43285 , n40677 );
buf ( n43286 , n35193 );
buf ( n43287 , n43286 );
buf ( n43288 , n35106 );
xor ( n43289 , n43285 , n43287 );
xor ( n43290 , n43289 , n43288 );
buf ( n43291 , n43290 );
xor ( n43292 , n43285 , n43287 );
and ( n43293 , n43292 , n43288 );
and ( n43294 , n43285 , n43287 );
or ( n43295 , n43293 , n43294 );
buf ( n43296 , n43295 );
buf ( n43297 , n35256 );
buf ( n43298 , n35273 );
buf ( n43299 , n43298 );
buf ( n43300 , n43299 );
buf ( n43301 , n40769 );
xor ( n43302 , n43297 , n43300 );
xor ( n43303 , n43302 , n43301 );
buf ( n43304 , n43303 );
xor ( n43305 , n43297 , n43300 );
and ( n43306 , n43305 , n43301 );
and ( n43307 , n43297 , n43300 );
or ( n43308 , n43306 , n43307 );
buf ( n43309 , n43308 );
buf ( n43310 , n35282 );
buf ( n43311 , n43310 );
not ( n43312 , n36277 );
buf ( n43313 , n43312 );
buf ( n43314 , n40529 );
xor ( n43315 , n43311 , n43313 );
xor ( n43316 , n43315 , n43314 );
buf ( n43317 , n43316 );
xor ( n43318 , n43311 , n43313 );
and ( n43319 , n43318 , n43314 );
and ( n43320 , n43311 , n43313 );
or ( n43321 , n43319 , n43320 );
buf ( n43322 , n43321 );
not ( n43323 , n33647 );
buf ( n43324 , n43323 );
buf ( n43325 , n27514 );
buf ( n43326 , n40628 );
xor ( n43327 , n43324 , n43325 );
xor ( n43328 , n43327 , n43326 );
buf ( n43329 , n43328 );
xor ( n43330 , n43324 , n43325 );
and ( n43331 , n43330 , n43326 );
and ( n43332 , n43324 , n43325 );
or ( n43333 , n43331 , n43332 );
buf ( n43334 , n43333 );
buf ( n43335 , n22526 );
buf ( n43336 , n33613 );
buf ( n43337 , n43336 );
buf ( n43338 , n40226 );
xor ( n43339 , n43335 , n43337 );
xor ( n43340 , n43339 , n43338 );
buf ( n43341 , n43340 );
xor ( n43342 , n43335 , n43337 );
and ( n43343 , n43342 , n43338 );
and ( n43344 , n43335 , n43337 );
or ( n43345 , n43343 , n43344 );
buf ( n43346 , n43345 );
buf ( n43347 , n24075 );
buf ( n43348 , n37510 );
buf ( n43349 , n40149 );
xor ( n43350 , n43347 , n43348 );
xor ( n43351 , n43350 , n43349 );
buf ( n43352 , n43351 );
xor ( n43353 , n43347 , n43348 );
and ( n43354 , n43353 , n43349 );
and ( n43355 , n43347 , n43348 );
or ( n43356 , n43354 , n43355 );
buf ( n43357 , n43356 );
buf ( n43358 , n33524 );
not ( n43359 , n33476 );
buf ( n43360 , n43359 );
buf ( n43361 , n40381 );
xor ( n43362 , n43358 , n43360 );
xor ( n43363 , n43362 , n43361 );
buf ( n43364 , n43363 );
xor ( n43365 , n43358 , n43360 );
and ( n43366 , n43365 , n43361 );
and ( n43367 , n43358 , n43360 );
or ( n43368 , n43366 , n43367 );
buf ( n43369 , n43368 );
buf ( n43370 , n32827 );
buf ( n43371 , n32810 );
buf ( n43372 , n39335 );
xor ( n43373 , n43370 , n43371 );
xor ( n43374 , n43373 , n43372 );
buf ( n43375 , n43374 );
xor ( n43376 , n43370 , n43371 );
and ( n43377 , n43376 , n43372 );
and ( n43378 , n43370 , n43371 );
or ( n43379 , n43377 , n43378 );
buf ( n43380 , n43379 );
buf ( n43381 , n33257 );
buf ( n43382 , n33312 );
buf ( n43383 , n39964 );
xor ( n43384 , n43381 , n43382 );
xor ( n43385 , n43384 , n43383 );
buf ( n43386 , n43385 );
xor ( n43387 , n43381 , n43382 );
and ( n43388 , n43387 , n43383 );
and ( n43389 , n43381 , n43382 );
or ( n43390 , n43388 , n43389 );
buf ( n43391 , n43390 );
buf ( n43392 , n33353 );
buf ( n43393 , n33347 );
buf ( n43394 , n43393 );
buf ( n43395 , n39847 );
xor ( n43396 , n43392 , n43394 );
xor ( n43397 , n43396 , n43395 );
buf ( n43398 , n43397 );
xor ( n43399 , n43392 , n43394 );
and ( n43400 , n43399 , n43395 );
and ( n43401 , n43392 , n43394 );
or ( n43402 , n43400 , n43401 );
buf ( n43403 , n43402 );
buf ( n43404 , n33386 );
buf ( n43405 , n33391 );
buf ( n43406 , n39779 );
xor ( n43407 , n43404 , n43405 );
xor ( n43408 , n43407 , n43406 );
buf ( n43409 , n43408 );
xor ( n43410 , n43404 , n43405 );
and ( n43411 , n43410 , n43406 );
and ( n43412 , n43404 , n43405 );
or ( n43413 , n43411 , n43412 );
buf ( n43414 , n43413 );
buf ( n43415 , n36523 );
buf ( n43416 , n36394 );
buf ( n43417 , n42460 );
xor ( n43418 , n43415 , n43416 );
xor ( n43419 , n43418 , n43417 );
buf ( n43420 , n43419 );
xor ( n43421 , n43415 , n43416 );
and ( n43422 , n43421 , n43417 );
and ( n43423 , n43415 , n43416 );
or ( n43424 , n43422 , n43423 );
buf ( n43425 , n43424 );
buf ( n43426 , n32764 );
buf ( n43427 , n32770 );
buf ( n43428 , n39056 );
xor ( n43429 , n43426 , n43427 );
xor ( n43430 , n43429 , n43428 );
buf ( n43431 , n43430 );
xor ( n43432 , n43426 , n43427 );
and ( n43433 , n43432 , n43428 );
and ( n43434 , n43426 , n43427 );
or ( n43435 , n43433 , n43434 );
buf ( n43436 , n43435 );
buf ( n43437 , n37293 );
buf ( n43438 , n37238 );
xor ( n43439 , n43437 , n43438 );
buf ( n43440 , n43439 );
and ( n43441 , n43437 , n43438 );
buf ( n43442 , n43441 );
buf ( n43443 , n37220 );
buf ( n43444 , n37158 );
xor ( n43445 , n43443 , n43444 );
buf ( n43446 , n43445 );
and ( n43447 , n43443 , n43444 );
buf ( n43448 , n43447 );
buf ( n43449 , n37345 );
buf ( n43450 , n37299 );
xor ( n43451 , n43449 , n43450 );
buf ( n43452 , n43451 );
and ( n43453 , n43449 , n43450 );
buf ( n43454 , n43453 );
buf ( n43455 , n37378 );
buf ( n43456 , n37352 );
xor ( n43457 , n43455 , n43456 );
buf ( n43458 , n43457 );
and ( n43459 , n43455 , n43456 );
buf ( n43460 , n43459 );
buf ( n43461 , n37633 );
buf ( n43462 , n37627 );
xor ( n43463 , n43461 , n43462 );
buf ( n43464 , n43463 );
buf ( n43465 , n43458 );
buf ( n43466 , n43454 );
buf ( n43467 , n43448 );
buf ( n43468 , n43440 );
or ( n43469 , n43467 , n43468 );
buf ( n43470 , n43469 );
buf ( n43471 , n43470 );
not ( n43472 , n43471 );
buf ( n43473 , n43442 );
buf ( n43474 , n43452 );
nor ( n43475 , n43473 , n43474 );
buf ( n43476 , n43475 );
buf ( n43477 , n43476 );
nor ( n43478 , n43472 , n43477 );
buf ( n43479 , n43478 );
buf ( n43480 , n43479 );
not ( n43481 , n43480 );
buf ( n43482 , n32688 );
buf ( n43483 , n32522 );
xor ( n43484 , n43482 , n43483 );
buf ( n43485 , n39575 );
xor ( n43486 , n43484 , n43485 );
buf ( n43487 , n43486 );
buf ( n43488 , n43487 );
not ( n43489 , n43488 );
xor ( n43490 , n32513 , n26379 );
and ( n43491 , n43490 , n39716 );
and ( n43492 , n32513 , n26379 );
nor ( n43493 , n43491 , n43492 );
buf ( n43494 , n43493 );
nand ( n43495 , n43489 , n43494 );
buf ( n43496 , n43495 );
buf ( n43497 , n43496 );
xor ( n43498 , n43482 , n43483 );
and ( n43499 , n43498 , n43485 );
and ( n43500 , n43482 , n43483 );
or ( n43501 , n43499 , n43500 );
buf ( n43502 , n43501 );
buf ( n43503 , n43502 );
buf ( n43504 , n43431 );
or ( n43505 , n43503 , n43504 );
buf ( n43506 , n43505 );
buf ( n43507 , n43506 );
and ( n43508 , n43497 , n43507 );
buf ( n43509 , n43508 );
buf ( n43510 , n43509 );
buf ( n43511 , n43414 );
xnor ( n43512 , n20096 , n32505 );
not ( n43513 , n39681 );
and ( n43514 , n43512 , n43513 );
not ( n43515 , n43512 );
and ( n43516 , n43515 , n39681 );
nor ( n43517 , n43514 , n43516 );
buf ( n43518 , n43517 );
nor ( n43519 , n43511 , n43518 );
buf ( n43520 , n43519 );
buf ( n43521 , n43520 );
xor ( n43522 , n32513 , n26379 );
xor ( n43523 , n43522 , n39716 );
or ( n43524 , n20096 , n32505 );
not ( n43525 , n43524 );
not ( n43526 , n39681 );
or ( n43527 , n43525 , n43526 );
nand ( n43528 , n20096 , n32505 );
nand ( n43529 , n43527 , n43528 );
nor ( n43530 , n43523 , n43529 );
buf ( n43531 , n43530 );
nor ( n43532 , n43521 , n43531 );
buf ( n43533 , n43532 );
buf ( n43534 , n43533 );
nand ( n43535 , n43510 , n43534 );
buf ( n43536 , n43535 );
buf ( n43537 , n43536 );
buf ( n43538 , n43436 );
buf ( n43539 , n32836 );
buf ( n43540 , n43539 );
buf ( n43541 , n32831 );
buf ( n43542 , n43541 );
xor ( n43543 , n43540 , n43542 );
buf ( n43544 , n38500 );
xor ( n43545 , n43543 , n43544 );
buf ( n43546 , n43545 );
buf ( n43547 , n43546 );
nor ( n43548 , n43538 , n43547 );
buf ( n43549 , n43548 );
buf ( n43550 , n43549 );
buf ( n43551 , n43375 );
xor ( n43552 , n43540 , n43542 );
and ( n43553 , n43552 , n43544 );
and ( n43554 , n43540 , n43542 );
or ( n43555 , n43553 , n43554 );
buf ( n43556 , n43555 );
buf ( n43557 , n43556 );
nor ( n43558 , n43551 , n43557 );
buf ( n43559 , n43558 );
buf ( n43560 , n43559 );
nor ( n43561 , n43550 , n43560 );
buf ( n43562 , n43561 );
buf ( n43563 , n43562 );
buf ( n43564 , n43420 );
buf ( n43565 , n43116 );
nor ( n43566 , n43564 , n43565 );
buf ( n43567 , n43566 );
buf ( n43568 , n43567 );
buf ( n43569 , n43111 );
buf ( n43570 , n43380 );
nor ( n43571 , n43569 , n43570 );
buf ( n43572 , n43571 );
buf ( n43573 , n43572 );
nor ( n43574 , n43568 , n43573 );
buf ( n43575 , n43574 );
buf ( n43576 , n43575 );
nand ( n43577 , n43563 , n43576 );
buf ( n43578 , n43577 );
buf ( n43579 , n43578 );
nor ( n43580 , n43537 , n43579 );
buf ( n43581 , n43580 );
buf ( n43582 , n43581 );
not ( n43583 , n43582 );
buf ( n43584 , n43398 );
buf ( n43585 , n43391 );
nor ( n43586 , n43584 , n43585 );
buf ( n43587 , n43586 );
buf ( n43588 , n43587 );
buf ( n43589 , n33419 );
buf ( n43590 , n33399 );
buf ( n43591 , n43590 );
xor ( n43592 , n43589 , n43591 );
buf ( n43593 , n40012 );
and ( n43594 , n43592 , n43593 );
and ( n43595 , n43589 , n43591 );
or ( n43596 , n43594 , n43595 );
buf ( n43597 , n43596 );
buf ( n43598 , n43597 );
buf ( n43599 , n43386 );
nor ( n43600 , n43598 , n43599 );
buf ( n43601 , n43600 );
buf ( n43602 , n43601 );
nor ( n43603 , n43588 , n43602 );
buf ( n43604 , n43603 );
buf ( n43605 , n43604 );
buf ( n43606 , n43409 );
not ( n43607 , n43606 );
xor ( n43608 , n33382 , n33361 );
not ( n43609 , n39895 );
and ( n43610 , n43608 , n43609 );
and ( n43611 , n33382 , n33361 );
or ( n43612 , n43610 , n43611 );
buf ( n43613 , n43612 );
not ( n43614 , n43613 );
buf ( n43615 , n43614 );
buf ( n43616 , n43615 );
nand ( n43617 , n43607 , n43616 );
buf ( n43618 , n43617 );
buf ( n43619 , n43618 );
xor ( n43620 , n33382 , n33361 );
xor ( n43621 , n43620 , n43609 );
buf ( n43622 , n43621 );
not ( n43623 , n43622 );
buf ( n43624 , n43403 );
not ( n43625 , n43624 );
buf ( n43626 , n43625 );
buf ( n43627 , n43626 );
nand ( n43628 , n43623 , n43627 );
buf ( n43629 , n43628 );
buf ( n43630 , n43629 );
and ( n43631 , n43605 , n43619 , n43630 );
buf ( n43632 , n43631 );
buf ( n43633 , n43632 );
not ( n43634 , n43633 );
xor ( n43635 , n43589 , n43591 );
xor ( n43636 , n43635 , n43593 );
buf ( n43637 , n43636 );
buf ( n43638 , n43637 );
not ( n43639 , n43638 );
xor ( n43640 , n26385 , n40515 );
not ( n43641 , n33426 );
and ( n43642 , n43640 , n43641 );
and ( n43643 , n26385 , n40515 );
or ( n43644 , n43642 , n43643 );
not ( n43645 , n43644 );
buf ( n43646 , n43645 );
nand ( n43647 , n43639 , n43646 );
buf ( n43648 , n43647 );
buf ( n43649 , n43648 );
not ( n43650 , n43649 );
buf ( n43651 , n43364 );
buf ( n43652 , n34044 );
buf ( n43653 , n34022 );
xor ( n43654 , n43652 , n43653 );
buf ( n43655 , n40389 );
and ( n43656 , n43654 , n43655 );
and ( n43657 , n43652 , n43653 );
or ( n43658 , n43656 , n43657 );
buf ( n43659 , n43658 );
buf ( n43660 , n43659 );
nand ( n43661 , n43651 , n43660 );
buf ( n43662 , n43661 );
buf ( n43663 , n43369 );
buf ( n43664 , n33533 );
xor ( n43665 , n43664 , n26183 );
xor ( n43666 , n43665 , n40452 );
buf ( n43667 , n43666 );
nor ( n43668 , n43663 , n43667 );
buf ( n43669 , n43668 );
or ( n43670 , n43662 , n43669 );
buf ( n43671 , n43369 );
buf ( n43672 , n43666 );
nand ( n43673 , n43671 , n43672 );
buf ( n43674 , n43673 );
nand ( n43675 , n43670 , n43674 );
not ( n43676 , n43675 );
xor ( n43677 , n26385 , n40515 );
not ( n43678 , n33426 );
xor ( n43679 , n43677 , n43678 );
xor ( n43680 , n43664 , n26183 );
and ( n43681 , n43680 , n40452 );
and ( n43682 , n43664 , n26183 );
nor ( n43683 , n43681 , n43682 );
not ( n43684 , n43683 );
or ( n43685 , n43679 , n43684 );
not ( n43686 , n43685 );
or ( n43687 , n43676 , n43686 );
not ( n43688 , n43683 );
nand ( n43689 , n43688 , n43679 );
nand ( n43690 , n43687 , n43689 );
buf ( n43691 , n43690 );
not ( n43692 , n43691 );
or ( n43693 , n43650 , n43692 );
buf ( n43694 , n43645 );
not ( n43695 , n43694 );
buf ( n43696 , n43637 );
nand ( n43697 , n43695 , n43696 );
buf ( n43698 , n43697 );
buf ( n43699 , n43698 );
nand ( n43700 , n43693 , n43699 );
buf ( n43701 , n43700 );
buf ( n43702 , n43701 );
not ( n43703 , n43702 );
or ( n43704 , n43634 , n43703 );
buf ( n43705 , n43629 );
not ( n43706 , n43705 );
buf ( n43707 , n43597 );
buf ( n43708 , n43386 );
and ( n43709 , n43707 , n43708 );
buf ( n43710 , n43709 );
buf ( n43711 , n43710 );
not ( n43712 , n43711 );
buf ( n43713 , n43587 );
not ( n43714 , n43713 );
buf ( n43715 , n43714 );
buf ( n43716 , n43715 );
not ( n43717 , n43716 );
or ( n43718 , n43712 , n43717 );
buf ( n43719 , n43398 );
buf ( n43720 , n43391 );
nand ( n43721 , n43719 , n43720 );
buf ( n43722 , n43721 );
buf ( n43723 , n43722 );
nand ( n43724 , n43718 , n43723 );
buf ( n43725 , n43724 );
buf ( n43726 , n43725 );
not ( n43727 , n43726 );
or ( n43728 , n43706 , n43727 );
buf ( n43729 , n43626 );
not ( n43730 , n43729 );
buf ( n43731 , n43621 );
nand ( n43732 , n43730 , n43731 );
buf ( n43733 , n43732 );
buf ( n43734 , n43733 );
nand ( n43735 , n43728 , n43734 );
buf ( n43736 , n43735 );
buf ( n43737 , n43736 );
buf ( n43738 , n43618 );
and ( n43739 , n43737 , n43738 );
buf ( n43740 , n43615 );
not ( n43741 , n43740 );
buf ( n43742 , n43409 );
nand ( n43743 , n43741 , n43742 );
buf ( n43744 , n43743 );
buf ( n43745 , n43744 );
not ( n43746 , n43745 );
buf ( n43747 , n43746 );
buf ( n43748 , n43747 );
nor ( n43749 , n43739 , n43748 );
buf ( n43750 , n43749 );
buf ( n43751 , n43750 );
nand ( n43752 , n43704 , n43751 );
buf ( n43753 , n43752 );
buf ( n43754 , n43753 );
not ( n43755 , n43754 );
buf ( n43756 , n43632 );
buf ( n43757 , n43685 );
or ( n43758 , n43659 , n43364 );
buf ( n43759 , n43758 );
buf ( n43760 , n43648 );
buf ( n43761 , n43669 );
not ( n43762 , n43761 );
buf ( n43763 , n43762 );
buf ( n43764 , n43763 );
and ( n43765 , n43757 , n43759 , n43760 , n43764 );
buf ( n43766 , n43765 );
buf ( n43767 , n43766 );
and ( n43768 , n43756 , n43767 );
buf ( n43769 , n43768 );
buf ( n43770 , n43769 );
buf ( n43771 , n35576 );
buf ( n43772 , n35570 );
buf ( n43773 , n43772 );
xor ( n43774 , n43771 , n43773 );
buf ( n43775 , n41286 );
xor ( n43776 , n43774 , n43775 );
buf ( n43777 , n43776 );
buf ( n43778 , n43777 );
buf ( n43779 , n28989 );
buf ( n43780 , n28900 );
xor ( n43781 , n43779 , n43780 );
buf ( n43782 , n41364 );
and ( n43783 , n43781 , n43782 );
and ( n43784 , n43779 , n43780 );
or ( n43785 , n43783 , n43784 );
buf ( n43786 , n43785 );
buf ( n43787 , n43786 );
nor ( n43788 , n43778 , n43787 );
buf ( n43789 , n43788 );
buf ( n43790 , n43789 );
xor ( n43791 , n43779 , n43780 );
xor ( n43792 , n43791 , n43782 );
buf ( n43793 , n43792 );
buf ( n43794 , n43793 );
buf ( n43795 , n43238 );
nor ( n43796 , n43794 , n43795 );
buf ( n43797 , n43796 );
buf ( n43798 , n43797 );
nor ( n43799 , n43790 , n43798 );
buf ( n43800 , n43799 );
buf ( n43801 , n43800 );
xor ( n43802 , n43771 , n43773 );
and ( n43803 , n43802 , n43775 );
and ( n43804 , n43771 , n43773 );
or ( n43805 , n43803 , n43804 );
buf ( n43806 , n43805 );
or ( n43807 , n43244 , n43806 );
buf ( n43808 , n43807 );
buf ( n43809 , n29873 );
not ( n43810 , n35694 );
buf ( n43811 , n43810 );
xor ( n43812 , n43809 , n43811 );
buf ( n43813 , n40856 );
xor ( n43814 , n43812 , n43813 );
buf ( n43815 , n43814 );
buf ( n43816 , n43815 );
buf ( n43817 , n43249 );
or ( n43818 , n43816 , n43817 );
buf ( n43819 , n43818 );
buf ( n43820 , n43819 );
and ( n43821 , n43801 , n43808 , n43820 );
buf ( n43822 , n43821 );
buf ( n43823 , n43822 );
buf ( n43824 , n43216 );
buf ( n43825 , n43222 );
or ( n43826 , n43824 , n43825 );
buf ( n43827 , n43826 );
buf ( n43828 , n43827 );
not ( n43829 , n43828 );
buf ( n43830 , n43205 );
buf ( n43831 , n43211 );
nor ( n43832 , n43830 , n43831 );
buf ( n43833 , n43832 );
buf ( n43834 , n43833 );
buf ( n43835 , n43200 );
buf ( n43836 , n43194 );
nand ( n43837 , n43835 , n43836 );
buf ( n43838 , n43837 );
buf ( n43839 , n43838 );
or ( n43840 , n43834 , n43839 );
buf ( n43841 , n43205 );
buf ( n43842 , n43211 );
nand ( n43843 , n43841 , n43842 );
buf ( n43844 , n43843 );
buf ( n43845 , n43844 );
nand ( n43846 , n43840 , n43845 );
buf ( n43847 , n43846 );
buf ( n43848 , n43847 );
not ( n43849 , n43848 );
or ( n43850 , n43829 , n43849 );
buf ( n43851 , n43216 );
buf ( n43852 , n43222 );
nand ( n43853 , n43851 , n43852 );
buf ( n43854 , n43853 );
buf ( n43855 , n43854 );
nand ( n43856 , n43850 , n43855 );
buf ( n43857 , n43856 );
buf ( n43858 , n43857 );
not ( n43859 , n43858 );
buf ( n43860 , n36192 );
buf ( n43861 , n27183 );
xor ( n43862 , n43860 , n43861 );
buf ( n43863 , n42127 );
xor ( n43864 , n43862 , n43863 );
buf ( n43865 , n43864 );
buf ( n43866 , n43865 );
buf ( n43867 , n43227 );
nor ( n43868 , n43866 , n43867 );
buf ( n43869 , n43868 );
buf ( n43870 , n43869 );
not ( n43871 , n43870 );
buf ( n43872 , n43871 );
buf ( n43873 , n43872 );
not ( n43874 , n43873 );
or ( n43875 , n43859 , n43874 );
buf ( n43876 , n43227 );
buf ( n43877 , n43865 );
nand ( n43878 , n43876 , n43877 );
buf ( n43879 , n43878 );
buf ( n43880 , n43879 );
nand ( n43881 , n43875 , n43880 );
buf ( n43882 , n43881 );
buf ( n43883 , n43882 );
not ( n43884 , n43883 );
buf ( n43885 , n43178 );
buf ( n43886 , n36165 );
buf ( n43887 , n36159 );
xor ( n43888 , n43886 , n43887 );
buf ( n43889 , n41860 );
and ( n43890 , n43888 , n43889 );
and ( n43891 , n43886 , n43887 );
or ( n43892 , n43890 , n43891 );
buf ( n43893 , n43892 );
buf ( n43894 , n43893 );
or ( n43895 , n43885 , n43894 );
buf ( n43896 , n43895 );
buf ( n43897 , n43896 );
not ( n43898 , n43897 );
buf ( n43899 , n36184 );
buf ( n43900 , n27468 );
xor ( n43901 , n43899 , n43900 );
buf ( n43902 , n41933 );
and ( n43903 , n43901 , n43902 );
and ( n43904 , n43899 , n43900 );
or ( n43905 , n43903 , n43904 );
buf ( n43906 , n43905 );
buf ( n43907 , n43906 );
xor ( n43908 , n43886 , n43887 );
xor ( n43909 , n43908 , n43889 );
buf ( n43910 , n43909 );
buf ( n43911 , n43910 );
nor ( n43912 , n43907 , n43911 );
buf ( n43913 , n43912 );
buf ( n43914 , n43913 );
xor ( n43915 , n43899 , n43900 );
xor ( n43916 , n43915 , n43902 );
buf ( n43917 , n43916 );
buf ( n43918 , n43917 );
buf ( n43919 , n43172 );
nand ( n43920 , n43918 , n43919 );
buf ( n43921 , n43920 );
buf ( n43922 , n43921 );
or ( n43923 , n43914 , n43922 );
buf ( n43924 , n43906 );
buf ( n43925 , n43910 );
nand ( n43926 , n43924 , n43925 );
buf ( n43927 , n43926 );
buf ( n43928 , n43927 );
nand ( n43929 , n43923 , n43928 );
buf ( n43930 , n43929 );
buf ( n43931 , n43930 );
not ( n43932 , n43931 );
or ( n43933 , n43898 , n43932 );
buf ( n43934 , n43178 );
buf ( n43935 , n43893 );
nand ( n43936 , n43934 , n43935 );
buf ( n43937 , n43936 );
buf ( n43938 , n43937 );
nand ( n43939 , n43933 , n43938 );
buf ( n43940 , n43939 );
buf ( n43941 , n43940 );
not ( n43942 , n43941 );
buf ( n43943 , n43189 );
buf ( n43944 , n43183 );
or ( n43945 , n43943 , n43944 );
buf ( n43946 , n43945 );
buf ( n43947 , n43946 );
not ( n43948 , n43947 );
or ( n43949 , n43942 , n43948 );
buf ( n43950 , n43189 );
buf ( n43951 , n43183 );
nand ( n43952 , n43950 , n43951 );
buf ( n43953 , n43952 );
buf ( n43954 , n43953 );
nand ( n43955 , n43949 , n43954 );
buf ( n43956 , n43955 );
buf ( n43957 , n43956 );
not ( n43958 , n43957 );
buf ( n43959 , n43161 );
buf ( n43960 , n43167 );
xor ( n43961 , n43959 , n43960 );
buf ( n43962 , n43156 );
buf ( n43963 , n35916 );
buf ( n43964 , n35922 );
xor ( n43965 , n43963 , n43964 );
buf ( n43966 , n41946 );
and ( n43967 , n43965 , n43966 );
and ( n43968 , n43963 , n43964 );
or ( n43969 , n43967 , n43968 );
buf ( n43970 , n43969 );
buf ( n43971 , n43970 );
xor ( n43972 , n43962 , n43971 );
xor ( n43973 , n43963 , n43964 );
xor ( n43974 , n43973 , n43966 );
buf ( n43975 , n43974 );
buf ( n43976 , n43975 );
buf ( n43977 , n43150 );
xor ( n43978 , n43976 , n43977 );
buf ( n43979 , n43139 );
buf ( n43980 , n43145 );
xor ( n43981 , n43979 , n43980 );
xor ( n43982 , n35959 , n35963 );
and ( n43983 , n43982 , n30465 );
and ( n43984 , n35959 , n35963 );
or ( n43985 , n43983 , n43984 );
buf ( n43986 , n43985 );
buf ( n43987 , n43134 );
xor ( n43988 , n43986 , n43987 );
buf ( n43989 , n29006 );
buf ( n43990 , n42006 );
xor ( n43991 , n43989 , n43990 );
buf ( n43992 , n43991 );
buf ( n43993 , n43992 );
not ( n43994 , n43993 );
buf ( n43995 , n43994 );
buf ( n43996 , n43995 );
buf ( n43997 , n35972 );
not ( n43998 , n43997 );
buf ( n43999 , n43998 );
buf ( n44000 , n43999 );
and ( n44001 , n43996 , n44000 );
buf ( n44002 , n42038 );
and ( n44003 , n863 , n895 );
buf ( n44004 , n44003 );
buf ( n44005 , n44004 );
nand ( n44006 , n44002 , n44005 );
buf ( n44007 , n44006 );
buf ( n44008 , n44007 );
nor ( n44009 , n44001 , n44008 );
buf ( n44010 , n44009 );
buf ( n44011 , n44010 );
buf ( n44012 , n43995 );
buf ( n44013 , n43999 );
nor ( n44014 , n44012 , n44013 );
buf ( n44015 , n44014 );
buf ( n44016 , n44015 );
nor ( n44017 , n44011 , n44016 );
buf ( n44018 , n44017 );
buf ( n44019 , n44018 );
xor ( n44020 , n35959 , n35963 );
xor ( n44021 , n44020 , n30465 );
buf ( n44022 , n44021 );
and ( n44023 , n43989 , n43990 );
buf ( n44024 , n44023 );
buf ( n44025 , n44024 );
nor ( n44026 , n44022 , n44025 );
buf ( n44027 , n44026 );
buf ( n44028 , n44027 );
or ( n44029 , n44019 , n44028 );
buf ( n44030 , n44021 );
buf ( n44031 , n44024 );
nand ( n44032 , n44030 , n44031 );
buf ( n44033 , n44032 );
buf ( n44034 , n44033 );
nand ( n44035 , n44029 , n44034 );
buf ( n44036 , n44035 );
buf ( n44037 , n44036 );
and ( n44038 , n43988 , n44037 );
and ( n44039 , n43986 , n43987 );
or ( n44040 , n44038 , n44039 );
buf ( n44041 , n44040 );
buf ( n44042 , n44041 );
and ( n44043 , n43981 , n44042 );
and ( n44044 , n43979 , n43980 );
or ( n44045 , n44043 , n44044 );
buf ( n44046 , n44045 );
buf ( n44047 , n44046 );
and ( n44048 , n43978 , n44047 );
and ( n44049 , n43976 , n43977 );
or ( n44050 , n44048 , n44049 );
buf ( n44051 , n44050 );
buf ( n44052 , n44051 );
and ( n44053 , n43972 , n44052 );
and ( n44054 , n43962 , n43971 );
or ( n44055 , n44053 , n44054 );
buf ( n44056 , n44055 );
buf ( n44057 , n44056 );
and ( n44058 , n43961 , n44057 );
and ( n44059 , n43959 , n43960 );
or ( n44060 , n44058 , n44059 );
buf ( n44061 , n44060 );
buf ( n44062 , n44061 );
buf ( n44063 , n43946 );
buf ( n44064 , n43913 );
buf ( n44065 , n43917 );
buf ( n44066 , n43172 );
nor ( n44067 , n44065 , n44066 );
buf ( n44068 , n44067 );
buf ( n44069 , n44068 );
nor ( n44070 , n44064 , n44069 );
buf ( n44071 , n44070 );
buf ( n44072 , n44071 );
buf ( n44073 , n43896 );
and ( n44074 , n44072 , n44073 );
buf ( n44075 , n44074 );
buf ( n44076 , n44075 );
nand ( n44077 , n44062 , n44063 , n44076 );
buf ( n44078 , n44077 );
buf ( n44079 , n44078 );
nand ( n44080 , n43958 , n44079 );
buf ( n44081 , n44080 );
buf ( n44082 , n44081 );
buf ( n44083 , n43869 );
buf ( n44084 , n43827 );
not ( n44085 , n44084 );
buf ( n44086 , n44085 );
buf ( n44087 , n44086 );
nor ( n44088 , n44083 , n44087 );
buf ( n44089 , n44088 );
buf ( n44090 , n44089 );
buf ( n44091 , n43833 );
not ( n44092 , n44091 );
buf ( n44093 , n44092 );
buf ( n44094 , n44093 );
buf ( n44095 , n43200 );
buf ( n44096 , n43194 );
or ( n44097 , n44095 , n44096 );
buf ( n44098 , n44097 );
buf ( n44099 , n44098 );
nand ( n44100 , n44082 , n44090 , n44094 , n44099 );
buf ( n44101 , n44100 );
buf ( n44102 , n44101 );
nand ( n44103 , n43884 , n44102 );
buf ( n44104 , n44103 );
buf ( n44105 , n44104 );
buf ( n44106 , n43233 );
not ( n44107 , n35628 );
buf ( n44108 , n35645 );
not ( n44109 , n44108 );
or ( n44110 , n44107 , n44109 );
or ( n44111 , n44108 , n35628 );
not ( n44112 , n41532 );
not ( n44113 , n44112 );
nand ( n44114 , n44111 , n44113 );
nand ( n44115 , n44110 , n44114 );
buf ( n44116 , n44115 );
or ( n44117 , n44106 , n44116 );
buf ( n44118 , n44117 );
buf ( n44119 , n44118 );
not ( n44120 , n44119 );
xor ( n44121 , n43860 , n43861 );
and ( n44122 , n44121 , n43863 );
and ( n44123 , n43860 , n43861 );
or ( n44124 , n44122 , n44123 );
buf ( n44125 , n44124 );
buf ( n44126 , n44125 );
buf ( n44127 , n35662 );
buf ( n44128 , n27054 );
xor ( n44129 , n44127 , n44128 );
buf ( n44130 , n41576 );
xor ( n44131 , n44129 , n44130 );
buf ( n44132 , n44131 );
buf ( n44133 , n44132 );
nor ( n44134 , n44126 , n44133 );
buf ( n44135 , n44134 );
buf ( n44136 , n44135 );
not ( n44137 , n44136 );
xor ( n44138 , n44108 , n35628 );
not ( n44139 , n35676 );
xor ( n44140 , n44139 , n35672 );
buf ( n44141 , n41667 );
and ( n44142 , n44140 , n44141 );
and ( n44143 , n44139 , n35672 );
or ( n44144 , n44142 , n44143 );
or ( n44145 , n44138 , n44144 , n44113 );
not ( n44146 , n44144 );
nand ( n44147 , n44146 , n44113 , n44138 );
nand ( n44148 , n44145 , n44147 );
not ( n44149 , n44148 );
buf ( n44150 , n44149 );
xor ( n44151 , n44127 , n44128 );
and ( n44152 , n44151 , n44130 );
and ( n44153 , n44127 , n44128 );
or ( n44154 , n44152 , n44153 );
buf ( n44155 , n44154 );
buf ( n44156 , n44155 );
xor ( n44157 , n44139 , n35672 );
xor ( n44158 , n44157 , n44141 );
buf ( n44159 , n44158 );
nor ( n44160 , n44156 , n44159 );
buf ( n44161 , n44160 );
buf ( n44162 , n44161 );
not ( n44163 , n44162 );
buf ( n44164 , n44163 );
buf ( n44165 , n44164 );
nand ( n44166 , n44137 , n44150 , n44165 );
buf ( n44167 , n44166 );
buf ( n44168 , n44167 );
nor ( n44169 , n44120 , n44168 );
buf ( n44170 , n44169 );
buf ( n44171 , n44170 );
and ( n44172 , n43823 , n44105 , n44171 );
buf ( n44173 , n44172 );
buf ( n44174 , n44173 );
buf ( n44175 , n43822 );
buf ( n44176 , n44118 );
not ( n44177 , n44176 );
not ( n44178 , n44161 );
buf ( n44179 , n44125 );
buf ( n44180 , n44132 );
nand ( n44181 , n44179 , n44180 );
buf ( n44182 , n44181 );
not ( n44183 , n44182 );
and ( n44184 , n44178 , n44183 );
buf ( n44185 , n44155 );
buf ( n44186 , n44158 );
and ( n44187 , n44185 , n44186 );
buf ( n44188 , n44187 );
nor ( n44189 , n44184 , n44188 );
buf ( n44190 , n44189 );
buf ( n44191 , n44148 );
or ( n44192 , n44190 , n44191 );
xor ( n44193 , n44113 , n44138 );
buf ( n44194 , n44193 );
buf ( n44195 , n44144 );
nand ( n44196 , n44194 , n44195 );
buf ( n44197 , n44196 );
buf ( n44198 , n44197 );
nand ( n44199 , n44192 , n44198 );
buf ( n44200 , n44199 );
buf ( n44201 , n44200 );
not ( n44202 , n44201 );
or ( n44203 , n44177 , n44202 );
buf ( n44204 , n43233 );
buf ( n44205 , n44115 );
nand ( n44206 , n44204 , n44205 );
buf ( n44207 , n44206 );
buf ( n44208 , n44207 );
nand ( n44209 , n44203 , n44208 );
buf ( n44210 , n44209 );
buf ( n44211 , n44210 );
nand ( n44212 , n44175 , n44211 );
buf ( n44213 , n44212 );
buf ( n44214 , n43807 );
not ( n44215 , n44214 );
buf ( n44216 , n43789 );
buf ( n44217 , n43793 );
buf ( n44218 , n43238 );
nand ( n44219 , n44217 , n44218 );
buf ( n44220 , n44219 );
buf ( n44221 , n44220 );
or ( n44222 , n44216 , n44221 );
buf ( n44223 , n43786 );
buf ( n44224 , n43777 );
nand ( n44225 , n44223 , n44224 );
buf ( n44226 , n44225 );
buf ( n44227 , n44226 );
nand ( n44228 , n44222 , n44227 );
buf ( n44229 , n44228 );
buf ( n44230 , n44229 );
not ( n44231 , n44230 );
or ( n44232 , n44215 , n44231 );
nand ( n44233 , n43244 , n43806 );
buf ( n44234 , n44233 );
nand ( n44235 , n44232 , n44234 );
buf ( n44236 , n44235 );
buf ( n44237 , n44236 );
buf ( n44238 , n43819 );
nand ( n44239 , n44237 , n44238 );
buf ( n44240 , n44239 );
buf ( n44241 , n43249 );
buf ( n44242 , n43815 );
nand ( n44243 , n44241 , n44242 );
buf ( n44244 , n44243 );
nand ( n44245 , n44213 , n44240 , n44244 );
buf ( n44246 , n44245 );
or ( n44247 , n44174 , n44246 );
buf ( n44248 , n43279 );
not ( n44249 , n44248 );
xor ( n44250 , n35506 , n41132 );
not ( n44251 , n36243 );
and ( n44252 , n44250 , n44251 );
and ( n44253 , n35506 , n41132 );
or ( n44254 , n44252 , n44253 );
not ( n44255 , n44254 );
buf ( n44256 , n44255 );
nand ( n44257 , n44249 , n44256 );
buf ( n44258 , n44257 );
buf ( n44259 , n44258 );
xor ( n44260 , n35506 , n41132 );
not ( n44261 , n36243 );
xor ( n44262 , n44260 , n44261 );
buf ( n44263 , n44262 );
buf ( n44264 , n43261 );
or ( n44265 , n44263 , n44264 );
buf ( n44266 , n44265 );
buf ( n44267 , n44266 );
not ( n44268 , n44267 );
buf ( n44269 , n43256 );
buf ( n44270 , n43272 );
nor ( n44271 , n44269 , n44270 );
buf ( n44272 , n44271 );
buf ( n44273 , n44272 );
not ( n44274 , n44273 );
buf ( n44275 , n44274 );
buf ( n44276 , n44275 );
buf ( n44277 , n43267 );
xor ( n44278 , n43809 , n43811 );
and ( n44279 , n44278 , n43813 );
and ( n44280 , n43809 , n43811 );
or ( n44281 , n44279 , n44280 );
buf ( n44282 , n44281 );
buf ( n44283 , n44282 );
or ( n44284 , n44277 , n44283 );
buf ( n44285 , n44284 );
buf ( n44286 , n44285 );
nand ( n44287 , n44276 , n44286 );
buf ( n44288 , n44287 );
buf ( n44289 , n44288 );
nor ( n44290 , n44268 , n44289 );
buf ( n44291 , n44290 );
buf ( n44292 , n44291 );
and ( n44293 , n44259 , n44292 );
buf ( n44294 , n44293 );
buf ( n44295 , n44294 );
nand ( n44296 , n44247 , n44295 );
buf ( n44297 , n44296 );
buf ( n44298 , n44297 );
not ( n44299 , n44298 );
buf ( n44300 , n44266 );
not ( n44301 , n44300 );
buf ( n44302 , n44272 );
buf ( n44303 , n43267 );
buf ( n44304 , n44282 );
nand ( n44305 , n44303 , n44304 );
buf ( n44306 , n44305 );
buf ( n44307 , n44306 );
or ( n44308 , n44302 , n44307 );
buf ( n44309 , n43272 );
buf ( n44310 , n43256 );
nand ( n44311 , n44309 , n44310 );
buf ( n44312 , n44311 );
buf ( n44313 , n44312 );
nand ( n44314 , n44308 , n44313 );
buf ( n44315 , n44314 );
buf ( n44316 , n44315 );
not ( n44317 , n44316 );
or ( n44318 , n44301 , n44317 );
buf ( n44319 , n44262 );
buf ( n44320 , n43261 );
nand ( n44321 , n44319 , n44320 );
buf ( n44322 , n44321 );
buf ( n44323 , n44322 );
nand ( n44324 , n44318 , n44323 );
buf ( n44325 , n44324 );
buf ( n44326 , n44325 );
not ( n44327 , n44326 );
buf ( n44328 , n44258 );
not ( n44329 , n44328 );
or ( n44330 , n44327 , n44329 );
buf ( n44331 , n44255 );
not ( n44332 , n44331 );
buf ( n44333 , n43279 );
nand ( n44334 , n44332 , n44333 );
buf ( n44335 , n44334 );
buf ( n44336 , n44335 );
nand ( n44337 , n44330 , n44336 );
buf ( n44338 , n44337 );
buf ( n44339 , n44338 );
not ( n44340 , n44339 );
buf ( n44341 , n44340 );
buf ( n44342 , n44341 );
not ( n44343 , n44342 );
or ( n44344 , n44299 , n44343 );
buf ( n44345 , n43309 );
not ( n44346 , n44345 );
buf ( n44347 , n43317 );
not ( n44348 , n44347 );
buf ( n44349 , n44348 );
buf ( n44350 , n44349 );
nand ( n44351 , n44346 , n44350 );
buf ( n44352 , n44351 );
buf ( n44353 , n44352 );
buf ( n44354 , n43304 );
buf ( n44355 , n35247 );
buf ( n44356 , n44355 );
buf ( n44357 , n44356 );
buf ( n44358 , n36271 );
buf ( n44359 , n44358 );
xor ( n44360 , n44357 , n44359 );
buf ( n44361 , n40734 );
and ( n44362 , n44360 , n44361 );
and ( n44363 , n44357 , n44359 );
or ( n44364 , n44362 , n44363 );
buf ( n44365 , n44364 );
buf ( n44366 , n44365 );
or ( n44367 , n44354 , n44366 );
buf ( n44368 , n44367 );
buf ( n44369 , n44368 );
nand ( n44370 , n44353 , n44369 );
buf ( n44371 , n44370 );
buf ( n44372 , n44371 );
buf ( n44373 , n43296 );
xor ( n44374 , n44357 , n44359 );
xor ( n44375 , n44374 , n44361 );
buf ( n44376 , n44375 );
buf ( n44377 , n44376 );
nor ( n44378 , n44373 , n44377 );
buf ( n44379 , n44378 );
buf ( n44380 , n44379 );
not ( n44381 , n44380 );
buf ( n44382 , n43291 );
buf ( n44383 , n43284 );
or ( n44384 , n44382 , n44383 );
buf ( n44385 , n44384 );
buf ( n44386 , n44385 );
nand ( n44387 , n44381 , n44386 );
buf ( n44388 , n44387 );
buf ( n44389 , n44388 );
nor ( n44390 , n44372 , n44389 );
buf ( n44391 , n44390 );
buf ( n44392 , n44391 );
nand ( n44393 , n44344 , n44392 );
buf ( n44394 , n44393 );
buf ( n44395 , n44394 );
buf ( n44396 , n44371 );
not ( n44397 , n44396 );
buf ( n44398 , n44397 );
buf ( n44399 , n44398 );
buf ( n44400 , n44379 );
buf ( n44401 , n43284 );
buf ( n44402 , n43291 );
nand ( n44403 , n44401 , n44402 );
buf ( n44404 , n44403 );
buf ( n44405 , n44404 );
or ( n44406 , n44400 , n44405 );
buf ( n44407 , n43296 );
buf ( n44408 , n44376 );
nand ( n44409 , n44407 , n44408 );
buf ( n44410 , n44409 );
buf ( n44411 , n44410 );
nand ( n44412 , n44406 , n44411 );
buf ( n44413 , n44412 );
buf ( n44414 , n44413 );
and ( n44415 , n44399 , n44414 );
buf ( n44416 , n44365 );
buf ( n44417 , n43304 );
and ( n44418 , n44416 , n44417 );
buf ( n44419 , n44418 );
buf ( n44420 , n44419 );
not ( n44421 , n44420 );
buf ( n44422 , n44352 );
not ( n44423 , n44422 );
or ( n44424 , n44421 , n44423 );
buf ( n44425 , n44349 );
not ( n44426 , n44425 );
buf ( n44427 , n43309 );
nand ( n44428 , n44426 , n44427 );
buf ( n44429 , n44428 );
buf ( n44430 , n44429 );
nand ( n44431 , n44424 , n44430 );
buf ( n44432 , n44431 );
buf ( n44433 , n44432 );
nor ( n44434 , n44415 , n44433 );
buf ( n44435 , n44434 );
buf ( n44436 , n44435 );
nand ( n44437 , n44395 , n44436 );
buf ( n44438 , n44437 );
buf ( n44439 , n44438 );
buf ( n44440 , n43341 );
buf ( n44441 , n34000 );
buf ( n44442 , n33995 );
buf ( n44443 , n44442 );
xor ( n44444 , n44441 , n44443 );
buf ( n44445 , n40377 );
and ( n44446 , n44444 , n44445 );
and ( n44447 , n44441 , n44443 );
or ( n44448 , n44446 , n44447 );
buf ( n44449 , n44448 );
buf ( n44450 , n44449 );
nor ( n44451 , n44440 , n44450 );
buf ( n44452 , n44451 );
buf ( n44453 , n44452 );
buf ( n44454 , n43346 );
xor ( n44455 , n33598 , n33604 );
xor ( n44456 , n44455 , n40364 );
buf ( n44457 , n44456 );
nor ( n44458 , n44454 , n44457 );
buf ( n44459 , n44458 );
buf ( n44460 , n44459 );
nor ( n44461 , n44453 , n44460 );
buf ( n44462 , n44461 );
buf ( n44463 , n44462 );
buf ( n44464 , n43352 );
not ( n44465 , n44464 );
xor ( n44466 , n33598 , n33604 );
and ( n44467 , n44466 , n40364 );
and ( n44468 , n33598 , n33604 );
nor ( n44469 , n44467 , n44468 );
buf ( n44470 , n44469 );
nand ( n44471 , n44465 , n44470 );
buf ( n44472 , n44471 );
buf ( n44473 , n44472 );
xor ( n44474 , n43652 , n43653 );
xor ( n44475 , n44474 , n43655 );
buf ( n44476 , n44475 );
buf ( n44477 , n44476 );
buf ( n44478 , n43357 );
or ( n44479 , n44477 , n44478 );
buf ( n44480 , n44479 );
buf ( n44481 , n44480 );
and ( n44482 , n44463 , n44473 , n44481 );
buf ( n44483 , n44482 );
buf ( n44484 , n44483 );
not ( n44485 , n44484 );
buf ( n44486 , n44485 );
buf ( n44487 , n44486 );
buf ( n44488 , n33985 );
buf ( n44489 , n23015 );
xor ( n44490 , n44488 , n44489 );
buf ( n44491 , n40636 );
and ( n44492 , n44490 , n44491 );
and ( n44493 , n44488 , n44489 );
or ( n44494 , n44492 , n44493 );
buf ( n44495 , n44494 );
buf ( n44496 , n44495 );
xor ( n44497 , n44441 , n44443 );
xor ( n44498 , n44497 , n44445 );
buf ( n44499 , n44498 );
buf ( n44500 , n44499 );
or ( n44501 , n44496 , n44500 );
buf ( n44502 , n44501 );
buf ( n44503 , n44502 );
xor ( n44504 , n44488 , n44489 );
xor ( n44505 , n44504 , n44491 );
buf ( n44506 , n44505 );
buf ( n44507 , n44506 );
buf ( n44508 , n43334 );
or ( n44509 , n44507 , n44508 );
buf ( n44510 , n44509 );
buf ( n44511 , n44510 );
and ( n44512 , n44503 , n44511 );
buf ( n44513 , n44512 );
buf ( n44514 , n44513 );
buf ( n44515 , n24855 );
buf ( n44516 , n33978 );
xor ( n44517 , n44515 , n44516 );
buf ( n44518 , n40592 );
xor ( n44519 , n44517 , n44518 );
buf ( n44520 , n44519 );
buf ( n44521 , n44520 );
buf ( n44522 , n43322 );
nor ( n44523 , n44521 , n44522 );
buf ( n44524 , n44523 );
buf ( n44525 , n44524 );
xor ( n44526 , n44515 , n44516 );
and ( n44527 , n44526 , n44518 );
and ( n44528 , n44515 , n44516 );
or ( n44529 , n44527 , n44528 );
buf ( n44530 , n44529 );
buf ( n44531 , n44530 );
buf ( n44532 , n43329 );
nor ( n44533 , n44531 , n44532 );
buf ( n44534 , n44533 );
buf ( n44535 , n44534 );
nor ( n44536 , n44525 , n44535 );
buf ( n44537 , n44536 );
buf ( n44538 , n44537 );
nand ( n44539 , n44514 , n44538 );
buf ( n44540 , n44539 );
buf ( n44541 , n44540 );
nor ( n44542 , n44487 , n44541 );
buf ( n44543 , n44542 );
buf ( n44544 , n44543 );
nand ( n44545 , n43770 , n44439 , n44544 );
buf ( n44546 , n44545 );
buf ( n44547 , n44546 );
buf ( n44548 , n43769 );
buf ( n44549 , n44513 );
not ( n44550 , n44549 );
buf ( n44551 , n44520 );
buf ( n44552 , n43322 );
nand ( n44553 , n44551 , n44552 );
buf ( n44554 , n44553 );
buf ( n44555 , n44554 );
buf ( n44556 , n44534 );
or ( n44557 , n44555 , n44556 );
buf ( n44558 , n44530 );
buf ( n44559 , n43329 );
nand ( n44560 , n44558 , n44559 );
buf ( n44561 , n44560 );
buf ( n44562 , n44561 );
nand ( n44563 , n44557 , n44562 );
buf ( n44564 , n44563 );
buf ( n44565 , n44564 );
not ( n44566 , n44565 );
or ( n44567 , n44550 , n44566 );
buf ( n44568 , n43334 );
buf ( n44569 , n44506 );
and ( n44570 , n44568 , n44569 );
buf ( n44571 , n44570 );
buf ( n44572 , n44571 );
not ( n44573 , n44572 );
buf ( n44574 , n44502 );
not ( n44575 , n44574 );
or ( n44576 , n44573 , n44575 );
buf ( n44577 , n44495 );
buf ( n44578 , n44499 );
nand ( n44579 , n44577 , n44578 );
buf ( n44580 , n44579 );
buf ( n44581 , n44580 );
nand ( n44582 , n44576 , n44581 );
buf ( n44583 , n44582 );
buf ( n44584 , n44583 );
not ( n44585 , n44584 );
buf ( n44586 , n44585 );
buf ( n44587 , n44586 );
nand ( n44588 , n44567 , n44587 );
buf ( n44589 , n44588 );
buf ( n44590 , n44589 );
buf ( n44591 , n44483 );
nand ( n44592 , n44590 , n44591 );
buf ( n44593 , n44592 );
buf ( n44594 , n44593 );
buf ( n44595 , n44472 );
not ( n44596 , n44595 );
buf ( n44597 , n44459 );
buf ( n44598 , n43341 );
buf ( n44599 , n44449 );
nand ( n44600 , n44598 , n44599 );
buf ( n44601 , n44600 );
buf ( n44602 , n44601 );
or ( n44603 , n44597 , n44602 );
buf ( n44604 , n43346 );
buf ( n44605 , n44456 );
nand ( n44606 , n44604 , n44605 );
buf ( n44607 , n44606 );
buf ( n44608 , n44607 );
nand ( n44609 , n44603 , n44608 );
buf ( n44610 , n44609 );
buf ( n44611 , n44610 );
not ( n44612 , n44611 );
or ( n44613 , n44596 , n44612 );
buf ( n44614 , n44469 );
not ( n44615 , n44614 );
buf ( n44616 , n43352 );
nand ( n44617 , n44615 , n44616 );
buf ( n44618 , n44617 );
buf ( n44619 , n44618 );
nand ( n44620 , n44613 , n44619 );
buf ( n44621 , n44620 );
buf ( n44622 , n44621 );
buf ( n44623 , n44480 );
nand ( n44624 , n44622 , n44623 );
buf ( n44625 , n44624 );
buf ( n44626 , n44625 );
buf ( n44627 , n43357 );
buf ( n44628 , n44476 );
nand ( n44629 , n44627 , n44628 );
buf ( n44630 , n44629 );
buf ( n44631 , n44630 );
nand ( n44632 , n44594 , n44626 , n44631 );
buf ( n44633 , n44632 );
buf ( n44634 , n44633 );
nand ( n44635 , n44548 , n44634 );
buf ( n44636 , n44635 );
buf ( n44637 , n44636 );
nand ( n44638 , n43755 , n44547 , n44637 );
buf ( n44639 , n44638 );
buf ( n44640 , n44639 );
not ( n44641 , n44640 );
or ( n44642 , n43583 , n44641 );
buf ( n44643 , n43506 );
not ( n44644 , n44643 );
buf ( n44645 , n43496 );
not ( n44646 , n44645 );
buf ( n44647 , n43414 );
buf ( n44648 , n43517 );
nand ( n44649 , n44647 , n44648 );
buf ( n44650 , n44649 );
buf ( n44651 , n44650 );
buf ( n44652 , n43530 );
or ( n44653 , n44651 , n44652 );
buf ( n44654 , n43523 );
buf ( n44655 , n43529 );
nand ( n44656 , n44654 , n44655 );
buf ( n44657 , n44656 );
buf ( n44658 , n44657 );
nand ( n44659 , n44653 , n44658 );
buf ( n44660 , n44659 );
buf ( n44661 , n44660 );
not ( n44662 , n44661 );
or ( n44663 , n44646 , n44662 );
buf ( n44664 , n43493 );
not ( n44665 , n44664 );
buf ( n44666 , n43487 );
nand ( n44667 , n44665 , n44666 );
buf ( n44668 , n44667 );
buf ( n44669 , n44668 );
nand ( n44670 , n44663 , n44669 );
buf ( n44671 , n44670 );
buf ( n44672 , n44671 );
not ( n44673 , n44672 );
or ( n44674 , n44644 , n44673 );
buf ( n44675 , n43502 );
buf ( n44676 , n43431 );
nand ( n44677 , n44675 , n44676 );
buf ( n44678 , n44677 );
buf ( n44679 , n44678 );
nand ( n44680 , n44674 , n44679 );
buf ( n44681 , n44680 );
buf ( n44682 , n43578 );
not ( n44683 , n44682 );
buf ( n44684 , n44683 );
and ( n44685 , n44681 , n44684 );
buf ( n44686 , n43572 );
not ( n44687 , n44686 );
buf ( n44688 , n44687 );
buf ( n44689 , n44688 );
not ( n44690 , n44689 );
buf ( n44691 , n43559 );
buf ( n44692 , n43436 );
buf ( n44693 , n43546 );
nand ( n44694 , n44692 , n44693 );
buf ( n44695 , n44694 );
buf ( n44696 , n44695 );
or ( n44697 , n44691 , n44696 );
buf ( n44698 , n43375 );
buf ( n44699 , n43556 );
nand ( n44700 , n44698 , n44699 );
buf ( n44701 , n44700 );
buf ( n44702 , n44701 );
nand ( n44703 , n44697 , n44702 );
buf ( n44704 , n44703 );
buf ( n44705 , n44704 );
not ( n44706 , n44705 );
or ( n44707 , n44690 , n44706 );
buf ( n44708 , n43380 );
buf ( n44709 , n43111 );
nand ( n44710 , n44708 , n44709 );
buf ( n44711 , n44710 );
buf ( n44712 , n44711 );
nand ( n44713 , n44707 , n44712 );
buf ( n44714 , n44713 );
buf ( n44715 , n43567 );
not ( n44716 , n44715 );
buf ( n44717 , n44716 );
and ( n44718 , n44714 , n44717 );
buf ( n44719 , n43420 );
buf ( n44720 , n43116 );
and ( n44721 , n44719 , n44720 );
buf ( n44722 , n44721 );
nor ( n44723 , n44685 , n44718 , n44722 );
buf ( n44724 , n44723 );
nand ( n44725 , n44642 , n44724 );
buf ( n44726 , n44725 );
buf ( n44727 , n44726 );
buf ( n44728 , n43100 );
buf ( n44729 , n43425 );
or ( n44730 , n44728 , n44729 );
buf ( n44731 , n44730 );
buf ( n44732 , n44731 );
nand ( n44733 , n44727 , n44732 );
buf ( n44734 , n44733 );
buf ( n44735 , n43089 );
buf ( n44736 , n43105 );
nor ( n44737 , n44735 , n44736 );
buf ( n44738 , n44737 );
not ( n44739 , n44738 );
buf ( n44740 , n43094 );
buf ( n44741 , n43123 );
or ( n44742 , n44740 , n44741 );
buf ( n44743 , n44742 );
buf ( n44744 , n43128 );
buf ( n44745 , n43446 );
or ( n44746 , n44744 , n44745 );
buf ( n44747 , n44746 );
nand ( n44748 , n44739 , n44743 , n44747 );
or ( n44749 , n44734 , n44748 );
buf ( n44750 , n44743 );
not ( n44751 , n44750 );
buf ( n44752 , n43100 );
buf ( n44753 , n43425 );
nand ( n44754 , n44752 , n44753 );
buf ( n44755 , n44754 );
or ( n44756 , n44738 , n44755 );
buf ( n44757 , n43089 );
buf ( n44758 , n43105 );
nand ( n44759 , n44757 , n44758 );
buf ( n44760 , n44759 );
nand ( n44761 , n44756 , n44760 );
buf ( n44762 , n44761 );
not ( n44763 , n44762 );
or ( n44764 , n44751 , n44763 );
buf ( n44765 , n43094 );
buf ( n44766 , n43123 );
nand ( n44767 , n44765 , n44766 );
buf ( n44768 , n44767 );
buf ( n44769 , n44768 );
nand ( n44770 , n44764 , n44769 );
buf ( n44771 , n44770 );
and ( n44772 , n44771 , n44747 );
buf ( n44773 , n43128 );
buf ( n44774 , n43446 );
and ( n44775 , n44773 , n44774 );
buf ( n44776 , n44775 );
nor ( n44777 , n44772 , n44776 );
nand ( n44778 , n44749 , n44777 );
buf ( n44779 , n44778 );
not ( n44780 , n44779 );
or ( n44781 , n43481 , n44780 );
buf ( n44782 , n43448 );
buf ( n44783 , n43440 );
nand ( n44784 , n44782 , n44783 );
buf ( n44785 , n44784 );
buf ( n44786 , n44785 );
not ( n44787 , n44786 );
buf ( n44788 , n43476 );
not ( n44789 , n44788 );
and ( n44790 , n44787 , n44789 );
buf ( n44791 , n43442 );
buf ( n44792 , n43452 );
and ( n44793 , n44791 , n44792 );
buf ( n44794 , n44793 );
buf ( n44795 , n44794 );
nor ( n44796 , n44790 , n44795 );
buf ( n44797 , n44796 );
buf ( n44798 , n44797 );
nand ( n44799 , n44781 , n44798 );
buf ( n44800 , n44799 );
buf ( n44801 , n44800 );
xor ( n44802 , n43465 , n43466 );
xor ( n44803 , n44802 , n44801 );
buf ( n44804 , n44803 );
xor ( n44805 , n43465 , n43466 );
and ( n44806 , n44805 , n44801 );
and ( n44807 , n43465 , n43466 );
or ( n44808 , n44806 , n44807 );
buf ( n44809 , n44808 );
buf ( n44810 , n44776 );
not ( n44811 , n44810 );
buf ( n44812 , n44747 );
nand ( n44813 , n44811 , n44812 );
buf ( n44814 , n44813 );
buf ( n44815 , n44814 );
buf ( n44816 , n44814 );
not ( n44817 , n44816 );
buf ( n44818 , n44817 );
buf ( n44819 , n44818 );
buf ( n44820 , n44743 );
not ( n44821 , n44820 );
or ( n44822 , n44734 , n44738 );
not ( n44823 , n44761 );
nand ( n44824 , n44822 , n44823 );
buf ( n44825 , n44824 );
not ( n44826 , n44825 );
or ( n44827 , n44821 , n44826 );
buf ( n44828 , n44768 );
nand ( n44829 , n44827 , n44828 );
buf ( n44830 , n44829 );
buf ( n44831 , n44830 );
and ( n44832 , n44831 , n44819 );
not ( n44833 , n44831 );
and ( n44834 , n44833 , n44815 );
nor ( n44835 , n44832 , n44834 );
buf ( n44836 , n44835 );
buf ( n44837 , n43629 );
buf ( n44838 , n43604 );
not ( n44839 , n44838 );
buf ( n44840 , n43766 );
not ( n44841 , n44840 );
buf ( n44842 , n44486 );
buf ( n44843 , n44540 );
not ( n44844 , n44843 );
buf ( n44845 , n44438 );
nand ( n44846 , n44844 , n44845 );
buf ( n44847 , n44846 );
buf ( n44848 , n44847 );
or ( n44849 , n44842 , n44848 );
buf ( n44850 , n44633 );
not ( n44851 , n44850 );
buf ( n44852 , n44851 );
buf ( n44853 , n44852 );
nand ( n44854 , n44849 , n44853 );
buf ( n44855 , n44854 );
buf ( n44856 , n44855 );
not ( n44857 , n44856 );
or ( n44858 , n44841 , n44857 );
buf ( n44859 , n43701 );
not ( n44860 , n44859 );
buf ( n44861 , n44860 );
buf ( n44862 , n44861 );
nand ( n44863 , n44858 , n44862 );
buf ( n44864 , n44863 );
buf ( n44865 , n44864 );
not ( n44866 , n44865 );
or ( n44867 , n44839 , n44866 );
buf ( n44868 , n43725 );
not ( n44869 , n44868 );
buf ( n44870 , n44869 );
buf ( n44871 , n44870 );
nand ( n44872 , n44867 , n44871 );
buf ( n44873 , n44872 );
buf ( n44874 , n44873 );
buf ( n44875 , n43733 );
not ( n44876 , n44837 );
not ( n44877 , n44874 );
or ( n44878 , n44876 , n44877 );
nand ( n44879 , n44878 , n44875 );
buf ( n44880 , n44879 );
buf ( n44881 , n43685 );
not ( n44882 , n43763 );
and ( n44883 , n44855 , n43758 );
not ( n44884 , n44883 );
or ( n44885 , n44882 , n44884 );
buf ( n44886 , n43675 );
not ( n44887 , n44886 );
buf ( n44888 , n44887 );
nand ( n44889 , n44885 , n44888 );
buf ( n44890 , n44889 );
buf ( n44891 , n43689 );
not ( n44892 , n44881 );
not ( n44893 , n44890 );
or ( n44894 , n44892 , n44893 );
nand ( n44895 , n44894 , n44891 );
buf ( n44896 , n44895 );
buf ( n44897 , n43549 );
not ( n44898 , n44897 );
buf ( n44899 , n44898 );
buf ( n44900 , n44899 );
buf ( n44901 , n43536 );
not ( n44902 , n44901 );
buf ( n44903 , n44902 );
buf ( n44904 , n44903 );
not ( n44905 , n44904 );
buf ( n44906 , n44639 );
not ( n44907 , n44906 );
or ( n44908 , n44905 , n44907 );
buf ( n44909 , n44681 );
not ( n44910 , n44909 );
buf ( n44911 , n44910 );
buf ( n44912 , n44911 );
nand ( n44913 , n44908 , n44912 );
buf ( n44914 , n44913 );
buf ( n44915 , n44914 );
buf ( n44916 , n44695 );
not ( n44917 , n44900 );
not ( n44918 , n44915 );
or ( n44919 , n44917 , n44918 );
nand ( n44920 , n44919 , n44916 );
buf ( n44921 , n44920 );
buf ( n44922 , n43601 );
not ( n44923 , n44922 );
buf ( n44924 , n44923 );
buf ( n44925 , n44924 );
buf ( n44926 , n44864 );
buf ( n44927 , n43710 );
not ( n44928 , n44927 );
buf ( n44929 , n44928 );
buf ( n44930 , n44929 );
not ( n44931 , n44925 );
not ( n44932 , n44926 );
or ( n44933 , n44931 , n44932 );
nand ( n44934 , n44933 , n44930 );
buf ( n44935 , n44934 );
buf ( n44936 , n43562 );
buf ( n44937 , n44914 );
buf ( n44938 , n44704 );
not ( n44939 , n44938 );
buf ( n44940 , n44939 );
buf ( n44941 , n44940 );
not ( n44942 , n44936 );
not ( n44943 , n44937 );
or ( n44944 , n44942 , n44943 );
nand ( n44945 , n44944 , n44941 );
buf ( n44946 , n44945 );
buf ( n44947 , n43496 );
buf ( n44948 , n43533 );
not ( n44949 , n44948 );
buf ( n44950 , n44639 );
not ( n44951 , n44950 );
or ( n44952 , n44949 , n44951 );
buf ( n44953 , n44660 );
not ( n44954 , n44953 );
buf ( n44955 , n44954 );
buf ( n44956 , n44955 );
nand ( n44957 , n44952 , n44956 );
buf ( n44958 , n44957 );
buf ( n44959 , n44958 );
buf ( n44960 , n44668 );
not ( n44961 , n44947 );
not ( n44962 , n44959 );
or ( n44963 , n44961 , n44962 );
nand ( n44964 , n44963 , n44960 );
buf ( n44965 , n44964 );
buf ( n44966 , n44472 );
buf ( n44967 , n44462 );
not ( n44968 , n44967 );
buf ( n44969 , n44589 );
not ( n44970 , n44969 );
buf ( n44971 , n44847 );
nand ( n44972 , n44970 , n44971 );
buf ( n44973 , n44972 );
buf ( n44974 , n44973 );
not ( n44975 , n44974 );
or ( n44976 , n44968 , n44975 );
buf ( n44977 , n44610 );
not ( n44978 , n44977 );
buf ( n44979 , n44978 );
buf ( n44980 , n44979 );
nand ( n44981 , n44976 , n44980 );
buf ( n44982 , n44981 );
buf ( n44983 , n44982 );
buf ( n44984 , n44618 );
not ( n44985 , n44966 );
not ( n44986 , n44983 );
or ( n44987 , n44985 , n44986 );
nand ( n44988 , n44987 , n44984 );
buf ( n44989 , n44988 );
buf ( n44990 , n43520 );
not ( n44991 , n44990 );
buf ( n44992 , n44991 );
buf ( n44993 , n44992 );
buf ( n44994 , n44639 );
buf ( n44995 , n44650 );
not ( n44996 , n44993 );
not ( n44997 , n44994 );
or ( n44998 , n44996 , n44997 );
nand ( n44999 , n44998 , n44995 );
buf ( n45000 , n44999 );
buf ( n45001 , n44452 );
not ( n45002 , n45001 );
buf ( n45003 , n45002 );
buf ( n45004 , n45003 );
buf ( n45005 , n44973 );
buf ( n45006 , n44601 );
not ( n45007 , n45004 );
not ( n45008 , n45005 );
or ( n45009 , n45007 , n45008 );
nand ( n45010 , n45009 , n45006 );
buf ( n45011 , n45010 );
buf ( n45012 , n44368 );
buf ( n45013 , n44294 );
not ( n45014 , n45013 );
buf ( n45015 , n43822 );
not ( n45016 , n45015 );
buf ( n45017 , n44170 );
not ( n45018 , n45017 );
buf ( n45019 , n44104 );
not ( n45020 , n45019 );
buf ( n45021 , n45020 );
buf ( n45022 , n45021 );
nor ( n45023 , n45018 , n45022 );
buf ( n45024 , n45023 );
buf ( n45025 , n45024 );
not ( n45026 , n45025 );
or ( n45027 , n45016 , n45026 );
not ( n45028 , n44245 );
buf ( n45029 , n45028 );
nand ( n45030 , n45027 , n45029 );
buf ( n45031 , n45030 );
buf ( n45032 , n45031 );
not ( n45033 , n45032 );
or ( n45034 , n45014 , n45033 );
buf ( n45035 , n44341 );
nand ( n45036 , n45034 , n45035 );
buf ( n45037 , n45036 );
buf ( n45038 , n45037 );
buf ( n45039 , n44385 );
nand ( n45040 , n45038 , n45039 );
buf ( n45041 , n45040 );
buf ( n45042 , n45041 );
buf ( n45043 , n44379 );
or ( n45044 , n45042 , n45043 );
buf ( n45045 , n44413 );
not ( n45046 , n45045 );
buf ( n45047 , n45046 );
buf ( n45048 , n45047 );
nand ( n45049 , n45044 , n45048 );
buf ( n45050 , n45049 );
buf ( n45051 , n45050 );
buf ( n45052 , n44419 );
not ( n45053 , n45052 );
buf ( n45054 , n45053 );
buf ( n45055 , n45054 );
not ( n45056 , n45012 );
not ( n45057 , n45051 );
or ( n45058 , n45056 , n45057 );
nand ( n45059 , n45058 , n45055 );
buf ( n45060 , n45059 );
buf ( n45061 , n44537 );
buf ( n45062 , n44438 );
buf ( n45063 , n44564 );
not ( n45064 , n45063 );
buf ( n45065 , n45064 );
buf ( n45066 , n45065 );
not ( n45067 , n45061 );
not ( n45068 , n45062 );
or ( n45069 , n45067 , n45068 );
nand ( n45070 , n45069 , n45066 );
buf ( n45071 , n45070 );
buf ( n45072 , n44524 );
not ( n45073 , n45072 );
buf ( n45074 , n45073 );
buf ( n45075 , n45074 );
buf ( n45076 , n44438 );
buf ( n45077 , n44554 );
not ( n45078 , n45075 );
not ( n45079 , n45076 );
or ( n45080 , n45078 , n45079 );
nand ( n45081 , n45080 , n45077 );
buf ( n45082 , n45081 );
buf ( n45083 , n45074 );
buf ( n45084 , n44554 );
nand ( n45085 , n45083 , n45084 );
buf ( n45086 , n45085 );
buf ( n45087 , n45086 );
buf ( n45088 , n44438 );
buf ( n45089 , n45086 );
buf ( n45090 , n44438 );
not ( n45091 , n45087 );
not ( n45092 , n45088 );
or ( n45093 , n45091 , n45092 );
or ( n45094 , n45089 , n45090 );
nand ( n45095 , n45093 , n45094 );
buf ( n45096 , n45095 );
buf ( n45097 , n44266 );
buf ( n45098 , n44288 );
not ( n45099 , n45098 );
buf ( n45100 , n45099 );
buf ( n45101 , n45100 );
not ( n45102 , n45101 );
buf ( n45103 , n45031 );
not ( n45104 , n45103 );
or ( n45105 , n45102 , n45104 );
buf ( n45106 , n44315 );
not ( n45107 , n45106 );
buf ( n45108 , n45107 );
buf ( n45109 , n45108 );
nand ( n45110 , n45105 , n45109 );
buf ( n45111 , n45110 );
buf ( n45112 , n45111 );
buf ( n45113 , n44322 );
not ( n45114 , n45097 );
not ( n45115 , n45112 );
or ( n45116 , n45114 , n45115 );
nand ( n45117 , n45116 , n45113 );
buf ( n45118 , n45117 );
buf ( n45119 , n44285 );
buf ( n45120 , n45031 );
buf ( n45121 , n44306 );
not ( n45122 , n45119 );
not ( n45123 , n45120 );
or ( n45124 , n45122 , n45123 );
nand ( n45125 , n45124 , n45121 );
buf ( n45126 , n45125 );
buf ( n45127 , n44285 );
buf ( n45128 , n44306 );
nand ( n45129 , n45127 , n45128 );
buf ( n45130 , n45129 );
buf ( n45131 , n45130 );
buf ( n45132 , n45031 );
buf ( n45133 , n45130 );
buf ( n45134 , n45031 );
not ( n45135 , n45131 );
not ( n45136 , n45132 );
or ( n45137 , n45135 , n45136 );
or ( n45138 , n45133 , n45134 );
nand ( n45139 , n45137 , n45138 );
buf ( n45140 , n45139 );
buf ( n45141 , n44164 );
not ( n45142 , n45141 );
buf ( n45143 , n45021 );
buf ( n45144 , n44135 );
nor ( n45145 , n45143 , n45144 );
buf ( n45146 , n45145 );
buf ( n45147 , n45146 );
not ( n45148 , n45147 );
or ( n45149 , n45142 , n45148 );
buf ( n45150 , n44189 );
nand ( n45151 , n45149 , n45150 );
buf ( n45152 , n45151 );
buf ( n45153 , n45152 );
buf ( n45154 , n44149 );
buf ( n45155 , n44197 );
nand ( n45156 , n45154 , n45155 );
buf ( n45157 , n45156 );
buf ( n45158 , n45157 );
buf ( n45159 , n45157 );
buf ( n45160 , n45152 );
not ( n45161 , n45153 );
not ( n45162 , n45158 );
or ( n45163 , n45161 , n45162 );
or ( n45164 , n45159 , n45160 );
nand ( n45165 , n45163 , n45164 );
buf ( n45166 , n45165 );
buf ( n45167 , n43797 );
not ( n45168 , n45167 );
buf ( n45169 , n45168 );
buf ( n45170 , n45169 );
buf ( n45171 , n45024 );
buf ( n45172 , n44210 );
or ( n45173 , n45171 , n45172 );
buf ( n45174 , n45173 );
buf ( n45175 , n45174 );
buf ( n45176 , n44220 );
not ( n45177 , n45170 );
not ( n45178 , n45175 );
or ( n45179 , n45177 , n45178 );
nand ( n45180 , n45179 , n45176 );
buf ( n45181 , n45180 );
buf ( n45182 , n45169 );
buf ( n45183 , n44220 );
nand ( n45184 , n45182 , n45183 );
buf ( n45185 , n45184 );
buf ( n45186 , n45185 );
buf ( n45187 , n45174 );
buf ( n45188 , n45185 );
buf ( n45189 , n45174 );
not ( n45190 , n45186 );
not ( n45191 , n45187 );
or ( n45192 , n45190 , n45191 );
or ( n45193 , n45188 , n45189 );
nand ( n45194 , n45192 , n45193 );
buf ( n45195 , n45194 );
buf ( n45196 , n45146 );
not ( n45197 , n45196 );
buf ( n45198 , n44182 );
nand ( n45199 , n45197 , n45198 );
buf ( n45200 , n45199 );
buf ( n45201 , n45200 );
buf ( n45202 , n44188 );
not ( n45203 , n45202 );
buf ( n45204 , n44164 );
nand ( n45205 , n45203 , n45204 );
buf ( n45206 , n45205 );
buf ( n45207 , n45206 );
buf ( n45208 , n45206 );
buf ( n45209 , n45200 );
not ( n45210 , n45201 );
not ( n45211 , n45207 );
or ( n45212 , n45210 , n45211 );
or ( n45213 , n45208 , n45209 );
nand ( n45214 , n45212 , n45213 );
buf ( n45215 , n45214 );
buf ( n45216 , n43872 );
buf ( n45217 , n43879 );
nand ( n45218 , n45216 , n45217 );
buf ( n45219 , n45218 );
buf ( n45220 , n45219 );
buf ( n45221 , n44081 );
buf ( n45222 , n44098 );
and ( n45223 , n45221 , n45222 );
buf ( n45224 , n45223 );
and ( n45225 , n45224 , n44093 );
nor ( n45226 , n45225 , n43847 );
buf ( n45227 , n45226 );
buf ( n45228 , n44086 );
or ( n45229 , n45227 , n45228 );
buf ( n45230 , n43854 );
nand ( n45231 , n45229 , n45230 );
buf ( n45232 , n45231 );
buf ( n45233 , n45232 );
buf ( n45234 , n45219 );
buf ( n45235 , n45232 );
not ( n45236 , n45220 );
not ( n45237 , n45233 );
or ( n45238 , n45236 , n45237 );
or ( n45239 , n45234 , n45235 );
nand ( n45240 , n45238 , n45239 );
buf ( n45241 , n45240 );
buf ( n45242 , n44182 );
not ( n45243 , n45242 );
buf ( n45244 , n44135 );
nor ( n45245 , n45243 , n45244 );
buf ( n45246 , n45245 );
buf ( n45247 , n45246 );
buf ( n45248 , n45021 );
buf ( n45249 , n45246 );
buf ( n45250 , n45021 );
not ( n45251 , n45247 );
not ( n45252 , n45248 );
or ( n45253 , n45251 , n45252 );
or ( n45254 , n45249 , n45250 );
nand ( n45255 , n45253 , n45254 );
buf ( n45256 , n45255 );
buf ( n45257 , n45226 );
buf ( n45258 , n43827 );
buf ( n45259 , n43854 );
and ( n45260 , n45258 , n45259 );
buf ( n45261 , n45260 );
buf ( n45262 , n45261 );
buf ( n45263 , n45261 );
buf ( n45264 , n45226 );
not ( n45265 , n45257 );
not ( n45266 , n45262 );
or ( n45267 , n45265 , n45266 );
or ( n45268 , n45263 , n45264 );
nand ( n45269 , n45267 , n45268 );
buf ( n45270 , n45269 );
buf ( n45271 , n44093 );
buf ( n45272 , n43844 );
nand ( n45273 , n45271 , n45272 );
buf ( n45274 , n45273 );
buf ( n45275 , n45274 );
buf ( n45276 , n45224 );
not ( n45277 , n45276 );
buf ( n45278 , n43838 );
nand ( n45279 , n45277 , n45278 );
buf ( n45280 , n45279 );
buf ( n45281 , n45280 );
buf ( n45282 , n45274 );
buf ( n45283 , n45280 );
not ( n45284 , n45275 );
not ( n45285 , n45281 );
or ( n45286 , n45284 , n45285 );
or ( n45287 , n45282 , n45283 );
nand ( n45288 , n45286 , n45287 );
buf ( n45289 , n45288 );
buf ( n45290 , n43946 );
buf ( n45291 , n43953 );
nand ( n45292 , n45290 , n45291 );
buf ( n45293 , n45292 );
buf ( n45294 , n45293 );
buf ( n45295 , n44061 );
buf ( n45296 , n44071 );
and ( n45297 , n45295 , n45296 );
buf ( n45298 , n43930 );
nor ( n45299 , n45297 , n45298 );
buf ( n45300 , n45299 );
buf ( n45301 , n45300 );
buf ( n45302 , n43896 );
not ( n45303 , n45302 );
buf ( n45304 , n45303 );
buf ( n45305 , n45304 );
or ( n45306 , n45301 , n45305 );
buf ( n45307 , n43937 );
nand ( n45308 , n45306 , n45307 );
buf ( n45309 , n45308 );
buf ( n45310 , n45309 );
buf ( n45311 , n45293 );
buf ( n45312 , n45309 );
not ( n45313 , n45294 );
not ( n45314 , n45310 );
or ( n45315 , n45313 , n45314 );
or ( n45316 , n45311 , n45312 );
nand ( n45317 , n45315 , n45316 );
buf ( n45318 , n45317 );
buf ( n45319 , n44098 );
buf ( n45320 , n43838 );
nand ( n45321 , n45319 , n45320 );
buf ( n45322 , n45321 );
buf ( n45323 , n45322 );
buf ( n45324 , n44081 );
buf ( n45325 , n45322 );
buf ( n45326 , n44081 );
not ( n45327 , n45323 );
not ( n45328 , n45324 );
or ( n45329 , n45327 , n45328 );
or ( n45330 , n45325 , n45326 );
nand ( n45331 , n45329 , n45330 );
buf ( n45332 , n45331 );
buf ( n45333 , n45300 );
buf ( n45334 , n43896 );
buf ( n45335 , n43937 );
and ( n45336 , n45334 , n45335 );
buf ( n45337 , n45336 );
buf ( n45338 , n45337 );
buf ( n45339 , n45337 );
buf ( n45340 , n45300 );
not ( n45341 , n45333 );
not ( n45342 , n45338 );
or ( n45343 , n45341 , n45342 );
or ( n45344 , n45339 , n45340 );
nand ( n45345 , n45343 , n45344 );
buf ( n45346 , n45345 );
buf ( n45347 , n43913 );
not ( n45348 , n45347 );
buf ( n45349 , n43927 );
nand ( n45350 , n45348 , n45349 );
buf ( n45351 , n45350 );
buf ( n45352 , n45351 );
buf ( n45353 , n44068 );
not ( n45354 , n45353 );
buf ( n45355 , n45354 );
buf ( n45356 , n45355 );
not ( n45357 , n45356 );
buf ( n45358 , n44061 );
not ( n45359 , n45358 );
or ( n45360 , n45357 , n45359 );
buf ( n45361 , n43921 );
nand ( n45362 , n45360 , n45361 );
buf ( n45363 , n45362 );
buf ( n45364 , n45363 );
buf ( n45365 , n45351 );
buf ( n45366 , n45363 );
not ( n45367 , n45352 );
not ( n45368 , n45364 );
or ( n45369 , n45367 , n45368 );
or ( n45370 , n45365 , n45366 );
nand ( n45371 , n45369 , n45370 );
buf ( n45372 , n45371 );
buf ( n45373 , n45355 );
buf ( n45374 , n43921 );
nand ( n45375 , n45373 , n45374 );
buf ( n45376 , n45375 );
buf ( n45377 , n45376 );
buf ( n45378 , n44061 );
buf ( n45379 , n45376 );
buf ( n45380 , n44061 );
not ( n45381 , n45377 );
not ( n45382 , n45378 );
or ( n45383 , n45381 , n45382 );
or ( n45384 , n45379 , n45380 );
nand ( n45385 , n45383 , n45384 );
buf ( n45386 , n45385 );
xor ( n45387 , n43959 , n43960 );
xor ( n45388 , n45387 , n44057 );
buf ( n45389 , n45388 );
xor ( n45390 , n43962 , n43971 );
xor ( n45391 , n45390 , n44052 );
buf ( n45392 , n45391 );
xor ( n45393 , n43976 , n43977 );
xor ( n45394 , n45393 , n44047 );
buf ( n45395 , n45394 );
xor ( n45396 , n43979 , n43980 );
xor ( n45397 , n45396 , n44042 );
buf ( n45398 , n45397 );
xor ( n45399 , n43986 , n43987 );
xor ( n45400 , n45399 , n44037 );
buf ( n45401 , n45400 );
buf ( n45402 , n44033 );
not ( n45403 , n45402 );
buf ( n45404 , n44027 );
nor ( n45405 , n45403 , n45404 );
buf ( n45406 , n45405 );
buf ( n45407 , n45406 );
buf ( n45408 , n44018 );
buf ( n45409 , n44018 );
buf ( n45410 , n45406 );
not ( n45411 , n45407 );
not ( n45412 , n45408 );
or ( n45413 , n45411 , n45412 );
or ( n45414 , n45409 , n45410 );
nand ( n45415 , n45413 , n45414 );
buf ( n45416 , n45415 );
buf ( n45417 , n44007 );
not ( n45418 , n45417 );
buf ( n45419 , n45418 );
buf ( n45420 , n45419 );
buf ( n45421 , n43995 );
buf ( n45422 , n43999 );
and ( n45423 , n45421 , n45422 );
buf ( n45424 , n44015 );
nor ( n45425 , n45423 , n45424 );
buf ( n45426 , n45425 );
buf ( n45427 , n45426 );
not ( n45428 , n45427 );
buf ( n45429 , n45428 );
buf ( n45430 , n45429 );
buf ( n45431 , n45419 );
buf ( n45432 , n45429 );
not ( n45433 , n45420 );
not ( n45434 , n45430 );
or ( n45435 , n45433 , n45434 );
or ( n45436 , n45431 , n45432 );
nand ( n45437 , n45435 , n45436 );
buf ( n45438 , n45437 );
buf ( n45439 , n44229 );
not ( n45440 , n45439 );
buf ( n45441 , n45440 );
buf ( n45442 , n44924 );
buf ( n45443 , n44929 );
nand ( n45444 , n45442 , n45443 );
buf ( n45445 , n45444 );
buf ( n45446 , n43648 );
buf ( n45447 , n43698 );
nand ( n45448 , n45446 , n45447 );
buf ( n45449 , n45448 );
buf ( n45450 , n43758 );
buf ( n45451 , n43662 );
nand ( n45452 , n45450 , n45451 );
buf ( n45453 , n45452 );
buf ( n45454 , n44480 );
buf ( n45455 , n44630 );
nand ( n45456 , n45454 , n45455 );
buf ( n45457 , n45456 );
buf ( n45458 , n44258 );
buf ( n45459 , n44335 );
nand ( n45460 , n45458 , n45459 );
buf ( n45461 , n45460 );
buf ( n45462 , n43789 );
buf ( n45463 , n44226 );
not ( n45464 , n45462 );
nand ( n45465 , n45464 , n45463 );
buf ( n45466 , n45465 );
buf ( n45467 , n45003 );
buf ( n45468 , n44601 );
nand ( n45469 , n45467 , n45468 );
buf ( n45470 , n45469 );
buf ( n45471 , n44510 );
buf ( n45472 , n44571 );
not ( n45473 , n45472 );
buf ( n45474 , n45473 );
buf ( n45475 , n45474 );
nand ( n45476 , n45471 , n45475 );
buf ( n45477 , n45476 );
buf ( n45478 , n44534 );
buf ( n45479 , n44561 );
not ( n45480 , n45478 );
nand ( n45481 , n45480 , n45479 );
buf ( n45482 , n45481 );
buf ( n45483 , n44385 );
buf ( n45484 , n44404 );
nand ( n45485 , n45483 , n45484 );
buf ( n45486 , n45485 );
buf ( n45487 , n43807 );
buf ( n45488 , n44233 );
nand ( n45489 , n45487 , n45488 );
buf ( n45490 , n45489 );
buf ( n45491 , n44472 );
buf ( n45492 , n44618 );
nand ( n45493 , n45491 , n45492 );
buf ( n45494 , n45493 );
buf ( n45495 , n44368 );
buf ( n45496 , n45054 );
nand ( n45497 , n45495 , n45496 );
buf ( n45498 , n45497 );
buf ( n45499 , n43618 );
buf ( n45500 , n43744 );
nand ( n45501 , n45499 , n45500 );
buf ( n45502 , n45501 );
buf ( n45503 , n43715 );
buf ( n45504 , n43722 );
nand ( n45505 , n45503 , n45504 );
buf ( n45506 , n45505 );
buf ( n45507 , n44266 );
buf ( n45508 , n44322 );
nand ( n45509 , n45507 , n45508 );
buf ( n45510 , n45509 );
buf ( n45511 , n44459 );
buf ( n45512 , n44607 );
not ( n45513 , n45511 );
nand ( n45514 , n45513 , n45512 );
buf ( n45515 , n45514 );
buf ( n45516 , n43763 );
buf ( n45517 , n43674 );
nand ( n45518 , n45516 , n45517 );
buf ( n45519 , n45518 );
buf ( n45520 , n44352 );
buf ( n45521 , n44429 );
nand ( n45522 , n45520 , n45521 );
buf ( n45523 , n45522 );
buf ( n45524 , n43629 );
buf ( n45525 , n43733 );
nand ( n45526 , n45524 , n45525 );
buf ( n45527 , n45526 );
buf ( n45528 , n43470 );
buf ( n45529 , n44785 );
nand ( n45530 , n45528 , n45529 );
buf ( n45531 , n45530 );
buf ( n45532 , n44743 );
buf ( n45533 , n44768 );
nand ( n45534 , n45532 , n45533 );
buf ( n45535 , n45534 );
buf ( n45536 , n44731 );
buf ( n45537 , n44755 );
nand ( n45538 , n45536 , n45537 );
buf ( n45539 , n45538 );
buf ( n45540 , n44688 );
buf ( n45541 , n44711 );
nand ( n45542 , n45540 , n45541 );
buf ( n45543 , n45542 );
buf ( n45544 , n43559 );
buf ( n45545 , n44701 );
not ( n45546 , n45544 );
nand ( n45547 , n45546 , n45545 );
buf ( n45548 , n45547 );
buf ( n45549 , n43819 );
buf ( n45550 , n44244 );
nand ( n45551 , n45549 , n45550 );
buf ( n45552 , n45551 );
buf ( n45553 , n44899 );
buf ( n45554 , n44695 );
nand ( n45555 , n45553 , n45554 );
buf ( n45556 , n45555 );
buf ( n45557 , n43506 );
buf ( n45558 , n44678 );
nand ( n45559 , n45557 , n45558 );
buf ( n45560 , n45559 );
buf ( n45561 , n43496 );
buf ( n45562 , n44668 );
nand ( n45563 , n45561 , n45562 );
buf ( n45564 , n45563 );
buf ( n45565 , n43530 );
buf ( n45566 , n44657 );
not ( n45567 , n45565 );
nand ( n45568 , n45567 , n45566 );
buf ( n45569 , n45568 );
buf ( n45570 , n44992 );
buf ( n45571 , n44650 );
nand ( n45572 , n45570 , n45571 );
buf ( n45573 , n45572 );
buf ( n45574 , n44275 );
buf ( n45575 , n44312 );
nand ( n45576 , n45574 , n45575 );
buf ( n45577 , n45576 );
buf ( n45578 , n43460 );
buf ( n45579 , n43464 );
buf ( n45580 , n43460 );
buf ( n45581 , n43464 );
not ( n45582 , n45578 );
not ( n45583 , n45579 );
and ( n45584 , n45582 , n45583 );
and ( n45585 , n45580 , n45581 );
nor ( n45586 , n45584 , n45585 );
buf ( n45587 , n45586 );
buf ( n45588 , n44824 );
buf ( n45589 , n45535 );
xnor ( n45590 , n45588 , n45589 );
buf ( n45591 , n45590 );
buf ( n45592 , n44883 );
buf ( n45593 , n43662 );
not ( n45594 , n45592 );
nand ( n45595 , n45594 , n45593 );
buf ( n45596 , n45595 );
buf ( n45597 , n45050 );
buf ( n45598 , n45498 );
xnor ( n45599 , n45597 , n45598 );
buf ( n45600 , n45599 );
buf ( n45601 , n44864 );
buf ( n45602 , n45445 );
xnor ( n45603 , n45601 , n45602 );
buf ( n45604 , n45603 );
buf ( n45605 , n44896 );
buf ( n45606 , n45449 );
xnor ( n45607 , n45605 , n45606 );
buf ( n45608 , n45607 );
buf ( n45609 , n44989 );
buf ( n45610 , n45457 );
xnor ( n45611 , n45609 , n45610 );
buf ( n45612 , n45611 );
buf ( n45613 , n45118 );
buf ( n45614 , n45461 );
xnor ( n45615 , n45613 , n45614 );
buf ( n45616 , n45615 );
buf ( n45617 , n45181 );
buf ( n45618 , n45466 );
xnor ( n45619 , n45617 , n45618 );
buf ( n45620 , n45619 );
buf ( n45621 , n44973 );
buf ( n45622 , n45470 );
xnor ( n45623 , n45621 , n45622 );
buf ( n45624 , n45623 );
buf ( n45625 , n45071 );
buf ( n45626 , n45477 );
xnor ( n45627 , n45625 , n45626 );
buf ( n45628 , n45627 );
buf ( n45629 , n45082 );
buf ( n45630 , n45482 );
xnor ( n45631 , n45629 , n45630 );
buf ( n45632 , n45631 );
buf ( n45633 , n45037 );
buf ( n45634 , n45486 );
xnor ( n45635 , n45633 , n45634 );
buf ( n45636 , n45635 );
not ( n45637 , n43800 );
not ( n45638 , n45174 );
or ( n45639 , n45637 , n45638 );
nand ( n45640 , n45639 , n45441 );
buf ( n45641 , n45640 );
buf ( n45642 , n45490 );
xnor ( n45643 , n45641 , n45642 );
buf ( n45644 , n45643 );
buf ( n45645 , n44982 );
buf ( n45646 , n45494 );
xnor ( n45647 , n45645 , n45646 );
buf ( n45648 , n45647 );
buf ( n45649 , n44880 );
buf ( n45650 , n45502 );
xnor ( n45651 , n45649 , n45650 );
buf ( n45652 , n45651 );
buf ( n45653 , n44935 );
buf ( n45654 , n45506 );
xnor ( n45655 , n45653 , n45654 );
buf ( n45656 , n45655 );
buf ( n45657 , n45111 );
buf ( n45658 , n45510 );
xnor ( n45659 , n45657 , n45658 );
buf ( n45660 , n45659 );
buf ( n45661 , n45011 );
buf ( n45662 , n45515 );
xnor ( n45663 , n45661 , n45662 );
buf ( n45664 , n45663 );
buf ( n45665 , n45596 );
buf ( n45666 , n45519 );
xnor ( n45667 , n45665 , n45666 );
buf ( n45668 , n45667 );
buf ( n45669 , n45060 );
buf ( n45670 , n45523 );
xnor ( n45671 , n45669 , n45670 );
buf ( n45672 , n45671 );
buf ( n45673 , n44873 );
buf ( n45674 , n45527 );
xnor ( n45675 , n45673 , n45674 );
buf ( n45676 , n45675 );
buf ( n45677 , n44778 );
buf ( n45678 , n45531 );
xnor ( n45679 , n45677 , n45678 );
buf ( n45680 , n45679 );
buf ( n45681 , n44726 );
buf ( n45682 , n45539 );
xnor ( n45683 , n45681 , n45682 );
buf ( n45684 , n45683 );
buf ( n45685 , n44946 );
buf ( n45686 , n45543 );
xnor ( n45687 , n45685 , n45686 );
buf ( n45688 , n45687 );
buf ( n45689 , n44921 );
buf ( n45690 , n45548 );
xnor ( n45691 , n45689 , n45690 );
buf ( n45692 , n45691 );
not ( n45693 , n43807 );
not ( n45694 , n45640 );
or ( n45695 , n45693 , n45694 );
nand ( n45696 , n45695 , n44233 );
buf ( n45697 , n45696 );
buf ( n45698 , n45552 );
xnor ( n45699 , n45697 , n45698 );
buf ( n45700 , n45699 );
buf ( n45701 , n44914 );
buf ( n45702 , n45556 );
xnor ( n45703 , n45701 , n45702 );
buf ( n45704 , n45703 );
buf ( n45705 , n44965 );
buf ( n45706 , n45560 );
xnor ( n45707 , n45705 , n45706 );
buf ( n45708 , n45707 );
buf ( n45709 , n44958 );
buf ( n45710 , n45564 );
xnor ( n45711 , n45709 , n45710 );
buf ( n45712 , n45711 );
buf ( n45713 , n45000 );
buf ( n45714 , n45569 );
xnor ( n45715 , n45713 , n45714 );
buf ( n45716 , n45715 );
buf ( n45717 , n44639 );
buf ( n45718 , n45573 );
xnor ( n45719 , n45717 , n45718 );
buf ( n45720 , n45719 );
buf ( n45721 , n45126 );
buf ( n45722 , n45577 );
xnor ( n45723 , n45721 , n45722 );
buf ( n45724 , n45723 );
not ( n45725 , n37536 );
not ( n45726 , n45725 );
not ( n45727 , n37533 );
not ( n45728 , n45727 );
or ( n45729 , n45726 , n45728 );
nand ( n45730 , n45729 , n37537 );
buf ( n45731 , n45730 );
not ( n45732 , n45731 );
or ( n45733 , n37469 , n37468 );
nand ( n45734 , n45733 , n37470 );
not ( n45735 , n45734 );
not ( n45736 , n45735 );
or ( n45737 , n45732 , n45736 );
not ( n45738 , n45731 );
nand ( n45739 , n45734 , n45738 );
nand ( n45740 , n45737 , n45739 );
buf ( n45741 , n42065 );
and ( n45742 , n45740 , n45741 );
not ( n45743 , n37665 );
and ( n45744 , n37651 , n45743 );
not ( n45745 , n37651 );
and ( n45746 , n45745 , n37665 );
nor ( n45747 , n45744 , n45746 );
not ( n45748 , n45747 );
not ( n45749 , n45748 );
buf ( n45750 , n45730 );
not ( n45751 , n45750 );
not ( n45752 , n30633 );
not ( n45753 , n45752 );
or ( n45754 , n45751 , n45753 );
not ( n45755 , n45730 );
nand ( n45756 , n45755 , n30633 );
nand ( n45757 , n45754 , n45756 );
not ( n45758 , n45757 );
or ( n45759 , n45749 , n45758 );
not ( n45760 , n45730 );
nand ( n45761 , n45760 , n45743 );
not ( n45762 , n45761 );
nand ( n45763 , n45730 , n37665 );
nand ( n45764 , n45763 , n45747 );
nor ( n45765 , n45762 , n45764 );
buf ( n45766 , n45765 );
not ( n45767 , n1212 );
or ( n45768 , n45730 , n45767 );
nand ( n45769 , n45767 , n45730 );
nand ( n45770 , n45768 , n45769 );
nand ( n45771 , n45766 , n45770 );
nand ( n45772 , n45759 , n45771 );
xor ( n45773 , n45742 , n45772 );
not ( n45774 , n42065 );
nand ( n45775 , n45743 , n45774 );
not ( n45776 , n37651 );
not ( n45777 , n45776 );
and ( n45778 , n45775 , n45777 );
and ( n45779 , n37665 , n45741 );
nor ( n45780 , n45778 , n45779 , n45755 );
xnor ( n45781 , n45774 , n45730 );
not ( n45782 , n45781 );
not ( n45783 , n45765 );
or ( n45784 , n45782 , n45783 );
not ( n45785 , n45747 );
nand ( n45786 , n45785 , n45770 );
nand ( n45787 , n45784 , n45786 );
and ( n45788 , n45780 , n45787 );
xor ( n45789 , n45773 , n45788 );
xor ( n45790 , n45742 , n45772 );
and ( n45791 , n45790 , n45788 );
and ( n45792 , n45742 , n45772 );
or ( n45793 , n45791 , n45792 );
not ( n45794 , n45741 );
xnor ( n45795 , n37463 , n37577 );
not ( n45796 , n45795 );
and ( n45797 , n45794 , n45796 );
not ( n45798 , n45794 );
not ( n45799 , n45796 );
and ( n45800 , n45798 , n45799 );
nor ( n45801 , n45797 , n45800 );
not ( n45802 , n45801 );
and ( n45803 , n45795 , n45734 );
not ( n45804 , n45795 );
and ( n45805 , n45804 , n45735 );
nor ( n45806 , n45803 , n45805 );
not ( n45807 , n45731 );
not ( n45808 , n45734 );
or ( n45809 , n45807 , n45808 );
nand ( n45810 , n45735 , n45738 );
nand ( n45811 , n45809 , n45810 );
and ( n45812 , n45806 , n45811 );
not ( n45813 , n45812 );
or ( n45814 , n45802 , n45813 );
not ( n45815 , n45811 );
not ( n45816 , n45767 );
not ( n45817 , n45816 );
not ( n45818 , n45796 );
or ( n45819 , n45817 , n45818 );
buf ( n45820 , n45795 );
nand ( n45821 , n45820 , n45767 );
nand ( n45822 , n45819 , n45821 );
nand ( n45823 , n45815 , n45822 );
nand ( n45824 , n45814 , n45823 );
not ( n45825 , n45735 );
or ( n45826 , n45825 , n45741 );
buf ( n45827 , n45750 );
nand ( n45828 , n45826 , n45827 );
not ( n45829 , n45794 );
nand ( n45830 , n45825 , n45829 );
and ( n45831 , n45799 , n45828 , n45830 );
not ( n45832 , n45747 );
not ( n45833 , n45832 );
not ( n45834 , n30610 );
and ( n45835 , n45834 , n45827 );
not ( n45836 , n45834 );
not ( n45837 , n45750 );
and ( n45838 , n45836 , n45837 );
or ( n45839 , n45835 , n45838 );
not ( n45840 , n45839 );
or ( n45841 , n45833 , n45840 );
buf ( n45842 , n45766 );
nand ( n45843 , n45757 , n45842 );
nand ( n45844 , n45841 , n45843 );
xor ( n45845 , n45831 , n45844 );
xor ( n45846 , n45824 , n45845 );
not ( n45847 , n44004 );
not ( n45848 , n42038 );
and ( n45849 , n45848 , n45777 );
not ( n45850 , n45848 );
and ( n45851 , n45850 , n45776 );
or ( n45852 , n45849 , n45851 );
not ( n45853 , n45852 );
or ( n45854 , n45847 , n45853 );
not ( n45855 , n45777 );
not ( n45856 , n42050 );
not ( n45857 , n45856 );
or ( n45858 , n45855 , n45857 );
nand ( n45859 , n42050 , n45776 );
nand ( n45860 , n45858 , n45859 );
not ( n45861 , n44004 );
nand ( n45862 , n45861 , n37651 );
not ( n45863 , n45862 );
nand ( n45864 , n45860 , n45863 );
nand ( n45865 , n45854 , n45864 );
xor ( n45866 , n45846 , n45865 );
xor ( n45867 , n45824 , n45845 );
and ( n45868 , n45867 , n45865 );
and ( n45869 , n45824 , n45845 );
or ( n45870 , n45868 , n45869 );
not ( n45871 , n45822 );
not ( n45872 , n45812 );
or ( n45873 , n45871 , n45872 );
not ( n45874 , n45796 );
not ( n45875 , n30633 );
or ( n45876 , n45874 , n45875 );
not ( n45877 , n45796 );
not ( n45878 , n30633 );
nand ( n45879 , n45877 , n45878 );
nand ( n45880 , n45876 , n45879 );
nand ( n45881 , n45880 , n45740 );
nand ( n45882 , n45873 , n45881 );
nand ( n45883 , n36116 , n36118 );
nand ( n45884 , n35981 , n37556 );
not ( n45885 , n45884 );
and ( n45886 , n45883 , n45885 );
not ( n45887 , n45883 );
and ( n45888 , n45887 , n45884 );
nor ( n45889 , n45886 , n45888 );
not ( n45890 , n45889 );
and ( n45891 , n45796 , n45890 );
not ( n45892 , n45796 );
and ( n45893 , n45892 , n45889 );
nor ( n45894 , n45891 , n45893 );
not ( n45895 , n45894 );
not ( n45896 , n45895 );
and ( n45897 , n45896 , n45741 );
xor ( n45898 , n45882 , n45897 );
not ( n45899 , n45748 );
not ( n45900 , n45827 );
not ( n45901 , n45856 );
or ( n45902 , n45900 , n45901 );
nand ( n45903 , n42050 , n45837 );
nand ( n45904 , n45902 , n45903 );
not ( n45905 , n45904 );
or ( n45906 , n45899 , n45905 );
buf ( n45907 , n45766 );
nand ( n45908 , n45839 , n45907 );
nand ( n45909 , n45906 , n45908 );
xor ( n45910 , n45898 , n45909 );
xor ( n45911 , n45882 , n45897 );
and ( n45912 , n45911 , n45909 );
and ( n45913 , n45882 , n45897 );
or ( n45914 , n45912 , n45913 );
and ( n45915 , n45831 , n45844 );
xor ( n45916 , n45915 , n45910 );
not ( n45917 , n44004 );
not ( n45918 , n45777 );
not ( n45919 , n42006 );
not ( n45920 , n45919 );
or ( n45921 , n45918 , n45920 );
not ( n45922 , n45919 );
nand ( n45923 , n45922 , n45776 );
nand ( n45924 , n45921 , n45923 );
not ( n45925 , n45924 );
or ( n45926 , n45917 , n45925 );
nand ( n45927 , n45852 , n45863 );
nand ( n45928 , n45926 , n45927 );
xor ( n45929 , n45916 , n45928 );
xor ( n45930 , n45915 , n45910 );
and ( n45931 , n45930 , n45928 );
and ( n45932 , n45915 , n45910 );
or ( n45933 , n45931 , n45932 );
not ( n45934 , n45829 );
not ( n45935 , n37595 );
and ( n45936 , n35930 , n35980 );
nand ( n45937 , n45936 , n37643 , n37469 );
not ( n45938 , n36115 );
not ( n45939 , n37642 );
or ( n45940 , n45938 , n45939 );
nand ( n45941 , n45940 , n35928 );
nand ( n45942 , n45937 , n45941 , n36118 );
not ( n45943 , n45942 );
not ( n45944 , n45943 );
or ( n45945 , n45935 , n45944 );
nand ( n45946 , n37594 , n45942 );
nand ( n45947 , n45945 , n45946 );
not ( n45948 , n45947 );
not ( n45949 , n45948 );
or ( n45950 , n45934 , n45949 );
buf ( n45951 , n45947 );
nand ( n45952 , n45951 , n45794 );
nand ( n45953 , n45950 , n45952 );
not ( n45954 , n45953 );
not ( n45955 , n45894 );
not ( n45956 , n45947 );
not ( n45957 , n45890 );
or ( n45958 , n45956 , n45957 );
or ( n45959 , n45947 , n45890 );
nand ( n45960 , n45958 , n45959 );
nand ( n45961 , n45955 , n45960 );
not ( n45962 , n45961 );
not ( n45963 , n45962 );
or ( n45964 , n45954 , n45963 );
not ( n45965 , n45816 );
not ( n45966 , n45948 );
or ( n45967 , n45965 , n45966 );
not ( n45968 , n45948 );
nand ( n45969 , n45968 , n45767 );
nand ( n45970 , n45967 , n45969 );
nand ( n45971 , n45896 , n45970 );
nand ( n45972 , n45964 , n45971 );
not ( n45973 , n45880 );
not ( n45974 , n45812 );
or ( n45975 , n45973 , n45974 );
not ( n45976 , n30610 );
not ( n45977 , n45796 );
or ( n45978 , n45976 , n45977 );
nand ( n45979 , n45834 , n45820 );
nand ( n45980 , n45978 , n45979 );
nand ( n45981 , n45980 , n45740 );
nand ( n45982 , n45975 , n45981 );
not ( n45983 , n45951 );
buf ( n45984 , n45889 );
nor ( n45985 , n45984 , n45829 );
or ( n45986 , n45985 , n45796 );
nand ( n45987 , n45984 , n45741 );
nand ( n45988 , n45986 , n45987 );
nor ( n45989 , n45983 , n45988 );
xor ( n45990 , n45982 , n45989 );
xor ( n45991 , n45972 , n45990 );
not ( n45992 , n45904 );
not ( n45993 , n45907 );
or ( n45994 , n45992 , n45993 );
not ( n45995 , n45837 );
not ( n45996 , n42038 );
and ( n45997 , n45995 , n45996 );
buf ( n45998 , n42038 );
and ( n45999 , n45998 , n45837 );
nor ( n46000 , n45997 , n45999 );
or ( n46001 , n46000 , n45747 );
nand ( n46002 , n45994 , n46001 );
xor ( n46003 , n45991 , n46002 );
xor ( n46004 , n45972 , n45990 );
and ( n46005 , n46004 , n46002 );
and ( n46006 , n45972 , n45990 );
or ( n46007 , n46005 , n46006 );
not ( n46008 , n44004 );
not ( n46009 , n45776 );
not ( n46010 , n30465 );
or ( n46011 , n46009 , n46010 );
not ( n46012 , n30465 );
nand ( n46013 , n46012 , n45777 );
nand ( n46014 , n46011 , n46013 );
not ( n46015 , n46014 );
or ( n46016 , n46008 , n46015 );
nand ( n46017 , n45924 , n45863 );
nand ( n46018 , n46016 , n46017 );
xor ( n46019 , n45914 , n46018 );
xor ( n46020 , n46019 , n46003 );
xor ( n46021 , n45914 , n46018 );
and ( n46022 , n46021 , n46003 );
and ( n46023 , n45914 , n46018 );
or ( n46024 , n46022 , n46023 );
not ( n46025 , n45740 );
and ( n46026 , n42049 , n45796 );
not ( n46027 , n42049 );
and ( n46028 , n46027 , n45820 );
or ( n46029 , n46026 , n46028 );
not ( n46030 , n46029 );
or ( n46031 , n46025 , n46030 );
nand ( n46032 , n45812 , n45980 );
nand ( n46033 , n46031 , n46032 );
not ( n46034 , n45970 );
not ( n46035 , n45962 );
or ( n46036 , n46034 , n46035 );
not ( n46037 , n45878 );
and ( n46038 , n45948 , n46037 );
not ( n46039 , n45948 );
and ( n46040 , n46039 , n45878 );
or ( n46041 , n46038 , n46040 );
nand ( n46042 , n46041 , n45896 );
nand ( n46043 , n46036 , n46042 );
xor ( n46044 , n46033 , n46043 );
xor ( n46045 , n36996 , n37641 );
xnor ( n46046 , n45968 , n46045 );
nor ( n46047 , n46046 , n45794 );
xor ( n46048 , n46044 , n46047 );
xor ( n46049 , n46033 , n46043 );
and ( n46050 , n46049 , n46047 );
and ( n46051 , n46033 , n46043 );
or ( n46052 , n46050 , n46051 );
and ( n46053 , n45982 , n45989 );
not ( n46054 , n45832 );
and ( n46055 , n45919 , n45827 );
not ( n46056 , n45919 );
and ( n46057 , n46056 , n45837 );
or ( n46058 , n46055 , n46057 );
not ( n46059 , n46058 );
or ( n46060 , n46054 , n46059 );
not ( n46061 , n46000 );
nand ( n46062 , n46061 , n45907 );
nand ( n46063 , n46060 , n46062 );
xor ( n46064 , n46053 , n46063 );
xor ( n46065 , n46064 , n46007 );
xor ( n46066 , n46053 , n46063 );
and ( n46067 , n46066 , n46007 );
and ( n46068 , n46053 , n46063 );
or ( n46069 , n46067 , n46068 );
not ( n46070 , n44004 );
buf ( n46071 , n45776 );
not ( n46072 , n46071 );
not ( n46073 , n46072 );
not ( n46074 , n30379 );
not ( n46075 , n46074 );
or ( n46076 , n46073 , n46075 );
nand ( n46077 , n30379 , n46071 );
nand ( n46078 , n46076 , n46077 );
not ( n46079 , n46078 );
or ( n46080 , n46070 , n46079 );
nand ( n46081 , n46014 , n45863 );
nand ( n46082 , n46080 , n46081 );
xor ( n46083 , n46048 , n46082 );
xor ( n46084 , n46083 , n46065 );
xor ( n46085 , n46048 , n46082 );
and ( n46086 , n46085 , n46065 );
and ( n46087 , n46048 , n46082 );
or ( n46088 , n46086 , n46087 );
buf ( n46089 , n37063 );
not ( n46090 , n46089 );
buf ( n46091 , n46045 );
nand ( n46092 , n46091 , n45829 );
not ( n46093 , n45951 );
and ( n46094 , n46092 , n46093 );
nor ( n46095 , n46091 , n45829 );
nor ( n46096 , n46094 , n46095 );
nor ( n46097 , n46090 , n46096 );
not ( n46098 , n45740 );
and ( n46099 , n42037 , n45796 );
not ( n46100 , n42037 );
and ( n46101 , n46100 , n45799 );
or ( n46102 , n46099 , n46101 );
not ( n46103 , n46102 );
or ( n46104 , n46098 , n46103 );
nand ( n46105 , n45812 , n46029 );
nand ( n46106 , n46104 , n46105 );
not ( n46107 , n46041 );
not ( n46108 , n45962 );
or ( n46109 , n46107 , n46108 );
not ( n46110 , n46093 );
buf ( n46111 , n30610 );
not ( n46112 , n46111 );
or ( n46113 , n46110 , n46112 );
not ( n46114 , n46111 );
nand ( n46115 , n45951 , n46114 );
nand ( n46116 , n46113 , n46115 );
nand ( n46117 , n46116 , n45896 );
nand ( n46118 , n46109 , n46117 );
xor ( n46119 , n46106 , n46118 );
xor ( n46120 , n46097 , n46119 );
xor ( n46121 , n46120 , n46052 );
xor ( n46122 , n46097 , n46119 );
and ( n46123 , n46122 , n46052 );
and ( n46124 , n46097 , n46119 );
or ( n46125 , n46123 , n46124 );
not ( n46126 , n45832 );
not ( n46127 , n45837 );
not ( n46128 , n30465 );
or ( n46129 , n46127 , n46128 );
nand ( n46130 , n46012 , n45827 );
nand ( n46131 , n46129 , n46130 );
not ( n46132 , n46131 );
or ( n46133 , n46126 , n46132 );
nand ( n46134 , n46058 , n45907 );
nand ( n46135 , n46133 , n46134 );
and ( n46136 , n45741 , n46089 );
not ( n46137 , n45741 );
not ( n46138 , n46089 );
and ( n46139 , n46137 , n46138 );
nor ( n46140 , n46136 , n46139 );
not ( n46141 , n46140 );
or ( n46142 , n46091 , n37063 );
nand ( n46143 , n46091 , n37063 );
and ( n46144 , n46142 , n46143 , n46046 );
not ( n46145 , n46144 );
or ( n46146 , n46141 , n46145 );
not ( n46147 , n45816 );
not ( n46148 , n37063 );
not ( n46149 , n46148 );
or ( n46150 , n46147 , n46149 );
nand ( n46151 , n46089 , n45767 );
nand ( n46152 , n46150 , n46151 );
not ( n46153 , n46046 );
nand ( n46154 , n46152 , n46153 );
nand ( n46155 , n46146 , n46154 );
xor ( n46156 , n46135 , n46155 );
xor ( n46157 , n46156 , n46121 );
xor ( n46158 , n46135 , n46155 );
and ( n46159 , n46158 , n46121 );
and ( n46160 , n46135 , n46155 );
or ( n46161 , n46159 , n46160 );
not ( n46162 , n44004 );
not ( n46163 , n30577 );
and ( n46164 , n46071 , n46163 );
not ( n46165 , n46071 );
and ( n46166 , n46165 , n41948 );
nor ( n46167 , n46164 , n46166 );
not ( n46168 , n46167 );
or ( n46169 , n46162 , n46168 );
nand ( n46170 , n46078 , n45863 );
nand ( n46171 , n46169 , n46170 );
xor ( n46172 , n46171 , n46069 );
xor ( n46173 , n46172 , n46157 );
xor ( n46174 , n46171 , n46069 );
and ( n46175 , n46174 , n46157 );
and ( n46176 , n46171 , n46069 );
or ( n46177 , n46175 , n46176 );
not ( n46178 , n46116 );
not ( n46179 , n45962 );
or ( n46180 , n46178 , n46179 );
not ( n46181 , n42050 );
not ( n46182 , n46093 );
or ( n46183 , n46181 , n46182 );
nand ( n46184 , n45968 , n45856 );
nand ( n46185 , n46183 , n46184 );
nand ( n46186 , n46185 , n45896 );
nand ( n46187 , n46180 , n46186 );
buf ( n46188 , n45740 );
not ( n46189 , n46188 );
and ( n46190 , n42006 , n45796 );
not ( n46191 , n42006 );
and ( n46192 , n46191 , n45799 );
or ( n46193 , n46190 , n46192 );
not ( n46194 , n46193 );
or ( n46195 , n46189 , n46194 );
nand ( n46196 , n46102 , n45812 );
nand ( n46197 , n46195 , n46196 );
xor ( n46198 , n46187 , n46197 );
not ( n46199 , n37051 );
not ( n46200 , n46199 );
not ( n46201 , n46089 );
and ( n46202 , n46200 , n46201 );
not ( n46203 , n46148 );
and ( n46204 , n46199 , n46203 );
nor ( n46205 , n46202 , n46204 );
nor ( n46206 , n46205 , n45794 );
xor ( n46207 , n46198 , n46206 );
xor ( n46208 , n46187 , n46197 );
and ( n46209 , n46208 , n46206 );
and ( n46210 , n46187 , n46197 );
or ( n46211 , n46209 , n46210 );
and ( n46212 , n46106 , n46118 );
not ( n46213 , n46152 );
not ( n46214 , n46144 );
or ( n46215 , n46213 , n46214 );
not ( n46216 , n46037 );
not ( n46217 , n46138 );
or ( n46218 , n46216 , n46217 );
nand ( n46219 , n46089 , n45878 );
nand ( n46220 , n46218 , n46219 );
nand ( n46221 , n46220 , n46153 );
nand ( n46222 , n46215 , n46221 );
xor ( n46223 , n46212 , n46222 );
not ( n46224 , n45832 );
not ( n46225 , n45750 );
not ( n46226 , n46074 );
or ( n46227 , n46225 , n46226 );
nand ( n46228 , n30379 , n45837 );
nand ( n46229 , n46227 , n46228 );
not ( n46230 , n46229 );
or ( n46231 , n46224 , n46230 );
nand ( n46232 , n46131 , n45907 );
nand ( n46233 , n46231 , n46232 );
xor ( n46234 , n46223 , n46233 );
xor ( n46235 , n46212 , n46222 );
and ( n46236 , n46235 , n46233 );
and ( n46237 , n46212 , n46222 );
or ( n46238 , n46236 , n46237 );
not ( n46239 , n44004 );
and ( n46240 , n41945 , n46071 );
not ( n46241 , n41945 );
and ( n46242 , n46241 , n46072 );
or ( n46243 , n46240 , n46242 );
not ( n46244 , n46243 );
or ( n46245 , n46239 , n46244 );
nand ( n46246 , n45863 , n46167 );
nand ( n46247 , n46245 , n46246 );
xor ( n46248 , n46207 , n46247 );
xor ( n46249 , n46248 , n46125 );
xor ( n46250 , n46207 , n46247 );
and ( n46251 , n46250 , n46125 );
and ( n46252 , n46207 , n46247 );
or ( n46253 , n46251 , n46252 );
xor ( n46254 , n46234 , n46161 );
xor ( n46255 , n46254 , n46249 );
xor ( n46256 , n46234 , n46161 );
and ( n46257 , n46256 , n46249 );
and ( n46258 , n46234 , n46161 );
or ( n46259 , n46257 , n46258 );
not ( n46260 , n46188 );
and ( n46261 , n30465 , n45796 );
not ( n46262 , n30465 );
and ( n46263 , n46262 , n45799 );
or ( n46264 , n46261 , n46263 );
not ( n46265 , n46264 );
or ( n46266 , n46260 , n46265 );
buf ( n46267 , n45812 );
nand ( n46268 , n46193 , n46267 );
nand ( n46269 , n46266 , n46268 );
not ( n46270 , n46220 );
not ( n46271 , n46144 );
or ( n46272 , n46270 , n46271 );
not ( n46273 , n46114 );
not ( n46274 , n46273 );
not ( n46275 , n46148 );
or ( n46276 , n46274 , n46275 );
nand ( n46277 , n46089 , n46114 );
nand ( n46278 , n46276 , n46277 );
nand ( n46279 , n46153 , n46278 );
nand ( n46280 , n46272 , n46279 );
xor ( n46281 , n46269 , n46280 );
not ( n46282 , n46185 );
not ( n46283 , n45962 );
or ( n46284 , n46282 , n46283 );
not ( n46285 , n45951 );
not ( n46286 , n45848 );
or ( n46287 , n46285 , n46286 );
nand ( n46288 , n45998 , n46093 );
nand ( n46289 , n46287 , n46288 );
nand ( n46290 , n45896 , n46289 );
nand ( n46291 , n46284 , n46290 );
nand ( n46292 , n46199 , n45794 );
nand ( n46293 , n46089 , n46292 );
not ( n46294 , n36229 );
nor ( n46295 , n46294 , n37573 );
and ( n46296 , n37393 , n46295 );
not ( n46297 , n37393 );
and ( n46298 , n46297 , n37575 );
nor ( n46299 , n46296 , n46298 );
not ( n46300 , n46299 );
not ( n46301 , n46300 );
nand ( n46302 , n37051 , n45741 );
and ( n46303 , n46293 , n46301 , n46302 );
xor ( n46304 , n46291 , n46303 );
xor ( n46305 , n46281 , n46304 );
xor ( n46306 , n46269 , n46280 );
and ( n46307 , n46306 , n46304 );
and ( n46308 , n46269 , n46280 );
or ( n46309 , n46307 , n46308 );
and ( n46310 , n45741 , n46301 );
not ( n46311 , n45741 );
buf ( n46312 , n46300 );
and ( n46313 , n46311 , n46312 );
nor ( n46314 , n46310 , n46313 );
not ( n46315 , n46314 );
not ( n46316 , n37051 );
not ( n46317 , n46300 );
or ( n46318 , n46316 , n46317 );
nand ( n46319 , n46299 , n46199 );
nand ( n46320 , n46318 , n46319 );
and ( n46321 , n46205 , n46320 );
not ( n46322 , n46321 );
or ( n46323 , n46315 , n46322 );
not ( n46324 , n45816 );
not ( n46325 , n46301 );
not ( n46326 , n46325 );
or ( n46327 , n46324 , n46326 );
nand ( n46328 , n46301 , n45767 );
nand ( n46329 , n46327 , n46328 );
and ( n46330 , n46199 , n46089 );
not ( n46331 , n46199 );
and ( n46332 , n46331 , n46138 );
nor ( n46333 , n46330 , n46332 );
not ( n46334 , n46333 );
nand ( n46335 , n46329 , n46334 );
nand ( n46336 , n46323 , n46335 );
xor ( n46337 , n46336 , n46211 );
not ( n46338 , n45832 );
not ( n46339 , n45750 );
not ( n46340 , n46163 );
or ( n46341 , n46339 , n46340 );
nand ( n46342 , n41948 , n45837 );
nand ( n46343 , n46341 , n46342 );
not ( n46344 , n46343 );
or ( n46345 , n46338 , n46344 );
nand ( n46346 , n46229 , n45907 );
nand ( n46347 , n46345 , n46346 );
xor ( n46348 , n46337 , n46347 );
xor ( n46349 , n46336 , n46211 );
and ( n46350 , n46349 , n46347 );
and ( n46351 , n46336 , n46211 );
or ( n46352 , n46350 , n46351 );
not ( n46353 , n45863 );
not ( n46354 , n46243 );
or ( n46355 , n46353 , n46354 );
or ( n46356 , n30351 , n46071 );
nand ( n46357 , n30351 , n46071 );
nand ( n46358 , n46356 , n46357 );
nand ( n46359 , n44004 , n46358 );
nand ( n46360 , n46355 , n46359 );
xor ( n46361 , n46360 , n46305 );
xor ( n46362 , n46361 , n46238 );
xor ( n46363 , n46360 , n46305 );
and ( n46364 , n46363 , n46238 );
and ( n46365 , n46360 , n46305 );
or ( n46366 , n46364 , n46365 );
xor ( n46367 , n46348 , n46253 );
xor ( n46368 , n46367 , n46362 );
xor ( n46369 , n46348 , n46253 );
and ( n46370 , n46369 , n46362 );
and ( n46371 , n46348 , n46253 );
or ( n46372 , n46370 , n46371 );
not ( n46373 , n45896 );
and ( n46374 , n45951 , n45919 );
not ( n46375 , n45951 );
and ( n46376 , n46375 , n45922 );
or ( n46377 , n46374 , n46376 );
not ( n46378 , n46377 );
or ( n46379 , n46373 , n46378 );
nand ( n46380 , n45962 , n46289 );
nand ( n46381 , n46379 , n46380 );
not ( n46382 , n46278 );
not ( n46383 , n46144 );
or ( n46384 , n46382 , n46383 );
not ( n46385 , n42050 );
not ( n46386 , n46148 );
or ( n46387 , n46385 , n46386 );
buf ( n46388 , n45856 );
nand ( n46389 , n46203 , n46388 );
nand ( n46390 , n46387 , n46389 );
nand ( n46391 , n46390 , n46153 );
nand ( n46392 , n46384 , n46391 );
xor ( n46393 , n46381 , n46392 );
and ( n46394 , n46291 , n46303 );
xor ( n46395 , n46393 , n46394 );
xor ( n46396 , n46381 , n46392 );
and ( n46397 , n46396 , n46394 );
and ( n46398 , n46381 , n46392 );
or ( n46399 , n46397 , n46398 );
not ( n46400 , n46329 );
nand ( n46401 , n46089 , n37051 );
not ( n46402 , n46401 );
not ( n46403 , n46089 );
nand ( n46404 , n46403 , n46199 );
not ( n46405 , n46404 );
or ( n46406 , n46402 , n46405 );
nand ( n46407 , n46406 , n46320 );
not ( n46408 , n46407 );
not ( n46409 , n46408 );
or ( n46410 , n46400 , n46409 );
not ( n46411 , n46037 );
buf ( n46412 , n46299 );
not ( n46413 , n46412 );
not ( n46414 , n46413 );
or ( n46415 , n46411 , n46414 );
not ( n46416 , n46312 );
nand ( n46417 , n46416 , n45878 );
nand ( n46418 , n46415 , n46417 );
nand ( n46419 , n46418 , n46334 );
nand ( n46420 , n46410 , n46419 );
not ( n46421 , n46188 );
buf ( n46422 , n45796 );
and ( n46423 , n30379 , n46422 );
not ( n46424 , n30379 );
not ( n46425 , n46422 );
and ( n46426 , n46424 , n46425 );
or ( n46427 , n46423 , n46426 );
not ( n46428 , n46427 );
or ( n46429 , n46421 , n46428 );
nand ( n46430 , n46264 , n46267 );
nand ( n46431 , n46429 , n46430 );
xor ( n46432 , n46420 , n46431 );
nor ( n46433 , n36993 , n36187 );
and ( n46434 , n46433 , n37581 );
not ( n46435 , n46433 );
and ( n46436 , n46435 , n37582 );
nor ( n46437 , n46434 , n46436 );
xnor ( n46438 , n46301 , n46437 );
buf ( n46439 , n46438 );
buf ( n46440 , n45741 );
not ( n46441 , n46440 );
nor ( n46442 , n46439 , n46441 );
xor ( n46443 , n46432 , n46442 );
xor ( n46444 , n46420 , n46431 );
and ( n46445 , n46444 , n46442 );
and ( n46446 , n46420 , n46431 );
or ( n46447 , n46445 , n46446 );
buf ( n46448 , n45766 );
not ( n46449 , n46448 );
not ( n46450 , n46343 );
or ( n46451 , n46449 , n46450 );
not ( n46452 , n45750 );
not ( n46453 , n41945 );
not ( n46454 , n46453 );
or ( n46455 , n46452 , n46454 );
nand ( n46456 , n41946 , n45837 );
nand ( n46457 , n46455 , n46456 );
nand ( n46458 , n45832 , n46457 );
nand ( n46459 , n46451 , n46458 );
xor ( n46460 , n46459 , n46309 );
xor ( n46461 , n46460 , n46395 );
xor ( n46462 , n46459 , n46309 );
and ( n46463 , n46462 , n46395 );
and ( n46464 , n46459 , n46309 );
or ( n46465 , n46463 , n46464 );
xor ( n46466 , n46352 , n46443 );
not ( n46467 , n44004 );
and ( n46468 , n30259 , n46071 );
not ( n46469 , n30259 );
and ( n46470 , n46469 , n46072 );
or ( n46471 , n46468 , n46470 );
not ( n46472 , n46471 );
or ( n46473 , n46467 , n46472 );
buf ( n46474 , n45863 );
nand ( n46475 , n46358 , n46474 );
nand ( n46476 , n46473 , n46475 );
xor ( n46477 , n46466 , n46476 );
xor ( n46478 , n46352 , n46443 );
and ( n46479 , n46478 , n46476 );
and ( n46480 , n46352 , n46443 );
or ( n46481 , n46479 , n46480 );
xor ( n46482 , n46366 , n46461 );
xor ( n46483 , n46482 , n46477 );
xor ( n46484 , n46366 , n46461 );
and ( n46485 , n46484 , n46477 );
and ( n46486 , n46366 , n46461 );
or ( n46487 , n46485 , n46486 );
not ( n46488 , n46418 );
not ( n46489 , n46408 );
or ( n46490 , n46488 , n46489 );
not ( n46491 , n46273 );
not ( n46492 , n46325 );
or ( n46493 , n46491 , n46492 );
nand ( n46494 , n46301 , n46114 );
nand ( n46495 , n46493 , n46494 );
nand ( n46496 , n46495 , n46334 );
nand ( n46497 , n46490 , n46496 );
buf ( n46498 , n46437 );
not ( n46499 , n46498 );
nand ( n46500 , n46499 , n45794 );
not ( n46501 , n46500 );
not ( n46502 , n45741 );
not ( n46503 , n46498 );
or ( n46504 , n46502 , n46503 );
buf ( n46505 , n46300 );
nand ( n46506 , n46504 , n46505 );
not ( n46507 , n46506 );
or ( n46508 , n46501 , n46507 );
not ( n46509 , n37006 );
buf ( n46510 , n46509 );
not ( n46511 , n46510 );
nand ( n46512 , n46508 , n46511 );
not ( n46513 , n46512 );
xor ( n46514 , n46497 , n46513 );
not ( n46515 , n46188 );
not ( n46516 , n46422 );
not ( n46517 , n41948 );
or ( n46518 , n46516 , n46517 );
nand ( n46519 , n46163 , n46425 );
nand ( n46520 , n46518 , n46519 );
not ( n46521 , n46520 );
or ( n46522 , n46515 , n46521 );
nand ( n46523 , n46427 , n46267 );
nand ( n46524 , n46522 , n46523 );
xor ( n46525 , n46514 , n46524 );
xor ( n46526 , n46497 , n46513 );
and ( n46527 , n46526 , n46524 );
and ( n46528 , n46497 , n46513 );
or ( n46529 , n46527 , n46528 );
not ( n46530 , n45896 );
not ( n46531 , n45951 );
not ( n46532 , n46012 );
or ( n46533 , n46531 , n46532 );
nand ( n46534 , n30465 , n46093 );
nand ( n46535 , n46533 , n46534 );
not ( n46536 , n46535 );
or ( n46537 , n46530 , n46536 );
nand ( n46538 , n46377 , n45962 );
nand ( n46539 , n46537 , n46538 );
not ( n46540 , n46390 );
not ( n46541 , n46144 );
or ( n46542 , n46540 , n46541 );
not ( n46543 , n46148 );
not ( n46544 , n45998 );
or ( n46545 , n46543 , n46544 );
not ( n46546 , n45998 );
nand ( n46547 , n46089 , n46546 );
nand ( n46548 , n46545 , n46547 );
nand ( n46549 , n46153 , n46548 );
nand ( n46550 , n46542 , n46549 );
xor ( n46551 , n46539 , n46550 );
xor ( n46552 , n46551 , n46399 );
not ( n46553 , n45832 );
buf ( n46554 , n45750 );
not ( n46555 , n46554 );
not ( n46556 , n30351 );
not ( n46557 , n46556 );
or ( n46558 , n46555 , n46557 );
buf ( n46559 , n45837 );
nand ( n46560 , n30351 , n46559 );
nand ( n46561 , n46558 , n46560 );
not ( n46562 , n46561 );
or ( n46563 , n46553 , n46562 );
buf ( n46564 , n46448 );
nand ( n46565 , n46564 , n46457 );
nand ( n46566 , n46563 , n46565 );
xor ( n46567 , n46552 , n46566 );
xor ( n46568 , n46551 , n46399 );
and ( n46569 , n46568 , n46566 );
and ( n46570 , n46551 , n46399 );
or ( n46571 , n46569 , n46570 );
not ( n46572 , n46440 );
not ( n46573 , n37006 );
not ( n46574 , n46573 );
or ( n46575 , n46572 , n46574 );
not ( n46576 , n46573 );
nand ( n46577 , n46576 , n46441 );
nand ( n46578 , n46575 , n46577 );
not ( n46579 , n46578 );
nand ( n46580 , n46573 , n46499 );
not ( n46581 , n46509 );
nand ( n46582 , n46581 , n46498 );
nand ( n46583 , n46580 , n46438 , n46582 );
not ( n46584 , n46583 );
not ( n46585 , n46584 );
or ( n46586 , n46579 , n46585 );
not ( n46587 , n45816 );
not ( n46588 , n46510 );
or ( n46589 , n46587 , n46588 );
nand ( n46590 , n46576 , n45767 );
nand ( n46591 , n46589 , n46590 );
not ( n46592 , n46439 );
nand ( n46593 , n46591 , n46592 );
nand ( n46594 , n46586 , n46593 );
xor ( n46595 , n46594 , n46447 );
xor ( n46596 , n46595 , n46525 );
xor ( n46597 , n46594 , n46447 );
and ( n46598 , n46597 , n46525 );
and ( n46599 , n46594 , n46447 );
or ( n46600 , n46598 , n46599 );
not ( n46601 , n44004 );
not ( n46602 , n46601 );
not ( n46603 , n46602 );
not ( n46604 , n46072 );
not ( n46605 , n41938 );
or ( n46606 , n46604 , n46605 );
not ( n46607 , n41933 );
not ( n46608 , n46607 );
nand ( n46609 , n46608 , n46071 );
nand ( n46610 , n46606 , n46609 );
not ( n46611 , n46610 );
or ( n46612 , n46603 , n46611 );
nand ( n46613 , n46471 , n46474 );
nand ( n46614 , n46612 , n46613 );
xor ( n46615 , n46614 , n46567 );
xor ( n46616 , n46615 , n46465 );
xor ( n46617 , n46614 , n46567 );
and ( n46618 , n46617 , n46465 );
and ( n46619 , n46614 , n46567 );
or ( n46620 , n46618 , n46619 );
xor ( n46621 , n46596 , n46481 );
xor ( n46622 , n46621 , n46616 );
xor ( n46623 , n46596 , n46481 );
and ( n46624 , n46623 , n46616 );
and ( n46625 , n46596 , n46481 );
or ( n46626 , n46624 , n46625 );
not ( n46627 , n46548 );
not ( n46628 , n46144 );
or ( n46629 , n46627 , n46628 );
not ( n46630 , n45922 );
not ( n46631 , n46138 );
or ( n46632 , n46630 , n46631 );
nand ( n46633 , n46203 , n45919 );
nand ( n46634 , n46632 , n46633 );
nand ( n46635 , n46634 , n46153 );
nand ( n46636 , n46629 , n46635 );
not ( n46637 , n46495 );
not ( n46638 , n46321 );
or ( n46639 , n46637 , n46638 );
not ( n46640 , n42050 );
buf ( n46641 , n46300 );
not ( n46642 , n46641 );
or ( n46643 , n46640 , n46642 );
nand ( n46644 , n46301 , n46388 );
nand ( n46645 , n46643 , n46644 );
nand ( n46646 , n46645 , n46334 );
nand ( n46647 , n46639 , n46646 );
xor ( n46648 , n46636 , n46647 );
not ( n46649 , n45896 );
buf ( n46650 , n45951 );
not ( n46651 , n46650 );
not ( n46652 , n46074 );
or ( n46653 , n46651 , n46652 );
not ( n46654 , n45951 );
nand ( n46655 , n30379 , n46654 );
nand ( n46656 , n46653 , n46655 );
not ( n46657 , n46656 );
or ( n46658 , n46649 , n46657 );
nand ( n46659 , n46535 , n45962 );
nand ( n46660 , n46658 , n46659 );
xor ( n46661 , n46648 , n46660 );
xor ( n46662 , n46636 , n46647 );
and ( n46663 , n46662 , n46660 );
and ( n46664 , n46636 , n46647 );
or ( n46665 , n46663 , n46664 );
not ( n46666 , n37006 );
and ( n46667 , n37039 , n46666 );
not ( n46668 , n37039 );
and ( n46669 , n46668 , n46581 );
nor ( n46670 , n46667 , n46669 );
nor ( n46671 , n46670 , n45794 );
and ( n46672 , n46550 , n46539 );
xor ( n46673 , n46671 , n46672 );
not ( n46674 , n46267 );
not ( n46675 , n46520 );
or ( n46676 , n46674 , n46675 );
not ( n46677 , n46425 );
not ( n46678 , n46453 );
or ( n46679 , n46677 , n46678 );
nand ( n46680 , n41945 , n46422 );
nand ( n46681 , n46679 , n46680 );
nand ( n46682 , n46681 , n46188 );
nand ( n46683 , n46676 , n46682 );
xor ( n46684 , n46673 , n46683 );
xor ( n46685 , n46671 , n46672 );
and ( n46686 , n46685 , n46683 );
and ( n46687 , n46671 , n46672 );
or ( n46688 , n46686 , n46687 );
not ( n46689 , n46591 );
and ( n46690 , n46580 , n46582 , n46438 );
not ( n46691 , n46690 );
or ( n46692 , n46689 , n46691 );
not ( n46693 , n46037 );
not ( n46694 , n46666 );
or ( n46695 , n46693 , n46694 );
nand ( n46696 , n46576 , n45878 );
nand ( n46697 , n46695 , n46696 );
nand ( n46698 , n46697 , n46592 );
nand ( n46699 , n46692 , n46698 );
xor ( n46700 , n46699 , n46661 );
not ( n46701 , n45832 );
and ( n46702 , n30259 , n46559 );
not ( n46703 , n30259 );
and ( n46704 , n46703 , n46554 );
or ( n46705 , n46702 , n46704 );
not ( n46706 , n46705 );
or ( n46707 , n46701 , n46706 );
nand ( n46708 , n46561 , n46448 );
nand ( n46709 , n46707 , n46708 );
xor ( n46710 , n46700 , n46709 );
xor ( n46711 , n46699 , n46661 );
and ( n46712 , n46711 , n46709 );
and ( n46713 , n46699 , n46661 );
or ( n46714 , n46712 , n46713 );
not ( n46715 , n46474 );
not ( n46716 , n46610 );
or ( n46717 , n46715 , n46716 );
not ( n46718 , n46072 );
not ( n46719 , n41861 );
not ( n46720 , n46719 );
or ( n46721 , n46718 , n46720 );
nand ( n46722 , n41861 , n46071 );
nand ( n46723 , n46721 , n46722 );
nand ( n46724 , n46723 , n46602 );
nand ( n46725 , n46717 , n46724 );
xor ( n46726 , n46529 , n46725 );
xor ( n46727 , n46726 , n46684 );
xor ( n46728 , n46529 , n46725 );
and ( n46729 , n46728 , n46684 );
and ( n46730 , n46529 , n46725 );
or ( n46731 , n46729 , n46730 );
xor ( n46732 , n46571 , n46710 );
xor ( n46733 , n46732 , n46600 );
xor ( n46734 , n46571 , n46710 );
and ( n46735 , n46734 , n46600 );
and ( n46736 , n46571 , n46710 );
or ( n46737 , n46735 , n46736 );
xor ( n46738 , n46620 , n46727 );
xor ( n46739 , n46738 , n46733 );
xor ( n46740 , n46620 , n46727 );
and ( n46741 , n46740 , n46733 );
and ( n46742 , n46620 , n46727 );
or ( n46743 , n46741 , n46742 );
or ( n46744 , n36993 , n36187 );
and ( n46745 , n46744 , n37667 );
not ( n46746 , n37032 );
not ( n46747 , n36205 );
or ( n46748 , n46746 , n46747 );
nand ( n46749 , n46748 , n37033 );
nor ( n46750 , n46745 , n46749 );
nand ( n46751 , n36193 , n36209 );
nor ( n46752 , n46750 , n46751 );
not ( n46753 , n46752 );
nand ( n46754 , n46744 , n37667 );
not ( n46755 , n46749 );
nand ( n46756 , n46754 , n46755 , n46751 );
nand ( n46757 , n46753 , n46756 );
not ( n46758 , n46757 );
not ( n46759 , n37039 );
nand ( n46760 , n46759 , n45794 );
not ( n46761 , n45741 );
not ( n46762 , n37039 );
or ( n46763 , n46761 , n46762 );
nand ( n46764 , n46763 , n46666 );
nand ( n46765 , n46760 , n46764 );
and ( n46766 , n46758 , n46765 );
not ( n46767 , n45896 );
not ( n46768 , n46650 );
not ( n46769 , n46163 );
or ( n46770 , n46768 , n46769 );
nand ( n46771 , n41948 , n46654 );
nand ( n46772 , n46770 , n46771 );
not ( n46773 , n46772 );
or ( n46774 , n46767 , n46773 );
not ( n46775 , n45962 );
not ( n46776 , n46775 );
nand ( n46777 , n46656 , n46776 );
nand ( n46778 , n46774 , n46777 );
xor ( n46779 , n46766 , n46778 );
not ( n46780 , n46634 );
not ( n46781 , n46144 );
or ( n46782 , n46780 , n46781 );
not ( n46783 , n41954 );
not ( n46784 , n46138 );
or ( n46785 , n46783 , n46784 );
nand ( n46786 , n46089 , n46012 );
nand ( n46787 , n46785 , n46786 );
nand ( n46788 , n46787 , n46153 );
nand ( n46789 , n46782 , n46788 );
not ( n46790 , n46645 );
not ( n46791 , n46321 );
or ( n46792 , n46790 , n46791 );
not ( n46793 , n45998 );
not ( n46794 , n46641 );
or ( n46795 , n46793 , n46794 );
nand ( n46796 , n46412 , n46546 );
nand ( n46797 , n46795 , n46796 );
nand ( n46798 , n46797 , n46334 );
nand ( n46799 , n46792 , n46798 );
xor ( n46800 , n46789 , n46799 );
xor ( n46801 , n46779 , n46800 );
xor ( n46802 , n46766 , n46778 );
and ( n46803 , n46802 , n46800 );
and ( n46804 , n46766 , n46778 );
or ( n46805 , n46803 , n46804 );
not ( n46806 , n46188 );
not ( n46807 , n46425 );
not ( n46808 , n46556 );
or ( n46809 , n46807 , n46808 );
nand ( n46810 , n30351 , n46422 );
nand ( n46811 , n46809 , n46810 );
not ( n46812 , n46811 );
or ( n46813 , n46806 , n46812 );
nand ( n46814 , n46681 , n46267 );
nand ( n46815 , n46813 , n46814 );
not ( n46816 , n46697 );
not ( n46817 , n46690 );
or ( n46818 , n46816 , n46817 );
not ( n46819 , n46273 );
not ( n46820 , n46666 );
not ( n46821 , n46820 );
not ( n46822 , n46821 );
or ( n46823 , n46819 , n46822 );
not ( n46824 , n46273 );
nand ( n46825 , n46576 , n46824 );
nand ( n46826 , n46823 , n46825 );
nand ( n46827 , n46826 , n46592 );
nand ( n46828 , n46818 , n46827 );
xor ( n46829 , n46815 , n46828 );
and ( n46830 , n45741 , n46757 );
not ( n46831 , n45741 );
not ( n46832 , n46752 );
nand ( n46833 , n46832 , n46756 );
not ( n46834 , n46833 );
buf ( n46835 , n46834 );
and ( n46836 , n46831 , n46835 );
or ( n46837 , n46830 , n46836 );
not ( n46838 , n46837 );
not ( n46839 , n46833 );
not ( n46840 , n37039 );
or ( n46841 , n46839 , n46840 );
nand ( n46842 , n46834 , n46759 );
nand ( n46843 , n46841 , n46842 );
buf ( n46844 , n46670 );
nand ( n46845 , n46843 , n46844 );
not ( n46846 , n46845 );
not ( n46847 , n46846 );
or ( n46848 , n46838 , n46847 );
not ( n46849 , n45816 );
not ( n46850 , n46833 );
or ( n46851 , n46849 , n46850 );
nand ( n46852 , n46758 , n45767 );
nand ( n46853 , n46851 , n46852 );
not ( n46854 , n46844 );
nand ( n46855 , n46853 , n46854 );
nand ( n46856 , n46848 , n46855 );
xor ( n46857 , n46829 , n46856 );
xor ( n46858 , n46815 , n46828 );
and ( n46859 , n46858 , n46856 );
and ( n46860 , n46815 , n46828 );
or ( n46861 , n46859 , n46860 );
xor ( n46862 , n46665 , n46688 );
xor ( n46863 , n46862 , n46801 );
xor ( n46864 , n46665 , n46688 );
and ( n46865 , n46864 , n46801 );
and ( n46866 , n46665 , n46688 );
or ( n46867 , n46865 , n46866 );
not ( n46868 , n45832 );
not ( n46869 , n46554 );
not ( n46870 , n46607 );
or ( n46871 , n46869 , n46870 );
nand ( n46872 , n41933 , n46559 );
nand ( n46873 , n46871 , n46872 );
not ( n46874 , n46873 );
or ( n46875 , n46868 , n46874 );
nand ( n46876 , n46705 , n46448 );
nand ( n46877 , n46875 , n46876 );
not ( n46878 , n46602 );
not ( n46879 , n46072 );
not ( n46880 , n41800 );
not ( n46881 , n46880 );
or ( n46882 , n46879 , n46881 );
nand ( n46883 , n41800 , n46071 );
nand ( n46884 , n46882 , n46883 );
not ( n46885 , n46884 );
or ( n46886 , n46878 , n46885 );
nand ( n46887 , n46723 , n46474 );
nand ( n46888 , n46886 , n46887 );
xor ( n46889 , n46877 , n46888 );
xor ( n46890 , n46889 , n46857 );
xor ( n46891 , n46877 , n46888 );
and ( n46892 , n46891 , n46857 );
and ( n46893 , n46877 , n46888 );
or ( n46894 , n46892 , n46893 );
xor ( n46895 , n46714 , n46863 );
xor ( n46896 , n46895 , n46731 );
xor ( n46897 , n46714 , n46863 );
and ( n46898 , n46897 , n46731 );
and ( n46899 , n46714 , n46863 );
or ( n46900 , n46898 , n46899 );
xor ( n46901 , n46737 , n46890 );
xor ( n46902 , n46901 , n46896 );
xor ( n46903 , n46737 , n46890 );
and ( n46904 , n46903 , n46896 );
and ( n46905 , n46737 , n46890 );
or ( n46906 , n46904 , n46905 );
not ( n46907 , n46797 );
not ( n46908 , n46321 );
or ( n46909 , n46907 , n46908 );
not ( n46910 , n45922 );
not ( n46911 , n46413 );
or ( n46912 , n46910 , n46911 );
nand ( n46913 , n46412 , n45919 );
nand ( n46914 , n46912 , n46913 );
nand ( n46915 , n46914 , n46334 );
nand ( n46916 , n46909 , n46915 );
not ( n46917 , n46153 );
not ( n46918 , n46089 );
not ( n46919 , n46074 );
or ( n46920 , n46918 , n46919 );
nand ( n46921 , n30379 , n46138 );
nand ( n46922 , n46920 , n46921 );
not ( n46923 , n46922 );
or ( n46924 , n46917 , n46923 );
buf ( n46925 , n46144 );
nand ( n46926 , n46925 , n46787 );
nand ( n46927 , n46924 , n46926 );
xor ( n46928 , n46916 , n46927 );
not ( n46929 , n45896 );
not ( n46930 , n46650 );
not ( n46931 , n46453 );
or ( n46932 , n46930 , n46931 );
nand ( n46933 , n41945 , n46654 );
nand ( n46934 , n46932 , n46933 );
not ( n46935 , n46934 );
or ( n46936 , n46929 , n46935 );
nand ( n46937 , n46772 , n46776 );
nand ( n46938 , n46936 , n46937 );
xor ( n46939 , n46928 , n46938 );
xor ( n46940 , n46916 , n46927 );
and ( n46941 , n46940 , n46938 );
and ( n46942 , n46916 , n46927 );
or ( n46943 , n46941 , n46942 );
and ( n46944 , n46789 , n46799 );
not ( n46945 , n46826 );
not ( n46946 , n46690 );
or ( n46947 , n46945 , n46946 );
not ( n46948 , n42050 );
not ( n46949 , n46510 );
or ( n46950 , n46948 , n46949 );
nand ( n46951 , n46820 , n45856 );
nand ( n46952 , n46950 , n46951 );
nand ( n46953 , n46952 , n46592 );
nand ( n46954 , n46947 , n46953 );
xor ( n46955 , n46944 , n46954 );
not ( n46956 , n46037 );
not ( n46957 , n46833 );
or ( n46958 , n46956 , n46957 );
nand ( n46959 , n46758 , n45878 );
nand ( n46960 , n46958 , n46959 );
not ( n46961 , n46960 );
not ( n46962 , n46854 );
or ( n46963 , n46961 , n46962 );
nand ( n46964 , n46846 , n46853 );
nand ( n46965 , n46963 , n46964 );
xor ( n46966 , n46955 , n46965 );
xor ( n46967 , n46944 , n46954 );
and ( n46968 , n46967 , n46965 );
and ( n46969 , n46944 , n46954 );
or ( n46970 , n46968 , n46969 );
not ( n46971 , n37013 );
and ( n46972 , n46757 , n46971 );
not ( n46973 , n46757 );
and ( n46974 , n46973 , n37013 );
nor ( n46975 , n46972 , n46974 );
and ( n46976 , n46975 , n46440 );
not ( n46977 , n46188 );
and ( n46978 , n30259 , n46422 );
not ( n46979 , n30259 );
and ( n46980 , n46979 , n46425 );
or ( n46981 , n46978 , n46980 );
not ( n46982 , n46981 );
or ( n46983 , n46977 , n46982 );
nand ( n46984 , n46811 , n46267 );
nand ( n46985 , n46983 , n46984 );
xor ( n46986 , n46976 , n46985 );
xor ( n46987 , n46986 , n46805 );
xor ( n46988 , n46976 , n46985 );
and ( n46989 , n46988 , n46805 );
and ( n46990 , n46976 , n46985 );
or ( n46991 , n46989 , n46990 );
not ( n46992 , n45832 );
not ( n46993 , n46554 );
not ( n46994 , n41861 );
not ( n46995 , n46994 );
or ( n46996 , n46993 , n46995 );
nand ( n46997 , n41861 , n46559 );
nand ( n46998 , n46996 , n46997 );
not ( n46999 , n46998 );
or ( n47000 , n46992 , n46999 );
nand ( n47001 , n46873 , n46448 );
nand ( n47002 , n47000 , n47001 );
xor ( n47003 , n46939 , n47002 );
xor ( n47004 , n47003 , n46861 );
xor ( n47005 , n46939 , n47002 );
and ( n47006 , n47005 , n46861 );
and ( n47007 , n46939 , n47002 );
or ( n47008 , n47006 , n47007 );
buf ( n47009 , n44004 );
not ( n47010 , n47009 );
xor ( n47011 , n46072 , n30964 );
not ( n47012 , n47011 );
or ( n47013 , n47010 , n47012 );
nand ( n47014 , n46884 , n46474 );
nand ( n47015 , n47013 , n47014 );
xor ( n47016 , n46966 , n47015 );
xor ( n47017 , n47016 , n46867 );
xor ( n47018 , n46966 , n47015 );
and ( n47019 , n47018 , n46867 );
and ( n47020 , n46966 , n47015 );
or ( n47021 , n47019 , n47020 );
xor ( n47022 , n46987 , n46894 );
xor ( n47023 , n47022 , n47004 );
xor ( n47024 , n46987 , n46894 );
and ( n47025 , n47024 , n47004 );
and ( n47026 , n46987 , n46894 );
or ( n47027 , n47025 , n47026 );
xor ( n47028 , n46900 , n47017 );
xor ( n47029 , n47028 , n47023 );
xor ( n47030 , n46900 , n47017 );
and ( n47031 , n47030 , n47023 );
and ( n47032 , n46900 , n47017 );
or ( n47033 , n47031 , n47032 );
not ( n47034 , n45896 );
not ( n47035 , n46650 );
not ( n47036 , n46556 );
or ( n47037 , n47035 , n47036 );
nand ( n47038 , n30351 , n46654 );
nand ( n47039 , n47037 , n47038 );
not ( n47040 , n47039 );
or ( n47041 , n47034 , n47040 );
nand ( n47042 , n46934 , n46776 );
nand ( n47043 , n47041 , n47042 );
not ( n47044 , n46952 );
not ( n47045 , n46584 );
or ( n47046 , n47044 , n47045 );
buf ( n47047 , n45998 );
xnor ( n47048 , n47047 , n46510 );
nand ( n47049 , n47048 , n46592 );
nand ( n47050 , n47046 , n47049 );
xor ( n47051 , n47043 , n47050 );
not ( n47052 , n46960 );
not ( n47053 , n46846 );
or ( n47054 , n47052 , n47053 );
not ( n47055 , n46273 );
not ( n47056 , n46757 );
or ( n47057 , n47055 , n47056 );
nand ( n47058 , n46835 , n46824 );
nand ( n47059 , n47057 , n47058 );
not ( n47060 , n46844 );
nand ( n47061 , n47059 , n47060 );
nand ( n47062 , n47054 , n47061 );
xor ( n47063 , n47051 , n47062 );
xor ( n47064 , n47043 , n47050 );
and ( n47065 , n47064 , n47062 );
and ( n47066 , n47043 , n47050 );
or ( n47067 , n47065 , n47066 );
not ( n47068 , n46153 );
not ( n47069 , n46203 );
not ( n47070 , n46163 );
or ( n47071 , n47069 , n47070 );
nand ( n47072 , n41948 , n46148 );
nand ( n47073 , n47071 , n47072 );
not ( n47074 , n47073 );
or ( n47075 , n47068 , n47074 );
nand ( n47076 , n46922 , n46925 );
nand ( n47077 , n47075 , n47076 );
not ( n47078 , n46914 );
not ( n47079 , n46408 );
or ( n47080 , n47078 , n47079 );
not ( n47081 , n41954 );
not ( n47082 , n46312 );
or ( n47083 , n47081 , n47082 );
nand ( n47084 , n46416 , n46012 );
nand ( n47085 , n47083 , n47084 );
nand ( n47086 , n47085 , n46334 );
nand ( n47087 , n47080 , n47086 );
xor ( n47088 , n47077 , n47087 );
nand ( n47089 , n46971 , n46441 );
not ( n47090 , n47089 );
not ( n47091 , n45741 );
not ( n47092 , n37013 );
or ( n47093 , n47091 , n47092 );
buf ( n47094 , n46833 );
nand ( n47095 , n47093 , n47094 );
not ( n47096 , n47095 );
or ( n47097 , n47090 , n47096 );
not ( n47098 , n37007 );
not ( n47099 , n36235 );
or ( n47100 , n47098 , n47099 );
nand ( n47101 , n47100 , n35663 );
and ( n47102 , n47101 , n37561 );
not ( n47103 , n47101 );
and ( n47104 , n47103 , n37560 );
nor ( n47105 , n47102 , n47104 );
buf ( n47106 , n47105 );
not ( n47107 , n47106 );
not ( n47108 , n47107 );
nand ( n47109 , n47097 , n47108 );
not ( n47110 , n47109 );
xor ( n47111 , n47088 , n47110 );
xor ( n47112 , n47111 , n46943 );
xor ( n47113 , n47088 , n47110 );
and ( n47114 , n47113 , n46943 );
and ( n47115 , n47088 , n47110 );
or ( n47116 , n47114 , n47115 );
not ( n47117 , n46188 );
not ( n47118 , n46425 );
not ( n47119 , n46607 );
or ( n47120 , n47118 , n47119 );
nand ( n47121 , n41939 , n46422 );
nand ( n47122 , n47120 , n47121 );
not ( n47123 , n47122 );
or ( n47124 , n47117 , n47123 );
nand ( n47125 , n46981 , n46267 );
nand ( n47126 , n47124 , n47125 );
not ( n47127 , n46440 );
not ( n47128 , n47107 );
or ( n47129 , n47127 , n47128 );
nand ( n47130 , n47108 , n46441 );
nand ( n47131 , n47129 , n47130 );
not ( n47132 , n47131 );
and ( n47133 , n47106 , n37013 );
not ( n47134 , n47106 );
and ( n47135 , n47134 , n46971 );
nor ( n47136 , n47133 , n47135 );
not ( n47137 , n46975 );
nand ( n47138 , n47136 , n47137 );
not ( n47139 , n47138 );
not ( n47140 , n47139 );
or ( n47141 , n47132 , n47140 );
not ( n47142 , n45816 );
not ( n47143 , n47107 );
or ( n47144 , n47142 , n47143 );
nand ( n47145 , n47108 , n45767 );
nand ( n47146 , n47144 , n47145 );
not ( n47147 , n47137 );
buf ( n47148 , n47147 );
nand ( n47149 , n47146 , n47148 );
nand ( n47150 , n47141 , n47149 );
xor ( n47151 , n47126 , n47150 );
not ( n47152 , n45832 );
not ( n47153 , n46554 );
not ( n47154 , n41801 );
not ( n47155 , n47154 );
or ( n47156 , n47153 , n47155 );
not ( n47157 , n41800 );
not ( n47158 , n47157 );
nand ( n47159 , n47158 , n46559 );
nand ( n47160 , n47156 , n47159 );
not ( n47161 , n47160 );
or ( n47162 , n47152 , n47161 );
nand ( n47163 , n46998 , n46448 );
nand ( n47164 , n47162 , n47163 );
xor ( n47165 , n47151 , n47164 );
xor ( n47166 , n47126 , n47150 );
and ( n47167 , n47166 , n47164 );
and ( n47168 , n47126 , n47150 );
or ( n47169 , n47167 , n47168 );
xor ( n47170 , n46970 , n47063 );
xor ( n47171 , n47170 , n47112 );
xor ( n47172 , n46970 , n47063 );
and ( n47173 , n47172 , n47112 );
and ( n47174 , n46970 , n47063 );
or ( n47175 , n47173 , n47174 );
not ( n47176 , n46602 );
not ( n47177 , n46072 );
not ( n47178 , n41692 );
not ( n47179 , n47178 );
or ( n47180 , n47177 , n47179 );
nand ( n47181 , n41692 , n46071 );
nand ( n47182 , n47180 , n47181 );
not ( n47183 , n47182 );
or ( n47184 , n47176 , n47183 );
nand ( n47185 , n47011 , n46474 );
nand ( n47186 , n47184 , n47185 );
xor ( n47187 , n46991 , n47186 );
xor ( n47188 , n47187 , n47008 );
xor ( n47189 , n46991 , n47186 );
and ( n47190 , n47189 , n47008 );
and ( n47191 , n46991 , n47186 );
or ( n47192 , n47190 , n47191 );
xor ( n47193 , n47171 , n47165 );
xor ( n47194 , n47193 , n47021 );
xor ( n47195 , n47171 , n47165 );
and ( n47196 , n47195 , n47021 );
and ( n47197 , n47171 , n47165 );
or ( n47198 , n47196 , n47197 );
xor ( n47199 , n47027 , n47188 );
xor ( n47200 , n47199 , n47194 );
xor ( n47201 , n47027 , n47188 );
and ( n47202 , n47201 , n47194 );
and ( n47203 , n47027 , n47188 );
or ( n47204 , n47202 , n47203 );
not ( n47205 , n46334 );
and ( n47206 , n30379 , n46641 );
not ( n47207 , n30379 );
and ( n47208 , n47207 , n46412 );
or ( n47209 , n47206 , n47208 );
not ( n47210 , n47209 );
or ( n47211 , n47205 , n47210 );
nand ( n47212 , n47085 , n46408 );
nand ( n47213 , n47211 , n47212 );
not ( n47214 , n46925 );
not ( n47215 , n47073 );
or ( n47216 , n47214 , n47215 );
and ( n47217 , n41945 , n46148 );
not ( n47218 , n41945 );
and ( n47219 , n47218 , n46203 );
or ( n47220 , n47217 , n47219 );
nand ( n47221 , n47220 , n46153 );
nand ( n47222 , n47216 , n47221 );
xor ( n47223 , n47213 , n47222 );
not ( n47224 , n47048 );
not ( n47225 , n46690 );
or ( n47226 , n47224 , n47225 );
buf ( n47227 , n45922 );
and ( n47228 , n47227 , n46510 );
not ( n47229 , n47227 );
and ( n47230 , n47229 , n46576 );
or ( n47231 , n47228 , n47230 );
nand ( n47232 , n47231 , n46592 );
nand ( n47233 , n47226 , n47232 );
xor ( n47234 , n47223 , n47233 );
xor ( n47235 , n47213 , n47222 );
and ( n47236 , n47235 , n47233 );
and ( n47237 , n47213 , n47222 );
or ( n47238 , n47236 , n47237 );
not ( n47239 , n47059 );
nand ( n47240 , n46843 , n46844 );
not ( n47241 , n47240 );
not ( n47242 , n47241 );
or ( n47243 , n47239 , n47242 );
not ( n47244 , n42050 );
not ( n47245 , n47094 );
or ( n47246 , n47244 , n47245 );
nand ( n47247 , n46835 , n45856 );
nand ( n47248 , n47246 , n47247 );
nand ( n47249 , n47248 , n47060 );
nand ( n47250 , n47243 , n47249 );
and ( n47251 , n47077 , n47087 );
xor ( n47252 , n47250 , n47251 );
not ( n47253 , n45896 );
not ( n47254 , n47253 );
not ( n47255 , n47254 );
not ( n47256 , n46650 );
not ( n47257 , n30259 );
not ( n47258 , n47257 );
or ( n47259 , n47256 , n47258 );
not ( n47260 , n46650 );
nand ( n47261 , n30259 , n47260 );
nand ( n47262 , n47259 , n47261 );
not ( n47263 , n47262 );
or ( n47264 , n47255 , n47263 );
nand ( n47265 , n47039 , n46776 );
nand ( n47266 , n47264 , n47265 );
xor ( n47267 , n47252 , n47266 );
xor ( n47268 , n47250 , n47251 );
and ( n47269 , n47268 , n47266 );
and ( n47270 , n47250 , n47251 );
or ( n47271 , n47269 , n47270 );
not ( n47272 , n47106 );
not ( n47273 , n36938 );
not ( n47274 , n47273 );
or ( n47275 , n47272 , n47274 );
not ( n47276 , n47106 );
nand ( n47277 , n36938 , n47276 );
nand ( n47278 , n47275 , n47277 );
and ( n47279 , n47278 , n46440 );
xor ( n47280 , n47234 , n47279 );
not ( n47281 , n46267 );
not ( n47282 , n47122 );
or ( n47283 , n47281 , n47282 );
not ( n47284 , n46425 );
not ( n47285 , n46719 );
or ( n47286 , n47284 , n47285 );
not ( n47287 , n41861 );
not ( n47288 , n47287 );
nand ( n47289 , n47288 , n46422 );
nand ( n47290 , n47286 , n47289 );
nand ( n47291 , n47290 , n46188 );
nand ( n47292 , n47283 , n47291 );
xor ( n47293 , n47280 , n47292 );
xor ( n47294 , n47234 , n47279 );
and ( n47295 , n47294 , n47292 );
and ( n47296 , n47234 , n47279 );
or ( n47297 , n47295 , n47296 );
not ( n47298 , n47146 );
buf ( n47299 , n47138 );
not ( n47300 , n47299 );
not ( n47301 , n47300 );
or ( n47302 , n47298 , n47301 );
not ( n47303 , n46037 );
not ( n47304 , n47107 );
or ( n47305 , n47303 , n47304 );
not ( n47306 , n46037 );
nand ( n47307 , n47108 , n47306 );
nand ( n47308 , n47305 , n47307 );
nand ( n47309 , n47308 , n47148 );
nand ( n47310 , n47302 , n47309 );
xor ( n47311 , n47310 , n47067 );
xor ( n47312 , n47311 , n47116 );
xor ( n47313 , n47310 , n47067 );
and ( n47314 , n47313 , n47116 );
and ( n47315 , n47310 , n47067 );
or ( n47316 , n47314 , n47315 );
not ( n47317 , n45832 );
not ( n47318 , n30964 );
and ( n47319 , n46559 , n47318 );
not ( n47320 , n46559 );
and ( n47321 , n47320 , n30964 );
nor ( n47322 , n47319 , n47321 );
not ( n47323 , n47322 );
or ( n47324 , n47317 , n47323 );
nand ( n47325 , n46448 , n47160 );
nand ( n47326 , n47324 , n47325 );
xor ( n47327 , n47267 , n47326 );
not ( n47328 , n46474 );
not ( n47329 , n47182 );
or ( n47330 , n47328 , n47329 );
not ( n47331 , n46072 );
not ( n47332 , n41683 );
not ( n47333 , n47332 );
or ( n47334 , n47331 , n47333 );
nand ( n47335 , n41683 , n46071 );
nand ( n47336 , n47334 , n47335 );
nand ( n47337 , n47336 , n46602 );
nand ( n47338 , n47330 , n47337 );
xor ( n47339 , n47327 , n47338 );
xor ( n47340 , n47267 , n47326 );
and ( n47341 , n47340 , n47338 );
and ( n47342 , n47267 , n47326 );
or ( n47343 , n47341 , n47342 );
xor ( n47344 , n47169 , n47293 );
xor ( n47345 , n47344 , n47312 );
xor ( n47346 , n47169 , n47293 );
and ( n47347 , n47346 , n47312 );
and ( n47348 , n47169 , n47293 );
or ( n47349 , n47347 , n47348 );
xor ( n47350 , n47175 , n47339 );
xor ( n47351 , n47350 , n47192 );
xor ( n47352 , n47175 , n47339 );
and ( n47353 , n47352 , n47192 );
and ( n47354 , n47175 , n47339 );
or ( n47355 , n47353 , n47354 );
xor ( n47356 , n47345 , n47198 );
xor ( n47357 , n47356 , n47351 );
xor ( n47358 , n47345 , n47198 );
and ( n47359 , n47358 , n47351 );
and ( n47360 , n47345 , n47198 );
or ( n47361 , n47359 , n47360 );
not ( n47362 , n47231 );
not ( n47363 , n46584 );
or ( n47364 , n47362 , n47363 );
not ( n47365 , n41954 );
not ( n47366 , n46510 );
or ( n47367 , n47365 , n47366 );
not ( n47368 , n41954 );
nand ( n47369 , n46576 , n47368 );
nand ( n47370 , n47367 , n47369 );
nand ( n47371 , n47370 , n46592 );
nand ( n47372 , n47364 , n47371 );
not ( n47373 , n47248 );
not ( n47374 , n47241 );
or ( n47375 , n47373 , n47374 );
and ( n47376 , n47047 , n47094 );
not ( n47377 , n47047 );
not ( n47378 , n47094 );
and ( n47379 , n47377 , n47378 );
or ( n47380 , n47376 , n47379 );
nand ( n47381 , n47380 , n46854 );
nand ( n47382 , n47375 , n47381 );
xor ( n47383 , n47372 , n47382 );
buf ( n47384 , n46334 );
not ( n47385 , n47384 );
not ( n47386 , n46412 );
not ( n47387 , n46163 );
or ( n47388 , n47386 , n47387 );
not ( n47389 , n41948 );
not ( n47390 , n47389 );
buf ( n47391 , n46325 );
nand ( n47392 , n47390 , n47391 );
nand ( n47393 , n47388 , n47392 );
not ( n47394 , n47393 );
or ( n47395 , n47385 , n47394 );
nand ( n47396 , n47209 , n46408 );
nand ( n47397 , n47395 , n47396 );
not ( n47398 , n46153 );
not ( n47399 , n46089 );
not ( n47400 , n46556 );
or ( n47401 , n47399 , n47400 );
not ( n47402 , n46089 );
nand ( n47403 , n30351 , n47402 );
nand ( n47404 , n47401 , n47403 );
not ( n47405 , n47404 );
or ( n47406 , n47398 , n47405 );
buf ( n47407 , n46925 );
nand ( n47408 , n47220 , n47407 );
nand ( n47409 , n47406 , n47408 );
xor ( n47410 , n47397 , n47409 );
xor ( n47411 , n47383 , n47410 );
xor ( n47412 , n47372 , n47382 );
and ( n47413 , n47412 , n47410 );
and ( n47414 , n47372 , n47382 );
or ( n47415 , n47413 , n47414 );
not ( n47416 , n47254 );
not ( n47417 , n46650 );
not ( n47418 , n41938 );
or ( n47419 , n47417 , n47418 );
nand ( n47420 , n46608 , n47260 );
nand ( n47421 , n47419 , n47420 );
not ( n47422 , n47421 );
or ( n47423 , n47416 , n47422 );
nand ( n47424 , n47262 , n46776 );
nand ( n47425 , n47423 , n47424 );
not ( n47426 , n47273 );
nand ( n47427 , n47426 , n46440 );
not ( n47428 , n47427 );
not ( n47429 , n47107 );
or ( n47430 , n47428 , n47429 );
nand ( n47431 , n47273 , n46441 );
nand ( n47432 , n47430 , n47431 );
and ( n47433 , n37022 , n37588 );
not ( n47434 , n37022 );
and ( n47435 , n47434 , n37589 );
nor ( n47436 , n47433 , n47435 );
buf ( n47437 , n47436 );
and ( n47438 , n47432 , n47437 );
xor ( n47439 , n47425 , n47438 );
xor ( n47440 , n47439 , n47238 );
xor ( n47441 , n47425 , n47438 );
and ( n47442 , n47441 , n47238 );
and ( n47443 , n47425 , n47438 );
or ( n47444 , n47442 , n47443 );
not ( n47445 , n47308 );
not ( n47446 , n47300 );
or ( n47447 , n47445 , n47446 );
not ( n47448 , n46273 );
buf ( n47449 , n47106 );
not ( n47450 , n47449 );
not ( n47451 , n47450 );
or ( n47452 , n47448 , n47451 );
nand ( n47453 , n47449 , n46824 );
nand ( n47454 , n47452 , n47453 );
nand ( n47455 , n47454 , n47148 );
nand ( n47456 , n47447 , n47455 );
not ( n47457 , n46188 );
not ( n47458 , n46425 );
not ( n47459 , n47154 );
or ( n47460 , n47458 , n47459 );
or ( n47461 , n47157 , n46425 );
nand ( n47462 , n47460 , n47461 );
not ( n47463 , n47462 );
or ( n47464 , n47457 , n47463 );
nand ( n47465 , n47290 , n46267 );
nand ( n47466 , n47464 , n47465 );
xor ( n47467 , n47456 , n47466 );
xor ( n47468 , n47467 , n47411 );
xor ( n47469 , n47456 , n47466 );
and ( n47470 , n47469 , n47411 );
and ( n47471 , n47456 , n47466 );
or ( n47472 , n47470 , n47471 );
not ( n47473 , n47437 );
and ( n47474 , n46441 , n47473 );
not ( n47475 , n46441 );
buf ( n47476 , n47437 );
and ( n47477 , n47475 , n47476 );
nor ( n47478 , n47474 , n47477 );
not ( n47479 , n47478 );
and ( n47480 , n47106 , n47273 );
not ( n47481 , n47106 );
and ( n47482 , n47481 , n47426 );
nor ( n47483 , n47480 , n47482 );
not ( n47484 , n47436 );
or ( n47485 , n47426 , n47484 );
nand ( n47486 , n47484 , n36938 );
nand ( n47487 , n47485 , n47486 );
nand ( n47488 , n47483 , n47487 );
not ( n47489 , n47488 );
not ( n47490 , n47489 );
or ( n47491 , n47479 , n47490 );
not ( n47492 , n45816 );
not ( n47493 , n47437 );
not ( n47494 , n47493 );
or ( n47495 , n47492 , n47494 );
nand ( n47496 , n47476 , n45767 );
nand ( n47497 , n47495 , n47496 );
buf ( n47498 , n47278 );
nand ( n47499 , n47497 , n47498 );
nand ( n47500 , n47491 , n47499 );
xor ( n47501 , n47500 , n47271 );
xor ( n47502 , n47501 , n47297 );
xor ( n47503 , n47500 , n47271 );
and ( n47504 , n47503 , n47297 );
and ( n47505 , n47500 , n47271 );
or ( n47506 , n47504 , n47505 );
not ( n47507 , n45748 );
not ( n47508 , n45837 );
not ( n47509 , n47508 );
not ( n47510 , n31958 );
buf ( n47511 , n47510 );
not ( n47512 , n47511 );
or ( n47513 , n47509 , n47512 );
not ( n47514 , n47508 );
nand ( n47515 , n41692 , n47514 );
nand ( n47516 , n47513 , n47515 );
not ( n47517 , n47516 );
or ( n47518 , n47507 , n47517 );
nand ( n47519 , n47322 , n46448 );
nand ( n47520 , n47518 , n47519 );
xor ( n47521 , n47440 , n47520 );
not ( n47522 , n46602 );
not ( n47523 , n46072 );
not ( n47524 , n30929 );
not ( n47525 , n47524 );
or ( n47526 , n47523 , n47525 );
buf ( n47527 , n30929 );
nand ( n47528 , n47527 , n46071 );
nand ( n47529 , n47526 , n47528 );
not ( n47530 , n47529 );
or ( n47531 , n47522 , n47530 );
nand ( n47532 , n46474 , n47336 );
nand ( n47533 , n47531 , n47532 );
xor ( n47534 , n47521 , n47533 );
xor ( n47535 , n47440 , n47520 );
and ( n47536 , n47535 , n47533 );
and ( n47537 , n47440 , n47520 );
or ( n47538 , n47536 , n47537 );
xor ( n47539 , n47316 , n47468 );
xor ( n47540 , n47539 , n47502 );
xor ( n47541 , n47316 , n47468 );
and ( n47542 , n47541 , n47502 );
and ( n47543 , n47316 , n47468 );
or ( n47544 , n47542 , n47543 );
xor ( n47545 , n47343 , n47349 );
xor ( n47546 , n47545 , n47534 );
xor ( n47547 , n47343 , n47349 );
and ( n47548 , n47547 , n47534 );
and ( n47549 , n47343 , n47349 );
or ( n47550 , n47548 , n47549 );
xor ( n47551 , n47540 , n47355 );
xor ( n47552 , n47551 , n47546 );
xor ( n47553 , n47540 , n47355 );
and ( n47554 , n47553 , n47546 );
and ( n47555 , n47540 , n47355 );
or ( n47556 , n47554 , n47555 );
not ( n47557 , n46408 );
not ( n47558 , n47393 );
or ( n47559 , n47557 , n47558 );
not ( n47560 , n47391 );
not ( n47561 , n47560 );
not ( n47562 , n46453 );
or ( n47563 , n47561 , n47562 );
nand ( n47564 , n47391 , n41946 );
nand ( n47565 , n47563 , n47564 );
nand ( n47566 , n47565 , n47384 );
nand ( n47567 , n47559 , n47566 );
not ( n47568 , n47370 );
not ( n47569 , n46584 );
or ( n47570 , n47568 , n47569 );
buf ( n47571 , n30379 );
not ( n47572 , n47571 );
not ( n47573 , n46510 );
or ( n47574 , n47572 , n47573 );
not ( n47575 , n47571 );
nand ( n47576 , n46511 , n47575 );
nand ( n47577 , n47574 , n47576 );
not ( n47578 , n46439 );
nand ( n47579 , n47577 , n47578 );
nand ( n47580 , n47570 , n47579 );
xor ( n47581 , n47567 , n47580 );
not ( n47582 , n47380 );
not ( n47583 , n47240 );
not ( n47584 , n47583 );
or ( n47585 , n47582 , n47584 );
not ( n47586 , n47227 );
not ( n47587 , n47094 );
or ( n47588 , n47586 , n47587 );
not ( n47589 , n47227 );
nand ( n47590 , n47378 , n47589 );
nand ( n47591 , n47588 , n47590 );
nand ( n47592 , n47591 , n46854 );
nand ( n47593 , n47585 , n47592 );
xor ( n47594 , n47581 , n47593 );
xor ( n47595 , n47567 , n47580 );
and ( n47596 , n47595 , n47593 );
and ( n47597 , n47567 , n47580 );
or ( n47598 , n47596 , n47597 );
and ( n47599 , n47409 , n47397 );
not ( n47600 , n46153 );
not ( n47601 , n46089 );
not ( n47602 , n47257 );
or ( n47603 , n47601 , n47602 );
nand ( n47604 , n30259 , n47402 );
nand ( n47605 , n47603 , n47604 );
not ( n47606 , n47605 );
or ( n47607 , n47600 , n47606 );
nand ( n47608 , n47404 , n47407 );
nand ( n47609 , n47607 , n47608 );
xor ( n47610 , n47599 , n47609 );
not ( n47611 , n46776 );
not ( n47612 , n47421 );
or ( n47613 , n47611 , n47612 );
not ( n47614 , n46650 );
not ( n47615 , n47287 );
or ( n47616 , n47614 , n47615 );
buf ( n47617 , n41861 );
nand ( n47618 , n47617 , n47260 );
nand ( n47619 , n47616 , n47618 );
nand ( n47620 , n47254 , n47619 );
nand ( n47621 , n47613 , n47620 );
xor ( n47622 , n47610 , n47621 );
xor ( n47623 , n47599 , n47609 );
and ( n47624 , n47623 , n47621 );
and ( n47625 , n47599 , n47609 );
or ( n47626 , n47624 , n47625 );
not ( n47627 , n47436 );
and ( n47628 , n37027 , n37571 );
not ( n47629 , n37027 );
not ( n47630 , n37571 );
and ( n47631 , n47629 , n47630 );
or ( n47632 , n47628 , n47631 );
not ( n47633 , n47632 );
or ( n47634 , n47627 , n47633 );
and ( n47635 , n37027 , n37571 );
not ( n47636 , n37027 );
and ( n47637 , n47636 , n47630 );
nor ( n47638 , n47635 , n47637 );
nand ( n47639 , n47638 , n47484 );
nand ( n47640 , n47634 , n47639 );
buf ( n47641 , n47640 );
nor ( n47642 , n47641 , n46441 );
not ( n47643 , n47454 );
not ( n47644 , n47300 );
or ( n47645 , n47643 , n47644 );
buf ( n47646 , n42050 );
not ( n47647 , n47646 );
not ( n47648 , n47107 );
or ( n47649 , n47647 , n47648 );
not ( n47650 , n47646 );
nand ( n47651 , n47449 , n47650 );
nand ( n47652 , n47649 , n47651 );
nand ( n47653 , n47652 , n47148 );
nand ( n47654 , n47645 , n47653 );
xor ( n47655 , n47642 , n47654 );
xor ( n47656 , n47655 , n47594 );
xor ( n47657 , n47642 , n47654 );
and ( n47658 , n47657 , n47594 );
and ( n47659 , n47642 , n47654 );
or ( n47660 , n47658 , n47659 );
not ( n47661 , n47497 );
not ( n47662 , n47489 );
or ( n47663 , n47661 , n47662 );
not ( n47664 , n46037 );
not ( n47665 , n47473 );
or ( n47666 , n47664 , n47665 );
nand ( n47667 , n47476 , n47306 );
nand ( n47668 , n47666 , n47667 );
nand ( n47669 , n47668 , n47498 );
nand ( n47670 , n47663 , n47669 );
xor ( n47671 , n47670 , n47415 );
xor ( n47672 , n47671 , n47622 );
xor ( n47673 , n47670 , n47415 );
and ( n47674 , n47673 , n47622 );
and ( n47675 , n47670 , n47415 );
or ( n47676 , n47674 , n47675 );
not ( n47677 , n46188 );
not ( n47678 , n46425 );
not ( n47679 , n30964 );
not ( n47680 , n47679 );
or ( n47681 , n47678 , n47680 );
nand ( n47682 , n30964 , n46422 );
nand ( n47683 , n47681 , n47682 );
not ( n47684 , n47683 );
or ( n47685 , n47677 , n47684 );
nand ( n47686 , n47462 , n46267 );
nand ( n47687 , n47685 , n47686 );
xor ( n47688 , n47687 , n47444 );
not ( n47689 , n46448 );
not ( n47690 , n47516 );
or ( n47691 , n47689 , n47690 );
not ( n47692 , n47508 );
not ( n47693 , n47332 );
or ( n47694 , n47692 , n47693 );
nand ( n47695 , n41683 , n45837 );
nand ( n47696 , n47694 , n47695 );
nand ( n47697 , n47696 , n45748 );
nand ( n47698 , n47691 , n47697 );
xor ( n47699 , n47688 , n47698 );
xor ( n47700 , n47687 , n47444 );
and ( n47701 , n47700 , n47698 );
and ( n47702 , n47687 , n47444 );
or ( n47703 , n47701 , n47702 );
not ( n47704 , n46474 );
not ( n47705 , n47529 );
or ( n47706 , n47704 , n47705 );
not ( n47707 , n46072 );
not ( n47708 , n41415 );
not ( n47709 , n47708 );
or ( n47710 , n47707 , n47709 );
nand ( n47711 , n41415 , n46071 );
nand ( n47712 , n47710 , n47711 );
nand ( n47713 , n47712 , n44004 );
nand ( n47714 , n47706 , n47713 );
xor ( n47715 , n47714 , n47472 );
xor ( n47716 , n47715 , n47656 );
xor ( n47717 , n47714 , n47472 );
and ( n47718 , n47717 , n47656 );
and ( n47719 , n47714 , n47472 );
or ( n47720 , n47718 , n47719 );
xor ( n47721 , n47506 , n47672 );
xor ( n47722 , n47721 , n47699 );
xor ( n47723 , n47506 , n47672 );
and ( n47724 , n47723 , n47699 );
and ( n47725 , n47506 , n47672 );
or ( n47726 , n47724 , n47725 );
xor ( n47727 , n47538 , n47716 );
xor ( n47728 , n47727 , n47544 );
xor ( n47729 , n47538 , n47716 );
and ( n47730 , n47729 , n47544 );
and ( n47731 , n47538 , n47716 );
or ( n47732 , n47730 , n47731 );
xor ( n47733 , n47722 , n47550 );
xor ( n47734 , n47733 , n47728 );
xor ( n47735 , n47722 , n47550 );
and ( n47736 , n47735 , n47728 );
and ( n47737 , n47722 , n47550 );
or ( n47738 , n47736 , n47737 );
not ( n47739 , n46854 );
buf ( n47740 , n41954 );
not ( n47741 , n47740 );
not ( n47742 , n47094 );
or ( n47743 , n47741 , n47742 );
buf ( n47744 , n46758 );
nand ( n47745 , n47744 , n47368 );
nand ( n47746 , n47743 , n47745 );
not ( n47747 , n47746 );
or ( n47748 , n47739 , n47747 );
nand ( n47749 , n47591 , n47583 );
nand ( n47750 , n47748 , n47749 );
not ( n47751 , n47384 );
not ( n47752 , n47560 );
not ( n47753 , n46556 );
or ( n47754 , n47752 , n47753 );
nand ( n47755 , n30351 , n47391 );
nand ( n47756 , n47754 , n47755 );
not ( n47757 , n47756 );
or ( n47758 , n47751 , n47757 );
nand ( n47759 , n47565 , n46408 );
nand ( n47760 , n47758 , n47759 );
not ( n47761 , n47760 );
not ( n47762 , n47577 );
not ( n47763 , n46584 );
or ( n47764 , n47762 , n47763 );
not ( n47765 , n46163 );
not ( n47766 , n47765 );
not ( n47767 , n46510 );
or ( n47768 , n47766 , n47767 );
not ( n47769 , n46510 );
nand ( n47770 , n47769 , n47389 );
nand ( n47771 , n47768 , n47770 );
nand ( n47772 , n47771 , n47578 );
nand ( n47773 , n47764 , n47772 );
not ( n47774 , n47773 );
not ( n47775 , n47774 );
or ( n47776 , n47761 , n47775 );
or ( n47777 , n47774 , n47760 );
nand ( n47778 , n47776 , n47777 );
xor ( n47779 , n47750 , n47778 );
nand ( n47780 , n47632 , n46440 );
nand ( n47781 , n47780 , n47473 );
not ( n47782 , n46440 );
nand ( n47783 , n47782 , n47638 );
and ( n47784 , n47781 , n47783 );
buf ( n47785 , n35578 );
nand ( n47786 , n35705 , n47785 );
not ( n47787 , n47786 );
not ( n47788 , n47787 );
not ( n47789 , n36984 );
not ( n47790 , n47789 );
or ( n47791 , n47788 , n47790 );
nand ( n47792 , n36984 , n47786 );
nand ( n47793 , n47791 , n47792 );
buf ( n47794 , n47793 );
not ( n47795 , n47794 );
nor ( n47796 , n47784 , n47795 );
xor ( n47797 , n47779 , n47796 );
xor ( n47798 , n47750 , n47778 );
and ( n47799 , n47798 , n47796 );
and ( n47800 , n47750 , n47778 );
or ( n47801 , n47799 , n47800 );
not ( n47802 , n46153 );
not ( n47803 , n47402 );
not ( n47804 , n47803 );
not ( n47805 , n41938 );
or ( n47806 , n47804 , n47805 );
not ( n47807 , n46607 );
buf ( n47808 , n47402 );
nand ( n47809 , n47807 , n47808 );
nand ( n47810 , n47806 , n47809 );
not ( n47811 , n47810 );
or ( n47812 , n47802 , n47811 );
nand ( n47813 , n47605 , n47407 );
nand ( n47814 , n47812 , n47813 );
not ( n47815 , n47652 );
not ( n47816 , n47300 );
or ( n47817 , n47815 , n47816 );
not ( n47818 , n47047 );
not ( n47819 , n47107 );
or ( n47820 , n47818 , n47819 );
not ( n47821 , n47047 );
nand ( n47822 , n47108 , n47821 );
nand ( n47823 , n47820 , n47822 );
nand ( n47824 , n47823 , n47148 );
nand ( n47825 , n47817 , n47824 );
xor ( n47826 , n47814 , n47825 );
not ( n47827 , n47253 );
not ( n47828 , n47827 );
not ( n47829 , n46650 );
not ( n47830 , n47154 );
or ( n47831 , n47829 , n47830 );
nand ( n47832 , n47260 , n47158 );
nand ( n47833 , n47831 , n47832 );
not ( n47834 , n47833 );
or ( n47835 , n47828 , n47834 );
nand ( n47836 , n47619 , n46776 );
nand ( n47837 , n47835 , n47836 );
xor ( n47838 , n47826 , n47837 );
xor ( n47839 , n47814 , n47825 );
and ( n47840 , n47839 , n47837 );
and ( n47841 , n47814 , n47825 );
or ( n47842 , n47840 , n47841 );
not ( n47843 , n47668 );
not ( n47844 , n47489 );
or ( n47845 , n47843 , n47844 );
not ( n47846 , n46273 );
not ( n47847 , n47473 );
or ( n47848 , n47846 , n47847 );
nand ( n47849 , n47476 , n46824 );
nand ( n47850 , n47848 , n47849 );
nand ( n47851 , n47850 , n47498 );
nand ( n47852 , n47845 , n47851 );
xor ( n47853 , n47598 , n47852 );
not ( n47854 , n47794 );
not ( n47855 , n47854 );
and ( n47856 , n46440 , n47855 );
not ( n47857 , n46440 );
and ( n47858 , n47857 , n47854 );
nor ( n47859 , n47856 , n47858 );
not ( n47860 , n47859 );
not ( n47861 , n47787 );
not ( n47862 , n47789 );
or ( n47863 , n47861 , n47862 );
nand ( n47864 , n47863 , n47792 );
nand ( n47865 , n47638 , n47864 );
not ( n47866 , n47865 );
not ( n47867 , n47864 );
nand ( n47868 , n47867 , n47632 );
not ( n47869 , n47868 );
or ( n47870 , n47866 , n47869 );
nand ( n47871 , n47870 , n47640 );
not ( n47872 , n47871 );
buf ( n47873 , n47872 );
not ( n47874 , n47873 );
or ( n47875 , n47860 , n47874 );
not ( n47876 , n45816 );
not ( n47877 , n47854 );
or ( n47878 , n47876 , n47877 );
nand ( n47879 , n47794 , n45767 );
nand ( n47880 , n47878 , n47879 );
not ( n47881 , n47641 );
nand ( n47882 , n47880 , n47881 );
nand ( n47883 , n47875 , n47882 );
xor ( n47884 , n47853 , n47883 );
xor ( n47885 , n47598 , n47852 );
and ( n47886 , n47885 , n47883 );
and ( n47887 , n47598 , n47852 );
or ( n47888 , n47886 , n47887 );
xor ( n47889 , n47797 , n47626 );
not ( n47890 , n46448 );
not ( n47891 , n47696 );
or ( n47892 , n47890 , n47891 );
not ( n47893 , n46554 );
not ( n47894 , n47524 );
or ( n47895 , n47893 , n47894 );
nand ( n47896 , n30929 , n46559 );
nand ( n47897 , n47895 , n47896 );
nand ( n47898 , n47897 , n45748 );
nand ( n47899 , n47892 , n47898 );
xor ( n47900 , n47889 , n47899 );
xor ( n47901 , n47797 , n47626 );
and ( n47902 , n47901 , n47899 );
and ( n47903 , n47797 , n47626 );
or ( n47904 , n47902 , n47903 );
not ( n47905 , n44004 );
and ( n47906 , n41575 , n46071 );
not ( n47907 , n41575 );
and ( n47908 , n47907 , n46072 );
or ( n47909 , n47906 , n47908 );
not ( n47910 , n47909 );
or ( n47911 , n47905 , n47910 );
nand ( n47912 , n47712 , n46474 );
nand ( n47913 , n47911 , n47912 );
not ( n47914 , n46188 );
not ( n47915 , n46425 );
not ( n47916 , n47178 );
or ( n47917 , n47915 , n47916 );
not ( n47918 , n47510 );
nand ( n47919 , n47918 , n46422 );
nand ( n47920 , n47917 , n47919 );
not ( n47921 , n47920 );
or ( n47922 , n47914 , n47921 );
nand ( n47923 , n47683 , n46267 );
nand ( n47924 , n47922 , n47923 );
xor ( n47925 , n47913 , n47924 );
xor ( n47926 , n47925 , n47660 );
xor ( n47927 , n47913 , n47924 );
and ( n47928 , n47927 , n47660 );
and ( n47929 , n47913 , n47924 );
or ( n47930 , n47928 , n47929 );
xor ( n47931 , n47838 , n47676 );
xor ( n47932 , n47931 , n47884 );
xor ( n47933 , n47838 , n47676 );
and ( n47934 , n47933 , n47884 );
and ( n47935 , n47838 , n47676 );
or ( n47936 , n47934 , n47935 );
xor ( n47937 , n47703 , n47900 );
xor ( n47938 , n47937 , n47720 );
xor ( n47939 , n47703 , n47900 );
and ( n47940 , n47939 , n47720 );
and ( n47941 , n47703 , n47900 );
or ( n47942 , n47940 , n47941 );
xor ( n47943 , n47926 , n47932 );
xor ( n47944 , n47943 , n47726 );
xor ( n47945 , n47926 , n47932 );
and ( n47946 , n47945 , n47726 );
and ( n47947 , n47926 , n47932 );
or ( n47948 , n47946 , n47947 );
xor ( n47949 , n47938 , n47732 );
xor ( n47950 , n47949 , n47944 );
xor ( n47951 , n47938 , n47732 );
and ( n47952 , n47951 , n47944 );
and ( n47953 , n47938 , n47732 );
or ( n47954 , n47952 , n47953 );
not ( n47955 , n47771 );
not ( n47956 , n46584 );
or ( n47957 , n47955 , n47956 );
not ( n47958 , n46453 );
not ( n47959 , n47958 );
not ( n47960 , n46510 );
or ( n47961 , n47959 , n47960 );
not ( n47962 , n46510 );
nand ( n47963 , n47962 , n46453 );
nand ( n47964 , n47961 , n47963 );
nand ( n47965 , n47964 , n47578 );
nand ( n47966 , n47957 , n47965 );
not ( n47967 , n47746 );
not ( n47968 , n47583 );
or ( n47969 , n47967 , n47968 );
not ( n47970 , n47571 );
not ( n47971 , n46757 );
or ( n47972 , n47970 , n47971 );
nand ( n47973 , n47575 , n46834 );
nand ( n47974 , n47972 , n47973 );
nand ( n47975 , n47974 , n46854 );
nand ( n47976 , n47969 , n47975 );
xor ( n47977 , n47966 , n47976 );
not ( n47978 , n47384 );
buf ( n47979 , n46505 );
not ( n47980 , n47979 );
not ( n47981 , n47980 );
not ( n47982 , n30259 );
not ( n47983 , n47982 );
or ( n47984 , n47981 , n47983 );
nand ( n47985 , n30259 , n47979 );
nand ( n47986 , n47984 , n47985 );
not ( n47987 , n47986 );
or ( n47988 , n47978 , n47987 );
nand ( n47989 , n47756 , n46408 );
nand ( n47990 , n47988 , n47989 );
xor ( n47991 , n47977 , n47990 );
xor ( n47992 , n47966 , n47976 );
and ( n47993 , n47992 , n47990 );
and ( n47994 , n47966 , n47976 );
or ( n47995 , n47993 , n47994 );
not ( n47996 , n47760 );
nor ( n47997 , n47996 , n47774 );
not ( n47998 , n47793 );
not ( n47999 , n47998 );
not ( n48000 , n36626 );
not ( n48001 , n35726 );
nor ( n48002 , n48001 , n36619 );
not ( n48003 , n48002 );
or ( n48004 , n48000 , n48003 );
nand ( n48005 , n48004 , n37649 );
nand ( n48006 , n36947 , n35592 );
and ( n48007 , n48005 , n48006 );
not ( n48008 , n48005 );
not ( n48009 , n48006 );
and ( n48010 , n48008 , n48009 );
nor ( n48011 , n48007 , n48010 );
not ( n48012 , n48011 );
or ( n48013 , n47999 , n48012 );
not ( n48014 , n48011 );
nand ( n48015 , n47793 , n48014 );
nand ( n48016 , n48013 , n48015 );
not ( n48017 , n48016 );
and ( n48018 , n48017 , n46440 );
xor ( n48019 , n47997 , n48018 );
not ( n48020 , n47407 );
not ( n48021 , n47810 );
or ( n48022 , n48020 , n48021 );
not ( n48023 , n47808 );
not ( n48024 , n48023 );
not ( n48025 , n46719 );
or ( n48026 , n48024 , n48025 );
not ( n48027 , n46994 );
nand ( n48028 , n48027 , n47808 );
nand ( n48029 , n48026 , n48028 );
nand ( n48030 , n48029 , n46153 );
nand ( n48031 , n48022 , n48030 );
xor ( n48032 , n48019 , n48031 );
xor ( n48033 , n47997 , n48018 );
and ( n48034 , n48033 , n48031 );
and ( n48035 , n47997 , n48018 );
or ( n48036 , n48034 , n48035 );
not ( n48037 , n47823 );
not ( n48038 , n47300 );
or ( n48039 , n48037 , n48038 );
not ( n48040 , n47227 );
not ( n48041 , n47276 );
or ( n48042 , n48040 , n48041 );
nand ( n48043 , n47108 , n47589 );
nand ( n48044 , n48042 , n48043 );
nand ( n48045 , n48044 , n47148 );
nand ( n48046 , n48039 , n48045 );
not ( n48047 , n47850 );
not ( n48048 , n47489 );
or ( n48049 , n48047 , n48048 );
not ( n48050 , n47646 );
not ( n48051 , n47493 );
or ( n48052 , n48050 , n48051 );
nand ( n48053 , n47476 , n47650 );
nand ( n48054 , n48052 , n48053 );
nand ( n48055 , n48054 , n47498 );
nand ( n48056 , n48049 , n48055 );
xor ( n48057 , n48046 , n48056 );
xor ( n48058 , n48057 , n47991 );
xor ( n48059 , n48046 , n48056 );
and ( n48060 , n48059 , n47991 );
and ( n48061 , n48046 , n48056 );
or ( n48062 , n48060 , n48061 );
not ( n48063 , n47880 );
not ( n48064 , n47873 );
or ( n48065 , n48063 , n48064 );
not ( n48066 , n46037 );
not ( n48067 , n47854 );
or ( n48068 , n48066 , n48067 );
nand ( n48069 , n47794 , n47306 );
nand ( n48070 , n48068 , n48069 );
nand ( n48071 , n48070 , n47881 );
nand ( n48072 , n48065 , n48071 );
buf ( n48073 , n45896 );
not ( n48074 , n48073 );
not ( n48075 , n46650 );
not ( n48076 , n47318 );
or ( n48077 , n48075 , n48076 );
not ( n48078 , n46650 );
nand ( n48079 , n30964 , n48078 );
nand ( n48080 , n48077 , n48079 );
not ( n48081 , n48080 );
or ( n48082 , n48074 , n48081 );
nand ( n48083 , n47833 , n46776 );
nand ( n48084 , n48082 , n48083 );
xor ( n48085 , n48072 , n48084 );
xor ( n48086 , n48085 , n47801 );
xor ( n48087 , n48072 , n48084 );
and ( n48088 , n48087 , n47801 );
and ( n48089 , n48072 , n48084 );
or ( n48090 , n48088 , n48089 );
not ( n48091 , n46448 );
not ( n48092 , n47897 );
or ( n48093 , n48091 , n48092 );
not ( n48094 , n46554 );
not ( n48095 , n47708 );
or ( n48096 , n48094 , n48095 );
nand ( n48097 , n41415 , n46559 );
nand ( n48098 , n48096 , n48097 );
nand ( n48099 , n48098 , n45832 );
nand ( n48100 , n48093 , n48099 );
xor ( n48101 , n48100 , n48032 );
xor ( n48102 , n48101 , n47842 );
xor ( n48103 , n48100 , n48032 );
and ( n48104 , n48103 , n47842 );
and ( n48105 , n48100 , n48032 );
or ( n48106 , n48104 , n48105 );
not ( n48107 , n46267 );
not ( n48108 , n47920 );
or ( n48109 , n48107 , n48108 );
and ( n48110 , n41683 , n46422 );
not ( n48111 , n41683 );
and ( n48112 , n48111 , n46425 );
or ( n48113 , n48110 , n48112 );
nand ( n48114 , n48113 , n46188 );
nand ( n48115 , n48109 , n48114 );
not ( n48116 , n44004 );
not ( n48117 , n46072 );
not ( n48118 , n44141 );
not ( n48119 , n48118 );
or ( n48120 , n48117 , n48119 );
nand ( n48121 , n41668 , n46071 );
nand ( n48122 , n48120 , n48121 );
not ( n48123 , n48122 );
or ( n48124 , n48116 , n48123 );
nand ( n48125 , n47909 , n46474 );
nand ( n48126 , n48124 , n48125 );
xor ( n48127 , n48115 , n48126 );
xor ( n48128 , n48127 , n47888 );
xor ( n48129 , n48115 , n48126 );
and ( n48130 , n48129 , n47888 );
and ( n48131 , n48115 , n48126 );
or ( n48132 , n48130 , n48131 );
xor ( n48133 , n48058 , n47930 );
xor ( n48134 , n48133 , n48086 );
xor ( n48135 , n48058 , n47930 );
and ( n48136 , n48135 , n48086 );
and ( n48137 , n48058 , n47930 );
or ( n48138 , n48136 , n48137 );
xor ( n48139 , n47904 , n48128 );
xor ( n48140 , n48139 , n48102 );
xor ( n48141 , n47904 , n48128 );
and ( n48142 , n48141 , n48102 );
and ( n48143 , n47904 , n48128 );
or ( n48144 , n48142 , n48143 );
xor ( n48145 , n47936 , n48134 );
xor ( n48146 , n48145 , n47942 );
xor ( n48147 , n47936 , n48134 );
and ( n48148 , n48147 , n47942 );
and ( n48149 , n47936 , n48134 );
or ( n48150 , n48148 , n48149 );
xor ( n48151 , n48140 , n47948 );
xor ( n48152 , n48151 , n48146 );
xor ( n48153 , n48140 , n47948 );
and ( n48154 , n48153 , n48146 );
and ( n48155 , n48140 , n47948 );
or ( n48156 , n48154 , n48155 );
not ( n48157 , n47384 );
not ( n48158 , n46608 );
not ( n48159 , n47979 );
or ( n48160 , n48158 , n48159 );
nand ( n48161 , n47980 , n41938 );
nand ( n48162 , n48160 , n48161 );
not ( n48163 , n48162 );
or ( n48164 , n48157 , n48163 );
nand ( n48165 , n47986 , n46408 );
nand ( n48166 , n48164 , n48165 );
not ( n48167 , n47964 );
not ( n48168 , n46584 );
or ( n48169 , n48167 , n48168 );
not ( n48170 , n46820 );
not ( n48171 , n30351 );
not ( n48172 , n48171 );
or ( n48173 , n48170 , n48172 );
nand ( n48174 , n30351 , n46573 );
nand ( n48175 , n48173 , n48174 );
nand ( n48176 , n48175 , n46592 );
nand ( n48177 , n48169 , n48176 );
not ( n48178 , n47974 );
not ( n48179 , n47241 );
or ( n48180 , n48178 , n48179 );
and ( n48181 , n46835 , n46163 );
not ( n48182 , n46835 );
and ( n48183 , n48182 , n47765 );
or ( n48184 , n48181 , n48183 );
nand ( n48185 , n48184 , n47060 );
nand ( n48186 , n48180 , n48185 );
xor ( n48187 , n48177 , n48186 );
xor ( n48188 , n48166 , n48187 );
not ( n48189 , n46440 );
not ( n48190 , n48011 );
not ( n48191 , n48190 );
or ( n48192 , n48189 , n48191 );
nand ( n48193 , n48192 , n47795 );
buf ( n48194 , n48011 );
nand ( n48195 , n48194 , n46441 );
and ( n48196 , n48193 , n48195 );
not ( n48197 , n37583 );
not ( n48198 , n36985 );
or ( n48199 , n48197 , n48198 );
nand ( n48200 , n48199 , n36952 );
buf ( n48201 , n48200 );
not ( n48202 , n48201 );
nor ( n48203 , n48196 , n48202 );
xor ( n48204 , n48188 , n48203 );
xor ( n48205 , n48166 , n48187 );
and ( n48206 , n48205 , n48203 );
and ( n48207 , n48166 , n48187 );
or ( n48208 , n48206 , n48207 );
not ( n48209 , n48044 );
not ( n48210 , n47139 );
or ( n48211 , n48209 , n48210 );
not ( n48212 , n47740 );
not ( n48213 , n47107 );
or ( n48214 , n48212 , n48213 );
nand ( n48215 , n47449 , n47368 );
nand ( n48216 , n48214 , n48215 );
nand ( n48217 , n48216 , n47147 );
nand ( n48218 , n48211 , n48217 );
not ( n48219 , n46153 );
not ( n48220 , n47803 );
not ( n48221 , n46880 );
or ( n48222 , n48220 , n48221 );
not ( n48223 , n47157 );
nand ( n48224 , n48223 , n47402 );
nand ( n48225 , n48222 , n48224 );
not ( n48226 , n48225 );
or ( n48227 , n48219 , n48226 );
nand ( n48228 , n48029 , n47407 );
nand ( n48229 , n48227 , n48228 );
xor ( n48230 , n48218 , n48229 );
not ( n48231 , n48070 );
not ( n48232 , n47872 );
or ( n48233 , n48231 , n48232 );
not ( n48234 , n46273 );
not ( n48235 , n47794 );
not ( n48236 , n48235 );
or ( n48237 , n48234 , n48236 );
nand ( n48238 , n47794 , n46824 );
nand ( n48239 , n48237 , n48238 );
not ( n48240 , n47641 );
nand ( n48241 , n48239 , n48240 );
nand ( n48242 , n48233 , n48241 );
xor ( n48243 , n48230 , n48242 );
xor ( n48244 , n48218 , n48229 );
and ( n48245 , n48244 , n48242 );
and ( n48246 , n48218 , n48229 );
or ( n48247 , n48245 , n48246 );
not ( n48248 , n48054 );
not ( n48249 , n47489 );
or ( n48250 , n48248 , n48249 );
not ( n48251 , n47047 );
not ( n48252 , n47493 );
or ( n48253 , n48251 , n48252 );
nand ( n48254 , n47476 , n47821 );
nand ( n48255 , n48253 , n48254 );
nand ( n48256 , n48255 , n47278 );
nand ( n48257 , n48250 , n48256 );
not ( n48258 , n46440 );
not ( n48259 , n48201 );
not ( n48260 , n48259 );
or ( n48261 , n48258 , n48260 );
not ( n48262 , n48259 );
nand ( n48263 , n48262 , n46441 );
nand ( n48264 , n48261 , n48263 );
not ( n48265 , n48264 );
xor ( n48266 , n48200 , n48190 );
nand ( n48267 , n48266 , n48016 );
not ( n48268 , n48267 );
not ( n48269 , n48268 );
or ( n48270 , n48265 , n48269 );
not ( n48271 , n45816 );
not ( n48272 , n48202 );
or ( n48273 , n48271 , n48272 );
nand ( n48274 , n48201 , n45767 );
nand ( n48275 , n48273 , n48274 );
not ( n48276 , n48017 );
not ( n48277 , n48276 );
nand ( n48278 , n48275 , n48277 );
nand ( n48279 , n48270 , n48278 );
xor ( n48280 , n48257 , n48279 );
xor ( n48281 , n48280 , n47995 );
xor ( n48282 , n48257 , n48279 );
and ( n48283 , n48282 , n47995 );
and ( n48284 , n48257 , n48279 );
or ( n48285 , n48283 , n48284 );
not ( n48286 , n47827 );
not ( n48287 , n46650 );
not ( n48288 , n47178 );
or ( n48289 , n48287 , n48288 );
not ( n48290 , n46650 );
nand ( n48291 , n47918 , n48290 );
nand ( n48292 , n48289 , n48291 );
not ( n48293 , n48292 );
or ( n48294 , n48286 , n48293 );
not ( n48295 , n46775 );
nand ( n48296 , n48080 , n48295 );
nand ( n48297 , n48294 , n48296 );
xor ( n48298 , n48036 , n48297 );
not ( n48299 , n46474 );
not ( n48300 , n48122 );
or ( n48301 , n48299 , n48300 );
not ( n48302 , n46072 );
not ( n48303 , n41531 );
not ( n48304 , n48303 );
or ( n48305 , n48302 , n48304 );
not ( n48306 , n41530 );
nand ( n48307 , n48306 , n46071 );
nand ( n48308 , n48305 , n48307 );
nand ( n48309 , n48308 , n44004 );
nand ( n48310 , n48301 , n48309 );
xor ( n48311 , n48298 , n48310 );
xor ( n48312 , n48036 , n48297 );
and ( n48313 , n48312 , n48310 );
and ( n48314 , n48036 , n48297 );
or ( n48315 , n48313 , n48314 );
not ( n48316 , n45832 );
not ( n48317 , n46554 );
not ( n48318 , n41575 );
not ( n48319 , n48318 );
or ( n48320 , n48317 , n48319 );
nand ( n48321 , n41575 , n46559 );
nand ( n48322 , n48320 , n48321 );
not ( n48323 , n48322 );
or ( n48324 , n48316 , n48323 );
nand ( n48325 , n48098 , n46448 );
nand ( n48326 , n48324 , n48325 );
xor ( n48327 , n48326 , n48204 );
not ( n48328 , n46188 );
not ( n48329 , n46425 );
not ( n48330 , n47524 );
or ( n48331 , n48329 , n48330 );
not ( n48332 , n47524 );
nand ( n48333 , n48332 , n46422 );
nand ( n48334 , n48331 , n48333 );
not ( n48335 , n48334 );
or ( n48336 , n48328 , n48335 );
nand ( n48337 , n48113 , n46267 );
nand ( n48338 , n48336 , n48337 );
xor ( n48339 , n48327 , n48338 );
xor ( n48340 , n48326 , n48204 );
and ( n48341 , n48340 , n48338 );
and ( n48342 , n48326 , n48204 );
or ( n48343 , n48341 , n48342 );
xor ( n48344 , n48062 , n48243 );
xor ( n48345 , n48344 , n48281 );
xor ( n48346 , n48062 , n48243 );
and ( n48347 , n48346 , n48281 );
and ( n48348 , n48062 , n48243 );
or ( n48349 , n48347 , n48348 );
xor ( n48350 , n48090 , n48106 );
xor ( n48351 , n48350 , n48339 );
xor ( n48352 , n48090 , n48106 );
and ( n48353 , n48352 , n48339 );
and ( n48354 , n48090 , n48106 );
or ( n48355 , n48353 , n48354 );
xor ( n48356 , n48132 , n48311 );
xor ( n48357 , n48356 , n48345 );
xor ( n48358 , n48132 , n48311 );
and ( n48359 , n48358 , n48345 );
and ( n48360 , n48132 , n48311 );
or ( n48361 , n48359 , n48360 );
xor ( n48362 , n48138 , n48351 );
xor ( n48363 , n48362 , n48144 );
xor ( n48364 , n48138 , n48351 );
and ( n48365 , n48364 , n48144 );
and ( n48366 , n48138 , n48351 );
or ( n48367 , n48365 , n48366 );
xor ( n48368 , n48357 , n48150 );
xor ( n48369 , n48368 , n48363 );
xor ( n48370 , n48357 , n48150 );
and ( n48371 , n48370 , n48363 );
and ( n48372 , n48357 , n48150 );
or ( n48373 , n48371 , n48372 );
not ( n48374 , n48184 );
not ( n48375 , n47241 );
or ( n48376 , n48374 , n48375 );
not ( n48377 , n47958 );
not ( n48378 , n46757 );
or ( n48379 , n48377 , n48378 );
nand ( n48380 , n46834 , n46453 );
nand ( n48381 , n48379 , n48380 );
nand ( n48382 , n47060 , n48381 );
nand ( n48383 , n48376 , n48382 );
not ( n48384 , n47578 );
not ( n48385 , n47962 );
not ( n48386 , n30259 );
not ( n48387 , n48386 );
or ( n48388 , n48385 , n48387 );
nand ( n48389 , n30259 , n46821 );
nand ( n48390 , n48388 , n48389 );
not ( n48391 , n48390 );
or ( n48392 , n48384 , n48391 );
nand ( n48393 , n48175 , n46584 );
nand ( n48394 , n48392 , n48393 );
xor ( n48395 , n48383 , n48394 );
not ( n48396 , n46408 );
not ( n48397 , n48162 );
or ( n48398 , n48396 , n48397 );
not ( n48399 , n47980 );
not ( n48400 , n46719 );
or ( n48401 , n48399 , n48400 );
nand ( n48402 , n41861 , n47979 );
nand ( n48403 , n48401 , n48402 );
nand ( n48404 , n48403 , n47384 );
nand ( n48405 , n48398 , n48404 );
xor ( n48406 , n48395 , n48405 );
xor ( n48407 , n48383 , n48394 );
and ( n48408 , n48407 , n48405 );
and ( n48409 , n48383 , n48394 );
or ( n48410 , n48408 , n48409 );
and ( n48411 , n48177 , n48186 );
not ( n48412 , n48216 );
not ( n48413 , n47300 );
or ( n48414 , n48412 , n48413 );
not ( n48415 , n47571 );
not ( n48416 , n47107 );
or ( n48417 , n48415 , n48416 );
nand ( n48418 , n47449 , n47575 );
nand ( n48419 , n48417 , n48418 );
nand ( n48420 , n48419 , n47148 );
nand ( n48421 , n48414 , n48420 );
xor ( n48422 , n48411 , n48421 );
not ( n48423 , n48255 );
not ( n48424 , n47489 );
or ( n48425 , n48423 , n48424 );
not ( n48426 , n47227 );
not ( n48427 , n47473 );
or ( n48428 , n48426 , n48427 );
nand ( n48429 , n47437 , n47589 );
nand ( n48430 , n48428 , n48429 );
nand ( n48431 , n47498 , n48430 );
nand ( n48432 , n48425 , n48431 );
xor ( n48433 , n48422 , n48432 );
xor ( n48434 , n48411 , n48421 );
and ( n48435 , n48434 , n48432 );
and ( n48436 , n48411 , n48421 );
or ( n48437 , n48435 , n48436 );
xor ( n48438 , n48247 , n48285 );
xor ( n48439 , n48438 , n48433 );
xor ( n48440 , n48439 , n48349 );
not ( n48441 , n48239 );
not ( n48442 , n47872 );
or ( n48443 , n48441 , n48442 );
not ( n48444 , n47646 );
not ( n48445 , n48235 );
or ( n48446 , n48444 , n48445 );
nand ( n48447 , n47794 , n47650 );
nand ( n48448 , n48446 , n48447 );
nand ( n48449 , n48448 , n48240 );
nand ( n48450 , n48443 , n48449 );
buf ( n48451 , n48016 );
not ( n48452 , n48451 );
not ( n48453 , n48452 );
not ( n48454 , n47306 );
not ( n48455 , n48200 );
not ( n48456 , n48455 );
not ( n48457 , n48456 );
or ( n48458 , n48454 , n48457 );
nand ( n48459 , n48259 , n46037 );
nand ( n48460 , n48458 , n48459 );
not ( n48461 , n48460 );
or ( n48462 , n48453 , n48461 );
not ( n48463 , n48267 );
nand ( n48464 , n48463 , n48275 );
nand ( n48465 , n48462 , n48464 );
xor ( n48466 , n48450 , n48465 );
and ( n48467 , n37457 , n36239 );
not ( n48468 , n48467 );
not ( n48469 , n36966 );
or ( n48470 , n48468 , n48469 );
or ( n48471 , n48467 , n36966 );
nand ( n48472 , n48470 , n48471 );
not ( n48473 , n48472 );
and ( n48474 , n48473 , n48201 );
not ( n48475 , n48473 );
and ( n48476 , n48475 , n48455 );
nor ( n48477 , n48474 , n48476 );
not ( n48478 , n48477 );
buf ( n48479 , n48478 );
nor ( n48480 , n48479 , n46441 );
xor ( n48481 , n48466 , n48480 );
not ( n48482 , n46072 );
not ( n48483 , n41407 );
not ( n48484 , n48483 );
or ( n48485 , n48482 , n48484 );
buf ( n48486 , n41407 );
nand ( n48487 , n48486 , n46071 );
nand ( n48488 , n48485 , n48487 );
not ( n48489 , n48488 );
not ( n48490 , n44004 );
or ( n48491 , n48489 , n48490 );
nand ( n48492 , n48308 , n46474 );
nand ( n48493 , n48491 , n48492 );
xor ( n48494 , n48481 , n48493 );
not ( n48495 , n46153 );
not ( n48496 , n30964 );
xor ( n48497 , n47402 , n48496 );
not ( n48498 , n48497 );
or ( n48499 , n48495 , n48498 );
nand ( n48500 , n48225 , n47407 );
nand ( n48501 , n48499 , n48500 );
xor ( n48502 , n48406 , n48501 );
xor ( n48503 , n48502 , n48208 );
xor ( n48504 , n48494 , n48503 );
xor ( n48505 , n48440 , n48504 );
xor ( n48506 , n48505 , n48367 );
xor ( n48507 , n48343 , n48315 );
not ( n48508 , n45832 );
not ( n48509 , n46554 );
not ( n48510 , n41667 );
not ( n48511 , n48510 );
or ( n48512 , n48509 , n48511 );
nand ( n48513 , n44141 , n46559 );
nand ( n48514 , n48512 , n48513 );
not ( n48515 , n48514 );
or ( n48516 , n48508 , n48515 );
nand ( n48517 , n48322 , n46448 );
nand ( n48518 , n48516 , n48517 );
not ( n48519 , n46776 );
not ( n48520 , n48292 );
or ( n48521 , n48519 , n48520 );
not ( n48522 , n46650 );
not ( n48523 , n41683 );
not ( n48524 , n48523 );
or ( n48525 , n48522 , n48524 );
nand ( n48526 , n41683 , n48290 );
nand ( n48527 , n48525 , n48526 );
nand ( n48528 , n48527 , n47827 );
nand ( n48529 , n48521 , n48528 );
xor ( n48530 , n48518 , n48529 );
not ( n48531 , n46267 );
not ( n48532 , n48334 );
or ( n48533 , n48531 , n48532 );
not ( n48534 , n46425 );
not ( n48535 , n41415 );
not ( n48536 , n48535 );
or ( n48537 , n48534 , n48536 );
nand ( n48538 , n41415 , n46422 );
nand ( n48539 , n48537 , n48538 );
nand ( n48540 , n48539 , n46188 );
nand ( n48541 , n48533 , n48540 );
xor ( n48542 , n48530 , n48541 );
xor ( n48543 , n48507 , n48542 );
xor ( n48544 , n48543 , n48355 );
xor ( n48545 , n48544 , n48361 );
xor ( n48546 , n48506 , n48545 );
xor ( n48547 , n48505 , n48367 );
and ( n48548 , n48547 , n48545 );
and ( n48549 , n48505 , n48367 );
or ( n48550 , n48548 , n48549 );
xor ( n48551 , n48450 , n48465 );
and ( n48552 , n48551 , n48480 );
and ( n48553 , n48450 , n48465 );
or ( n48554 , n48552 , n48553 );
xor ( n48555 , n48406 , n48501 );
and ( n48556 , n48555 , n48208 );
and ( n48557 , n48406 , n48501 );
or ( n48558 , n48556 , n48557 );
xor ( n48559 , n48518 , n48529 );
and ( n48560 , n48559 , n48541 );
and ( n48561 , n48518 , n48529 );
or ( n48562 , n48560 , n48561 );
xor ( n48563 , n48247 , n48285 );
and ( n48564 , n48563 , n48433 );
and ( n48565 , n48247 , n48285 );
or ( n48566 , n48564 , n48565 );
xor ( n48567 , n48481 , n48493 );
and ( n48568 , n48567 , n48503 );
and ( n48569 , n48481 , n48493 );
or ( n48570 , n48568 , n48569 );
xor ( n48571 , n48343 , n48315 );
and ( n48572 , n48571 , n48542 );
and ( n48573 , n48343 , n48315 );
or ( n48574 , n48572 , n48573 );
xor ( n48575 , n48439 , n48349 );
and ( n48576 , n48575 , n48504 );
and ( n48577 , n48439 , n48349 );
or ( n48578 , n48576 , n48577 );
xor ( n48579 , n48543 , n48355 );
and ( n48580 , n48579 , n48361 );
and ( n48581 , n48543 , n48355 );
or ( n48582 , n48580 , n48581 );
not ( n48583 , n48419 );
not ( n48584 , n47300 );
or ( n48585 , n48583 , n48584 );
not ( n48586 , n47765 );
not ( n48587 , n47107 );
or ( n48588 , n48586 , n48587 );
not ( n48589 , n47765 );
nand ( n48590 , n47108 , n48589 );
nand ( n48591 , n48588 , n48590 );
nand ( n48592 , n48591 , n47148 );
nand ( n48593 , n48585 , n48592 );
not ( n48594 , n47384 );
not ( n48595 , n47980 );
not ( n48596 , n46880 );
or ( n48597 , n48595 , n48596 );
nand ( n48598 , n47979 , n47158 );
nand ( n48599 , n48597 , n48598 );
not ( n48600 , n48599 );
or ( n48601 , n48594 , n48600 );
nand ( n48602 , n48403 , n46408 );
nand ( n48603 , n48601 , n48602 );
xor ( n48604 , n48593 , n48603 );
not ( n48605 , n48430 );
not ( n48606 , n47489 );
or ( n48607 , n48605 , n48606 );
not ( n48608 , n47740 );
not ( n48609 , n47493 );
or ( n48610 , n48608 , n48609 );
not ( n48611 , n47473 );
nand ( n48612 , n48611 , n47368 );
nand ( n48613 , n48610 , n48612 );
nand ( n48614 , n48613 , n47498 );
nand ( n48615 , n48607 , n48614 );
xor ( n48616 , n48604 , n48615 );
xor ( n48617 , n48593 , n48603 );
and ( n48618 , n48617 , n48615 );
and ( n48619 , n48593 , n48603 );
or ( n48620 , n48618 , n48619 );
not ( n48621 , n48448 );
not ( n48622 , n47872 );
or ( n48623 , n48621 , n48622 );
not ( n48624 , n47047 );
not ( n48625 , n47854 );
or ( n48626 , n48624 , n48625 );
nand ( n48627 , n47794 , n47821 );
nand ( n48628 , n48626 , n48627 );
nand ( n48629 , n48628 , n48240 );
nand ( n48630 , n48623 , n48629 );
not ( n48631 , n48460 );
not ( n48632 , n48268 );
or ( n48633 , n48631 , n48632 );
not ( n48634 , n46273 );
not ( n48635 , n48202 );
or ( n48636 , n48634 , n48635 );
nand ( n48637 , n48201 , n46824 );
nand ( n48638 , n48636 , n48637 );
nand ( n48639 , n48638 , n48452 );
nand ( n48640 , n48633 , n48639 );
xor ( n48641 , n48630 , n48640 );
not ( n48642 , n46854 );
not ( n48643 , n48171 );
not ( n48644 , n48643 );
buf ( n48645 , n47378 );
not ( n48646 , n48645 );
not ( n48647 , n48646 );
or ( n48648 , n48644 , n48647 );
nand ( n48649 , n48645 , n48171 );
nand ( n48650 , n48648 , n48649 );
not ( n48651 , n48650 );
or ( n48652 , n48642 , n48651 );
not ( n48653 , n47240 );
nand ( n48654 , n48653 , n48381 );
nand ( n48655 , n48652 , n48654 );
not ( n48656 , n46439 );
not ( n48657 , n48656 );
not ( n48658 , n47962 );
not ( n48659 , n41938 );
or ( n48660 , n48658 , n48659 );
not ( n48661 , n47962 );
nand ( n48662 , n41939 , n48661 );
nand ( n48663 , n48660 , n48662 );
not ( n48664 , n48663 );
or ( n48665 , n48657 , n48664 );
nand ( n48666 , n48390 , n46584 );
nand ( n48667 , n48665 , n48666 );
xor ( n48668 , n48655 , n48667 );
xor ( n48669 , n48641 , n48668 );
xor ( n48670 , n48630 , n48640 );
and ( n48671 , n48670 , n48668 );
and ( n48672 , n48630 , n48640 );
or ( n48673 , n48671 , n48672 );
xor ( n48674 , n48616 , n48558 );
xor ( n48675 , n48674 , n48669 );
xor ( n48676 , n48675 , n48570 );
not ( n48677 , n44004 );
not ( n48678 , n46072 );
not ( n48679 , n41363 );
not ( n48680 , n48679 );
or ( n48681 , n48678 , n48680 );
nand ( n48682 , n41364 , n46071 );
nand ( n48683 , n48681 , n48682 );
not ( n48684 , n48683 );
or ( n48685 , n48677 , n48684 );
nand ( n48686 , n48488 , n46474 );
nand ( n48687 , n48685 , n48686 );
xor ( n48688 , n48687 , n48562 );
not ( n48689 , n46441 );
and ( n48690 , n48473 , n48689 );
nor ( n48691 , n48690 , n48456 );
nor ( n48692 , n48473 , n46440 );
or ( n48693 , n48691 , n48692 );
not ( n48694 , n37640 );
buf ( n48695 , n36239 );
nand ( n48696 , n37458 , n36989 , n48695 );
not ( n48697 , n48696 );
or ( n48698 , n48694 , n48697 );
not ( n48699 , n48695 );
nor ( n48700 , n48699 , n37640 );
nand ( n48701 , n37458 , n36989 , n48700 );
nand ( n48702 , n48698 , n48701 );
not ( n48703 , n48702 );
buf ( n48704 , n48703 );
not ( n48705 , n48704 );
nand ( n48706 , n48693 , n48705 );
not ( n48707 , n48706 );
xor ( n48708 , n48707 , n48410 );
not ( n48709 , n48073 );
not ( n48710 , n46650 );
not ( n48711 , n47524 );
or ( n48712 , n48710 , n48711 );
nand ( n48713 , n30929 , n48078 );
nand ( n48714 , n48712 , n48713 );
not ( n48715 , n48714 );
or ( n48716 , n48709 , n48715 );
nand ( n48717 , n48527 , n46776 );
nand ( n48718 , n48716 , n48717 );
xor ( n48719 , n48708 , n48718 );
xor ( n48720 , n48688 , n48719 );
xor ( n48721 , n48676 , n48720 );
xor ( n48722 , n48721 , n48582 );
not ( n48723 , n46153 );
not ( n48724 , n48023 );
not ( n48725 , n47510 );
or ( n48726 , n48724 , n48725 );
not ( n48727 , n47803 );
nand ( n48728 , n41692 , n48727 );
nand ( n48729 , n48726 , n48728 );
not ( n48730 , n48729 );
or ( n48731 , n48723 , n48730 );
nand ( n48732 , n48497 , n47407 );
nand ( n48733 , n48731 , n48732 );
not ( n48734 , n46188 );
not ( n48735 , n46425 );
not ( n48736 , n41575 );
not ( n48737 , n48736 );
or ( n48738 , n48735 , n48737 );
not ( n48739 , n48318 );
nand ( n48740 , n48739 , n46422 );
nand ( n48741 , n48738 , n48740 );
not ( n48742 , n48741 );
or ( n48743 , n48734 , n48742 );
nand ( n48744 , n48539 , n46267 );
nand ( n48745 , n48743 , n48744 );
xor ( n48746 , n48733 , n48745 );
not ( n48747 , n48473 );
buf ( n48748 , n48702 );
not ( n48749 , n48748 );
not ( n48750 , n48749 );
or ( n48751 , n48747 , n48750 );
nand ( n48752 , n48748 , n48472 );
nand ( n48753 , n48751 , n48752 );
nand ( n48754 , n48753 , n48478 );
not ( n48755 , n48754 );
not ( n48756 , n48755 );
not ( n48757 , n48748 );
not ( n48758 , n48757 );
and ( n48759 , n48758 , n46441 );
not ( n48760 , n48758 );
and ( n48761 , n48760 , n46440 );
nor ( n48762 , n48759 , n48761 );
or ( n48763 , n48756 , n48762 );
not ( n48764 , n48757 );
not ( n48765 , n48764 );
buf ( n48766 , n45767 );
not ( n48767 , n48766 );
and ( n48768 , n48765 , n48767 );
and ( n48769 , n48705 , n45767 );
nor ( n48770 , n48768 , n48769 );
or ( n48771 , n48770 , n48479 );
nand ( n48772 , n48763 , n48771 );
xor ( n48773 , n48746 , n48772 );
xor ( n48774 , n48773 , n48566 );
not ( n48775 , n45832 );
not ( n48776 , n46554 );
not ( n48777 , n41530 );
or ( n48778 , n48776 , n48777 );
not ( n48779 , n41530 );
nand ( n48780 , n48779 , n46559 );
nand ( n48781 , n48778 , n48780 );
not ( n48782 , n48781 );
or ( n48783 , n48775 , n48782 );
nand ( n48784 , n48514 , n46448 );
nand ( n48785 , n48783 , n48784 );
xor ( n48786 , n48785 , n48437 );
xor ( n48787 , n48786 , n48554 );
xor ( n48788 , n48774 , n48787 );
xor ( n48789 , n48574 , n48788 );
xor ( n48790 , n48789 , n48578 );
xor ( n48791 , n48722 , n48790 );
xor ( n48792 , n48721 , n48582 );
and ( n48793 , n48792 , n48790 );
and ( n48794 , n48721 , n48582 );
or ( n48795 , n48793 , n48794 );
xor ( n48796 , n48707 , n48410 );
and ( n48797 , n48796 , n48718 );
and ( n48798 , n48707 , n48410 );
or ( n48799 , n48797 , n48798 );
xor ( n48800 , n48733 , n48745 );
and ( n48801 , n48800 , n48772 );
and ( n48802 , n48733 , n48745 );
or ( n48803 , n48801 , n48802 );
xor ( n48804 , n48785 , n48437 );
and ( n48805 , n48804 , n48554 );
and ( n48806 , n48785 , n48437 );
or ( n48807 , n48805 , n48806 );
xor ( n48808 , n48616 , n48558 );
and ( n48809 , n48808 , n48669 );
and ( n48810 , n48616 , n48558 );
or ( n48811 , n48809 , n48810 );
xor ( n48812 , n48687 , n48562 );
and ( n48813 , n48812 , n48719 );
and ( n48814 , n48687 , n48562 );
or ( n48815 , n48813 , n48814 );
xor ( n48816 , n48773 , n48566 );
and ( n48817 , n48816 , n48787 );
and ( n48818 , n48773 , n48566 );
or ( n48819 , n48817 , n48818 );
xor ( n48820 , n48675 , n48570 );
and ( n48821 , n48820 , n48720 );
and ( n48822 , n48675 , n48570 );
or ( n48823 , n48821 , n48822 );
xor ( n48824 , n48574 , n48788 );
and ( n48825 , n48824 , n48578 );
and ( n48826 , n48574 , n48788 );
or ( n48827 , n48825 , n48826 );
not ( n48828 , n46854 );
not ( n48829 , n30259 );
and ( n48830 , n47744 , n48829 );
not ( n48831 , n47744 );
not ( n48832 , n48829 );
and ( n48833 , n48831 , n48832 );
or ( n48834 , n48830 , n48833 );
not ( n48835 , n48834 );
or ( n48836 , n48828 , n48835 );
nand ( n48837 , n47583 , n48650 );
nand ( n48838 , n48836 , n48837 );
not ( n48839 , n46584 );
not ( n48840 , n48663 );
or ( n48841 , n48839 , n48840 );
not ( n48842 , n46994 );
not ( n48843 , n48842 );
not ( n48844 , n46821 );
and ( n48845 , n48843 , n48844 );
and ( n48846 , n47617 , n48661 );
nor ( n48847 , n48845 , n48846 );
not ( n48848 , n48847 );
nand ( n48849 , n48848 , n48656 );
nand ( n48850 , n48841 , n48849 );
xor ( n48851 , n48838 , n48850 );
not ( n48852 , n48591 );
not ( n48853 , n47300 );
or ( n48854 , n48852 , n48853 );
not ( n48855 , n47958 );
buf ( n48856 , n47108 );
not ( n48857 , n48856 );
not ( n48858 , n48857 );
or ( n48859 , n48855 , n48858 );
not ( n48860 , n47958 );
nand ( n48861 , n48856 , n48860 );
nand ( n48862 , n48859 , n48861 );
nand ( n48863 , n48862 , n47148 );
nand ( n48864 , n48854 , n48863 );
xor ( n48865 , n48851 , n48864 );
xor ( n48866 , n48838 , n48850 );
and ( n48867 , n48866 , n48864 );
and ( n48868 , n48838 , n48850 );
or ( n48869 , n48867 , n48868 );
not ( n48870 , n37673 );
not ( n48871 , n48870 );
not ( n48872 , n36986 );
buf ( n48873 , n35565 );
nand ( n48874 , n48872 , n36625 , n48873 );
not ( n48875 , n36614 );
nand ( n48876 , n48875 , n48873 );
not ( n48877 , n36960 );
nand ( n48878 , n48874 , n48876 , n48877 );
not ( n48879 , n48878 );
or ( n48880 , n48871 , n48879 );
nand ( n48881 , n48874 , n48876 , n48877 , n37673 );
nand ( n48882 , n48880 , n48881 );
not ( n48883 , n48882 );
and ( n48884 , n48883 , n48703 );
not ( n48885 , n48883 );
not ( n48886 , n48702 );
not ( n48887 , n48886 );
and ( n48888 , n48885 , n48887 );
nor ( n48889 , n48884 , n48888 );
buf ( n48890 , n48889 );
not ( n48891 , n48890 );
and ( n48892 , n48891 , n46440 );
not ( n48893 , n48613 );
buf ( n48894 , n47489 );
not ( n48895 , n48894 );
or ( n48896 , n48893 , n48895 );
buf ( n48897 , n47575 );
not ( n48898 , n48897 );
and ( n48899 , n48898 , n47476 );
not ( n48900 , n48898 );
and ( n48901 , n48900 , n47473 );
nor ( n48902 , n48899 , n48901 );
nand ( n48903 , n47498 , n48902 );
nand ( n48904 , n48896 , n48903 );
xor ( n48905 , n48892 , n48904 );
not ( n48906 , n48628 );
not ( n48907 , n47873 );
or ( n48908 , n48906 , n48907 );
nand ( n48909 , n47794 , n47589 );
nand ( n48910 , n47227 , n47795 );
nand ( n48911 , n48909 , n48910 );
nand ( n48912 , n48240 , n48911 );
nand ( n48913 , n48908 , n48912 );
xor ( n48914 , n48905 , n48913 );
xor ( n48915 , n48892 , n48904 );
and ( n48916 , n48915 , n48913 );
and ( n48917 , n48892 , n48904 );
or ( n48918 , n48916 , n48917 );
not ( n48919 , n46776 );
not ( n48920 , n48714 );
or ( n48921 , n48919 , n48920 );
not ( n48922 , n46650 );
not ( n48923 , n41416 );
or ( n48924 , n48922 , n48923 );
nand ( n48925 , n41415 , n48078 );
nand ( n48926 , n48924 , n48925 );
nand ( n48927 , n48926 , n47827 );
nand ( n48928 , n48921 , n48927 );
buf ( n48929 , n46153 );
not ( n48930 , n48929 );
not ( n48931 , n48023 );
not ( n48932 , n48523 );
or ( n48933 , n48931 , n48932 );
nand ( n48934 , n41683 , n48727 );
nand ( n48935 , n48933 , n48934 );
not ( n48936 , n48935 );
or ( n48937 , n48930 , n48936 );
nand ( n48938 , n48729 , n47407 );
nand ( n48939 , n48937 , n48938 );
xor ( n48940 , n48928 , n48939 );
xor ( n48941 , n48940 , n48865 );
xor ( n48942 , n48941 , n48811 );
xor ( n48943 , n48942 , n48815 );
xor ( n48944 , n48819 , n48943 );
xor ( n48945 , n48944 , n48823 );
xor ( n48946 , n48819 , n48943 );
and ( n48947 , n48946 , n48823 );
and ( n48948 , n48819 , n48943 );
or ( n48949 , n48947 , n48948 );
not ( n48950 , n45748 );
not ( n48951 , n41407 );
buf ( n48952 , n45750 );
and ( n48953 , n48951 , n48952 );
not ( n48954 , n48951 );
buf ( n48955 , n45837 );
and ( n48956 , n48954 , n48955 );
or ( n48957 , n48953 , n48956 );
not ( n48958 , n48957 );
or ( n48959 , n48950 , n48958 );
nand ( n48960 , n48781 , n46564 );
nand ( n48961 , n48959 , n48960 );
xor ( n48962 , n48673 , n48961 );
not ( n48963 , n48638 );
not ( n48964 , n48463 );
or ( n48965 , n48963 , n48964 );
not ( n48966 , n47646 );
not ( n48967 , n48456 );
not ( n48968 , n48967 );
or ( n48969 , n48966 , n48968 );
not ( n48970 , n48201 );
not ( n48971 , n48970 );
nand ( n48972 , n48971 , n47650 );
nand ( n48973 , n48969 , n48972 );
nand ( n48974 , n48973 , n48452 );
nand ( n48975 , n48965 , n48974 );
and ( n48976 , n48655 , n48667 );
xor ( n48977 , n48975 , n48976 );
not ( n48978 , n47384 );
not ( n48979 , n47980 );
not ( n48980 , n30964 );
not ( n48981 , n48980 );
or ( n48982 , n48979 , n48981 );
buf ( n48983 , n30964 );
nand ( n48984 , n48983 , n47979 );
nand ( n48985 , n48982 , n48984 );
not ( n48986 , n48985 );
or ( n48987 , n48978 , n48986 );
not ( n48988 , n46408 );
not ( n48989 , n48988 );
nand ( n48990 , n48599 , n48989 );
nand ( n48991 , n48987 , n48990 );
xor ( n48992 , n48977 , n48991 );
xor ( n48993 , n48962 , n48992 );
not ( n48994 , n46602 );
not ( n48995 , n46072 );
not ( n48996 , n41284 );
not ( n48997 , n48996 );
not ( n48998 , n48997 );
or ( n48999 , n48995 , n48998 );
not ( n49000 , n41283 );
buf ( n49001 , n49000 );
nand ( n49002 , n49001 , n46071 );
nand ( n49003 , n48999 , n49002 );
not ( n49004 , n49003 );
or ( n49005 , n48994 , n49004 );
nand ( n49006 , n48683 , n46474 );
nand ( n49007 , n49005 , n49006 );
xor ( n49008 , n48914 , n49007 );
xor ( n49009 , n49008 , n48799 );
xor ( n49010 , n48993 , n49009 );
xor ( n49011 , n48803 , n48807 );
not ( n49012 , n48770 );
not ( n49013 , n49012 );
not ( n49014 , n48754 );
not ( n49015 , n49014 );
or ( n49016 , n49013 , n49015 );
not ( n49017 , n48749 );
and ( n49018 , n46037 , n49017 );
not ( n49019 , n46037 );
and ( n49020 , n49019 , n48704 );
nor ( n49021 , n49018 , n49020 );
not ( n49022 , n48479 );
nand ( n49023 , n49021 , n49022 );
nand ( n49024 , n49016 , n49023 );
buf ( n49025 , n45811 );
not ( n49026 , n49025 );
not ( n49027 , n49026 );
not ( n49028 , n46425 );
not ( n49029 , n44141 );
not ( n49030 , n49029 );
or ( n49031 , n49028 , n49030 );
nand ( n49032 , n44141 , n46422 );
nand ( n49033 , n49031 , n49032 );
not ( n49034 , n49033 );
or ( n49035 , n49027 , n49034 );
nand ( n49036 , n48741 , n46267 );
nand ( n49037 , n49035 , n49036 );
xor ( n49038 , n49024 , n49037 );
xor ( n49039 , n49038 , n48620 );
xor ( n49040 , n49011 , n49039 );
xor ( n49041 , n49010 , n49040 );
xor ( n49042 , n49041 , n48827 );
xor ( n49043 , n49042 , n48945 );
xor ( n49044 , n49041 , n48827 );
and ( n49045 , n49044 , n48945 );
and ( n49046 , n49041 , n48827 );
or ( n49047 , n49045 , n49046 );
xor ( n49048 , n48975 , n48976 );
and ( n49049 , n49048 , n48991 );
and ( n49050 , n48975 , n48976 );
or ( n49051 , n49049 , n49050 );
xor ( n49052 , n48928 , n48939 );
and ( n49053 , n49052 , n48865 );
and ( n49054 , n48928 , n48939 );
or ( n49055 , n49053 , n49054 );
xor ( n49056 , n49024 , n49037 );
and ( n49057 , n49056 , n48620 );
and ( n49058 , n49024 , n49037 );
or ( n49059 , n49057 , n49058 );
xor ( n49060 , n48673 , n48961 );
and ( n49061 , n49060 , n48992 );
and ( n49062 , n48673 , n48961 );
or ( n49063 , n49061 , n49062 );
xor ( n49064 , n48914 , n49007 );
and ( n49065 , n49064 , n48799 );
and ( n49066 , n48914 , n49007 );
or ( n49067 , n49065 , n49066 );
xor ( n49068 , n48803 , n48807 );
and ( n49069 , n49068 , n49039 );
and ( n49070 , n48803 , n48807 );
or ( n49071 , n49069 , n49070 );
xor ( n49072 , n48941 , n48811 );
and ( n49073 , n49072 , n48815 );
and ( n49074 , n48941 , n48811 );
or ( n49075 , n49073 , n49074 );
xor ( n49076 , n48993 , n49009 );
and ( n49077 , n49076 , n49040 );
and ( n49078 , n48993 , n49009 );
or ( n49079 , n49077 , n49078 );
not ( n49080 , n48862 );
not ( n49081 , n47300 );
or ( n49082 , n49080 , n49081 );
not ( n49083 , n48643 );
not ( n49084 , n47107 );
or ( n49085 , n49083 , n49084 );
nand ( n49086 , n47106 , n48171 );
nand ( n49087 , n49085 , n49086 );
nand ( n49088 , n49087 , n47148 );
nand ( n49089 , n49082 , n49088 );
nand ( n49090 , n48883 , n46440 );
not ( n49091 , n49090 );
buf ( n49092 , n48886 );
not ( n49093 , n49092 );
not ( n49094 , n49093 );
not ( n49095 , n49094 );
or ( n49096 , n49091 , n49095 );
not ( n49097 , n48883 );
nand ( n49098 , n49097 , n46441 );
nand ( n49099 , n49096 , n49098 );
buf ( n49100 , n36256 );
nand ( n49101 , n49100 , n36259 );
not ( n49102 , n49101 );
not ( n49103 , n49102 );
not ( n49104 , n36964 );
not ( n49105 , n49104 );
or ( n49106 , n49103 , n49105 );
nand ( n49107 , n36964 , n49101 );
nand ( n49108 , n49106 , n49107 );
buf ( n49109 , n49108 );
not ( n49110 , n49109 );
not ( n49111 , n49110 );
buf ( n49112 , n49111 );
and ( n49113 , n49099 , n49112 );
xor ( n49114 , n49089 , n49113 );
not ( n49115 , n48902 );
not ( n49116 , n47488 );
not ( n49117 , n49116 );
or ( n49118 , n49115 , n49117 );
and ( n49119 , n47493 , n47765 );
not ( n49120 , n47493 );
and ( n49121 , n49120 , n48589 );
or ( n49122 , n49119 , n49121 );
nand ( n49123 , n47498 , n49122 );
nand ( n49124 , n49118 , n49123 );
xor ( n49125 , n49114 , n49124 );
xor ( n49126 , n49089 , n49113 );
and ( n49127 , n49126 , n49124 );
and ( n49128 , n49089 , n49113 );
or ( n49129 , n49127 , n49128 );
not ( n49130 , n48911 );
not ( n49131 , n47872 );
or ( n49132 , n49130 , n49131 );
not ( n49133 , n47740 );
not ( n49134 , n48235 );
or ( n49135 , n49133 , n49134 );
nand ( n49136 , n47794 , n47368 );
nand ( n49137 , n49135 , n49136 );
nand ( n49138 , n49137 , n47881 );
nand ( n49139 , n49132 , n49138 );
not ( n49140 , n48973 );
not ( n49141 , n48463 );
or ( n49142 , n49140 , n49141 );
not ( n49143 , n47047 );
not ( n49144 , n48202 );
or ( n49145 , n49143 , n49144 );
nand ( n49146 , n48201 , n47821 );
nand ( n49147 , n49145 , n49146 );
buf ( n49148 , n48017 );
nand ( n49149 , n49147 , n49148 );
nand ( n49150 , n49142 , n49149 );
xor ( n49151 , n49139 , n49150 );
not ( n49152 , n46854 );
not ( n49153 , n46607 );
not ( n49154 , n46835 );
and ( n49155 , n49153 , n49154 );
and ( n49156 , n41938 , n47744 );
nor ( n49157 , n49155 , n49156 );
not ( n49158 , n49157 );
not ( n49159 , n49158 );
or ( n49160 , n49152 , n49159 );
nand ( n49161 , n48834 , n47583 );
nand ( n49162 , n49160 , n49161 );
not ( n49163 , n49162 );
not ( n49164 , n49163 );
not ( n49165 , n47962 );
not ( n49166 , n46880 );
or ( n49167 , n49165 , n49166 );
nand ( n49168 , n47158 , n46821 );
nand ( n49169 , n49167 , n49168 );
and ( n49170 , n49169 , n48656 );
not ( n49171 , n46584 );
nor ( n49172 , n49171 , n48847 );
nor ( n49173 , n49170 , n49172 );
not ( n49174 , n49173 );
not ( n49175 , n49174 );
or ( n49176 , n49164 , n49175 );
or ( n49177 , n49163 , n49174 );
nand ( n49178 , n49176 , n49177 );
xor ( n49179 , n49151 , n49178 );
xor ( n49180 , n49139 , n49150 );
and ( n49181 , n49180 , n49178 );
and ( n49182 , n49139 , n49150 );
or ( n49183 , n49181 , n49182 );
xor ( n49184 , n49063 , n49067 );
xor ( n49185 , n49051 , n49179 );
not ( n49186 , n46564 );
not ( n49187 , n48957 );
or ( n49188 , n49186 , n49187 );
not ( n49189 , n48952 );
not ( n49190 , n41363 );
not ( n49191 , n49190 );
or ( n49192 , n49189 , n49191 );
nand ( n49193 , n41363 , n48955 );
nand ( n49194 , n49192 , n49193 );
nand ( n49195 , n49194 , n45748 );
nand ( n49196 , n49188 , n49195 );
xor ( n49197 , n49185 , n49196 );
xor ( n49198 , n49184 , n49197 );
xor ( n49199 , n49075 , n49198 );
xor ( n49200 , n49199 , n49079 );
xor ( n49201 , n49075 , n49198 );
and ( n49202 , n49201 , n49079 );
and ( n49203 , n49075 , n49198 );
or ( n49204 , n49202 , n49203 );
not ( n49205 , n46474 );
not ( n49206 , n49003 );
or ( n49207 , n49205 , n49206 );
not ( n49208 , n46072 );
not ( n49209 , n41216 );
not ( n49210 , n49209 );
not ( n49211 , n49210 );
or ( n49212 , n49208 , n49211 );
nand ( n49213 , n49209 , n46071 );
nand ( n49214 , n49212 , n49213 );
nand ( n49215 , n49214 , n46602 );
nand ( n49216 , n49207 , n49215 );
xor ( n49217 , n49055 , n49216 );
not ( n49218 , n48929 );
not ( n49219 , n48023 );
not ( n49220 , n30929 );
not ( n49221 , n49220 );
or ( n49222 , n49219 , n49221 );
nand ( n49223 , n30929 , n48727 );
nand ( n49224 , n49222 , n49223 );
not ( n49225 , n49224 );
or ( n49226 , n49218 , n49225 );
nand ( n49227 , n48935 , n47407 );
nand ( n49228 , n49226 , n49227 );
not ( n49229 , n46188 );
not ( n49230 , n46425 );
not ( n49231 , n41529 );
buf ( n49232 , n49231 );
not ( n49233 , n49232 );
not ( n49234 , n49233 );
or ( n49235 , n49230 , n49234 );
nand ( n49236 , n48306 , n46422 );
nand ( n49237 , n49235 , n49236 );
not ( n49238 , n49237 );
or ( n49239 , n49229 , n49238 );
nand ( n49240 , n49033 , n46267 );
nand ( n49241 , n49239 , n49240 );
xor ( n49242 , n49228 , n49241 );
not ( n49243 , n47384 );
not ( n49244 , n47980 );
not ( n49245 , n47918 );
not ( n49246 , n49245 );
or ( n49247 , n49244 , n49246 );
nand ( n49248 , n47918 , n47979 );
nand ( n49249 , n49247 , n49248 );
not ( n49250 , n49249 );
or ( n49251 , n49243 , n49250 );
not ( n49252 , n48988 );
nand ( n49253 , n48985 , n49252 );
nand ( n49254 , n49251 , n49253 );
xor ( n49255 , n49242 , n49254 );
xor ( n49256 , n49217 , n49255 );
xor ( n49257 , n49071 , n49256 );
not ( n49258 , n49108 );
buf ( n49259 , n49258 );
and ( n49260 , n46441 , n49259 );
not ( n49261 , n46441 );
buf ( n49262 , n49109 );
and ( n49263 , n49261 , n49262 );
nor ( n49264 , n49260 , n49263 );
not ( n49265 , n49264 );
not ( n49266 , n49102 );
not ( n49267 , n49104 );
or ( n49268 , n49266 , n49267 );
nand ( n49269 , n49268 , n49107 );
and ( n49270 , n48883 , n49269 );
not ( n49271 , n48883 );
and ( n49272 , n49271 , n49258 );
nor ( n49273 , n49270 , n49272 );
nand ( n49274 , n48889 , n49273 );
buf ( n49275 , n49274 );
not ( n49276 , n49275 );
not ( n49277 , n49276 );
or ( n49278 , n49265 , n49277 );
and ( n49279 , n45816 , n49259 );
not ( n49280 , n45816 );
buf ( n49281 , n49269 );
not ( n49282 , n49281 );
buf ( n49283 , n49282 );
not ( n49284 , n49283 );
and ( n49285 , n49280 , n49284 );
nor ( n49286 , n49279 , n49285 );
not ( n49287 , n49286 );
not ( n49288 , n48890 );
nand ( n49289 , n49287 , n49288 );
nand ( n49290 , n49278 , n49289 );
xor ( n49291 , n49290 , n48869 );
not ( n49292 , n45896 );
not ( n49293 , n48736 );
not ( n49294 , n49293 );
not ( n49295 , n48078 );
and ( n49296 , n49294 , n49295 );
not ( n49297 , n41575 );
not ( n49298 , n49297 );
and ( n49299 , n49298 , n48290 );
nor ( n49300 , n49296 , n49299 );
not ( n49301 , n49300 );
not ( n49302 , n49301 );
or ( n49303 , n49292 , n49302 );
nand ( n49304 , n48926 , n48295 );
nand ( n49305 , n49303 , n49304 );
xor ( n49306 , n49291 , n49305 );
xor ( n49307 , n49059 , n49306 );
not ( n49308 , n49021 );
not ( n49309 , n48756 );
not ( n49310 , n49309 );
or ( n49311 , n49308 , n49310 );
not ( n49312 , n46273 );
not ( n49313 , n48757 );
not ( n49314 , n49313 );
not ( n49315 , n49314 );
or ( n49316 , n49312 , n49315 );
not ( n49317 , n48704 );
nand ( n49318 , n49317 , n46824 );
nand ( n49319 , n49316 , n49318 );
not ( n49320 , n48478 );
nand ( n49321 , n49319 , n49320 );
nand ( n49322 , n49311 , n49321 );
xor ( n49323 , n49322 , n48918 );
xor ( n49324 , n49323 , n49125 );
xor ( n49325 , n49307 , n49324 );
xor ( n49326 , n49257 , n49325 );
xor ( n49327 , n49326 , n48949 );
xor ( n49328 , n49327 , n49200 );
xor ( n49329 , n49326 , n48949 );
and ( n49330 , n49329 , n49200 );
and ( n49331 , n49326 , n48949 );
or ( n49332 , n49330 , n49331 );
xor ( n49333 , n49290 , n48869 );
and ( n49334 , n49333 , n49305 );
and ( n49335 , n49290 , n48869 );
or ( n49336 , n49334 , n49335 );
xor ( n49337 , n49228 , n49241 );
and ( n49338 , n49337 , n49254 );
and ( n49339 , n49228 , n49241 );
or ( n49340 , n49338 , n49339 );
xor ( n49341 , n49322 , n48918 );
and ( n49342 , n49341 , n49125 );
and ( n49343 , n49322 , n48918 );
or ( n49344 , n49342 , n49343 );
xor ( n49345 , n49051 , n49179 );
and ( n49346 , n49345 , n49196 );
and ( n49347 , n49051 , n49179 );
or ( n49348 , n49346 , n49347 );
xor ( n49349 , n49055 , n49216 );
and ( n49350 , n49349 , n49255 );
and ( n49351 , n49055 , n49216 );
or ( n49352 , n49350 , n49351 );
xor ( n49353 , n49059 , n49306 );
and ( n49354 , n49353 , n49324 );
and ( n49355 , n49059 , n49306 );
or ( n49356 , n49354 , n49355 );
xor ( n49357 , n49063 , n49067 );
and ( n49358 , n49357 , n49197 );
and ( n49359 , n49063 , n49067 );
or ( n49360 , n49358 , n49359 );
xor ( n49361 , n49071 , n49256 );
and ( n49362 , n49361 , n49325 );
and ( n49363 , n49071 , n49256 );
or ( n49364 , n49362 , n49363 );
not ( n49365 , n47060 );
and ( n49366 , n41861 , n47094 );
not ( n49367 , n41861 );
and ( n49368 , n49367 , n47378 );
or ( n49369 , n49366 , n49368 );
not ( n49370 , n49369 );
or ( n49371 , n49365 , n49370 );
not ( n49372 , n47241 );
or ( n49373 , n49157 , n49372 );
nand ( n49374 , n49371 , n49373 );
not ( n49375 , n49087 );
not ( n49376 , n47139 );
or ( n49377 , n49375 , n49376 );
and ( n49378 , n30259 , n47276 );
not ( n49379 , n30259 );
and ( n49380 , n49379 , n47449 );
or ( n49381 , n49378 , n49380 );
nand ( n49382 , n49381 , n47147 );
nand ( n49383 , n49377 , n49382 );
xor ( n49384 , n49374 , n49383 );
not ( n49385 , n46440 );
and ( n49386 , n49108 , n36637 );
not ( n49387 , n49108 );
not ( n49388 , n36637 );
and ( n49389 , n49387 , n49388 );
nor ( n49390 , n49386 , n49389 );
not ( n49391 , n49390 );
nor ( n49392 , n49385 , n49391 );
xor ( n49393 , n49384 , n49392 );
xor ( n49394 , n49374 , n49383 );
and ( n49395 , n49394 , n49392 );
and ( n49396 , n49374 , n49383 );
or ( n49397 , n49395 , n49396 );
not ( n49398 , n49122 );
not ( n49399 , n47489 );
or ( n49400 , n49398 , n49399 );
not ( n49401 , n47958 );
not ( n49402 , n47473 );
or ( n49403 , n49401 , n49402 );
nand ( n49404 , n47476 , n48860 );
nand ( n49405 , n49403 , n49404 );
nand ( n49406 , n47498 , n49405 );
nand ( n49407 , n49400 , n49406 );
not ( n49408 , n49137 );
not ( n49409 , n47873 );
or ( n49410 , n49408 , n49409 );
not ( n49411 , n48898 );
not ( n49412 , n47854 );
or ( n49413 , n49411 , n49412 );
nand ( n49414 , n47794 , n48897 );
nand ( n49415 , n49413 , n49414 );
nand ( n49416 , n49415 , n47881 );
nand ( n49417 , n49410 , n49416 );
xor ( n49418 , n49407 , n49417 );
not ( n49419 , n49147 );
not ( n49420 , n48463 );
not ( n49421 , n49420 );
not ( n49422 , n49421 );
or ( n49423 , n49419 , n49422 );
not ( n49424 , n47227 );
not ( n49425 , n48455 );
or ( n49426 , n49424 , n49425 );
nand ( n49427 , n48456 , n47589 );
nand ( n49428 , n49426 , n49427 );
nand ( n49429 , n49428 , n48452 );
nand ( n49430 , n49423 , n49429 );
xor ( n49431 , n49418 , n49430 );
xor ( n49432 , n49407 , n49417 );
and ( n49433 , n49432 , n49430 );
and ( n49434 , n49407 , n49417 );
or ( n49435 , n49433 , n49434 );
not ( n49436 , n48656 );
and ( n49437 , n30964 , n46821 );
not ( n49438 , n30964 );
and ( n49439 , n49438 , n47962 );
or ( n49440 , n49437 , n49439 );
not ( n49441 , n49440 );
or ( n49442 , n49436 , n49441 );
nand ( n49443 , n49169 , n46584 );
nand ( n49444 , n49442 , n49443 );
not ( n49445 , n49162 );
nor ( n49446 , n49445 , n49173 );
xor ( n49447 , n49444 , n49446 );
or ( n49448 , n49275 , n49286 );
not ( n49449 , n46037 );
not ( n49450 , n49110 );
or ( n49451 , n49449 , n49450 );
not ( n49452 , n49259 );
nand ( n49453 , n49452 , n47306 );
nand ( n49454 , n49451 , n49453 );
not ( n49455 , n49454 );
or ( n49456 , n49455 , n48890 );
nand ( n49457 , n49448 , n49456 );
xor ( n49458 , n49447 , n49457 );
xor ( n49459 , n49340 , n49458 );
not ( n49460 , n47407 );
not ( n49461 , n49224 );
or ( n49462 , n49460 , n49461 );
not ( n49463 , n47803 );
not ( n49464 , n48535 );
or ( n49465 , n49463 , n49464 );
nand ( n49466 , n41415 , n48727 );
nand ( n49467 , n49465 , n49466 );
nand ( n49468 , n49467 , n48929 );
nand ( n49469 , n49462 , n49468 );
not ( n49470 , n47254 );
not ( n49471 , n46650 );
not ( n49472 , n41667 );
not ( n49473 , n49472 );
or ( n49474 , n49471 , n49473 );
nand ( n49475 , n41667 , n47260 );
nand ( n49476 , n49474 , n49475 );
not ( n49477 , n49476 );
or ( n49478 , n49470 , n49477 );
or ( n49479 , n49300 , n46775 );
nand ( n49480 , n49478 , n49479 );
xor ( n49481 , n49469 , n49480 );
not ( n49482 , n49319 );
not ( n49483 , n49014 );
or ( n49484 , n49482 , n49483 );
not ( n49485 , n49320 );
not ( n49486 , n49485 );
not ( n49487 , n47650 );
not ( n49488 , n48758 );
or ( n49489 , n49487 , n49488 );
nand ( n49490 , n48704 , n47646 );
nand ( n49491 , n49489 , n49490 );
nand ( n49492 , n49486 , n49491 );
nand ( n49493 , n49484 , n49492 );
xor ( n49494 , n49481 , n49493 );
xor ( n49495 , n49459 , n49494 );
xor ( n49496 , n49495 , n49356 );
not ( n49497 , n48989 );
not ( n49498 , n49249 );
or ( n49499 , n49497 , n49498 );
not ( n49500 , n47979 );
not ( n49501 , n49500 );
not ( n49502 , n48523 );
or ( n49503 , n49501 , n49502 );
nand ( n49504 , n41683 , n47979 );
nand ( n49505 , n49503 , n49504 );
nand ( n49506 , n49505 , n47384 );
nand ( n49507 , n49499 , n49506 );
xor ( n49508 , n49507 , n49393 );
xor ( n49509 , n49508 , n49129 );
xor ( n49510 , n49344 , n49509 );
not ( n49511 , n46188 );
not ( n49512 , n46425 );
not ( n49513 , n48951 );
or ( n49514 , n49512 , n49513 );
nand ( n49515 , n48486 , n46422 );
nand ( n49516 , n49514 , n49515 );
not ( n49517 , n49516 );
or ( n49518 , n49511 , n49517 );
nand ( n49519 , n49237 , n46267 );
nand ( n49520 , n49518 , n49519 );
xor ( n49521 , n49183 , n49520 );
xor ( n49522 , n49521 , n49431 );
xor ( n49523 , n49510 , n49522 );
xor ( n49524 , n49496 , n49523 );
xor ( n49525 , n49495 , n49356 );
and ( n49526 , n49525 , n49523 );
and ( n49527 , n49495 , n49356 );
or ( n49528 , n49526 , n49527 );
xor ( n49529 , n49360 , n49364 );
xor ( n49530 , n49348 , n49352 );
not ( n49531 , n45748 );
not ( n49532 , n48952 );
not ( n49533 , n48997 );
or ( n49534 , n49532 , n49533 );
nand ( n49535 , n49001 , n48955 );
nand ( n49536 , n49534 , n49535 );
not ( n49537 , n49536 );
or ( n49538 , n49531 , n49537 );
nand ( n49539 , n49194 , n46564 );
nand ( n49540 , n49538 , n49539 );
not ( n49541 , n46474 );
not ( n49542 , n49214 );
or ( n49543 , n49541 , n49542 );
not ( n49544 , n46072 );
not ( n49545 , n40854 );
not ( n49546 , n49545 );
or ( n49547 , n49544 , n49546 );
not ( n49548 , n40853 );
not ( n49549 , n49548 );
nand ( n49550 , n49549 , n46071 );
nand ( n49551 , n49547 , n49550 );
nand ( n49552 , n49551 , n46602 );
nand ( n49553 , n49543 , n49552 );
xor ( n49554 , n49540 , n49553 );
xor ( n49555 , n49554 , n49336 );
xor ( n49556 , n49530 , n49555 );
xor ( n49557 , n49529 , n49556 );
xor ( n49558 , n49360 , n49364 );
and ( n49559 , n49558 , n49556 );
and ( n49560 , n49360 , n49364 );
or ( n49561 , n49559 , n49560 );
xor ( n49562 , n49524 , n49204 );
xor ( n49563 , n49562 , n49557 );
xor ( n49564 , n49524 , n49204 );
and ( n49565 , n49564 , n49557 );
and ( n49566 , n49524 , n49204 );
or ( n49567 , n49565 , n49566 );
xor ( n49568 , n49444 , n49446 );
and ( n49569 , n49568 , n49457 );
and ( n49570 , n49444 , n49446 );
or ( n49571 , n49569 , n49570 );
xor ( n49572 , n49469 , n49480 );
and ( n49573 , n49572 , n49493 );
and ( n49574 , n49469 , n49480 );
or ( n49575 , n49573 , n49574 );
xor ( n49576 , n49507 , n49393 );
and ( n49577 , n49576 , n49129 );
and ( n49578 , n49507 , n49393 );
or ( n49579 , n49577 , n49578 );
xor ( n49580 , n49183 , n49520 );
and ( n49581 , n49580 , n49431 );
and ( n49582 , n49183 , n49520 );
or ( n49583 , n49581 , n49582 );
xor ( n49584 , n49540 , n49553 );
and ( n49585 , n49584 , n49336 );
and ( n49586 , n49540 , n49553 );
or ( n49587 , n49585 , n49586 );
xor ( n49588 , n49340 , n49458 );
and ( n49589 , n49588 , n49494 );
and ( n49590 , n49340 , n49458 );
or ( n49591 , n49589 , n49590 );
xor ( n49592 , n49344 , n49509 );
and ( n49593 , n49592 , n49522 );
and ( n49594 , n49344 , n49509 );
or ( n49595 , n49593 , n49594 );
xor ( n49596 , n49348 , n49352 );
and ( n49597 , n49596 , n49555 );
and ( n49598 , n49348 , n49352 );
or ( n49599 , n49597 , n49598 );
not ( n49600 , n49388 );
nand ( n49601 , n49600 , n46440 );
not ( n49602 , n49601 );
not ( n49603 , n49259 );
or ( n49604 , n49602 , n49603 );
nand ( n49605 , n49388 , n46441 );
nand ( n49606 , n49604 , n49605 );
not ( n49607 , n37467 );
nand ( n49608 , n49607 , n37459 , n36971 );
buf ( n49609 , n36272 );
buf ( n49610 , n35249 );
nand ( n49611 , n49609 , n49610 );
not ( n49612 , n49611 );
and ( n49613 , n49608 , n49612 );
not ( n49614 , n49608 );
and ( n49615 , n49614 , n49611 );
nor ( n49616 , n49613 , n49615 );
buf ( n49617 , n49616 );
buf ( n49618 , n49617 );
buf ( n49619 , n49618 );
and ( n49620 , n49606 , n49619 );
not ( n49621 , n49405 );
not ( n49622 , n48894 );
or ( n49623 , n49621 , n49622 );
buf ( n49624 , n48643 );
not ( n49625 , n49624 );
not ( n49626 , n47473 );
or ( n49627 , n49625 , n49626 );
buf ( n49628 , n47493 );
not ( n49629 , n49628 );
not ( n49630 , n49624 );
nand ( n49631 , n49629 , n49630 );
nand ( n49632 , n49627 , n49631 );
nand ( n49633 , n47498 , n49632 );
nand ( n49634 , n49623 , n49633 );
xor ( n49635 , n49620 , n49634 );
not ( n49636 , n49415 );
not ( n49637 , n47873 );
or ( n49638 , n49636 , n49637 );
not ( n49639 , n47765 );
not ( n49640 , n47795 );
or ( n49641 , n49639 , n49640 );
nand ( n49642 , n47794 , n48589 );
nand ( n49643 , n49641 , n49642 );
nand ( n49644 , n48240 , n49643 );
nand ( n49645 , n49638 , n49644 );
xor ( n49646 , n49635 , n49645 );
xor ( n49647 , n49620 , n49634 );
and ( n49648 , n49647 , n49645 );
and ( n49649 , n49620 , n49634 );
or ( n49650 , n49648 , n49649 );
not ( n49651 , n49428 );
not ( n49652 , n48463 );
or ( n49653 , n49651 , n49652 );
not ( n49654 , n47368 );
not ( n49655 , n49654 );
not ( n49656 , n48259 );
or ( n49657 , n49655 , n49656 );
not ( n49658 , n48455 );
nand ( n49659 , n49658 , n47368 );
nand ( n49660 , n49657 , n49659 );
nand ( n49661 , n48017 , n49660 );
nand ( n49662 , n49653 , n49661 );
not ( n49663 , n49454 );
not ( n49664 , n49276 );
or ( n49665 , n49663 , n49664 );
not ( n49666 , n46273 );
not ( n49667 , n49110 );
or ( n49668 , n49666 , n49667 );
nand ( n49669 , n49281 , n46824 );
nand ( n49670 , n49668 , n49669 );
nand ( n49671 , n49670 , n48891 );
nand ( n49672 , n49665 , n49671 );
xor ( n49673 , n49662 , n49672 );
not ( n49674 , n46854 );
buf ( n49675 , n47744 );
not ( n49676 , n49675 );
not ( n49677 , n47154 );
or ( n49678 , n49676 , n49677 );
not ( n49679 , n48645 );
nand ( n49680 , n47158 , n49679 );
nand ( n49681 , n49678 , n49680 );
not ( n49682 , n49681 );
or ( n49683 , n49674 , n49682 );
nand ( n49684 , n49369 , n48653 );
nand ( n49685 , n49683 , n49684 );
not ( n49686 , n49381 );
not ( n49687 , n47139 );
or ( n49688 , n49686 , n49687 );
not ( n49689 , n47807 );
not ( n49690 , n47107 );
or ( n49691 , n49689 , n49690 );
not ( n49692 , n47450 );
nand ( n49693 , n49692 , n46607 );
nand ( n49694 , n49691 , n49693 );
nand ( n49695 , n49694 , n47148 );
nand ( n49696 , n49688 , n49695 );
xor ( n49697 , n49685 , n49696 );
xor ( n49698 , n49673 , n49697 );
xor ( n49699 , n49662 , n49672 );
and ( n49700 , n49699 , n49697 );
and ( n49701 , n49662 , n49672 );
or ( n49702 , n49700 , n49701 );
not ( n49703 , n48656 );
not ( n49704 , n47510 );
not ( n49705 , n46820 );
or ( n49706 , n49704 , n49705 );
not ( n49707 , n48661 );
not ( n49708 , n49707 );
nand ( n49709 , n49708 , n47918 );
nand ( n49710 , n49706 , n49709 );
not ( n49711 , n49710 );
or ( n49712 , n49703 , n49711 );
buf ( n49713 , n46584 );
nand ( n49714 , n49440 , n49713 );
nand ( n49715 , n49712 , n49714 );
not ( n49716 , n47384 );
not ( n49717 , n49500 );
not ( n49718 , n49220 );
or ( n49719 , n49717 , n49718 );
nand ( n49720 , n30929 , n47979 );
nand ( n49721 , n49719 , n49720 );
not ( n49722 , n49721 );
or ( n49723 , n49716 , n49722 );
nand ( n49724 , n49505 , n46408 );
nand ( n49725 , n49723 , n49724 );
xor ( n49726 , n49715 , n49725 );
not ( n49727 , n49491 );
not ( n49728 , n49014 );
or ( n49729 , n49727 , n49728 );
not ( n49730 , n47821 );
not ( n49731 , n48758 );
or ( n49732 , n49730 , n49731 );
not ( n49733 , n49093 );
not ( n49734 , n47821 );
nand ( n49735 , n49733 , n49734 );
nand ( n49736 , n49732 , n49735 );
not ( n49737 , n48478 );
nand ( n49738 , n49736 , n49737 );
nand ( n49739 , n49729 , n49738 );
xor ( n49740 , n49726 , n49739 );
not ( n49741 , n47827 );
not ( n49742 , n46650 );
not ( n49743 , n41530 );
or ( n49744 , n49742 , n49743 );
nand ( n49745 , n49231 , n47260 );
nand ( n49746 , n49744 , n49745 );
not ( n49747 , n49746 );
or ( n49748 , n49741 , n49747 );
nand ( n49749 , n49476 , n46776 );
nand ( n49750 , n49748 , n49749 );
xor ( n49751 , n49750 , n49397 );
not ( n49752 , n47407 );
not ( n49753 , n49467 );
or ( n49754 , n49752 , n49753 );
not ( n49755 , n48023 );
not ( n49756 , n41575 );
not ( n49757 , n49756 );
or ( n49758 , n49755 , n49757 );
nand ( n49759 , n49298 , n48727 );
nand ( n49760 , n49758 , n49759 );
nand ( n49761 , n49760 , n48929 );
nand ( n49762 , n49754 , n49761 );
xor ( n49763 , n49751 , n49762 );
xor ( n49764 , n49740 , n49763 );
xor ( n49765 , n49764 , n49579 );
not ( n49766 , n49618 );
and ( n49767 , n46441 , n49766 );
not ( n49768 , n46441 );
not ( n49769 , n49617 );
not ( n49770 , n49769 );
and ( n49771 , n49768 , n49770 );
nor ( n49772 , n49767 , n49771 );
not ( n49773 , n49772 );
not ( n49774 , n49617 );
nand ( n49775 , n49774 , n49388 );
nand ( n49776 , n49617 , n49600 );
nand ( n49777 , n49775 , n49776 , n49391 );
buf ( n49778 , n49777 );
not ( n49779 , n49778 );
not ( n49780 , n49779 );
or ( n49781 , n49773 , n49780 );
not ( n49782 , n45816 );
buf ( n49783 , n49774 );
not ( n49784 , n49783 );
or ( n49785 , n49782 , n49784 );
nand ( n49786 , n49618 , n48766 );
nand ( n49787 , n49785 , n49786 );
buf ( n49788 , n49391 );
not ( n49789 , n49788 );
nand ( n49790 , n49787 , n49789 );
nand ( n49791 , n49781 , n49790 );
xor ( n49792 , n49791 , n49435 );
xor ( n49793 , n49792 , n49571 );
xor ( n49794 , n49793 , n49583 );
xor ( n49795 , n49794 , n49587 );
xor ( n49796 , n49765 , n49795 );
xor ( n49797 , n49796 , n49595 );
xor ( n49798 , n49765 , n49795 );
and ( n49799 , n49798 , n49595 );
and ( n49800 , n49765 , n49795 );
or ( n49801 , n49799 , n49800 );
not ( n49802 , n46602 );
not ( n49803 , n46072 );
not ( n49804 , n40948 );
not ( n49805 , n49804 );
buf ( n49806 , n49805 );
not ( n49807 , n49806 );
or ( n49808 , n49803 , n49807 );
not ( n49809 , n49804 );
not ( n49810 , n49809 );
nand ( n49811 , n49810 , n46071 );
nand ( n49812 , n49808 , n49811 );
not ( n49813 , n49812 );
or ( n49814 , n49802 , n49813 );
nand ( n49815 , n49551 , n46474 );
nand ( n49816 , n49814 , n49815 );
xor ( n49817 , n49816 , n49575 );
not ( n49818 , n49026 );
not ( n49819 , n46425 );
not ( n49820 , n41364 );
not ( n49821 , n49820 );
or ( n49822 , n49819 , n49821 );
not ( n49823 , n48679 );
nand ( n49824 , n49823 , n46422 );
nand ( n49825 , n49822 , n49824 );
not ( n49826 , n49825 );
or ( n49827 , n49818 , n49826 );
nand ( n49828 , n49516 , n46267 );
nand ( n49829 , n49827 , n49828 );
xor ( n49830 , n49817 , n49829 );
xor ( n49831 , n49830 , n49591 );
buf ( n49832 , n45748 );
not ( n49833 , n49832 );
not ( n49834 , n48952 );
not ( n49835 , n41216 );
or ( n49836 , n49834 , n49835 );
buf ( n49837 , n41216 );
not ( n49838 , n49837 );
nand ( n49839 , n49838 , n48955 );
nand ( n49840 , n49836 , n49839 );
not ( n49841 , n49840 );
or ( n49842 , n49833 , n49841 );
nand ( n49843 , n49536 , n46564 );
nand ( n49844 , n49842 , n49843 );
xor ( n49845 , n49646 , n49844 );
xor ( n49846 , n49845 , n49698 );
xor ( n49847 , n49831 , n49846 );
xor ( n49848 , n49599 , n49847 );
xor ( n49849 , n49848 , n49528 );
xor ( n49850 , n49599 , n49847 );
and ( n49851 , n49850 , n49528 );
and ( n49852 , n49599 , n49847 );
or ( n49853 , n49851 , n49852 );
xor ( n49854 , n49797 , n49561 );
xor ( n49855 , n49854 , n49849 );
xor ( n49856 , n49797 , n49561 );
and ( n49857 , n49856 , n49849 );
and ( n49858 , n49797 , n49561 );
or ( n49859 , n49857 , n49858 );
xor ( n49860 , n49750 , n49397 );
and ( n49861 , n49860 , n49762 );
and ( n49862 , n49750 , n49397 );
or ( n49863 , n49861 , n49862 );
xor ( n49864 , n49715 , n49725 );
and ( n49865 , n49864 , n49739 );
and ( n49866 , n49715 , n49725 );
or ( n49867 , n49865 , n49866 );
xor ( n49868 , n49791 , n49435 );
and ( n49869 , n49868 , n49571 );
and ( n49870 , n49791 , n49435 );
or ( n49871 , n49869 , n49870 );
xor ( n49872 , n49646 , n49844 );
and ( n49873 , n49872 , n49698 );
and ( n49874 , n49646 , n49844 );
or ( n49875 , n49873 , n49874 );
xor ( n49876 , n49816 , n49575 );
and ( n49877 , n49876 , n49829 );
and ( n49878 , n49816 , n49575 );
or ( n49879 , n49877 , n49878 );
xor ( n49880 , n49740 , n49763 );
and ( n49881 , n49880 , n49579 );
and ( n49882 , n49740 , n49763 );
or ( n49883 , n49881 , n49882 );
xor ( n49884 , n49793 , n49583 );
and ( n49885 , n49884 , n49587 );
and ( n49886 , n49793 , n49583 );
or ( n49887 , n49885 , n49886 );
xor ( n49888 , n49830 , n49591 );
and ( n49889 , n49888 , n49846 );
and ( n49890 , n49830 , n49591 );
or ( n49891 , n49889 , n49890 );
not ( n49892 , n49694 );
not ( n49893 , n47300 );
or ( n49894 , n49892 , n49893 );
and ( n49895 , n41861 , n47108 );
not ( n49896 , n41861 );
and ( n49897 , n49896 , n47107 );
nor ( n49898 , n49895 , n49897 );
nand ( n49899 , n47148 , n49898 );
nand ( n49900 , n49894 , n49899 );
not ( n49901 , n49632 );
not ( n49902 , n49116 );
or ( n49903 , n49901 , n49902 );
not ( n49904 , n30259 );
not ( n49905 , n47473 );
or ( n49906 , n49904 , n49905 );
nand ( n49907 , n47476 , n48829 );
nand ( n49908 , n49906 , n49907 );
nand ( n49909 , n47498 , n49908 );
nand ( n49910 , n49903 , n49909 );
xor ( n49911 , n49900 , n49910 );
and ( n49912 , n37653 , n37567 );
not ( n49913 , n37653 );
and ( n49914 , n49913 , n37566 );
nor ( n49915 , n49912 , n49914 );
and ( n49916 , n49915 , n49774 );
not ( n49917 , n49915 );
and ( n49918 , n49917 , n49617 );
nor ( n49919 , n49916 , n49918 );
not ( n49920 , n49919 );
and ( n49921 , n49920 , n46440 );
xor ( n49922 , n49911 , n49921 );
xor ( n49923 , n49900 , n49910 );
and ( n49924 , n49923 , n49921 );
and ( n49925 , n49900 , n49910 );
or ( n49926 , n49924 , n49925 );
not ( n49927 , n49643 );
not ( n49928 , n47873 );
or ( n49929 , n49927 , n49928 );
not ( n49930 , n47958 );
not ( n49931 , n47795 );
or ( n49932 , n49930 , n49931 );
nand ( n49933 , n47855 , n48860 );
nand ( n49934 , n49932 , n49933 );
nand ( n49935 , n49934 , n47881 );
nand ( n49936 , n49929 , n49935 );
not ( n49937 , n49660 );
not ( n49938 , n48463 );
or ( n49939 , n49937 , n49938 );
and ( n49940 , n48898 , n49658 );
not ( n49941 , n48898 );
and ( n49942 , n49941 , n48202 );
nor ( n49943 , n49940 , n49942 );
nand ( n49944 , n49148 , n49943 );
nand ( n49945 , n49939 , n49944 );
xor ( n49946 , n49936 , n49945 );
and ( n49947 , n49685 , n49696 );
xor ( n49948 , n49946 , n49947 );
xor ( n49949 , n49936 , n49945 );
and ( n49950 , n49949 , n49947 );
and ( n49951 , n49936 , n49945 );
or ( n49952 , n49950 , n49951 );
not ( n49953 , n49026 );
not ( n49954 , n46425 );
not ( n49955 , n48997 );
or ( n49956 , n49954 , n49955 );
nand ( n49957 , n49001 , n46422 );
nand ( n49958 , n49956 , n49957 );
not ( n49959 , n49958 );
or ( n49960 , n49953 , n49959 );
nand ( n49961 , n49825 , n46267 );
nand ( n49962 , n49960 , n49961 );
xor ( n49963 , n49863 , n49962 );
not ( n49964 , n46854 );
not ( n49965 , n48645 );
not ( n49966 , n48980 );
or ( n49967 , n49965 , n49966 );
not ( n49968 , n30964 );
not ( n49969 , n49968 );
not ( n49970 , n49675 );
nand ( n49971 , n49969 , n49970 );
nand ( n49972 , n49967 , n49971 );
not ( n49973 , n49972 );
or ( n49974 , n49964 , n49973 );
nand ( n49975 , n49681 , n48653 );
nand ( n49976 , n49974 , n49975 );
not ( n49977 , n49670 );
not ( n49978 , n49274 );
buf ( n49979 , n49978 );
not ( n49980 , n49979 );
or ( n49981 , n49977 , n49980 );
not ( n49982 , n47646 );
not ( n49983 , n49110 );
or ( n49984 , n49982 , n49983 );
nand ( n49985 , n49109 , n47650 );
nand ( n49986 , n49984 , n49985 );
nand ( n49987 , n49288 , n49986 );
nand ( n49988 , n49981 , n49987 );
xor ( n49989 , n49976 , n49988 );
not ( n49990 , n47407 );
not ( n49991 , n49760 );
or ( n49992 , n49990 , n49991 );
not ( n49993 , n48023 );
not ( n49994 , n48510 );
or ( n49995 , n49993 , n49994 );
nand ( n49996 , n41668 , n48727 );
nand ( n49997 , n49995 , n49996 );
nand ( n49998 , n49997 , n48929 );
nand ( n49999 , n49992 , n49998 );
xor ( n50000 , n49989 , n49999 );
xor ( n50001 , n49963 , n50000 );
not ( n50002 , n49832 );
not ( n50003 , n48952 );
not ( n50004 , n49549 );
not ( n50005 , n50004 );
or ( n50006 , n50003 , n50005 );
not ( n50007 , n40854 );
not ( n50008 , n50007 );
nand ( n50009 , n50008 , n48955 );
nand ( n50010 , n50006 , n50009 );
not ( n50011 , n50010 );
or ( n50012 , n50002 , n50011 );
nand ( n50013 , n49840 , n46564 );
nand ( n50014 , n50012 , n50013 );
xor ( n50015 , n49867 , n50014 );
not ( n50016 , n46474 );
not ( n50017 , n49812 );
or ( n50018 , n50016 , n50017 );
not ( n50019 , n46071 );
not ( n50020 , n41036 );
not ( n50021 , n50020 );
not ( n50022 , n50021 );
or ( n50023 , n50019 , n50022 );
nand ( n50024 , n50020 , n46072 );
nand ( n50025 , n50023 , n50024 );
nand ( n50026 , n50025 , n46602 );
nand ( n50027 , n50018 , n50026 );
xor ( n50028 , n50015 , n50027 );
xor ( n50029 , n50001 , n50028 );
xor ( n50030 , n50029 , n49883 );
xor ( n50031 , n50001 , n50028 );
and ( n50032 , n50031 , n49883 );
and ( n50033 , n50001 , n50028 );
or ( n50034 , n50032 , n50033 );
not ( n50035 , n47384 );
not ( n50036 , n49500 );
not ( n50037 , n41416 );
or ( n50038 , n50036 , n50037 );
nand ( n50039 , n41415 , n47979 );
nand ( n50040 , n50038 , n50039 );
not ( n50041 , n50040 );
or ( n50042 , n50035 , n50041 );
nand ( n50043 , n49721 , n46408 );
nand ( n50044 , n50042 , n50043 );
not ( n50045 , n49736 );
not ( n50046 , n48755 );
or ( n50047 , n50045 , n50046 );
not ( n50048 , n47227 );
not ( n50049 , n49314 );
or ( n50050 , n50048 , n50049 );
nand ( n50051 , n48705 , n47589 );
nand ( n50052 , n50050 , n50051 );
nand ( n50053 , n49022 , n50052 );
nand ( n50054 , n50047 , n50053 );
xor ( n50055 , n50044 , n50054 );
not ( n50056 , n49710 );
not ( n50057 , n49713 );
or ( n50058 , n50056 , n50057 );
not ( n50059 , n49707 );
not ( n50060 , n47332 );
or ( n50061 , n50059 , n50060 );
nand ( n50062 , n41683 , n48661 );
nand ( n50063 , n50061 , n50062 );
not ( n50064 , n50063 );
or ( n50065 , n50064 , n46439 );
nand ( n50066 , n50058 , n50065 );
xor ( n50067 , n50055 , n50066 );
xor ( n50068 , n50067 , n49871 );
not ( n50069 , n49787 );
not ( n50070 , n49778 );
not ( n50071 , n50070 );
or ( n50072 , n50069 , n50071 );
not ( n50073 , n46037 );
not ( n50074 , n49783 );
or ( n50075 , n50073 , n50074 );
nand ( n50076 , n49619 , n47306 );
nand ( n50077 , n50075 , n50076 );
buf ( n50078 , n49789 );
nand ( n50079 , n50077 , n50078 );
nand ( n50080 , n50072 , n50079 );
xor ( n50081 , n50080 , n49650 );
not ( n50082 , n45896 );
not ( n50083 , n46650 );
not ( n50084 , n48486 );
not ( n50085 , n50084 );
or ( n50086 , n50083 , n50085 );
not ( n50087 , n45951 );
nand ( n50088 , n48486 , n50087 );
nand ( n50089 , n50086 , n50088 );
not ( n50090 , n50089 );
or ( n50091 , n50082 , n50090 );
nand ( n50092 , n49746 , n48295 );
nand ( n50093 , n50091 , n50092 );
xor ( n50094 , n50081 , n50093 );
xor ( n50095 , n50068 , n50094 );
xor ( n50096 , n49887 , n50095 );
xor ( n50097 , n50096 , n49891 );
xor ( n50098 , n49887 , n50095 );
and ( n50099 , n50098 , n49891 );
and ( n50100 , n49887 , n50095 );
or ( n50101 , n50099 , n50100 );
xor ( n50102 , n49702 , n49948 );
xor ( n50103 , n50102 , n49922 );
xor ( n50104 , n50103 , n49879 );
xor ( n50105 , n50104 , n49875 );
xor ( n50106 , n50105 , n50030 );
xor ( n50107 , n50106 , n49801 );
xor ( n50108 , n50105 , n50030 );
and ( n50109 , n50108 , n49801 );
and ( n50110 , n50105 , n50030 );
or ( n50111 , n50109 , n50110 );
xor ( n50112 , n50097 , n50107 );
xor ( n50113 , n50112 , n49853 );
xor ( n50114 , n50097 , n50107 );
and ( n50115 , n50114 , n49853 );
and ( n50116 , n50097 , n50107 );
or ( n50117 , n50115 , n50116 );
xor ( n50118 , n49976 , n49988 );
and ( n50119 , n50118 , n49999 );
and ( n50120 , n49976 , n49988 );
or ( n50121 , n50119 , n50120 );
xor ( n50122 , n50044 , n50054 );
and ( n50123 , n50122 , n50066 );
and ( n50124 , n50044 , n50054 );
or ( n50125 , n50123 , n50124 );
xor ( n50126 , n50080 , n49650 );
and ( n50127 , n50126 , n50093 );
and ( n50128 , n50080 , n49650 );
or ( n50129 , n50127 , n50128 );
xor ( n50130 , n49702 , n49948 );
and ( n50131 , n50130 , n49922 );
and ( n50132 , n49702 , n49948 );
or ( n50133 , n50131 , n50132 );
xor ( n50134 , n49867 , n50014 );
and ( n50135 , n50134 , n50027 );
and ( n50136 , n49867 , n50014 );
or ( n50137 , n50135 , n50136 );
xor ( n50138 , n49863 , n49962 );
and ( n50139 , n50138 , n50000 );
and ( n50140 , n49863 , n49962 );
or ( n50141 , n50139 , n50140 );
xor ( n50142 , n50067 , n49871 );
and ( n50143 , n50142 , n50094 );
and ( n50144 , n50067 , n49871 );
or ( n50145 , n50143 , n50144 );
xor ( n50146 , n50103 , n49879 );
and ( n50147 , n50146 , n49875 );
and ( n50148 , n50103 , n49879 );
or ( n50149 , n50147 , n50148 );
not ( n50150 , n46440 );
not ( n50151 , n49915 );
or ( n50152 , n50150 , n50151 );
nand ( n50153 , n50152 , n49774 );
not ( n50154 , n49915 );
nand ( n50155 , n50154 , n46441 );
and ( n50156 , n50153 , n50155 );
not ( n50157 , n37580 );
not ( n50158 , n36696 );
or ( n50159 , n50157 , n50158 );
nand ( n50160 , n36695 , n37579 );
nand ( n50161 , n50159 , n50160 );
buf ( n50162 , n50161 );
not ( n50163 , n50162 );
nor ( n50164 , n50156 , n50163 );
not ( n50165 , n49934 );
not ( n50166 , n47873 );
or ( n50167 , n50165 , n50166 );
not ( n50168 , n49624 );
and ( n50169 , n47794 , n50168 );
not ( n50170 , n47794 );
and ( n50171 , n50170 , n49624 );
or ( n50172 , n50169 , n50171 );
nand ( n50173 , n50172 , n47881 );
nand ( n50174 , n50167 , n50173 );
xor ( n50175 , n50164 , n50174 );
buf ( n50176 , n48463 );
not ( n50177 , n50176 );
not ( n50178 , n49943 );
or ( n50179 , n50177 , n50178 );
not ( n50180 , n47765 );
not ( n50181 , n48967 );
or ( n50182 , n50180 , n50181 );
not ( n50183 , n47765 );
nand ( n50184 , n50183 , n48971 );
nand ( n50185 , n50182 , n50184 );
not ( n50186 , n50185 );
or ( n50187 , n50186 , n48276 );
nand ( n50188 , n50179 , n50187 );
xor ( n50189 , n50175 , n50188 );
xor ( n50190 , n50164 , n50174 );
and ( n50191 , n50190 , n50188 );
and ( n50192 , n50164 , n50174 );
or ( n50193 , n50191 , n50192 );
not ( n50194 , n49986 );
buf ( n50195 , n49979 );
not ( n50196 , n50195 );
or ( n50197 , n50194 , n50196 );
not ( n50198 , n49734 );
not ( n50199 , n49283 );
or ( n50200 , n50198 , n50199 );
not ( n50201 , n49259 );
nand ( n50202 , n50201 , n47821 );
nand ( n50203 , n50200 , n50202 );
nand ( n50204 , n49288 , n50203 );
nand ( n50205 , n50197 , n50204 );
not ( n50206 , n49898 );
not ( n50207 , n47139 );
or ( n50208 , n50206 , n50207 );
not ( n50209 , n47449 );
not ( n50210 , n47157 );
or ( n50211 , n50209 , n50210 );
nand ( n50212 , n41801 , n47107 );
nand ( n50213 , n50211 , n50212 );
nand ( n50214 , n50213 , n47147 );
nand ( n50215 , n50208 , n50214 );
not ( n50216 , n50215 );
not ( n50217 , n50216 );
not ( n50218 , n50217 );
and ( n50219 , n47489 , n49908 );
not ( n50220 , n47807 );
not ( n50221 , n47493 );
or ( n50222 , n50220 , n50221 );
nand ( n50223 , n46607 , n47476 );
nand ( n50224 , n50222 , n50223 );
and ( n50225 , n50224 , n47278 );
nor ( n50226 , n50219 , n50225 );
not ( n50227 , n50226 );
or ( n50228 , n50218 , n50227 );
or ( n50229 , n50217 , n50226 );
nand ( n50230 , n50228 , n50229 );
xor ( n50231 , n50205 , n50230 );
not ( n50232 , n49679 );
not ( n50233 , n50232 );
not ( n50234 , n47178 );
or ( n50235 , n50233 , n50234 );
nand ( n50236 , n47918 , n49679 );
nand ( n50237 , n50235 , n50236 );
not ( n50238 , n50237 );
not ( n50239 , n46854 );
or ( n50240 , n50238 , n50239 );
not ( n50241 , n48653 );
not ( n50242 , n50241 );
nand ( n50243 , n49972 , n50242 );
nand ( n50244 , n50240 , n50243 );
xor ( n50245 , n50231 , n50244 );
xor ( n50246 , n50205 , n50230 );
and ( n50247 , n50246 , n50244 );
and ( n50248 , n50205 , n50230 );
or ( n50249 , n50247 , n50248 );
not ( n50250 , n49832 );
not ( n50251 , n48952 );
not ( n50252 , n49809 );
or ( n50253 , n50251 , n50252 );
not ( n50254 , n49806 );
nand ( n50255 , n50254 , n47514 );
nand ( n50256 , n50253 , n50255 );
not ( n50257 , n50256 );
or ( n50258 , n50250 , n50257 );
nand ( n50259 , n50010 , n46564 );
nand ( n50260 , n50258 , n50259 );
buf ( n50261 , n45896 );
not ( n50262 , n50261 );
not ( n50263 , n50087 );
not ( n50264 , n50263 );
not ( n50265 , n48679 );
or ( n50266 , n50264 , n50265 );
not ( n50267 , n46650 );
nand ( n50268 , n50267 , n49823 );
nand ( n50269 , n50266 , n50268 );
not ( n50270 , n50269 );
or ( n50271 , n50262 , n50270 );
nand ( n50272 , n50089 , n48295 );
nand ( n50273 , n50271 , n50272 );
xor ( n50274 , n50260 , n50273 );
xor ( n50275 , n50274 , n50121 );
xor ( n50276 , n50275 , n50145 );
not ( n50277 , n48656 );
not ( n50278 , n49707 );
not ( n50279 , n47524 );
or ( n50280 , n50278 , n50279 );
nand ( n50281 , n30929 , n48661 );
nand ( n50282 , n50280 , n50281 );
not ( n50283 , n50282 );
or ( n50284 , n50277 , n50283 );
nand ( n50285 , n50063 , n49713 );
nand ( n50286 , n50284 , n50285 );
not ( n50287 , n50077 );
not ( n50288 , n50070 );
or ( n50289 , n50287 , n50288 );
not ( n50290 , n49788 );
not ( n50291 , n46273 );
not ( n50292 , n49618 );
not ( n50293 , n50292 );
or ( n50294 , n50291 , n50293 );
not ( n50295 , n49774 );
nand ( n50296 , n50295 , n46824 );
nand ( n50297 , n50294 , n50296 );
nand ( n50298 , n50290 , n50297 );
nand ( n50299 , n50289 , n50298 );
xor ( n50300 , n50286 , n50299 );
not ( n50301 , n50162 );
and ( n50302 , n46441 , n50301 );
not ( n50303 , n46441 );
buf ( n50304 , n50162 );
not ( n50305 , n50304 );
not ( n50306 , n50305 );
and ( n50307 , n50303 , n50306 );
nor ( n50308 , n50302 , n50307 );
not ( n50309 , n50308 );
not ( n50310 , n50154 );
not ( n50311 , n49617 );
and ( n50312 , n50310 , n50311 );
and ( n50313 , n50154 , n49617 );
nor ( n50314 , n50312 , n50313 );
and ( n50315 , n50162 , n49915 );
not ( n50316 , n50162 );
and ( n50317 , n50316 , n50154 );
nor ( n50318 , n50315 , n50317 );
nand ( n50319 , n50314 , n50318 );
buf ( n50320 , n50319 );
not ( n50321 , n50320 );
not ( n50322 , n50321 );
or ( n50323 , n50309 , n50322 );
not ( n50324 , n50163 );
and ( n50325 , n48766 , n50324 );
not ( n50326 , n48766 );
not ( n50327 , n50304 );
and ( n50328 , n50326 , n50327 );
or ( n50329 , n50325 , n50328 );
buf ( n50330 , n49919 );
not ( n50331 , n50330 );
nand ( n50332 , n50329 , n50331 );
nand ( n50333 , n50323 , n50332 );
xor ( n50334 , n50300 , n50333 );
not ( n50335 , n48929 );
not ( n50336 , n47803 );
not ( n50337 , n41530 );
or ( n50338 , n50336 , n50337 );
nand ( n50339 , n48779 , n47808 );
nand ( n50340 , n50338 , n50339 );
not ( n50341 , n50340 );
or ( n50342 , n50335 , n50341 );
nand ( n50343 , n49997 , n47407 );
nand ( n50344 , n50342 , n50343 );
not ( n50345 , n49252 );
not ( n50346 , n50040 );
or ( n50347 , n50345 , n50346 );
not ( n50348 , n47980 );
not ( n50349 , n48318 );
or ( n50350 , n50348 , n50349 );
nand ( n50351 , n41575 , n47979 );
nand ( n50352 , n50350 , n50351 );
nand ( n50353 , n50352 , n47384 );
nand ( n50354 , n50347 , n50353 );
xor ( n50355 , n50344 , n50354 );
not ( n50356 , n50052 );
not ( n50357 , n49309 );
or ( n50358 , n50356 , n50357 );
not ( n50359 , n49654 );
not ( n50360 , n48704 );
or ( n50361 , n50359 , n50360 );
nand ( n50362 , n48758 , n47368 );
nand ( n50363 , n50361 , n50362 );
nand ( n50364 , n50363 , n49320 );
nand ( n50365 , n50358 , n50364 );
xor ( n50366 , n50355 , n50365 );
xor ( n50367 , n50334 , n50366 );
xor ( n50368 , n50367 , n50245 );
xor ( n50369 , n50276 , n50368 );
xor ( n50370 , n50275 , n50145 );
and ( n50371 , n50370 , n50368 );
and ( n50372 , n50275 , n50145 );
or ( n50373 , n50371 , n50372 );
xor ( n50374 , n50129 , n50133 );
xor ( n50375 , n49926 , n49952 );
xor ( n50376 , n50375 , n50189 );
xor ( n50377 , n50374 , n50376 );
xor ( n50378 , n50149 , n50377 );
xor ( n50379 , n50378 , n50034 );
xor ( n50380 , n50149 , n50377 );
and ( n50381 , n50380 , n50034 );
and ( n50382 , n50149 , n50377 );
or ( n50383 , n50381 , n50382 );
xor ( n50384 , n50141 , n50137 );
not ( n50385 , n49026 );
not ( n50386 , n46425 );
not ( n50387 , n41217 );
not ( n50388 , n50387 );
or ( n50389 , n50386 , n50388 );
not ( n50390 , n49837 );
nand ( n50391 , n50390 , n46422 );
nand ( n50392 , n50389 , n50391 );
not ( n50393 , n50392 );
or ( n50394 , n50385 , n50393 );
nand ( n50395 , n49958 , n46267 );
nand ( n50396 , n50394 , n50395 );
xor ( n50397 , n50125 , n50396 );
not ( n50398 , n46602 );
not ( n50399 , n46072 );
not ( n50400 , n41132 );
not ( n50401 , n50400 );
or ( n50402 , n50399 , n50401 );
not ( n50403 , n41131 );
not ( n50404 , n50403 );
not ( n50405 , n46072 );
nand ( n50406 , n50404 , n50405 );
nand ( n50407 , n50402 , n50406 );
not ( n50408 , n50407 );
or ( n50409 , n50398 , n50408 );
nand ( n50410 , n50025 , n46474 );
nand ( n50411 , n50409 , n50410 );
xor ( n50412 , n50397 , n50411 );
xor ( n50413 , n50384 , n50412 );
xor ( n50414 , n50413 , n50369 );
xor ( n50415 , n50414 , n50379 );
xor ( n50416 , n50413 , n50369 );
and ( n50417 , n50416 , n50379 );
and ( n50418 , n50413 , n50369 );
or ( n50419 , n50417 , n50418 );
xor ( n50420 , n50101 , n50111 );
xor ( n50421 , n50420 , n50415 );
xor ( n50422 , n50101 , n50111 );
and ( n50423 , n50422 , n50415 );
and ( n50424 , n50101 , n50111 );
or ( n50425 , n50423 , n50424 );
xor ( n50426 , n50344 , n50354 );
and ( n50427 , n50426 , n50365 );
and ( n50428 , n50344 , n50354 );
or ( n50429 , n50427 , n50428 );
xor ( n50430 , n50286 , n50299 );
and ( n50431 , n50430 , n50333 );
and ( n50432 , n50286 , n50299 );
or ( n50433 , n50431 , n50432 );
xor ( n50434 , n49926 , n49952 );
and ( n50435 , n50434 , n50189 );
and ( n50436 , n49926 , n49952 );
or ( n50437 , n50435 , n50436 );
xor ( n50438 , n50260 , n50273 );
and ( n50439 , n50438 , n50121 );
and ( n50440 , n50260 , n50273 );
or ( n50441 , n50439 , n50440 );
xor ( n50442 , n50125 , n50396 );
and ( n50443 , n50442 , n50411 );
and ( n50444 , n50125 , n50396 );
or ( n50445 , n50443 , n50444 );
xor ( n50446 , n50334 , n50366 );
and ( n50447 , n50446 , n50245 );
and ( n50448 , n50334 , n50366 );
or ( n50449 , n50447 , n50448 );
xor ( n50450 , n50129 , n50133 );
and ( n50451 , n50450 , n50376 );
and ( n50452 , n50129 , n50133 );
or ( n50453 , n50451 , n50452 );
xor ( n50454 , n50141 , n50137 );
and ( n50455 , n50454 , n50412 );
and ( n50456 , n50141 , n50137 );
or ( n50457 , n50455 , n50456 );
not ( n50458 , n50224 );
not ( n50459 , n47489 );
or ( n50460 , n50458 , n50459 );
not ( n50461 , n47288 );
not ( n50462 , n47473 );
or ( n50463 , n50461 , n50462 );
nand ( n50464 , n47476 , n46994 );
nand ( n50465 , n50463 , n50464 );
nand ( n50466 , n47278 , n50465 );
nand ( n50467 , n50460 , n50466 );
not ( n50468 , n50172 );
not ( n50469 , n47873 );
or ( n50470 , n50468 , n50469 );
not ( n50471 , n48832 );
not ( n50472 , n48235 );
or ( n50473 , n50471 , n50472 );
nand ( n50474 , n47794 , n47982 );
nand ( n50475 , n50473 , n50474 );
nand ( n50476 , n50475 , n47881 );
nand ( n50477 , n50470 , n50476 );
xor ( n50478 , n50467 , n50477 );
not ( n50479 , n50185 );
not ( n50480 , n49421 );
or ( n50481 , n50479 , n50480 );
not ( n50482 , n47958 );
not ( n50483 , n48970 );
or ( n50484 , n50482 , n50483 );
nand ( n50485 , n49658 , n48860 );
nand ( n50486 , n50484 , n50485 );
nand ( n50487 , n50486 , n48452 );
nand ( n50488 , n50481 , n50487 );
xor ( n50489 , n50478 , n50488 );
xor ( n50490 , n50467 , n50477 );
and ( n50491 , n50490 , n50488 );
and ( n50492 , n50467 , n50477 );
or ( n50493 , n50491 , n50492 );
not ( n50494 , n47148 );
not ( n50495 , n48856 );
not ( n50496 , n47679 );
or ( n50497 , n50495 , n50496 );
not ( n50498 , n48856 );
nand ( n50499 , n50498 , n30964 );
nand ( n50500 , n50497 , n50499 );
not ( n50501 , n50500 );
or ( n50502 , n50494 , n50501 );
nand ( n50503 , n47300 , n50213 );
nand ( n50504 , n50502 , n50503 );
not ( n50505 , n50203 );
not ( n50506 , n49979 );
or ( n50507 , n50505 , n50506 );
not ( n50508 , n47227 );
not ( n50509 , n49282 );
or ( n50510 , n50508 , n50509 );
nand ( n50511 , n49109 , n47589 );
nand ( n50512 , n50510 , n50511 );
not ( n50513 , n48889 );
buf ( n50514 , n50513 );
nand ( n50515 , n50512 , n50514 );
nand ( n50516 , n50507 , n50515 );
xor ( n50517 , n50504 , n50516 );
not ( n50518 , n46854 );
not ( n50519 , n48645 );
not ( n50520 , n48523 );
or ( n50521 , n50519 , n50520 );
nand ( n50522 , n41683 , n49970 );
nand ( n50523 , n50521 , n50522 );
not ( n50524 , n50523 );
or ( n50525 , n50518 , n50524 );
nand ( n50526 , n50237 , n48653 );
nand ( n50527 , n50525 , n50526 );
xor ( n50528 , n50517 , n50527 );
xor ( n50529 , n50504 , n50516 );
and ( n50530 , n50529 , n50527 );
and ( n50531 , n50504 , n50516 );
or ( n50532 , n50530 , n50531 );
xor ( n50533 , n50489 , n50528 );
xor ( n50534 , n50533 , n50429 );
xor ( n50535 , n50534 , n50445 );
xor ( n50536 , n50535 , n50449 );
xor ( n50537 , n50534 , n50445 );
and ( n50538 , n50537 , n50449 );
and ( n50539 , n50534 , n50445 );
or ( n50540 , n50538 , n50539 );
not ( n50541 , n46267 );
not ( n50542 , n50392 );
or ( n50543 , n50541 , n50542 );
and ( n50544 , n46425 , n40854 );
not ( n50545 , n46425 );
not ( n50546 , n40854 );
and ( n50547 , n50545 , n50546 );
nor ( n50548 , n50544 , n50547 );
nand ( n50549 , n50548 , n49026 );
nand ( n50550 , n50543 , n50549 );
xor ( n50551 , n50550 , n50433 );
not ( n50552 , n50363 );
nand ( n50553 , n48753 , n48478 );
not ( n50554 , n50553 );
not ( n50555 , n50554 );
or ( n50556 , n50552 , n50555 );
not ( n50557 , n48898 );
not ( n50558 , n48704 );
or ( n50559 , n50557 , n50558 );
nand ( n50560 , n49093 , n48897 );
nand ( n50561 , n50559 , n50560 );
nand ( n50562 , n49320 , n50561 );
nand ( n50563 , n50556 , n50562 );
not ( n50564 , n50297 );
not ( n50565 , n49777 );
not ( n50566 , n50565 );
not ( n50567 , n50566 );
not ( n50568 , n50567 );
or ( n50569 , n50564 , n50568 );
not ( n50570 , n47646 );
not ( n50571 , n49774 );
or ( n50572 , n50570 , n50571 );
nand ( n50573 , n49618 , n47650 );
nand ( n50574 , n50572 , n50573 );
not ( n50575 , n49788 );
nand ( n50576 , n50574 , n50575 );
nand ( n50577 , n50569 , n50576 );
xor ( n50578 , n50563 , n50577 );
not ( n50579 , n50329 );
not ( n50580 , n50320 );
not ( n50581 , n50580 );
or ( n50582 , n50579 , n50581 );
not ( n50583 , n46037 );
not ( n50584 , n50163 );
or ( n50585 , n50583 , n50584 );
nand ( n50586 , n50304 , n47306 );
nand ( n50587 , n50585 , n50586 );
nand ( n50588 , n50587 , n50331 );
nand ( n50589 , n50582 , n50588 );
xor ( n50590 , n50578 , n50589 );
xor ( n50591 , n50551 , n50590 );
nor ( n50592 , n50226 , n50216 );
not ( n50593 , n47384 );
not ( n50594 , n47980 );
not ( n50595 , n49472 );
or ( n50596 , n50594 , n50595 );
nand ( n50597 , n46505 , n41667 );
nand ( n50598 , n50596 , n50597 );
not ( n50599 , n50598 );
or ( n50600 , n50593 , n50599 );
nand ( n50601 , n50352 , n46408 );
nand ( n50602 , n50600 , n50601 );
xor ( n50603 , n50592 , n50602 );
not ( n50604 , n49713 );
not ( n50605 , n50282 );
or ( n50606 , n50604 , n50605 );
and ( n50607 , n41415 , n48661 );
not ( n50608 , n41415 );
and ( n50609 , n50608 , n49707 );
or ( n50610 , n50607 , n50609 );
nand ( n50611 , n50610 , n48656 );
nand ( n50612 , n50606 , n50611 );
xor ( n50613 , n50603 , n50612 );
not ( n50614 , n37597 );
not ( n50615 , n50614 );
not ( n50616 , n36287 );
not ( n50617 , n50616 );
or ( n50618 , n50615 , n50617 );
nand ( n50619 , n36287 , n37597 );
nand ( n50620 , n50618 , n50619 );
not ( n50621 , n50620 );
and ( n50622 , n50162 , n50621 );
not ( n50623 , n50162 );
and ( n50624 , n50623 , n50620 );
nor ( n50625 , n50622 , n50624 );
buf ( n50626 , n50625 );
nor ( n50627 , n50626 , n46441 );
xor ( n50628 , n50627 , n50193 );
not ( n50629 , n48929 );
not ( n50630 , n47803 );
not ( n50631 , n41407 );
not ( n50632 , n50631 );
or ( n50633 , n50630 , n50632 );
buf ( n50634 , n48727 );
nand ( n50635 , n41407 , n50634 );
nand ( n50636 , n50633 , n50635 );
not ( n50637 , n50636 );
or ( n50638 , n50629 , n50637 );
nand ( n50639 , n50340 , n47407 );
nand ( n50640 , n50638 , n50639 );
xor ( n50641 , n50628 , n50640 );
xor ( n50642 , n50613 , n50641 );
xor ( n50643 , n50642 , n50437 );
xor ( n50644 , n50591 , n50643 );
xor ( n50645 , n50644 , n50453 );
xor ( n50646 , n50591 , n50643 );
and ( n50647 , n50646 , n50453 );
and ( n50648 , n50591 , n50643 );
or ( n50649 , n50647 , n50648 );
not ( n50650 , n46602 );
not ( n50651 , n46071 );
not ( n50652 , n40691 );
or ( n50653 , n50651 , n50652 );
not ( n50654 , n40691 );
nand ( n50655 , n50654 , n46072 );
nand ( n50656 , n50653 , n50655 );
not ( n50657 , n50656 );
or ( n50658 , n50650 , n50657 );
buf ( n50659 , n46474 );
nand ( n50660 , n50407 , n50659 );
nand ( n50661 , n50658 , n50660 );
xor ( n50662 , n50661 , n50441 );
not ( n50663 , n46564 );
not ( n50664 , n50256 );
or ( n50665 , n50663 , n50664 );
not ( n50666 , n47508 );
not ( n50667 , n41036 );
not ( n50668 , n50667 );
or ( n50669 , n50666 , n50668 );
or ( n50670 , n50667 , n47508 );
nand ( n50671 , n50669 , n50670 );
nand ( n50672 , n50671 , n45748 );
nand ( n50673 , n50665 , n50672 );
not ( n50674 , n45896 );
not ( n50675 , n46650 );
not ( n50676 , n41285 );
or ( n50677 , n50675 , n50676 );
nand ( n50678 , n49001 , n50087 );
nand ( n50679 , n50677 , n50678 );
not ( n50680 , n50679 );
or ( n50681 , n50674 , n50680 );
nand ( n50682 , n50269 , n48295 );
nand ( n50683 , n50681 , n50682 );
xor ( n50684 , n50673 , n50683 );
xor ( n50685 , n50684 , n50249 );
xor ( n50686 , n50662 , n50685 );
xor ( n50687 , n50457 , n50686 );
xor ( n50688 , n50687 , n50536 );
xor ( n50689 , n50457 , n50686 );
and ( n50690 , n50689 , n50536 );
and ( n50691 , n50457 , n50686 );
or ( n50692 , n50690 , n50691 );
xor ( n50693 , n50373 , n50383 );
xor ( n50694 , n50693 , n50645 );
xor ( n50695 , n50373 , n50383 );
and ( n50696 , n50695 , n50645 );
and ( n50697 , n50373 , n50383 );
or ( n50698 , n50696 , n50697 );
xor ( n50699 , n50688 , n50419 );
xor ( n50700 , n50699 , n50694 );
xor ( n50701 , n50688 , n50419 );
and ( n50702 , n50701 , n50694 );
and ( n50703 , n50688 , n50419 );
or ( n50704 , n50702 , n50703 );
xor ( n50705 , n50592 , n50602 );
and ( n50706 , n50705 , n50612 );
and ( n50707 , n50592 , n50602 );
or ( n50708 , n50706 , n50707 );
xor ( n50709 , n50563 , n50577 );
and ( n50710 , n50709 , n50589 );
and ( n50711 , n50563 , n50577 );
or ( n50712 , n50710 , n50711 );
xor ( n50713 , n50627 , n50193 );
and ( n50714 , n50713 , n50640 );
and ( n50715 , n50627 , n50193 );
or ( n50716 , n50714 , n50715 );
xor ( n50717 , n50489 , n50528 );
and ( n50718 , n50717 , n50429 );
and ( n50719 , n50489 , n50528 );
or ( n50720 , n50718 , n50719 );
xor ( n50721 , n50673 , n50683 );
and ( n50722 , n50721 , n50249 );
and ( n50723 , n50673 , n50683 );
or ( n50724 , n50722 , n50723 );
xor ( n50725 , n50550 , n50433 );
and ( n50726 , n50725 , n50590 );
and ( n50727 , n50550 , n50433 );
or ( n50728 , n50726 , n50727 );
xor ( n50729 , n50613 , n50641 );
and ( n50730 , n50729 , n50437 );
and ( n50731 , n50613 , n50641 );
or ( n50732 , n50730 , n50731 );
xor ( n50733 , n50661 , n50441 );
and ( n50734 , n50733 , n50685 );
and ( n50735 , n50661 , n50441 );
or ( n50736 , n50734 , n50735 );
not ( n50737 , n50486 );
nand ( n50738 , n48016 , n48266 );
not ( n50739 , n50738 );
not ( n50740 , n50739 );
or ( n50741 , n50737 , n50740 );
not ( n50742 , n48643 );
not ( n50743 , n48970 );
or ( n50744 , n50742 , n50743 );
nand ( n50745 , n48201 , n48171 );
nand ( n50746 , n50744 , n50745 );
nand ( n50747 , n50746 , n48277 );
nand ( n50748 , n50741 , n50747 );
not ( n50749 , n50512 );
not ( n50750 , n49978 );
or ( n50751 , n50749 , n50750 );
not ( n50752 , n49654 );
not ( n50753 , n49282 );
or ( n50754 , n50752 , n50753 );
not ( n50755 , n47740 );
nand ( n50756 , n50755 , n49281 );
nand ( n50757 , n50754 , n50756 );
nand ( n50758 , n50757 , n50513 );
nand ( n50759 , n50751 , n50758 );
xor ( n50760 , n50748 , n50759 );
not ( n50761 , n48856 );
not ( n50762 , n47510 );
or ( n50763 , n50761 , n50762 );
nand ( n50764 , n41692 , n50498 );
nand ( n50765 , n50763 , n50764 );
not ( n50766 , n50765 );
buf ( n50767 , n46975 );
not ( n50768 , n50767 );
or ( n50769 , n50766 , n50768 );
nand ( n50770 , n50500 , n47300 );
nand ( n50771 , n50769 , n50770 );
xor ( n50772 , n50760 , n50771 );
xor ( n50773 , n50748 , n50759 );
and ( n50774 , n50773 , n50771 );
and ( n50775 , n50748 , n50759 );
or ( n50776 , n50774 , n50775 );
not ( n50777 , n50475 );
not ( n50778 , n47872 );
or ( n50779 , n50777 , n50778 );
not ( n50780 , n46608 );
not ( n50781 , n48235 );
or ( n50782 , n50780 , n50781 );
nand ( n50783 , n47794 , n41938 );
nand ( n50784 , n50782 , n50783 );
nand ( n50785 , n50784 , n47881 );
nand ( n50786 , n50779 , n50785 );
not ( n50787 , n50465 );
not ( n50788 , n47489 );
or ( n50789 , n50787 , n50788 );
not ( n50790 , n47476 );
not ( n50791 , n47157 );
or ( n50792 , n50790 , n50791 );
nand ( n50793 , n41801 , n47473 );
nand ( n50794 , n50792 , n50793 );
nand ( n50795 , n50794 , n47278 );
nand ( n50796 , n50789 , n50795 );
xor ( n50797 , n50786 , n50796 );
not ( n50798 , n47384 );
not ( n50799 , n47979 );
not ( n50800 , n41531 );
or ( n50801 , n50799 , n50800 );
nand ( n50802 , n41530 , n49500 );
nand ( n50803 , n50801 , n50802 );
not ( n50804 , n50803 );
or ( n50805 , n50798 , n50804 );
nand ( n50806 , n46408 , n50598 );
nand ( n50807 , n50805 , n50806 );
xor ( n50808 , n50797 , n50807 );
not ( n50809 , n50523 );
or ( n50810 , n50809 , n50241 );
and ( n50811 , n47524 , n50232 );
not ( n50812 , n47524 );
and ( n50813 , n50812 , n48646 );
or ( n50814 , n50811 , n50813 );
not ( n50815 , n50814 );
or ( n50816 , n50815 , n50239 );
nand ( n50817 , n50810 , n50816 );
xor ( n50818 , n50808 , n50817 );
xor ( n50819 , n50797 , n50807 );
and ( n50820 , n50819 , n50817 );
and ( n50821 , n50797 , n50807 );
or ( n50822 , n50820 , n50821 );
not ( n50823 , n46188 );
not ( n50824 , n46425 );
not ( n50825 , n49805 );
or ( n50826 , n50824 , n50825 );
not ( n50827 , n49809 );
nand ( n50828 , n50827 , n46422 );
nand ( n50829 , n50826 , n50828 );
not ( n50830 , n50829 );
or ( n50831 , n50823 , n50830 );
nand ( n50832 , n50548 , n46267 );
nand ( n50833 , n50831 , n50832 );
xor ( n50834 , n50708 , n50833 );
xor ( n50835 , n50834 , n50772 );
not ( n50836 , n50671 );
not ( n50837 , n46564 );
or ( n50838 , n50836 , n50837 );
xor ( n50839 , n50400 , n47508 );
not ( n50840 , n49832 );
or ( n50841 , n50839 , n50840 );
nand ( n50842 , n50838 , n50841 );
xor ( n50843 , n50712 , n50842 );
not ( n50844 , n49713 );
not ( n50845 , n50610 );
or ( n50846 , n50844 , n50845 );
not ( n50847 , n47962 );
not ( n50848 , n48318 );
or ( n50849 , n50847 , n50848 );
not ( n50850 , n47962 );
nand ( n50851 , n50850 , n41575 );
nand ( n50852 , n50849 , n50851 );
nand ( n50853 , n50852 , n48656 );
nand ( n50854 , n50846 , n50853 );
not ( n50855 , n50561 );
not ( n50856 , n50554 );
or ( n50857 , n50855 , n50856 );
not ( n50858 , n47765 );
not ( n50859 , n48704 );
or ( n50860 , n50858 , n50859 );
nand ( n50861 , n48758 , n48589 );
nand ( n50862 , n50860 , n50861 );
nand ( n50863 , n50862 , n49320 );
nand ( n50864 , n50857 , n50863 );
xor ( n50865 , n50854 , n50864 );
not ( n50866 , n50574 );
not ( n50867 , n50567 );
or ( n50868 , n50866 , n50867 );
not ( n50869 , n49734 );
not ( n50870 , n49769 );
or ( n50871 , n50869 , n50870 );
nand ( n50872 , n49770 , n47821 );
nand ( n50873 , n50871 , n50872 );
nand ( n50874 , n50873 , n50575 );
nand ( n50875 , n50868 , n50874 );
xor ( n50876 , n50865 , n50875 );
xor ( n50877 , n50843 , n50876 );
xor ( n50878 , n50835 , n50877 );
xor ( n50879 , n50878 , n50732 );
xor ( n50880 , n50835 , n50877 );
and ( n50881 , n50880 , n50732 );
and ( n50882 , n50835 , n50877 );
or ( n50883 , n50881 , n50882 );
buf ( n50884 , n33649 );
buf ( n50885 , n50884 );
nand ( n50886 , n50885 , n36365 );
not ( n50887 , n50886 );
not ( n50888 , n50887 );
not ( n50889 , n36556 );
not ( n50890 , n50889 );
or ( n50891 , n50888 , n50890 );
nand ( n50892 , n36556 , n50886 );
nand ( n50893 , n50891 , n50892 );
not ( n50894 , n50893 );
not ( n50895 , n50894 );
and ( n50896 , n48689 , n50895 );
not ( n50897 , n48689 );
not ( n50898 , n50894 );
not ( n50899 , n50898 );
and ( n50900 , n50897 , n50899 );
nor ( n50901 , n50896 , n50900 );
not ( n50902 , n50901 );
nand ( n50903 , n50621 , n50894 );
not ( n50904 , n50887 );
not ( n50905 , n50889 );
or ( n50906 , n50904 , n50905 );
nand ( n50907 , n50906 , n50892 );
nand ( n50908 , n50907 , n50620 );
nand ( n50909 , n50903 , n50908 , n50625 );
buf ( n50910 , n50909 );
not ( n50911 , n50910 );
not ( n50912 , n50911 );
or ( n50913 , n50902 , n50912 );
not ( n50914 , n48766 );
not ( n50915 , n50914 );
not ( n50916 , n50893 );
not ( n50917 , n50916 );
or ( n50918 , n50915 , n50917 );
nand ( n50919 , n50898 , n48766 );
nand ( n50920 , n50918 , n50919 );
not ( n50921 , n50626 );
buf ( n50922 , n50921 );
nand ( n50923 , n50920 , n50922 );
nand ( n50924 , n50913 , n50923 );
xor ( n50925 , n50818 , n50924 );
xor ( n50926 , n50925 , n50716 );
xor ( n50927 , n50926 , n50540 );
not ( n50928 , n50587 );
not ( n50929 , n50319 );
not ( n50930 , n50929 );
or ( n50931 , n50928 , n50930 );
not ( n50932 , n46273 );
not ( n50933 , n50301 );
or ( n50934 , n50932 , n50933 );
nand ( n50935 , n50304 , n46824 );
nand ( n50936 , n50934 , n50935 );
nand ( n50937 , n50936 , n49920 );
nand ( n50938 , n50931 , n50937 );
not ( n50939 , n50620 );
not ( n50940 , n46440 );
and ( n50941 , n50939 , n50940 );
nand ( n50942 , n50620 , n46440 );
not ( n50943 , n50304 );
and ( n50944 , n50942 , n50943 );
nor ( n50945 , n50941 , n50944 );
buf ( n50946 , n50894 );
nor ( n50947 , n50945 , n50946 );
xor ( n50948 , n50938 , n50947 );
xor ( n50949 , n50948 , n50493 );
xor ( n50950 , n50949 , n50724 );
xor ( n50951 , n50950 , n50720 );
xor ( n50952 , n50927 , n50951 );
xor ( n50953 , n50926 , n50540 );
and ( n50954 , n50953 , n50951 );
and ( n50955 , n50926 , n50540 );
or ( n50956 , n50954 , n50955 );
not ( n50957 , n47009 );
not ( n50958 , n40677 );
and ( n50959 , n46072 , n50958 );
not ( n50960 , n46072 );
and ( n50961 , n50960 , n40677 );
or ( n50962 , n50959 , n50961 );
not ( n50963 , n50962 );
or ( n50964 , n50957 , n50963 );
nand ( n50965 , n50656 , n50659 );
nand ( n50966 , n50964 , n50965 );
not ( n50967 , n48295 );
not ( n50968 , n50679 );
or ( n50969 , n50967 , n50968 );
not ( n50970 , n46650 );
not ( n50971 , n41216 );
or ( n50972 , n50970 , n50971 );
not ( n50973 , n41216 );
nand ( n50974 , n50973 , n50087 );
nand ( n50975 , n50972 , n50974 );
nand ( n50976 , n50975 , n45896 );
nand ( n50977 , n50969 , n50976 );
not ( n50978 , n48929 );
not ( n50979 , n47803 );
not ( n50980 , n41363 );
not ( n50981 , n50980 );
or ( n50982 , n50979 , n50981 );
nand ( n50983 , n41363 , n50634 );
nand ( n50984 , n50982 , n50983 );
not ( n50985 , n50984 );
or ( n50986 , n50978 , n50985 );
nand ( n50987 , n50636 , n47407 );
nand ( n50988 , n50986 , n50987 );
xor ( n50989 , n50977 , n50988 );
xor ( n50990 , n50989 , n50532 );
xor ( n50991 , n50966 , n50990 );
xor ( n50992 , n50991 , n50728 );
xor ( n50993 , n50736 , n50992 );
xor ( n50994 , n50993 , n50879 );
xor ( n50995 , n50736 , n50992 );
and ( n50996 , n50995 , n50879 );
and ( n50997 , n50736 , n50992 );
or ( n50998 , n50996 , n50997 );
xor ( n50999 , n50649 , n50692 );
xor ( n51000 , n50999 , n50952 );
xor ( n51001 , n50649 , n50692 );
and ( n51002 , n51001 , n50952 );
and ( n51003 , n50649 , n50692 );
or ( n51004 , n51002 , n51003 );
xor ( n51005 , n50994 , n50698 );
xor ( n51006 , n51005 , n51000 );
xor ( n51007 , n50994 , n50698 );
and ( n51008 , n51007 , n51000 );
and ( n51009 , n50994 , n50698 );
or ( n51010 , n51008 , n51009 );
xor ( n51011 , n50854 , n50864 );
and ( n51012 , n51011 , n50875 );
and ( n51013 , n50854 , n50864 );
or ( n51014 , n51012 , n51013 );
xor ( n51015 , n50938 , n50947 );
and ( n51016 , n51015 , n50493 );
and ( n51017 , n50938 , n50947 );
or ( n51018 , n51016 , n51017 );
xor ( n51019 , n50977 , n50988 );
and ( n51020 , n51019 , n50532 );
and ( n51021 , n50977 , n50988 );
or ( n51022 , n51020 , n51021 );
xor ( n51023 , n50708 , n50833 );
and ( n51024 , n51023 , n50772 );
and ( n51025 , n50708 , n50833 );
or ( n51026 , n51024 , n51025 );
xor ( n51027 , n50712 , n50842 );
and ( n51028 , n51027 , n50876 );
and ( n51029 , n50712 , n50842 );
or ( n51030 , n51028 , n51029 );
xor ( n51031 , n50818 , n50924 );
and ( n51032 , n51031 , n50716 );
and ( n51033 , n50818 , n50924 );
or ( n51034 , n51032 , n51033 );
xor ( n51035 , n50949 , n50724 );
and ( n51036 , n51035 , n50720 );
and ( n51037 , n50949 , n50724 );
or ( n51038 , n51036 , n51037 );
xor ( n51039 , n50966 , n50990 );
and ( n51040 , n51039 , n50728 );
and ( n51041 , n50966 , n50990 );
or ( n51042 , n51040 , n51041 );
not ( n51043 , n50784 );
not ( n51044 , n47872 );
or ( n51045 , n51043 , n51044 );
not ( n51046 , n47617 );
not ( n51047 , n47795 );
or ( n51048 , n51046 , n51047 );
nand ( n51049 , n47794 , n46994 );
nand ( n51050 , n51048 , n51049 );
nand ( n51051 , n51050 , n47881 );
nand ( n51052 , n51045 , n51051 );
not ( n51053 , n50746 );
or ( n51054 , n50738 , n51053 );
not ( n51055 , n48832 );
not ( n51056 , n48455 );
or ( n51057 , n51055 , n51056 );
nand ( n51058 , n48201 , n47982 );
nand ( n51059 , n51057 , n51058 );
not ( n51060 , n51059 );
or ( n51061 , n51060 , n48276 );
nand ( n51062 , n51054 , n51061 );
xor ( n51063 , n51052 , n51062 );
not ( n51064 , n47498 );
not ( n51065 , n47476 );
not ( n51066 , n47318 );
or ( n51067 , n51065 , n51066 );
not ( n51068 , n47476 );
nand ( n51069 , n51068 , n30964 );
nand ( n51070 , n51067 , n51069 );
not ( n51071 , n51070 );
or ( n51072 , n51064 , n51071 );
nand ( n51073 , n47489 , n50794 );
nand ( n51074 , n51072 , n51073 );
xor ( n51075 , n51063 , n51074 );
xor ( n51076 , n51052 , n51062 );
and ( n51077 , n51076 , n51074 );
and ( n51078 , n51052 , n51062 );
or ( n51079 , n51077 , n51078 );
not ( n51080 , n50757 );
not ( n51081 , n49978 );
or ( n51082 , n51080 , n51081 );
not ( n51083 , n48898 );
not ( n51084 , n49259 );
or ( n51085 , n51083 , n51084 );
nand ( n51086 , n48897 , n49109 );
nand ( n51087 , n51085 , n51086 );
nand ( n51088 , n51087 , n50513 );
nand ( n51089 , n51082 , n51088 );
not ( n51090 , n47148 );
and ( n51091 , n41683 , n48857 );
not ( n51092 , n41683 );
and ( n51093 , n51092 , n48856 );
or ( n51094 , n51091 , n51093 );
not ( n51095 , n51094 );
or ( n51096 , n51090 , n51095 );
nand ( n51097 , n50765 , n47300 );
nand ( n51098 , n51096 , n51097 );
xor ( n51099 , n51089 , n51098 );
and ( n51100 , n50786 , n50796 );
xor ( n51101 , n51099 , n51100 );
xor ( n51102 , n51089 , n51098 );
and ( n51103 , n51102 , n51100 );
and ( n51104 , n51089 , n51098 );
or ( n51105 , n51103 , n51104 );
not ( n51106 , n46267 );
not ( n51107 , n50829 );
or ( n51108 , n51106 , n51107 );
not ( n51109 , n46425 );
not ( n51110 , n41036 );
not ( n51111 , n51110 );
or ( n51112 , n51109 , n51111 );
nand ( n51113 , n41036 , n46422 );
nand ( n51114 , n51112 , n51113 );
nand ( n51115 , n51114 , n46188 );
nand ( n51116 , n51108 , n51115 );
xor ( n51117 , n51014 , n51116 );
xor ( n51118 , n51117 , n51018 );
not ( n51119 , n47384 );
not ( n51120 , n47980 );
not ( n51121 , n50631 );
or ( n51122 , n51120 , n51121 );
not ( n51123 , n48483 );
nand ( n51124 , n51123 , n47979 );
nand ( n51125 , n51122 , n51124 );
not ( n51126 , n51125 );
or ( n51127 , n51119 , n51126 );
nand ( n51128 , n50803 , n49252 );
nand ( n51129 , n51127 , n51128 );
not ( n51130 , n37568 );
not ( n51131 , n36341 );
or ( n51132 , n51130 , n51131 );
nand ( n51133 , n51132 , n37553 );
nand ( n51134 , n36362 , n36369 );
not ( n51135 , n51134 );
and ( n51136 , n51133 , n51135 );
not ( n51137 , n51133 );
and ( n51138 , n51137 , n51134 );
nor ( n51139 , n51136 , n51138 );
and ( n51140 , n50907 , n51139 );
not ( n51141 , n50907 );
not ( n51142 , n51139 );
and ( n51143 , n51141 , n51142 );
nor ( n51144 , n51140 , n51143 );
buf ( n51145 , n51144 );
not ( n51146 , n51145 );
nor ( n51147 , n51146 , n46441 );
xor ( n51148 , n51129 , n51147 );
not ( n51149 , n50261 );
not ( n51150 , n46650 );
not ( n51151 , n49545 );
or ( n51152 , n51150 , n51151 );
nand ( n51153 , n49549 , n50087 );
nand ( n51154 , n51152 , n51153 );
not ( n51155 , n51154 );
or ( n51156 , n51149 , n51155 );
not ( n51157 , n46775 );
nand ( n51158 , n50975 , n51157 );
nand ( n51159 , n51156 , n51158 );
xor ( n51160 , n51148 , n51159 );
xor ( n51161 , n51118 , n51160 );
not ( n51162 , n50984 );
not ( n51163 , n47407 );
or ( n51164 , n51162 , n51163 );
not ( n51165 , n47803 );
not ( n51166 , n41284 );
or ( n51167 , n51165 , n51166 );
nand ( n51168 , n49000 , n48727 );
nand ( n51169 , n51167 , n51168 );
nand ( n51170 , n51169 , n48929 );
nand ( n51171 , n51164 , n51170 );
xor ( n51172 , n51171 , n50776 );
xor ( n51173 , n51172 , n50822 );
xor ( n51174 , n51161 , n51173 );
xor ( n51175 , n51118 , n51160 );
and ( n51176 , n51175 , n51173 );
and ( n51177 , n51118 , n51160 );
or ( n51178 , n51176 , n51177 );
not ( n51179 , n48656 );
not ( n51180 , n46820 );
not ( n51181 , n48510 );
or ( n51182 , n51180 , n51181 );
nand ( n51183 , n41667 , n48661 );
nand ( n51184 , n51182 , n51183 );
not ( n51185 , n51184 );
or ( n51186 , n51179 , n51185 );
nand ( n51187 , n50852 , n46584 );
nand ( n51188 , n51186 , n51187 );
not ( n51189 , n48653 );
not ( n51190 , n50814 );
or ( n51191 , n51189 , n51190 );
not ( n51192 , n49675 );
not ( n51193 , n41415 );
not ( n51194 , n51193 );
or ( n51195 , n51192 , n51194 );
nand ( n51196 , n48646 , n41415 );
nand ( n51197 , n51195 , n51196 );
nand ( n51198 , n51197 , n46854 );
nand ( n51199 , n51191 , n51198 );
xor ( n51200 , n51188 , n51199 );
not ( n51201 , n50862 );
not ( n51202 , n48755 );
or ( n51203 , n51201 , n51202 );
not ( n51204 , n48860 );
not ( n51205 , n51204 );
not ( n51206 , n48704 );
or ( n51207 , n51205 , n51206 );
nand ( n51208 , n49017 , n48860 );
nand ( n51209 , n51207 , n51208 );
nand ( n51210 , n49737 , n51209 );
nand ( n51211 , n51203 , n51210 );
xor ( n51212 , n51200 , n51211 );
xor ( n51213 , n51212 , n51101 );
not ( n51214 , n50920 );
not ( n51215 , n50910 );
not ( n51216 , n51215 );
or ( n51217 , n51214 , n51216 );
not ( n51218 , n46037 );
not ( n51219 , n50916 );
or ( n51220 , n51218 , n51219 );
nand ( n51221 , n50898 , n47306 );
nand ( n51222 , n51220 , n51221 );
not ( n51223 , n50626 );
nand ( n51224 , n51222 , n51223 );
nand ( n51225 , n51217 , n51224 );
xor ( n51226 , n51213 , n51225 );
xor ( n51227 , n51226 , n51034 );
xor ( n51228 , n51227 , n51038 );
xor ( n51229 , n51226 , n51034 );
and ( n51230 , n51229 , n51038 );
and ( n51231 , n51226 , n51034 );
or ( n51232 , n51230 , n51231 );
not ( n51233 , n50873 );
not ( n51234 , n49778 );
not ( n51235 , n51234 );
or ( n51236 , n51233 , n51235 );
not ( n51237 , n47227 );
not ( n51238 , n50292 );
or ( n51239 , n51237 , n51238 );
nand ( n51240 , n49770 , n47589 );
nand ( n51241 , n51239 , n51240 );
nand ( n51242 , n51241 , n50575 );
nand ( n51243 , n51236 , n51242 );
not ( n51244 , n50936 );
not ( n51245 , n50580 );
or ( n51246 , n51244 , n51245 );
not ( n51247 , n47646 );
not ( n51248 , n50301 );
or ( n51249 , n51247 , n51248 );
not ( n51250 , n50301 );
nand ( n51251 , n51250 , n47650 );
nand ( n51252 , n51249 , n51251 );
nand ( n51253 , n51252 , n49920 );
nand ( n51254 , n51246 , n51253 );
xor ( n51255 , n51243 , n51254 );
xor ( n51256 , n51255 , n51075 );
xor ( n51257 , n51256 , n51026 );
xor ( n51258 , n51257 , n51022 );
xor ( n51259 , n51258 , n51042 );
xor ( n51260 , n51259 , n51174 );
xor ( n51261 , n51258 , n51042 );
and ( n51262 , n51261 , n51174 );
and ( n51263 , n51258 , n51042 );
or ( n51264 , n51262 , n51263 );
not ( n51265 , n49832 );
not ( n51266 , n47514 );
not ( n51267 , n40691 );
or ( n51268 , n51266 , n51267 );
nand ( n51269 , n50654 , n48952 );
nand ( n51270 , n51268 , n51269 );
not ( n51271 , n51270 );
or ( n51272 , n51265 , n51271 );
not ( n51273 , n50839 );
nand ( n51274 , n51273 , n46564 );
nand ( n51275 , n51272 , n51274 );
xor ( n51276 , n51275 , n51030 );
not ( n51277 , n50962 );
not ( n51278 , n50659 );
or ( n51279 , n51277 , n51278 );
not ( n51280 , n40732 );
xor ( n51281 , n51280 , n46072 );
not ( n51282 , n51281 );
or ( n51283 , n51282 , n45861 );
nand ( n51284 , n51279 , n51283 );
xor ( n51285 , n51276 , n51284 );
xor ( n51286 , n50883 , n51285 );
xor ( n51287 , n51286 , n51228 );
xor ( n51288 , n50883 , n51285 );
and ( n51289 , n51288 , n51228 );
and ( n51290 , n50883 , n51285 );
or ( n51291 , n51289 , n51290 );
xor ( n51292 , n50956 , n51260 );
xor ( n51293 , n51292 , n50998 );
xor ( n51294 , n50956 , n51260 );
and ( n51295 , n51294 , n50998 );
and ( n51296 , n50956 , n51260 );
or ( n51297 , n51295 , n51296 );
xor ( n51298 , n51287 , n51004 );
xor ( n51299 , n51298 , n51293 );
xor ( n51300 , n51287 , n51004 );
and ( n51301 , n51300 , n51293 );
and ( n51302 , n51287 , n51004 );
or ( n51303 , n51301 , n51302 );
xor ( n51304 , n51188 , n51199 );
and ( n51305 , n51304 , n51211 );
and ( n51306 , n51188 , n51199 );
or ( n51307 , n51305 , n51306 );
xor ( n51308 , n51243 , n51254 );
and ( n51309 , n51308 , n51075 );
and ( n51310 , n51243 , n51254 );
or ( n51311 , n51309 , n51310 );
xor ( n51312 , n51129 , n51147 );
and ( n51313 , n51312 , n51159 );
and ( n51314 , n51129 , n51147 );
or ( n51315 , n51313 , n51314 );
xor ( n51316 , n51171 , n50776 );
and ( n51317 , n51316 , n50822 );
and ( n51318 , n51171 , n50776 );
or ( n51319 , n51317 , n51318 );
xor ( n51320 , n51014 , n51116 );
and ( n51321 , n51320 , n51018 );
and ( n51322 , n51014 , n51116 );
or ( n51323 , n51321 , n51322 );
xor ( n51324 , n51212 , n51101 );
and ( n51325 , n51324 , n51225 );
and ( n51326 , n51212 , n51101 );
or ( n51327 , n51325 , n51326 );
xor ( n51328 , n51256 , n51026 );
and ( n51329 , n51328 , n51022 );
and ( n51330 , n51256 , n51026 );
or ( n51331 , n51329 , n51330 );
xor ( n51332 , n51275 , n51030 );
and ( n51333 , n51332 , n51284 );
and ( n51334 , n51275 , n51030 );
or ( n51335 , n51333 , n51334 );
not ( n51336 , n51087 );
not ( n51337 , n49275 );
not ( n51338 , n51337 );
or ( n51339 , n51336 , n51338 );
not ( n51340 , n47765 );
not ( n51341 , n49283 );
or ( n51342 , n51340 , n51341 );
nand ( n51343 , n49262 , n48589 );
nand ( n51344 , n51342 , n51343 );
nand ( n51345 , n51344 , n50514 );
nand ( n51346 , n51339 , n51345 );
not ( n51347 , n48656 );
not ( n51348 , n49707 );
not ( n51349 , n41530 );
or ( n51350 , n51348 , n51349 );
buf ( n51351 , n48661 );
nand ( n51352 , n41531 , n51351 );
nand ( n51353 , n51350 , n51352 );
not ( n51354 , n51353 );
or ( n51355 , n51347 , n51354 );
nand ( n51356 , n51184 , n49713 );
nand ( n51357 , n51355 , n51356 );
xor ( n51358 , n51346 , n51357 );
not ( n51359 , n50767 );
not ( n51360 , n47527 );
and ( n51361 , n48856 , n51360 );
not ( n51362 , n48856 );
and ( n51363 , n51362 , n47527 );
or ( n51364 , n51361 , n51363 );
not ( n51365 , n51364 );
or ( n51366 , n51359 , n51365 );
buf ( n51367 , n47299 );
not ( n51368 , n51367 );
nand ( n51369 , n51094 , n51368 );
nand ( n51370 , n51366 , n51369 );
xor ( n51371 , n51358 , n51370 );
xor ( n51372 , n51346 , n51357 );
and ( n51373 , n51372 , n51370 );
and ( n51374 , n51346 , n51357 );
or ( n51375 , n51373 , n51374 );
not ( n51376 , n51059 );
not ( n51377 , n50739 );
or ( n51378 , n51376 , n51377 );
not ( n51379 , n47807 );
not ( n51380 , n48259 );
or ( n51381 , n51379 , n51380 );
nand ( n51382 , n49658 , n46607 );
nand ( n51383 , n51381 , n51382 );
nand ( n51384 , n51383 , n48017 );
nand ( n51385 , n51378 , n51384 );
not ( n51386 , n47881 );
not ( n51387 , n47794 );
not ( n51388 , n47157 );
or ( n51389 , n51387 , n51388 );
nand ( n51390 , n48235 , n47158 );
nand ( n51391 , n51389 , n51390 );
not ( n51392 , n51391 );
or ( n51393 , n51386 , n51392 );
nand ( n51394 , n51050 , n47872 );
nand ( n51395 , n51393 , n51394 );
xor ( n51396 , n51385 , n51395 );
not ( n51397 , n46854 );
and ( n51398 , n41575 , n48646 );
not ( n51399 , n41575 );
and ( n51400 , n51399 , n49675 );
or ( n51401 , n51398 , n51400 );
not ( n51402 , n51401 );
or ( n51403 , n51397 , n51402 );
nand ( n51404 , n51197 , n48653 );
nand ( n51405 , n51403 , n51404 );
xor ( n51406 , n51396 , n51405 );
not ( n51407 , n47498 );
not ( n51408 , n47437 );
not ( n51409 , n47178 );
or ( n51410 , n51408 , n51409 );
nand ( n51411 , n41692 , n49628 );
nand ( n51412 , n51410 , n51411 );
not ( n51413 , n51412 );
or ( n51414 , n51407 , n51413 );
nand ( n51415 , n51070 , n49116 );
nand ( n51416 , n51414 , n51415 );
xor ( n51417 , n51406 , n51416 );
xor ( n51418 , n51396 , n51405 );
and ( n51419 , n51418 , n51416 );
and ( n51420 , n51396 , n51405 );
or ( n51421 , n51419 , n51420 );
not ( n51422 , n51209 );
not ( n51423 , n48755 );
or ( n51424 , n51422 , n51423 );
not ( n51425 , n49624 );
not ( n51426 , n48764 );
not ( n51427 , n51426 );
or ( n51428 , n51425 , n51427 );
nand ( n51429 , n49093 , n50168 );
nand ( n51430 , n51428 , n51429 );
nand ( n51431 , n49022 , n51430 );
nand ( n51432 , n51424 , n51431 );
not ( n51433 , n51241 );
not ( n51434 , n50070 );
or ( n51435 , n51433 , n51434 );
not ( n51436 , n49654 );
not ( n51437 , n49766 );
or ( n51438 , n51436 , n51437 );
nand ( n51439 , n49619 , n47368 );
nand ( n51440 , n51438 , n51439 );
nand ( n51441 , n51440 , n49789 );
nand ( n51442 , n51435 , n51441 );
xor ( n51443 , n51432 , n51442 );
not ( n51444 , n51252 );
not ( n51445 , n50580 );
or ( n51446 , n51444 , n51445 );
not ( n51447 , n49734 );
not ( n51448 , n50301 );
or ( n51449 , n51447 , n51448 );
nand ( n51450 , n50324 , n47821 );
nand ( n51451 , n51449 , n51450 );
not ( n51452 , n49919 );
nand ( n51453 , n51451 , n51452 );
nand ( n51454 , n51446 , n51453 );
xor ( n51455 , n51443 , n51454 );
xor ( n51456 , n51455 , n51417 );
not ( n51457 , n51222 );
not ( n51458 , n50911 );
or ( n51459 , n51457 , n51458 );
not ( n51460 , n46273 );
buf ( n51461 , n50907 );
not ( n51462 , n51461 );
not ( n51463 , n51462 );
or ( n51464 , n51460 , n51463 );
not ( n51465 , n50916 );
nand ( n51466 , n51465 , n46824 );
nand ( n51467 , n51464 , n51466 );
nand ( n51468 , n51467 , n50922 );
nand ( n51469 , n51459 , n51468 );
xor ( n51470 , n51456 , n51469 );
xor ( n51471 , n51327 , n51470 );
not ( n51472 , n47384 );
not ( n51473 , n49500 );
not ( n51474 , n49820 );
or ( n51475 , n51473 , n51474 );
not ( n51476 , n49190 );
nand ( n51477 , n51476 , n47979 );
nand ( n51478 , n51475 , n51477 );
not ( n51479 , n51478 );
or ( n51480 , n51472 , n51479 );
nand ( n51481 , n48989 , n51125 );
nand ( n51482 , n51480 , n51481 );
xor ( n51483 , n51482 , n51371 );
not ( n51484 , n49026 );
not ( n51485 , n46425 );
not ( n51486 , n50400 );
or ( n51487 , n51485 , n51486 );
nand ( n51488 , n41132 , n46422 );
nand ( n51489 , n51487 , n51488 );
not ( n51490 , n51489 );
or ( n51491 , n51484 , n51490 );
nand ( n51492 , n51114 , n46267 );
nand ( n51493 , n51491 , n51492 );
xor ( n51494 , n51483 , n51493 );
xor ( n51495 , n51471 , n51494 );
xor ( n51496 , n51327 , n51470 );
and ( n51497 , n51496 , n51494 );
and ( n51498 , n51327 , n51470 );
or ( n51499 , n51497 , n51498 );
not ( n51500 , n37590 );
not ( n51501 , n36608 );
or ( n51502 , n51500 , n51501 );
nand ( n51503 , n51502 , n36375 );
not ( n51504 , n51503 );
not ( n51505 , n51504 );
and ( n51506 , n48689 , n51505 );
not ( n51507 , n48689 );
buf ( n51508 , n51504 );
and ( n51509 , n51507 , n51508 );
nor ( n51510 , n51506 , n51509 );
not ( n51511 , n51510 );
not ( n51512 , n50907 );
not ( n51513 , n51142 );
or ( n51514 , n51512 , n51513 );
nand ( n51515 , n50894 , n51139 );
nand ( n51516 , n51514 , n51515 );
not ( n51517 , n51139 );
not ( n51518 , n51503 );
or ( n51519 , n51517 , n51518 );
not ( n51520 , n51503 );
nand ( n51521 , n51520 , n51142 );
nand ( n51522 , n51519 , n51521 );
nor ( n51523 , n51516 , n51522 );
not ( n51524 , n51523 );
not ( n51525 , n51524 );
not ( n51526 , n51525 );
or ( n51527 , n51511 , n51526 );
not ( n51528 , n50914 );
not ( n51529 , n51504 );
or ( n51530 , n51528 , n51529 );
nand ( n51531 , n51505 , n48766 );
nand ( n51532 , n51530 , n51531 );
buf ( n51533 , n51145 );
nand ( n51534 , n51532 , n51533 );
nand ( n51535 , n51527 , n51534 );
xor ( n51536 , n51535 , n51311 );
xor ( n51537 , n51536 , n51315 );
xor ( n51538 , n51331 , n51537 );
xor ( n51539 , n51538 , n51335 );
xor ( n51540 , n51331 , n51537 );
and ( n51541 , n51540 , n51335 );
and ( n51542 , n51331 , n51537 );
or ( n51543 , n51541 , n51542 );
not ( n51544 , n48929 );
not ( n51545 , n50634 );
not ( n51546 , n51545 );
not ( n51547 , n49210 );
or ( n51548 , n51546 , n51547 );
nand ( n51549 , n49209 , n50634 );
nand ( n51550 , n51548 , n51549 );
not ( n51551 , n51550 );
or ( n51552 , n51544 , n51551 );
nand ( n51553 , n51169 , n47407 );
nand ( n51554 , n51552 , n51553 );
xor ( n51555 , n51079 , n51554 );
not ( n51556 , n50898 );
nand ( n51557 , n51139 , n48689 );
nand ( n51558 , n51556 , n51557 );
nand ( n51559 , n51142 , n46441 );
and ( n51560 , n51558 , n51559 );
not ( n51561 , n37590 );
not ( n51562 , n36608 );
or ( n51563 , n51561 , n51562 );
nand ( n51564 , n51563 , n36375 );
not ( n51565 , n51564 );
buf ( n51566 , n51565 );
nor ( n51567 , n51560 , n51566 );
xor ( n51568 , n51555 , n51567 );
xor ( n51569 , n51319 , n51568 );
not ( n51570 , n49832 );
not ( n51571 , n47508 );
buf ( n51572 , n40676 );
not ( n51573 , n51572 );
buf ( n51574 , n51573 );
not ( n51575 , n51574 );
or ( n51576 , n51571 , n51575 );
not ( n51577 , n48952 );
nand ( n51578 , n40677 , n51577 );
nand ( n51579 , n51576 , n51578 );
not ( n51580 , n51579 );
or ( n51581 , n51570 , n51580 );
nand ( n51582 , n51270 , n46564 );
nand ( n51583 , n51581 , n51582 );
xor ( n51584 , n51569 , n51583 );
xor ( n51585 , n51178 , n51584 );
xor ( n51586 , n51105 , n51307 );
not ( n51587 , n50261 );
not ( n51588 , n46650 );
not ( n51589 , n49809 );
or ( n51590 , n51588 , n51589 );
nand ( n51591 , n50827 , n48290 );
nand ( n51592 , n51590 , n51591 );
not ( n51593 , n51592 );
or ( n51594 , n51587 , n51593 );
nand ( n51595 , n51154 , n48295 );
nand ( n51596 , n51594 , n51595 );
xor ( n51597 , n51586 , n51596 );
xor ( n51598 , n51597 , n51323 );
not ( n51599 , n47009 );
not ( n51600 , n46072 );
buf ( n51601 , n40768 );
not ( n51602 , n51601 );
not ( n51603 , n51602 );
or ( n51604 , n51600 , n51603 );
nand ( n51605 , n51601 , n50405 );
nand ( n51606 , n51604 , n51605 );
not ( n51607 , n51606 );
or ( n51608 , n51599 , n51607 );
nand ( n51609 , n51281 , n50659 );
nand ( n51610 , n51608 , n51609 );
xor ( n51611 , n51598 , n51610 );
xor ( n51612 , n51585 , n51611 );
xor ( n51613 , n51178 , n51584 );
and ( n51614 , n51613 , n51611 );
and ( n51615 , n51178 , n51584 );
or ( n51616 , n51614 , n51615 );
xor ( n51617 , n51495 , n51232 );
xor ( n51618 , n51617 , n51539 );
xor ( n51619 , n51495 , n51232 );
and ( n51620 , n51619 , n51539 );
and ( n51621 , n51495 , n51232 );
or ( n51622 , n51620 , n51621 );
xor ( n51623 , n51264 , n51612 );
xor ( n51624 , n51623 , n51291 );
xor ( n51625 , n51264 , n51612 );
and ( n51626 , n51625 , n51291 );
and ( n51627 , n51264 , n51612 );
or ( n51628 , n51626 , n51627 );
xor ( n51629 , n51618 , n51297 );
xor ( n51630 , n51629 , n51624 );
xor ( n51631 , n51618 , n51297 );
and ( n51632 , n51631 , n51624 );
and ( n51633 , n51618 , n51297 );
or ( n51634 , n51632 , n51633 );
xor ( n51635 , n51432 , n51442 );
and ( n51636 , n51635 , n51454 );
and ( n51637 , n51432 , n51442 );
or ( n51638 , n51636 , n51637 );
xor ( n51639 , n51079 , n51554 );
and ( n51640 , n51639 , n51567 );
and ( n51641 , n51079 , n51554 );
or ( n51642 , n51640 , n51641 );
xor ( n51643 , n51105 , n51307 );
and ( n51644 , n51643 , n51596 );
and ( n51645 , n51105 , n51307 );
or ( n51646 , n51644 , n51645 );
xor ( n51647 , n51482 , n51371 );
and ( n51648 , n51647 , n51493 );
and ( n51649 , n51482 , n51371 );
or ( n51650 , n51648 , n51649 );
xor ( n51651 , n51455 , n51417 );
and ( n51652 , n51651 , n51469 );
and ( n51653 , n51455 , n51417 );
or ( n51654 , n51652 , n51653 );
xor ( n51655 , n51535 , n51311 );
and ( n51656 , n51655 , n51315 );
and ( n51657 , n51535 , n51311 );
or ( n51658 , n51656 , n51657 );
xor ( n51659 , n51319 , n51568 );
and ( n51660 , n51659 , n51583 );
and ( n51661 , n51319 , n51568 );
or ( n51662 , n51660 , n51661 );
xor ( n51663 , n51597 , n51323 );
and ( n51664 , n51663 , n51610 );
and ( n51665 , n51597 , n51323 );
or ( n51666 , n51664 , n51665 );
not ( n51667 , n48268 );
not ( n51668 , n51383 );
or ( n51669 , n51667 , n51668 );
buf ( n51670 , n47287 );
not ( n51671 , n51670 );
not ( n51672 , n51671 );
not ( n51673 , n48202 );
or ( n51674 , n51672 , n51673 );
nand ( n51675 , n49658 , n51670 );
nand ( n51676 , n51674 , n51675 );
nand ( n51677 , n51676 , n49148 );
nand ( n51678 , n51669 , n51677 );
not ( n51679 , n48240 );
buf ( n51680 , n47794 );
not ( n51681 , n51680 );
not ( n51682 , n48980 );
or ( n51683 , n51681 , n51682 );
not ( n51684 , n51680 );
nand ( n51685 , n30964 , n51684 );
nand ( n51686 , n51683 , n51685 );
not ( n51687 , n51686 );
or ( n51688 , n51679 , n51687 );
nand ( n51689 , n47873 , n51391 );
nand ( n51690 , n51688 , n51689 );
xor ( n51691 , n51678 , n51690 );
not ( n51692 , n51344 );
not ( n51693 , n50195 );
or ( n51694 , n51692 , n51693 );
not ( n51695 , n51204 );
not ( n51696 , n49283 );
or ( n51697 , n51695 , n51696 );
nand ( n51698 , n49111 , n48860 );
nand ( n51699 , n51697 , n51698 );
nand ( n51700 , n51699 , n48891 );
nand ( n51701 , n51694 , n51700 );
xor ( n51702 , n51691 , n51701 );
xor ( n51703 , n51678 , n51690 );
and ( n51704 , n51703 , n51701 );
and ( n51705 , n51678 , n51690 );
or ( n51706 , n51704 , n51705 );
not ( n51707 , n46854 );
not ( n51708 , n50232 );
not ( n51709 , n48510 );
or ( n51710 , n51708 , n51709 );
nand ( n51711 , n44141 , n49679 );
nand ( n51712 , n51710 , n51711 );
not ( n51713 , n51712 );
or ( n51714 , n51707 , n51713 );
nand ( n51715 , n51401 , n48653 );
nand ( n51716 , n51714 , n51715 );
not ( n51717 , n51368 );
not ( n51718 , n51364 );
or ( n51719 , n51717 , n51718 );
not ( n51720 , n48856 );
not ( n51721 , n41416 );
or ( n51722 , n51720 , n51721 );
buf ( n51723 , n47106 );
not ( n51724 , n51723 );
nand ( n51725 , n51724 , n41415 );
nand ( n51726 , n51722 , n51725 );
nand ( n51727 , n51726 , n47148 );
nand ( n51728 , n51719 , n51727 );
xor ( n51729 , n51716 , n51728 );
and ( n51730 , n51385 , n51395 );
xor ( n51731 , n51729 , n51730 );
xor ( n51732 , n51716 , n51728 );
and ( n51733 , n51732 , n51730 );
and ( n51734 , n51716 , n51728 );
or ( n51735 , n51733 , n51734 );
not ( n51736 , n47407 );
not ( n51737 , n51550 );
or ( n51738 , n51736 , n51737 );
not ( n51739 , n51545 );
not ( n51740 , n49548 );
not ( n51741 , n51740 );
not ( n51742 , n51741 );
or ( n51743 , n51739 , n51742 );
nand ( n51744 , n40854 , n50634 );
nand ( n51745 , n51743 , n51744 );
nand ( n51746 , n51745 , n48929 );
nand ( n51747 , n51738 , n51746 );
buf ( n51748 , n34054 );
not ( n51749 , n51748 );
buf ( n51750 , n33614 );
nor ( n51751 , n51749 , n51750 );
and ( n51752 , n37538 , n51751 );
not ( n51753 , n51752 );
buf ( n51754 , n36286 );
nand ( n51755 , n51754 , n37550 );
not ( n51756 , n51755 );
or ( n51757 , n51753 , n51756 );
not ( n51758 , n51755 );
not ( n51759 , n37538 );
or ( n51760 , n51758 , n51759 );
not ( n51761 , n51751 );
nand ( n51762 , n51760 , n51761 );
nand ( n51763 , n51757 , n51762 );
xnor ( n51764 , n51503 , n51763 );
not ( n51765 , n51764 );
buf ( n51766 , n51765 );
not ( n51767 , n51766 );
nor ( n51768 , n51767 , n46441 );
xor ( n51769 , n51747 , n51768 );
xor ( n51770 , n51769 , n51375 );
xor ( n51771 , n51650 , n51770 );
xor ( n51772 , n51771 , n51654 );
xor ( n51773 , n51650 , n51770 );
and ( n51774 , n51773 , n51654 );
and ( n51775 , n51650 , n51770 );
or ( n51776 , n51774 , n51775 );
xor ( n51777 , n51731 , n51638 );
not ( n51778 , n47498 );
not ( n51779 , n47437 );
not ( n51780 , n47332 );
or ( n51781 , n51779 , n51780 );
not ( n51782 , n47476 );
nand ( n51783 , n41683 , n51782 );
nand ( n51784 , n51781 , n51783 );
not ( n51785 , n51784 );
or ( n51786 , n51778 , n51785 );
nand ( n51787 , n51412 , n47489 );
nand ( n51788 , n51786 , n51787 );
not ( n51789 , n51430 );
not ( n51790 , n48755 );
or ( n51791 , n51789 , n51790 );
not ( n51792 , n48829 );
not ( n51793 , n51792 );
not ( n51794 , n48704 );
or ( n51795 , n51793 , n51794 );
nand ( n51796 , n49313 , n48829 );
nand ( n51797 , n51795 , n51796 );
nand ( n51798 , n51797 , n49737 );
nand ( n51799 , n51791 , n51798 );
xor ( n51800 , n51788 , n51799 );
not ( n51801 , n51440 );
not ( n51802 , n49779 );
or ( n51803 , n51801 , n51802 );
not ( n51804 , n48898 );
not ( n51805 , n50292 );
or ( n51806 , n51804 , n51805 );
nand ( n51807 , n49619 , n48897 );
nand ( n51808 , n51806 , n51807 );
not ( n51809 , n49788 );
nand ( n51810 , n51808 , n51809 );
nand ( n51811 , n51803 , n51810 );
xor ( n51812 , n51800 , n51811 );
xor ( n51813 , n51777 , n51812 );
xor ( n51814 , n51813 , n51658 );
not ( n51815 , n51532 );
not ( n51816 , n51525 );
or ( n51817 , n51815 , n51816 );
not ( n51818 , n51566 );
and ( n51819 , n46037 , n51818 );
not ( n51820 , n46037 );
and ( n51821 , n51820 , n51566 );
nor ( n51822 , n51819 , n51821 );
nand ( n51823 , n51822 , n51533 );
nand ( n51824 , n51817 , n51823 );
not ( n51825 , n51467 );
not ( n51826 , n50911 );
or ( n51827 , n51825 , n51826 );
not ( n51828 , n47646 );
not ( n51829 , n50899 );
or ( n51830 , n51828 , n51829 );
not ( n51831 , n50916 );
nand ( n51832 , n51831 , n47650 );
nand ( n51833 , n51830 , n51832 );
nand ( n51834 , n51833 , n50921 );
nand ( n51835 , n51827 , n51834 );
xor ( n51836 , n51824 , n51835 );
not ( n51837 , n49026 );
not ( n51838 , n46422 );
not ( n51839 , n40692 );
or ( n51840 , n51838 , n51839 );
not ( n51841 , n40691 );
nand ( n51842 , n51841 , n46425 );
nand ( n51843 , n51840 , n51842 );
not ( n51844 , n51843 );
or ( n51845 , n51837 , n51844 );
nand ( n51846 , n51489 , n46267 );
nand ( n51847 , n51845 , n51846 );
xor ( n51848 , n51836 , n51847 );
xor ( n51849 , n51814 , n51848 );
xor ( n51850 , n51813 , n51658 );
and ( n51851 , n51850 , n51848 );
and ( n51852 , n51813 , n51658 );
or ( n51853 , n51851 , n51852 );
xor ( n51854 , n51642 , n51646 );
not ( n51855 , n51451 );
not ( n51856 , n50321 );
or ( n51857 , n51855 , n51856 );
not ( n51858 , n47227 );
not ( n51859 , n50327 );
or ( n51860 , n51858 , n51859 );
nand ( n51861 , n50324 , n47589 );
nand ( n51862 , n51860 , n51861 );
nand ( n51863 , n51862 , n50331 );
nand ( n51864 , n51857 , n51863 );
buf ( n51865 , n48656 );
not ( n51866 , n51865 );
not ( n51867 , n49707 );
not ( n51868 , n50631 );
or ( n51869 , n51867 , n51868 );
nand ( n51870 , n48486 , n48661 );
nand ( n51871 , n51869 , n51870 );
not ( n51872 , n51871 );
or ( n51873 , n51866 , n51872 );
nand ( n51874 , n51353 , n49713 );
nand ( n51875 , n51873 , n51874 );
xor ( n51876 , n51864 , n51875 );
xor ( n51877 , n51876 , n51702 );
xor ( n51878 , n51854 , n51877 );
xor ( n51879 , n51662 , n51878 );
xor ( n51880 , n51879 , n51666 );
xor ( n51881 , n51662 , n51878 );
and ( n51882 , n51881 , n51666 );
and ( n51883 , n51662 , n51878 );
or ( n51884 , n51882 , n51883 );
not ( n51885 , n46776 );
not ( n51886 , n51592 );
or ( n51887 , n51885 , n51886 );
not ( n51888 , n46650 );
not ( n51889 , n41037 );
or ( n51890 , n51888 , n51889 );
buf ( n51891 , n41036 );
nand ( n51892 , n51891 , n48290 );
nand ( n51893 , n51890 , n51892 );
nand ( n51894 , n51893 , n50261 );
nand ( n51895 , n51887 , n51894 );
xor ( n51896 , n51421 , n51895 );
not ( n51897 , n47384 );
not ( n51898 , n49500 );
not ( n51899 , n48997 );
or ( n51900 , n51898 , n51899 );
nand ( n51901 , n49001 , n47979 );
nand ( n51902 , n51900 , n51901 );
not ( n51903 , n51902 );
or ( n51904 , n51897 , n51903 );
nand ( n51905 , n51478 , n48989 );
nand ( n51906 , n51904 , n51905 );
xor ( n51907 , n51896 , n51906 );
not ( n51908 , n50659 );
not ( n51909 , n51606 );
or ( n51910 , n51908 , n51909 );
not ( n51911 , n46072 );
buf ( n51912 , n40526 );
not ( n51913 , n51912 );
not ( n51914 , n51913 );
or ( n51915 , n51911 , n51914 );
buf ( n51916 , n40525 );
nand ( n51917 , n51916 , n46071 );
nand ( n51918 , n51915 , n51917 );
nand ( n51919 , n51918 , n44004 );
nand ( n51920 , n51910 , n51919 );
xor ( n51921 , n51907 , n51920 );
not ( n51922 , n49832 );
not ( n51923 , n47508 );
not ( n51924 , n51280 );
buf ( n51925 , n51924 );
not ( n51926 , n51925 );
or ( n51927 , n51923 , n51926 );
not ( n51928 , n40731 );
not ( n51929 , n51928 );
nand ( n51930 , n51929 , n47514 );
nand ( n51931 , n51927 , n51930 );
not ( n51932 , n51931 );
or ( n51933 , n51922 , n51932 );
nand ( n51934 , n51579 , n46564 );
nand ( n51935 , n51933 , n51934 );
xor ( n51936 , n51921 , n51935 );
xor ( n51937 , n51772 , n51936 );
xor ( n51938 , n51937 , n51499 );
xor ( n51939 , n51772 , n51936 );
and ( n51940 , n51939 , n51499 );
and ( n51941 , n51772 , n51936 );
or ( n51942 , n51940 , n51941 );
xor ( n51943 , n51543 , n51849 );
xor ( n51944 , n51943 , n51616 );
xor ( n51945 , n51543 , n51849 );
and ( n51946 , n51945 , n51616 );
and ( n51947 , n51543 , n51849 );
or ( n51948 , n51946 , n51947 );
xor ( n51949 , n51880 , n51938 );
xor ( n51950 , n51949 , n51622 );
xor ( n51951 , n51880 , n51938 );
and ( n51952 , n51951 , n51622 );
and ( n51953 , n51880 , n51938 );
or ( n51954 , n51952 , n51953 );
xor ( n51955 , n51944 , n51628 );
xor ( n51956 , n51955 , n51950 );
xor ( n51957 , n51944 , n51628 );
and ( n51958 , n51957 , n51950 );
and ( n51959 , n51944 , n51628 );
or ( n51960 , n51958 , n51959 );
xor ( n51961 , n51788 , n51799 );
and ( n51962 , n51961 , n51811 );
and ( n51963 , n51788 , n51799 );
or ( n51964 , n51962 , n51963 );
xor ( n51965 , n51864 , n51875 );
and ( n51966 , n51965 , n51702 );
and ( n51967 , n51864 , n51875 );
or ( n51968 , n51966 , n51967 );
xor ( n51969 , n51747 , n51768 );
and ( n51970 , n51969 , n51375 );
and ( n51971 , n51747 , n51768 );
or ( n51972 , n51970 , n51971 );
xor ( n51973 , n51421 , n51895 );
and ( n51974 , n51973 , n51906 );
and ( n51975 , n51421 , n51895 );
or ( n51976 , n51974 , n51975 );
xor ( n51977 , n51731 , n51638 );
and ( n51978 , n51977 , n51812 );
and ( n51979 , n51731 , n51638 );
or ( n51980 , n51978 , n51979 );
xor ( n51981 , n51824 , n51835 );
and ( n51982 , n51981 , n51847 );
and ( n51983 , n51824 , n51835 );
or ( n51984 , n51982 , n51983 );
xor ( n51985 , n51642 , n51646 );
and ( n51986 , n51985 , n51877 );
and ( n51987 , n51642 , n51646 );
or ( n51988 , n51986 , n51987 );
xor ( n51989 , n51907 , n51920 );
and ( n51990 , n51989 , n51935 );
and ( n51991 , n51907 , n51920 );
or ( n51992 , n51990 , n51991 );
not ( n51993 , n50767 );
not ( n51994 , n48856 );
not ( n51995 , n49298 );
not ( n51996 , n51995 );
or ( n51997 , n51994 , n51996 );
nand ( n51998 , n49293 , n51724 );
nand ( n51999 , n51997 , n51998 );
not ( n52000 , n51999 );
or ( n52001 , n51993 , n52000 );
nand ( n52002 , n51726 , n47139 );
nand ( n52003 , n52001 , n52002 );
buf ( n52004 , n47498 );
not ( n52005 , n52004 );
xor ( n52006 , n49628 , n49220 );
not ( n52007 , n52006 );
or ( n52008 , n52005 , n52007 );
nand ( n52009 , n49116 , n51784 );
nand ( n52010 , n52008 , n52009 );
xor ( n52011 , n52003 , n52010 );
not ( n52012 , n48240 );
not ( n52013 , n47855 );
not ( n52014 , n47510 );
or ( n52015 , n52013 , n52014 );
not ( n52016 , n47855 );
nand ( n52017 , n41692 , n52016 );
nand ( n52018 , n52015 , n52017 );
not ( n52019 , n52018 );
or ( n52020 , n52012 , n52019 );
not ( n52021 , n47872 );
not ( n52022 , n52021 );
nand ( n52023 , n51686 , n52022 );
nand ( n52024 , n52020 , n52023 );
xor ( n52025 , n52011 , n52024 );
xor ( n52026 , n52003 , n52010 );
and ( n52027 , n52026 , n52024 );
and ( n52028 , n52003 , n52010 );
or ( n52029 , n52027 , n52028 );
not ( n52030 , n51797 );
not ( n52031 , n49014 );
or ( n52032 , n52030 , n52031 );
buf ( n52033 , n47807 );
not ( n52034 , n52033 );
not ( n52035 , n51426 );
or ( n52036 , n52034 , n52035 );
not ( n52037 , n48704 );
not ( n52038 , n52033 );
nand ( n52039 , n52037 , n52038 );
nand ( n52040 , n52036 , n52039 );
nand ( n52041 , n49737 , n52040 );
nand ( n52042 , n52032 , n52041 );
not ( n52043 , n50239 );
not ( n52044 , n52043 );
not ( n52045 , n50232 );
not ( n52046 , n49233 );
or ( n52047 , n52045 , n52046 );
not ( n52048 , n48645 );
nand ( n52049 , n41531 , n52048 );
nand ( n52050 , n52047 , n52049 );
not ( n52051 , n52050 );
or ( n52052 , n52044 , n52051 );
nand ( n52053 , n51712 , n48653 );
nand ( n52054 , n52052 , n52053 );
xor ( n52055 , n52042 , n52054 );
not ( n52056 , n51808 );
buf ( n52057 , n50565 );
buf ( n52058 , n52057 );
not ( n52059 , n52058 );
or ( n52060 , n52056 , n52059 );
not ( n52061 , n47765 );
not ( n52062 , n50292 );
or ( n52063 , n52061 , n52062 );
nand ( n52064 , n49770 , n48589 );
nand ( n52065 , n52063 , n52064 );
nand ( n52066 , n52065 , n50078 );
nand ( n52067 , n52060 , n52066 );
xor ( n52068 , n52055 , n52067 );
xor ( n52069 , n52042 , n52054 );
and ( n52070 , n52069 , n52067 );
and ( n52071 , n52042 , n52054 );
or ( n52072 , n52070 , n52071 );
xor ( n52073 , n52025 , n52068 );
not ( n52074 , n47827 );
not ( n52075 , n50263 );
not ( n52076 , n41132 );
not ( n52077 , n52076 );
or ( n52078 , n52075 , n52077 );
buf ( n52079 , n50404 );
not ( n52080 , n46650 );
nand ( n52081 , n52079 , n52080 );
nand ( n52082 , n52078 , n52081 );
not ( n52083 , n52082 );
or ( n52084 , n52074 , n52083 );
nand ( n52085 , n51893 , n51157 );
nand ( n52086 , n52084 , n52085 );
xor ( n52087 , n52073 , n52086 );
xor ( n52088 , n51980 , n52087 );
xor ( n52089 , n52088 , n51984 );
xor ( n52090 , n51980 , n52087 );
and ( n52091 , n52090 , n51984 );
and ( n52092 , n51980 , n52087 );
or ( n52093 , n52091 , n52092 );
not ( n52094 , n46440 );
and ( n52095 , n37550 , n51748 );
not ( n52096 , n52095 );
not ( n52097 , n51754 );
or ( n52098 , n52096 , n52097 );
and ( n52099 , n37515 , n51748 );
nor ( n52100 , n52099 , n51750 );
nand ( n52101 , n52098 , n52100 );
and ( n52102 , n52101 , n37558 );
not ( n52103 , n52101 );
and ( n52104 , n52103 , n37559 );
nor ( n52105 , n52102 , n52104 );
buf ( n52106 , n52105 );
not ( n52107 , n52106 );
not ( n52108 , n52107 );
not ( n52109 , n52108 );
buf ( n52110 , n52109 );
not ( n52111 , n52110 );
or ( n52112 , n52094 , n52111 );
buf ( n52113 , n52107 );
not ( n52114 , n52113 );
nand ( n52115 , n52114 , n46441 );
nand ( n52116 , n52112 , n52115 );
not ( n52117 , n52116 );
and ( n52118 , n51763 , n52106 );
not ( n52119 , n51763 );
not ( n52120 , n52105 );
and ( n52121 , n52119 , n52120 );
nor ( n52122 , n52118 , n52121 );
nand ( n52123 , n52122 , n51764 );
buf ( n52124 , n52123 );
not ( n52125 , n52124 );
not ( n52126 , n52125 );
or ( n52127 , n52117 , n52126 );
not ( n52128 , n50914 );
buf ( n52129 , n52120 );
buf ( n52130 , n52129 );
not ( n52131 , n52130 );
or ( n52132 , n52128 , n52131 );
not ( n52133 , n52130 );
nand ( n52134 , n52133 , n48766 );
nand ( n52135 , n52132 , n52134 );
nand ( n52136 , n52135 , n51766 );
nand ( n52137 , n52127 , n52136 );
not ( n52138 , n51822 );
not ( n52139 , n51524 );
not ( n52140 , n52139 );
or ( n52141 , n52138 , n52140 );
not ( n52142 , n46273 );
not ( n52143 , n51508 );
or ( n52144 , n52142 , n52143 );
nand ( n52145 , n51505 , n46824 );
nand ( n52146 , n52144 , n52145 );
nand ( n52147 , n52146 , n51533 );
nand ( n52148 , n52141 , n52147 );
xor ( n52149 , n52137 , n52148 );
not ( n52150 , n51833 );
buf ( n52151 , n51215 );
not ( n52152 , n52151 );
or ( n52153 , n52150 , n52152 );
and ( n52154 , n47047 , n51461 );
not ( n52155 , n47047 );
and ( n52156 , n52155 , n51462 );
nor ( n52157 , n52154 , n52156 );
nand ( n52158 , n52157 , n51223 );
nand ( n52159 , n52153 , n52158 );
xor ( n52160 , n52149 , n52159 );
xor ( n52161 , n52160 , n51988 );
not ( n52162 , n51862 );
not ( n52163 , n50321 );
or ( n52164 , n52162 , n52163 );
not ( n52165 , n47368 );
not ( n52166 , n52165 );
not ( n52167 , n50327 );
or ( n52168 , n52166 , n52167 );
nand ( n52169 , n50304 , n47368 );
nand ( n52170 , n52168 , n52169 );
nand ( n52171 , n52170 , n49920 );
nand ( n52172 , n52164 , n52171 );
not ( n52173 , n51676 );
not ( n52174 , n48463 );
or ( n52175 , n52173 , n52174 );
not ( n52176 , n46880 );
and ( n52177 , n48970 , n52176 );
not ( n52178 , n48970 );
and ( n52179 , n52178 , n47157 );
or ( n52180 , n52177 , n52179 );
nand ( n52181 , n52180 , n48452 );
nand ( n52182 , n52175 , n52181 );
not ( n52183 , n51699 );
not ( n52184 , n49276 );
or ( n52185 , n52183 , n52184 );
not ( n52186 , n49624 );
not ( n52187 , n49259 );
or ( n52188 , n52186 , n52187 );
nand ( n52189 , n49284 , n50168 );
nand ( n52190 , n52188 , n52189 );
not ( n52191 , n48890 );
nand ( n52192 , n52190 , n52191 );
nand ( n52193 , n52185 , n52192 );
xor ( n52194 , n52182 , n52193 );
xor ( n52195 , n52172 , n52194 );
xor ( n52196 , n52195 , n51706 );
xor ( n52197 , n52196 , n51968 );
xor ( n52198 , n52197 , n51972 );
xor ( n52199 , n52161 , n52198 );
xor ( n52200 , n52160 , n51988 );
and ( n52201 , n52200 , n52198 );
and ( n52202 , n52160 , n51988 );
or ( n52203 , n52201 , n52202 );
not ( n52204 , n50659 );
not ( n52205 , n51918 );
or ( n52206 , n52204 , n52205 );
not ( n52207 , n46072 );
not ( n52208 , n40592 );
not ( n52209 , n52208 );
or ( n52210 , n52207 , n52209 );
not ( n52211 , n40590 );
not ( n52212 , n52211 );
nand ( n52213 , n52212 , n46071 );
nand ( n52214 , n52210 , n52213 );
nand ( n52215 , n52214 , n46602 );
nand ( n52216 , n52206 , n52215 );
not ( n52217 , n46564 );
not ( n52218 , n51931 );
or ( n52219 , n52217 , n52218 );
and ( n52220 , n48952 , n51602 );
not ( n52221 , n48952 );
not ( n52222 , n40768 );
not ( n52223 , n52222 );
and ( n52224 , n52221 , n52223 );
or ( n52225 , n52220 , n52224 );
nand ( n52226 , n52225 , n49832 );
nand ( n52227 , n52219 , n52226 );
xor ( n52228 , n52216 , n52227 );
not ( n52229 , n48929 );
not ( n52230 , n51545 );
not ( n52231 , n49809 );
or ( n52232 , n52230 , n52231 );
nand ( n52233 , n50254 , n48727 );
nand ( n52234 , n52232 , n52233 );
not ( n52235 , n52234 );
or ( n52236 , n52229 , n52235 );
nand ( n52237 , n51745 , n47407 );
nand ( n52238 , n52236 , n52237 );
and ( n52239 , n51763 , n46440 );
nor ( n52240 , n52239 , n51505 );
not ( n52241 , n46441 );
nor ( n52242 , n52241 , n51763 );
or ( n52243 , n52240 , n52242 );
nand ( n52244 , n52243 , n52114 );
not ( n52245 , n52244 );
xor ( n52246 , n52238 , n52245 );
xor ( n52247 , n52246 , n51735 );
xor ( n52248 , n52228 , n52247 );
xor ( n52249 , n51992 , n52248 );
xor ( n52250 , n52249 , n51776 );
xor ( n52251 , n51992 , n52248 );
and ( n52252 , n52251 , n51776 );
and ( n52253 , n51992 , n52248 );
or ( n52254 , n52252 , n52253 );
not ( n52255 , n48989 );
not ( n52256 , n51902 );
or ( n52257 , n52255 , n52256 );
not ( n52258 , n49500 );
not ( n52259 , n49837 );
or ( n52260 , n52258 , n52259 );
nand ( n52261 , n50973 , n47979 );
nand ( n52262 , n52260 , n52261 );
nand ( n52263 , n52262 , n47384 );
nand ( n52264 , n52257 , n52263 );
xor ( n52265 , n51964 , n52264 );
not ( n52266 , n51865 );
not ( n52267 , n51351 );
not ( n52268 , n52267 );
not ( n52269 , n48679 );
or ( n52270 , n52268 , n52269 );
not ( n52271 , n41363 );
not ( n52272 , n52271 );
not ( n52273 , n49707 );
nand ( n52274 , n52272 , n52273 );
nand ( n52275 , n52270 , n52274 );
not ( n52276 , n52275 );
or ( n52277 , n52266 , n52276 );
nand ( n52278 , n51871 , n49713 );
nand ( n52279 , n52277 , n52278 );
xor ( n52280 , n52265 , n52279 );
xor ( n52281 , n51976 , n52280 );
not ( n52282 , n49026 );
not ( n52283 , n46425 );
buf ( n52284 , n51572 );
not ( n52285 , n52284 );
buf ( n52286 , n52285 );
not ( n52287 , n52286 );
or ( n52288 , n52283 , n52287 );
buf ( n52289 , n40677 );
nand ( n52290 , n52289 , n46422 );
nand ( n52291 , n52288 , n52290 );
not ( n52292 , n52291 );
or ( n52293 , n52282 , n52292 );
nand ( n52294 , n51843 , n46267 );
nand ( n52295 , n52293 , n52294 );
xor ( n52296 , n52281 , n52295 );
xor ( n52297 , n52296 , n52089 );
xor ( n52298 , n52297 , n51853 );
xor ( n52299 , n52296 , n52089 );
and ( n52300 , n52299 , n51853 );
and ( n52301 , n52296 , n52089 );
or ( n52302 , n52300 , n52301 );
xor ( n52303 , n51884 , n52199 );
xor ( n52304 , n52303 , n51942 );
xor ( n52305 , n51884 , n52199 );
and ( n52306 , n52305 , n51942 );
and ( n52307 , n51884 , n52199 );
or ( n52308 , n52306 , n52307 );
xor ( n52309 , n52250 , n52298 );
xor ( n52310 , n52309 , n51948 );
xor ( n52311 , n52250 , n52298 );
and ( n52312 , n52311 , n51948 );
and ( n52313 , n52250 , n52298 );
or ( n52314 , n52312 , n52313 );
xor ( n52315 , n52304 , n51954 );
xor ( n52316 , n52315 , n52310 );
xor ( n52317 , n52304 , n51954 );
and ( n52318 , n52317 , n52310 );
and ( n52319 , n52304 , n51954 );
or ( n52320 , n52318 , n52319 );
xor ( n52321 , n52172 , n52194 );
and ( n52322 , n52321 , n51706 );
and ( n52323 , n52172 , n52194 );
or ( n52324 , n52322 , n52323 );
xor ( n52325 , n52238 , n52245 );
and ( n52326 , n52325 , n51735 );
and ( n52327 , n52238 , n52245 );
or ( n52328 , n52326 , n52327 );
xor ( n52329 , n51964 , n52264 );
and ( n52330 , n52329 , n52279 );
and ( n52331 , n51964 , n52264 );
or ( n52332 , n52330 , n52331 );
xor ( n52333 , n52025 , n52068 );
and ( n52334 , n52333 , n52086 );
and ( n52335 , n52025 , n52068 );
or ( n52336 , n52334 , n52335 );
xor ( n52337 , n52137 , n52148 );
and ( n52338 , n52337 , n52159 );
and ( n52339 , n52137 , n52148 );
or ( n52340 , n52338 , n52339 );
xor ( n52341 , n52196 , n51968 );
and ( n52342 , n52341 , n51972 );
and ( n52343 , n52196 , n51968 );
or ( n52344 , n52342 , n52343 );
xor ( n52345 , n51976 , n52280 );
and ( n52346 , n52345 , n52295 );
and ( n52347 , n51976 , n52280 );
or ( n52348 , n52346 , n52347 );
xor ( n52349 , n52216 , n52227 );
and ( n52350 , n52349 , n52247 );
and ( n52351 , n52216 , n52227 );
or ( n52352 , n52350 , n52351 );
not ( n52353 , n48277 );
not ( n52354 , n48456 );
not ( n52355 , n48980 );
or ( n52356 , n52354 , n52355 );
nand ( n52357 , n48983 , n48970 );
nand ( n52358 , n52356 , n52357 );
not ( n52359 , n52358 );
or ( n52360 , n52353 , n52359 );
nand ( n52361 , n49421 , n52180 );
nand ( n52362 , n52360 , n52361 );
not ( n52363 , n52190 );
not ( n52364 , n49979 );
or ( n52365 , n52363 , n52364 );
not ( n52366 , n51792 );
not ( n52367 , n49110 );
or ( n52368 , n52366 , n52367 );
nand ( n52369 , n49111 , n48829 );
nand ( n52370 , n52368 , n52369 );
nand ( n52371 , n52370 , n49288 );
nand ( n52372 , n52365 , n52371 );
xor ( n52373 , n52362 , n52372 );
not ( n52374 , n49116 );
not ( n52375 , n52006 );
or ( n52376 , n52374 , n52375 );
buf ( n52377 , n47476 );
not ( n52378 , n52377 );
not ( n52379 , n51193 );
not ( n52380 , n52379 );
not ( n52381 , n52380 );
or ( n52382 , n52378 , n52381 );
nand ( n52383 , n41415 , n49628 );
nand ( n52384 , n52382 , n52383 );
nand ( n52385 , n52384 , n52004 );
nand ( n52386 , n52376 , n52385 );
xor ( n52387 , n52373 , n52386 );
xor ( n52388 , n52362 , n52372 );
and ( n52389 , n52388 , n52386 );
and ( n52390 , n52362 , n52372 );
or ( n52391 , n52389 , n52390 );
not ( n52392 , n47873 );
not ( n52393 , n52018 );
or ( n52394 , n52392 , n52393 );
and ( n52395 , n41683 , n48235 );
not ( n52396 , n41683 );
and ( n52397 , n52396 , n47794 );
or ( n52398 , n52395 , n52397 );
nand ( n52399 , n48240 , n52398 );
nand ( n52400 , n52394 , n52399 );
not ( n52401 , n52040 );
not ( n52402 , n49014 );
or ( n52403 , n52401 , n52402 );
not ( n52404 , n51671 );
not ( n52405 , n49092 );
or ( n52406 , n52404 , n52405 );
nand ( n52407 , n48705 , n51670 );
nand ( n52408 , n52406 , n52407 );
nand ( n52409 , n49737 , n52408 );
nand ( n52410 , n52403 , n52409 );
xor ( n52411 , n52400 , n52410 );
not ( n52412 , n47148 );
not ( n52413 , n48856 );
not ( n52414 , n41667 );
not ( n52415 , n52414 );
or ( n52416 , n52413 , n52415 );
nand ( n52417 , n41668 , n51724 );
nand ( n52418 , n52416 , n52417 );
not ( n52419 , n52418 );
or ( n52420 , n52412 , n52419 );
buf ( n52421 , n51368 );
nand ( n52422 , n51999 , n52421 );
nand ( n52423 , n52420 , n52422 );
xor ( n52424 , n52411 , n52423 );
xor ( n52425 , n52400 , n52410 );
and ( n52426 , n52425 , n52423 );
and ( n52427 , n52400 , n52410 );
or ( n52428 , n52426 , n52427 );
not ( n52429 , n50659 );
not ( n52430 , n52214 );
or ( n52431 , n52429 , n52430 );
not ( n52432 , n40628 );
and ( n52433 , n46072 , n52432 );
not ( n52434 , n46072 );
and ( n52435 , n52434 , n40626 );
or ( n52436 , n52433 , n52435 );
nand ( n52437 , n52436 , n44004 );
nand ( n52438 , n52431 , n52437 );
not ( n52439 , n46267 );
not ( n52440 , n52291 );
or ( n52441 , n52439 , n52440 );
not ( n52442 , n46425 );
not ( n52443 , n40733 );
or ( n52444 , n52442 , n52443 );
nand ( n52445 , n51929 , n46422 );
nand ( n52446 , n52444 , n52445 );
nand ( n52447 , n52446 , n49026 );
nand ( n52448 , n52441 , n52447 );
xor ( n52449 , n52438 , n52448 );
not ( n52450 , n37552 );
not ( n52451 , n36286 );
or ( n52452 , n52450 , n52451 );
and ( n52453 , n37512 , n37515 );
nor ( n52454 , n52453 , n37518 );
nand ( n52455 , n52452 , n52454 );
nand ( n52456 , n37511 , n34041 );
not ( n52457 , n52456 );
and ( n52458 , n52455 , n52457 );
not ( n52459 , n52455 );
and ( n52460 , n52459 , n52456 );
nor ( n52461 , n52458 , n52460 );
not ( n52462 , n52461 );
not ( n52463 , n52120 );
or ( n52464 , n52462 , n52463 );
not ( n52465 , n52461 );
nand ( n52466 , n52106 , n52465 );
nand ( n52467 , n52464 , n52466 );
buf ( n52468 , n52467 );
buf ( n52469 , n52468 );
not ( n52470 , n52469 );
nor ( n52471 , n52470 , n46441 );
xor ( n52472 , n52471 , n52029 );
xor ( n52473 , n52472 , n52072 );
xor ( n52474 , n52449 , n52473 );
xor ( n52475 , n52438 , n52448 );
and ( n52476 , n52475 , n52473 );
and ( n52477 , n52438 , n52448 );
or ( n52478 , n52476 , n52477 );
xor ( n52479 , n52340 , n52344 );
not ( n52480 , n52135 );
buf ( n52481 , n52124 );
not ( n52482 , n52481 );
not ( n52483 , n52482 );
or ( n52484 , n52480 , n52483 );
not ( n52485 , n46037 );
not ( n52486 , n52109 );
not ( n52487 , n52486 );
not ( n52488 , n52487 );
or ( n52489 , n52485 , n52488 );
not ( n52490 , n52110 );
nand ( n52491 , n52490 , n47306 );
nand ( n52492 , n52489 , n52491 );
nand ( n52493 , n52492 , n51766 );
nand ( n52494 , n52484 , n52493 );
xor ( n52495 , n52494 , n52324 );
xor ( n52496 , n52495 , n52328 );
xor ( n52497 , n52479 , n52496 );
xor ( n52498 , n52340 , n52344 );
and ( n52499 , n52498 , n52496 );
and ( n52500 , n52340 , n52344 );
or ( n52501 , n52499 , n52500 );
not ( n52502 , n52065 );
not ( n52503 , n51234 );
or ( n52504 , n52502 , n52503 );
not ( n52505 , n51204 );
not ( n52506 , n50292 );
or ( n52507 , n52505 , n52506 );
nand ( n52508 , n49618 , n48860 );
nand ( n52509 , n52507 , n52508 );
nand ( n52510 , n52509 , n49789 );
nand ( n52511 , n52504 , n52510 );
not ( n52512 , n52170 );
not ( n52513 , n50580 );
or ( n52514 , n52512 , n52513 );
not ( n52515 , n48898 );
not ( n52516 , n50163 );
or ( n52517 , n52515 , n52516 );
nand ( n52518 , n50304 , n48897 );
nand ( n52519 , n52517 , n52518 );
nand ( n52520 , n52519 , n51452 );
nand ( n52521 , n52514 , n52520 );
xor ( n52522 , n52511 , n52521 );
and ( n52523 , n52182 , n52193 );
xor ( n52524 , n52522 , n52523 );
not ( n52525 , n52157 );
not ( n52526 , n50910 );
not ( n52527 , n52526 );
or ( n52528 , n52525 , n52527 );
not ( n52529 , n47227 );
not ( n52530 , n50899 );
or ( n52531 , n52529 , n52530 );
nand ( n52532 , n50898 , n47589 );
nand ( n52533 , n52531 , n52532 );
nand ( n52534 , n52533 , n51223 );
nand ( n52535 , n52528 , n52534 );
xor ( n52536 , n52524 , n52535 );
not ( n52537 , n52146 );
not ( n52538 , n52139 );
or ( n52539 , n52537 , n52538 );
not ( n52540 , n47646 );
not ( n52541 , n51504 );
or ( n52542 , n52540 , n52541 );
nand ( n52543 , n51818 , n47650 );
nand ( n52544 , n52542 , n52543 );
nand ( n52545 , n51533 , n52544 );
nand ( n52546 , n52539 , n52545 );
xor ( n52547 , n52536 , n52546 );
not ( n52548 , n47827 );
not ( n52549 , n46650 );
not ( n52550 , n51841 );
or ( n52551 , n52549 , n52550 );
nand ( n52552 , n40691 , n48078 );
nand ( n52553 , n52551 , n52552 );
not ( n52554 , n52553 );
or ( n52555 , n52548 , n52554 );
nand ( n52556 , n52082 , n51157 );
nand ( n52557 , n52555 , n52556 );
xor ( n52558 , n52332 , n52557 );
xor ( n52559 , n52558 , n52336 );
xor ( n52560 , n52547 , n52559 );
xor ( n52561 , n52560 , n52352 );
xor ( n52562 , n52547 , n52559 );
and ( n52563 , n52562 , n52352 );
and ( n52564 , n52547 , n52559 );
or ( n52565 , n52563 , n52564 );
not ( n52566 , n46564 );
not ( n52567 , n52225 );
or ( n52568 , n52566 , n52567 );
not ( n52569 , n47508 );
not ( n52570 , n51916 );
not ( n52571 , n52570 );
or ( n52572 , n52569 , n52571 );
nand ( n52573 , n40526 , n51577 );
nand ( n52574 , n52572 , n52573 );
nand ( n52575 , n52574 , n49832 );
nand ( n52576 , n52568 , n52575 );
not ( n52577 , n48989 );
not ( n52578 , n52262 );
or ( n52579 , n52577 , n52578 );
not ( n52580 , n49500 );
not ( n52581 , n49545 );
or ( n52582 , n52580 , n52581 );
nand ( n52583 , n49549 , n47979 );
nand ( n52584 , n52582 , n52583 );
nand ( n52585 , n52584 , n47384 );
nand ( n52586 , n52579 , n52585 );
not ( n52587 , n51865 );
not ( n52588 , n49707 );
not ( n52589 , n49001 );
not ( n52590 , n52589 );
or ( n52591 , n52588 , n52590 );
not ( n52592 , n48997 );
nand ( n52593 , n52592 , n51351 );
nand ( n52594 , n52591 , n52593 );
not ( n52595 , n52594 );
or ( n52596 , n52587 , n52595 );
nand ( n52597 , n52275 , n49713 );
nand ( n52598 , n52596 , n52597 );
xor ( n52599 , n52586 , n52598 );
xor ( n52600 , n52599 , n52424 );
xor ( n52601 , n52576 , n52600 );
not ( n52602 , n52043 );
not ( n52603 , n50232 );
not ( n52604 , n48951 );
or ( n52605 , n52603 , n52604 );
nand ( n52606 , n41407 , n52048 );
nand ( n52607 , n52605 , n52606 );
not ( n52608 , n52607 );
or ( n52609 , n52602 , n52608 );
nand ( n52610 , n52050 , n50242 );
nand ( n52611 , n52609 , n52610 );
not ( n52612 , n47407 );
not ( n52613 , n52234 );
or ( n52614 , n52612 , n52613 );
not ( n52615 , n51545 );
not ( n52616 , n41037 );
or ( n52617 , n52615 , n52616 );
nand ( n52618 , n41036 , n48727 );
nand ( n52619 , n52617 , n52618 );
nand ( n52620 , n52619 , n48929 );
nand ( n52621 , n52614 , n52620 );
xor ( n52622 , n52611 , n52621 );
xor ( n52623 , n52622 , n52387 );
xor ( n52624 , n52601 , n52623 );
xor ( n52625 , n52348 , n52624 );
xor ( n52626 , n52625 , n52474 );
xor ( n52627 , n52348 , n52624 );
and ( n52628 , n52627 , n52474 );
and ( n52629 , n52348 , n52624 );
or ( n52630 , n52628 , n52629 );
xor ( n52631 , n52093 , n52497 );
xor ( n52632 , n52631 , n52203 );
xor ( n52633 , n52093 , n52497 );
and ( n52634 , n52633 , n52203 );
and ( n52635 , n52093 , n52497 );
or ( n52636 , n52634 , n52635 );
xor ( n52637 , n52561 , n52254 );
xor ( n52638 , n52637 , n52626 );
xor ( n52639 , n52561 , n52254 );
and ( n52640 , n52639 , n52626 );
and ( n52641 , n52561 , n52254 );
or ( n52642 , n52640 , n52641 );
xor ( n52643 , n52302 , n52308 );
xor ( n52644 , n52643 , n52632 );
xor ( n52645 , n52302 , n52308 );
and ( n52646 , n52645 , n52632 );
and ( n52647 , n52302 , n52308 );
or ( n52648 , n52646 , n52647 );
xor ( n52649 , n52638 , n52314 );
xor ( n52650 , n52649 , n52644 );
xor ( n52651 , n52638 , n52314 );
and ( n52652 , n52651 , n52644 );
and ( n52653 , n52638 , n52314 );
or ( n52654 , n52652 , n52653 );
xor ( n52655 , n52511 , n52521 );
and ( n52656 , n52655 , n52523 );
and ( n52657 , n52511 , n52521 );
or ( n52658 , n52656 , n52657 );
xor ( n52659 , n52611 , n52621 );
and ( n52660 , n52659 , n52387 );
and ( n52661 , n52611 , n52621 );
or ( n52662 , n52660 , n52661 );
xor ( n52663 , n52471 , n52029 );
and ( n52664 , n52663 , n52072 );
and ( n52665 , n52471 , n52029 );
or ( n52666 , n52664 , n52665 );
xor ( n52667 , n52586 , n52598 );
and ( n52668 , n52667 , n52424 );
and ( n52669 , n52586 , n52598 );
or ( n52670 , n52668 , n52669 );
xor ( n52671 , n52524 , n52535 );
and ( n52672 , n52671 , n52546 );
and ( n52673 , n52524 , n52535 );
or ( n52674 , n52672 , n52673 );
xor ( n52675 , n52494 , n52324 );
and ( n52676 , n52675 , n52328 );
and ( n52677 , n52494 , n52324 );
or ( n52678 , n52676 , n52677 );
xor ( n52679 , n52332 , n52557 );
and ( n52680 , n52679 , n52336 );
and ( n52681 , n52332 , n52557 );
or ( n52682 , n52680 , n52681 );
xor ( n52683 , n52576 , n52600 );
and ( n52684 , n52683 , n52623 );
and ( n52685 , n52576 , n52600 );
or ( n52686 , n52684 , n52685 );
not ( n52687 , n47873 );
not ( n52688 , n52398 );
or ( n52689 , n52687 , n52688 );
or ( n52690 , n30929 , n47795 );
nand ( n52691 , n30929 , n48235 );
nand ( n52692 , n52690 , n52691 );
nand ( n52693 , n52692 , n47881 );
nand ( n52694 , n52689 , n52693 );
not ( n52695 , n47139 );
not ( n52696 , n52418 );
or ( n52697 , n52695 , n52696 );
not ( n52698 , n51723 );
not ( n52699 , n41530 );
or ( n52700 , n52698 , n52699 );
nand ( n52701 , n48779 , n48857 );
nand ( n52702 , n52700 , n52701 );
nand ( n52703 , n52702 , n47148 );
nand ( n52704 , n52697 , n52703 );
xor ( n52705 , n52694 , n52704 );
not ( n52706 , n52408 );
not ( n52707 , n48755 );
or ( n52708 , n52706 , n52707 );
not ( n52709 , n48223 );
not ( n52710 , n49092 );
or ( n52711 , n52709 , n52710 );
not ( n52712 , n48223 );
nand ( n52713 , n49093 , n52712 );
nand ( n52714 , n52711 , n52713 );
nand ( n52715 , n49022 , n52714 );
nand ( n52716 , n52708 , n52715 );
xor ( n52717 , n52705 , n52716 );
xor ( n52718 , n52694 , n52704 );
and ( n52719 , n52718 , n52716 );
and ( n52720 , n52694 , n52704 );
or ( n52721 , n52719 , n52720 );
buf ( n52722 , n48451 );
not ( n52723 , n52722 );
not ( n52724 , n52723 );
not ( n52725 , n48971 );
not ( n52726 , n47510 );
or ( n52727 , n52725 , n52726 );
buf ( n52728 , n48967 );
nand ( n52729 , n47918 , n52728 );
nand ( n52730 , n52727 , n52729 );
not ( n52731 , n52730 );
or ( n52732 , n52724 , n52731 );
nand ( n52733 , n52358 , n50176 );
nand ( n52734 , n52732 , n52733 );
not ( n52735 , n52509 );
buf ( n52736 , n49779 );
not ( n52737 , n52736 );
or ( n52738 , n52735 , n52737 );
not ( n52739 , n49624 );
not ( n52740 , n49618 );
not ( n52741 , n52740 );
or ( n52742 , n52739 , n52741 );
nand ( n52743 , n49619 , n49630 );
nand ( n52744 , n52742 , n52743 );
nand ( n52745 , n52744 , n50078 );
nand ( n52746 , n52738 , n52745 );
xor ( n52747 , n52734 , n52746 );
not ( n52748 , n52519 );
not ( n52749 , n50320 );
not ( n52750 , n52749 );
or ( n52751 , n52748 , n52750 );
not ( n52752 , n47765 );
not ( n52753 , n50943 );
or ( n52754 , n52752 , n52753 );
nand ( n52755 , n51250 , n48589 );
nand ( n52756 , n52754 , n52755 );
buf ( n52757 , n49920 );
nand ( n52758 , n52756 , n52757 );
nand ( n52759 , n52751 , n52758 );
xor ( n52760 , n52747 , n52759 );
xor ( n52761 , n52734 , n52746 );
and ( n52762 , n52761 , n52759 );
and ( n52763 , n52734 , n52746 );
or ( n52764 , n52762 , n52763 );
not ( n52765 , n48929 );
not ( n52766 , n47803 );
not ( n52767 , n41131 );
not ( n52768 , n52767 );
or ( n52769 , n52766 , n52768 );
nand ( n52770 , n41132 , n50634 );
nand ( n52771 , n52769 , n52770 );
not ( n52772 , n52771 );
or ( n52773 , n52765 , n52772 );
nand ( n52774 , n52619 , n47407 );
nand ( n52775 , n52773 , n52774 );
xor ( n52776 , n52658 , n52775 );
not ( n52777 , n52533 );
not ( n52778 , n52526 );
or ( n52779 , n52777 , n52778 );
not ( n52780 , n49654 );
not ( n52781 , n51465 );
not ( n52782 , n52781 );
or ( n52783 , n52780 , n52782 );
not ( n52784 , n52165 );
nand ( n52785 , n52784 , n50898 );
nand ( n52786 , n52783 , n52785 );
nand ( n52787 , n52786 , n50921 );
nand ( n52788 , n52779 , n52787 );
xor ( n52789 , n52776 , n52788 );
not ( n52790 , n49713 );
not ( n52791 , n52594 );
or ( n52792 , n52790 , n52791 );
not ( n52793 , n52267 );
not ( n52794 , n49837 );
or ( n52795 , n52793 , n52794 );
not ( n52796 , n49209 );
not ( n52797 , n52796 );
nand ( n52798 , n52797 , n48661 );
nand ( n52799 , n52795 , n52798 );
nand ( n52800 , n52799 , n51865 );
nand ( n52801 , n52792 , n52800 );
xor ( n52802 , n52801 , n52717 );
xor ( n52803 , n52802 , n52760 );
xor ( n52804 , n52789 , n52803 );
xor ( n52805 , n52804 , n52674 );
xor ( n52806 , n52789 , n52803 );
and ( n52807 , n52806 , n52674 );
and ( n52808 , n52789 , n52803 );
or ( n52809 , n52807 , n52808 );
not ( n52810 , n52544 );
not ( n52811 , n51525 );
or ( n52812 , n52810 , n52811 );
not ( n52813 , n49734 );
not ( n52814 , n51566 );
or ( n52815 , n52813 , n52814 );
not ( n52816 , n51566 );
nand ( n52817 , n52816 , n47821 );
nand ( n52818 , n52815 , n52817 );
nand ( n52819 , n52818 , n51533 );
nand ( n52820 , n52812 , n52819 );
nor ( n52821 , n37513 , n37551 );
not ( n52822 , n52821 );
not ( n52823 , n36286 );
or ( n52824 , n52822 , n52823 );
nand ( n52825 , n52824 , n37522 );
not ( n52826 , n34023 );
not ( n52827 , n34028 );
or ( n52828 , n52826 , n52827 );
nand ( n52829 , n52828 , n34045 );
and ( n52830 , n52825 , n52829 );
not ( n52831 , n52825 );
not ( n52832 , n52829 );
and ( n52833 , n52831 , n52832 );
nor ( n52834 , n52830 , n52833 );
not ( n52835 , n52834 );
buf ( n52836 , n52835 );
not ( n52837 , n52836 );
and ( n52838 , n46441 , n52837 );
not ( n52839 , n46441 );
not ( n52840 , n52837 );
buf ( n52841 , n52840 );
and ( n52842 , n52839 , n52841 );
nor ( n52843 , n52838 , n52842 );
not ( n52844 , n52843 );
not ( n52845 , n52835 );
nand ( n52846 , n52845 , n52465 );
nand ( n52847 , n52835 , n52461 );
nand ( n52848 , n52846 , n52847 );
not ( n52849 , n52848 );
xor ( n52850 , n52106 , n52465 );
nand ( n52851 , n52849 , n52850 );
not ( n52852 , n52851 );
buf ( n52853 , n52852 );
buf ( n52854 , n52853 );
not ( n52855 , n52854 );
or ( n52856 , n52844 , n52855 );
and ( n52857 , n52841 , n48766 );
not ( n52858 , n52841 );
and ( n52859 , n52858 , n50914 );
or ( n52860 , n52857 , n52859 );
nand ( n52861 , n52860 , n52469 );
nand ( n52862 , n52856 , n52861 );
xor ( n52863 , n52820 , n52862 );
not ( n52864 , n52492 );
not ( n52865 , n52482 );
or ( n52866 , n52864 , n52865 );
not ( n52867 , n46273 );
not ( n52868 , n52130 );
or ( n52869 , n52867 , n52868 );
not ( n52870 , n52129 );
not ( n52871 , n52870 );
or ( n52872 , n52871 , n46273 );
nand ( n52873 , n52869 , n52872 );
nand ( n52874 , n52873 , n51766 );
nand ( n52875 , n52866 , n52874 );
xor ( n52876 , n52863 , n52875 );
xor ( n52877 , n52678 , n52876 );
xor ( n52878 , n52877 , n52682 );
xor ( n52879 , n52678 , n52876 );
and ( n52880 , n52879 , n52682 );
and ( n52881 , n52678 , n52876 );
or ( n52882 , n52880 , n52881 );
xor ( n52883 , n52662 , n52666 );
xor ( n52884 , n52883 , n52670 );
xor ( n52885 , n52686 , n52884 );
xor ( n52886 , n52885 , n52478 );
xor ( n52887 , n52686 , n52884 );
and ( n52888 , n52887 , n52478 );
and ( n52889 , n52686 , n52884 );
or ( n52890 , n52888 , n52889 );
not ( n52891 , n46188 );
not ( n52892 , n46425 );
buf ( n52893 , n40768 );
not ( n52894 , n52893 );
not ( n52895 , n52894 );
or ( n52896 , n52892 , n52895 );
nand ( n52897 , n52893 , n46422 );
nand ( n52898 , n52896 , n52897 );
not ( n52899 , n52898 );
or ( n52900 , n52891 , n52899 );
nand ( n52901 , n52446 , n46267 );
nand ( n52902 , n52900 , n52901 );
not ( n52903 , n50659 );
not ( n52904 , n52436 );
or ( n52905 , n52903 , n52904 );
not ( n52906 , n40635 );
not ( n52907 , n52906 );
not ( n52908 , n52907 );
nand ( n52909 , n52908 , n46071 );
not ( n52910 , n52906 );
nand ( n52911 , n52910 , n46072 );
nand ( n52912 , n52909 , n52911 , n44004 );
nand ( n52913 , n52905 , n52912 );
xor ( n52914 , n52902 , n52913 );
not ( n52915 , n47384 );
not ( n52916 , n49805 );
not ( n52917 , n52916 );
not ( n52918 , n52917 );
not ( n52919 , n49500 );
or ( n52920 , n52918 , n52919 );
or ( n52921 , n52917 , n49500 );
nand ( n52922 , n52920 , n52921 );
not ( n52923 , n52922 );
or ( n52924 , n52915 , n52923 );
nand ( n52925 , n52584 , n49252 );
nand ( n52926 , n52924 , n52925 );
xor ( n52927 , n52926 , n52391 );
xor ( n52928 , n52927 , n52428 );
xor ( n52929 , n52914 , n52928 );
not ( n52930 , n48073 );
not ( n52931 , n50263 );
not ( n52932 , n50958 );
or ( n52933 , n52931 , n52932 );
nand ( n52934 , n40677 , n50087 );
nand ( n52935 , n52933 , n52934 );
not ( n52936 , n52935 );
or ( n52937 , n52930 , n52936 );
nand ( n52938 , n52553 , n48295 );
nand ( n52939 , n52937 , n52938 );
not ( n52940 , n52370 );
not ( n52941 , n51337 );
or ( n52942 , n52940 , n52941 );
not ( n52943 , n52033 );
not ( n52944 , n49283 );
or ( n52945 , n52943 , n52944 );
nand ( n52946 , n49452 , n52038 );
nand ( n52947 , n52945 , n52946 );
nand ( n52948 , n52191 , n52947 );
nand ( n52949 , n52942 , n52948 );
not ( n52950 , n52004 );
not ( n52951 , n52377 );
not ( n52952 , n49756 );
or ( n52953 , n52951 , n52952 );
not ( n52954 , n51995 );
nand ( n52955 , n52954 , n49628 );
nand ( n52956 , n52953 , n52955 );
not ( n52957 , n52956 );
or ( n52958 , n52950 , n52957 );
nand ( n52959 , n52384 , n48894 );
nand ( n52960 , n52958 , n52959 );
xor ( n52961 , n52949 , n52960 );
not ( n52962 , n50239 );
not ( n52963 , n52962 );
and ( n52964 , n49820 , n48645 );
not ( n52965 , n49820 );
and ( n52966 , n52965 , n52048 );
or ( n52967 , n52964 , n52966 );
not ( n52968 , n52967 );
or ( n52969 , n52963 , n52968 );
not ( n52970 , n50241 );
nand ( n52971 , n52607 , n52970 );
nand ( n52972 , n52969 , n52971 );
xor ( n52973 , n52961 , n52972 );
not ( n52974 , n46440 );
not ( n52975 , n52461 );
or ( n52976 , n52974 , n52975 );
nand ( n52977 , n52976 , n52871 );
nand ( n52978 , n52465 , n46441 );
and ( n52979 , n52977 , n52978 );
not ( n52980 , n52841 );
nor ( n52981 , n52979 , n52980 );
xor ( n52982 , n52973 , n52981 );
xor ( n52983 , n52939 , n52982 );
not ( n52984 , n46564 );
not ( n52985 , n52574 );
or ( n52986 , n52984 , n52985 );
not ( n52987 , n47508 );
not ( n52988 , n52208 );
or ( n52989 , n52987 , n52988 );
not ( n52990 , n47508 );
nand ( n52991 , n52212 , n52990 );
nand ( n52992 , n52989 , n52991 );
not ( n52993 , n52992 );
or ( n52994 , n52993 , n50840 );
nand ( n52995 , n52986 , n52994 );
xor ( n52996 , n52983 , n52995 );
xor ( n52997 , n52929 , n52996 );
xor ( n52998 , n52997 , n52501 );
xor ( n52999 , n52929 , n52996 );
and ( n53000 , n52999 , n52501 );
and ( n53001 , n52929 , n52996 );
or ( n53002 , n53000 , n53001 );
xor ( n53003 , n52805 , n52878 );
xor ( n53004 , n53003 , n52565 );
xor ( n53005 , n52805 , n52878 );
and ( n53006 , n53005 , n52565 );
and ( n53007 , n52805 , n52878 );
or ( n53008 , n53006 , n53007 );
xor ( n53009 , n52630 , n52886 );
xor ( n53010 , n53009 , n52998 );
xor ( n53011 , n52630 , n52886 );
and ( n53012 , n53011 , n52998 );
and ( n53013 , n52630 , n52886 );
or ( n53014 , n53012 , n53013 );
xor ( n53015 , n52636 , n53004 );
xor ( n53016 , n53015 , n52642 );
xor ( n53017 , n52636 , n53004 );
and ( n53018 , n53017 , n52642 );
and ( n53019 , n52636 , n53004 );
or ( n53020 , n53018 , n53019 );
xor ( n53021 , n53010 , n52648 );
xor ( n53022 , n53021 , n53016 );
xor ( n53023 , n53010 , n52648 );
and ( n53024 , n53023 , n53016 );
and ( n53025 , n53010 , n52648 );
or ( n53026 , n53024 , n53025 );
xor ( n53027 , n52961 , n52972 );
and ( n53028 , n53027 , n52981 );
and ( n53029 , n52961 , n52972 );
or ( n53030 , n53028 , n53029 );
xor ( n53031 , n52926 , n52391 );
and ( n53032 , n53031 , n52428 );
and ( n53033 , n52926 , n52391 );
or ( n53034 , n53032 , n53033 );
xor ( n53035 , n52801 , n52717 );
and ( n53036 , n53035 , n52760 );
and ( n53037 , n52801 , n52717 );
or ( n53038 , n53036 , n53037 );
xor ( n53039 , n52658 , n52775 );
and ( n53040 , n53039 , n52788 );
and ( n53041 , n52658 , n52775 );
or ( n53042 , n53040 , n53041 );
xor ( n53043 , n52820 , n52862 );
and ( n53044 , n53043 , n52875 );
and ( n53045 , n52820 , n52862 );
or ( n53046 , n53044 , n53045 );
xor ( n53047 , n52662 , n52666 );
and ( n53048 , n53047 , n52670 );
and ( n53049 , n52662 , n52666 );
or ( n53050 , n53048 , n53049 );
xor ( n53051 , n52939 , n52982 );
and ( n53052 , n53051 , n52995 );
and ( n53053 , n52939 , n52982 );
or ( n53054 , n53052 , n53053 );
xor ( n53055 , n52902 , n52913 );
and ( n53056 , n53055 , n52928 );
and ( n53057 , n52902 , n52913 );
or ( n53058 , n53056 , n53057 );
not ( n53059 , n52947 );
not ( n53060 , n49276 );
or ( n53061 , n53059 , n53060 );
not ( n53062 , n51671 );
not ( n53063 , n49259 );
or ( n53064 , n53062 , n53063 );
nand ( n53065 , n49111 , n51670 );
nand ( n53066 , n53064 , n53065 );
nand ( n53067 , n53066 , n52191 );
nand ( n53068 , n53061 , n53067 );
not ( n53069 , n48240 );
not ( n53070 , n47855 );
not ( n53071 , n51193 );
or ( n53072 , n53070 , n53071 );
nand ( n53073 , n52016 , n41415 );
nand ( n53074 , n53072 , n53073 );
not ( n53075 , n53074 );
or ( n53076 , n53069 , n53075 );
nand ( n53077 , n52692 , n47873 );
nand ( n53078 , n53076 , n53077 );
xor ( n53079 , n53068 , n53078 );
not ( n53080 , n52004 );
not ( n53081 , n52377 );
not ( n53082 , n48118 );
or ( n53083 , n53081 , n53082 );
nand ( n53084 , n41668 , n51782 );
nand ( n53085 , n53083 , n53084 );
not ( n53086 , n53085 );
or ( n53087 , n53080 , n53086 );
nand ( n53088 , n52956 , n49116 );
nand ( n53089 , n53087 , n53088 );
xor ( n53090 , n53079 , n53089 );
xor ( n53091 , n53068 , n53078 );
and ( n53092 , n53091 , n53089 );
and ( n53093 , n53068 , n53078 );
or ( n53094 , n53092 , n53093 );
not ( n53095 , n52714 );
or ( n53096 , n48756 , n53095 );
and ( n53097 , n48758 , n47318 );
not ( n53098 , n48758 );
and ( n53099 , n53098 , n30964 );
or ( n53100 , n53097 , n53099 );
not ( n53101 , n53100 );
or ( n53102 , n53101 , n49485 );
nand ( n53103 , n53096 , n53102 );
not ( n53104 , n49420 );
not ( n53105 , n53104 );
not ( n53106 , n52730 );
or ( n53107 , n53105 , n53106 );
not ( n53108 , n48456 );
not ( n53109 , n48523 );
or ( n53110 , n53108 , n53109 );
not ( n53111 , n831 );
not ( n53112 , n18833 );
or ( n53113 , n53111 , n53112 );
nand ( n53114 , n53113 , n32079 );
nand ( n53115 , n53114 , n48967 );
nand ( n53116 , n53110 , n53115 );
nand ( n53117 , n53116 , n52723 );
nand ( n53118 , n53107 , n53117 );
xor ( n53119 , n53103 , n53118 );
not ( n53120 , n52744 );
not ( n53121 , n52058 );
or ( n53122 , n53120 , n53121 );
not ( n53123 , n51792 );
not ( n53124 , n52740 );
or ( n53125 , n53123 , n53124 );
not ( n53126 , n51792 );
nand ( n53127 , n49619 , n53126 );
nand ( n53128 , n53125 , n53127 );
nand ( n53129 , n53128 , n50078 );
nand ( n53130 , n53122 , n53129 );
xor ( n53131 , n53119 , n53130 );
xor ( n53132 , n53103 , n53118 );
and ( n53133 , n53132 , n53130 );
and ( n53134 , n53103 , n53118 );
or ( n53135 , n53133 , n53134 );
not ( n53136 , n49713 );
not ( n53137 , n52799 );
or ( n53138 , n53136 , n53137 );
not ( n53139 , n49707 );
not ( n53140 , n50007 );
or ( n53141 , n53139 , n53140 );
nand ( n53142 , n49549 , n52273 );
nand ( n53143 , n53141 , n53142 );
nand ( n53144 , n53143 , n51865 );
nand ( n53145 , n53138 , n53144 );
xor ( n53146 , n52721 , n53145 );
xor ( n53147 , n53146 , n53090 );
xor ( n53148 , n53038 , n53147 );
xor ( n53149 , n53131 , n52764 );
not ( n53150 , n52786 );
not ( n53151 , n52526 );
or ( n53152 , n53150 , n53151 );
not ( n53153 , n48898 );
not ( n53154 , n52781 );
or ( n53155 , n53153 , n53154 );
not ( n53156 , n50916 );
nand ( n53157 , n53156 , n48897 );
nand ( n53158 , n53155 , n53157 );
nand ( n53159 , n53158 , n51223 );
nand ( n53160 , n53152 , n53159 );
xor ( n53161 , n53149 , n53160 );
xor ( n53162 , n53148 , n53161 );
xor ( n53163 , n53038 , n53147 );
and ( n53164 , n53163 , n53161 );
and ( n53165 , n53038 , n53147 );
or ( n53166 , n53164 , n53165 );
xor ( n53167 , n53046 , n53042 );
not ( n53168 , n52818 );
not ( n53169 , n51524 );
buf ( n53170 , n53169 );
not ( n53171 , n53170 );
or ( n53172 , n53168 , n53171 );
not ( n53173 , n47227 );
not ( n53174 , n51566 );
or ( n53175 , n53173 , n53174 );
not ( n53176 , n47227 );
nand ( n53177 , n53176 , n51505 );
nand ( n53178 , n53175 , n53177 );
nand ( n53179 , n53178 , n51533 );
nand ( n53180 , n53172 , n53179 );
not ( n53181 , n52860 );
buf ( n53182 , n52853 );
not ( n53183 , n53182 );
or ( n53184 , n53181 , n53183 );
not ( n53185 , n46037 );
not ( n53186 , n52841 );
not ( n53187 , n53186 );
or ( n53188 , n53185 , n53187 );
buf ( n53189 , n52837 );
not ( n53190 , n53189 );
nand ( n53191 , n53190 , n47306 );
nand ( n53192 , n53188 , n53191 );
nand ( n53193 , n53192 , n52469 );
nand ( n53194 , n53184 , n53193 );
xor ( n53195 , n53180 , n53194 );
not ( n53196 , n52873 );
not ( n53197 , n52481 );
not ( n53198 , n53197 );
or ( n53199 , n53196 , n53198 );
not ( n53200 , n47646 );
not ( n53201 , n52487 );
or ( n53202 , n53200 , n53201 );
nand ( n53203 , n52490 , n47650 );
nand ( n53204 , n53202 , n53203 );
nand ( n53205 , n53204 , n51766 );
nand ( n53206 , n53199 , n53205 );
xor ( n53207 , n53195 , n53206 );
xor ( n53208 , n53167 , n53207 );
xor ( n53209 , n53046 , n53042 );
and ( n53210 , n53209 , n53207 );
and ( n53211 , n53046 , n53042 );
or ( n53212 , n53210 , n53211 );
xor ( n53213 , n53054 , n53058 );
not ( n53214 , n52756 );
not ( n53215 , n50580 );
or ( n53216 , n53214 , n53215 );
not ( n53217 , n51204 );
not ( n53218 , n50327 );
or ( n53219 , n53217 , n53218 );
nand ( n53220 , n50304 , n48860 );
nand ( n53221 , n53219 , n53220 );
nand ( n53222 , n53221 , n52757 );
nand ( n53223 , n53216 , n53222 );
not ( n53224 , n47148 );
not ( n53225 , n48856 );
not ( n53226 , n48951 );
or ( n53227 , n53225 , n53226 );
not ( n53228 , n47106 );
nand ( n53229 , n41407 , n53228 );
nand ( n53230 , n53227 , n53229 );
not ( n53231 , n53230 );
or ( n53232 , n53224 , n53231 );
nand ( n53233 , n52702 , n52421 );
nand ( n53234 , n53232 , n53233 );
xor ( n53235 , n53223 , n53234 );
and ( n53236 , n52949 , n52960 );
xor ( n53237 , n53235 , n53236 );
xor ( n53238 , n53237 , n53030 );
xor ( n53239 , n53238 , n53034 );
xor ( n53240 , n53213 , n53239 );
xor ( n53241 , n53054 , n53058 );
and ( n53242 , n53241 , n53239 );
and ( n53243 , n53054 , n53058 );
or ( n53244 , n53242 , n53243 );
xor ( n53245 , n53050 , n53162 );
not ( n53246 , n48929 );
not ( n53247 , n50634 );
not ( n53248 , n40691 );
or ( n53249 , n53247 , n53248 );
nand ( n53250 , n50654 , n47803 );
nand ( n53251 , n53249 , n53250 );
not ( n53252 , n53251 );
or ( n53253 , n53246 , n53252 );
nand ( n53254 , n52771 , n47407 );
nand ( n53255 , n53253 , n53254 );
not ( n53256 , n47827 );
not ( n53257 , n50263 );
not ( n53258 , n51928 );
not ( n53259 , n53258 );
not ( n53260 , n53259 );
or ( n53261 , n53257 , n53260 );
nand ( n53262 , n40734 , n48078 );
nand ( n53263 , n53261 , n53262 );
not ( n53264 , n53263 );
or ( n53265 , n53256 , n53264 );
nand ( n53266 , n52935 , n46776 );
nand ( n53267 , n53265 , n53266 );
xor ( n53268 , n53255 , n53267 );
not ( n53269 , n49832 );
not ( n53270 , n48952 );
not ( n53271 , n40626 );
not ( n53272 , n53271 );
or ( n53273 , n53270 , n53272 );
nand ( n53274 , n40628 , n52990 );
nand ( n53275 , n53273 , n53274 );
not ( n53276 , n53275 );
or ( n53277 , n53269 , n53276 );
nand ( n53278 , n52992 , n46564 );
nand ( n53279 , n53277 , n53278 );
xor ( n53280 , n53268 , n53279 );
xor ( n53281 , n53245 , n53280 );
xor ( n53282 , n53050 , n53162 );
and ( n53283 , n53282 , n53280 );
and ( n53284 , n53050 , n53162 );
or ( n53285 , n53283 , n53284 );
not ( n53286 , n40377 );
and ( n53287 , n46072 , n53286 );
not ( n53288 , n46072 );
not ( n53289 , n40376 );
not ( n53290 , n53289 );
and ( n53291 , n53288 , n53290 );
nor ( n53292 , n53287 , n53291 );
or ( n53293 , n53292 , n45861 );
nand ( n53294 , n52909 , n52911 , n50659 );
nand ( n53295 , n53293 , n53294 );
not ( n53296 , n52043 );
not ( n53297 , n48645 );
not ( n53298 , n52589 );
or ( n53299 , n53297 , n53298 );
nand ( n53300 , n48996 , n52048 );
nand ( n53301 , n53299 , n53300 );
not ( n53302 , n53301 );
or ( n53303 , n53296 , n53302 );
nand ( n53304 , n52967 , n50242 );
nand ( n53305 , n53303 , n53304 );
not ( n53306 , n36617 );
not ( n53307 , n36965 );
or ( n53308 , n53306 , n53307 );
nor ( n53309 , n36612 , n36283 );
nand ( n53310 , n53308 , n53309 );
not ( n53311 , n53310 );
buf ( n53312 , n35286 );
buf ( n53313 , n36283 );
nor ( n53314 , n53312 , n53313 );
nor ( n53315 , n53314 , n34091 );
not ( n53316 , n53315 );
or ( n53317 , n53311 , n53316 );
nand ( n53318 , n53317 , n37502 );
not ( n53319 , n37576 );
and ( n53320 , n53318 , n53319 );
not ( n53321 , n53318 );
and ( n53322 , n53321 , n37576 );
nor ( n53323 , n53320 , n53322 );
xnor ( n53324 , n53323 , n52835 );
not ( n53325 , n53324 );
buf ( n53326 , n53325 );
not ( n53327 , n53326 );
nor ( n53328 , n53327 , n46441 );
xor ( n53329 , n53305 , n53328 );
not ( n53330 , n48989 );
not ( n53331 , n52922 );
or ( n53332 , n53330 , n53331 );
not ( n53333 , n47980 );
not ( n53334 , n50667 );
or ( n53335 , n53333 , n53334 );
nand ( n53336 , n51891 , n47979 );
nand ( n53337 , n53335 , n53336 );
nand ( n53338 , n53337 , n47384 );
nand ( n53339 , n53332 , n53338 );
xor ( n53340 , n53329 , n53339 );
xor ( n53341 , n53295 , n53340 );
not ( n53342 , n52898 );
not ( n53343 , n46267 );
or ( n53344 , n53342 , n53343 );
and ( n53345 , n46425 , n40528 );
not ( n53346 , n46425 );
not ( n53347 , n51913 );
and ( n53348 , n53346 , n53347 );
or ( n53349 , n53345 , n53348 );
not ( n53350 , n53349 );
or ( n53351 , n53350 , n49025 );
nand ( n53352 , n53344 , n53351 );
xor ( n53353 , n53341 , n53352 );
xor ( n53354 , n53353 , n52809 );
xor ( n53355 , n53354 , n53208 );
xor ( n53356 , n53353 , n52809 );
and ( n53357 , n53356 , n53208 );
and ( n53358 , n53353 , n52809 );
or ( n53359 , n53357 , n53358 );
xor ( n53360 , n52882 , n52890 );
xor ( n53361 , n53360 , n53240 );
xor ( n53362 , n52882 , n52890 );
and ( n53363 , n53362 , n53240 );
and ( n53364 , n52882 , n52890 );
or ( n53365 , n53363 , n53364 );
xor ( n53366 , n53002 , n53355 );
xor ( n53367 , n53366 , n53281 );
xor ( n53368 , n53002 , n53355 );
and ( n53369 , n53368 , n53281 );
and ( n53370 , n53002 , n53355 );
or ( n53371 , n53369 , n53370 );
xor ( n53372 , n53008 , n53361 );
xor ( n53373 , n53372 , n53014 );
xor ( n53374 , n53008 , n53361 );
and ( n53375 , n53374 , n53014 );
and ( n53376 , n53008 , n53361 );
or ( n53377 , n53375 , n53376 );
xor ( n53378 , n53367 , n53373 );
xor ( n53379 , n53378 , n53020 );
xor ( n53380 , n53367 , n53373 );
and ( n53381 , n53380 , n53020 );
and ( n53382 , n53367 , n53373 );
or ( n53383 , n53381 , n53382 );
xor ( n53384 , n53223 , n53234 );
and ( n53385 , n53384 , n53236 );
and ( n53386 , n53223 , n53234 );
or ( n53387 , n53385 , n53386 );
xor ( n53388 , n53305 , n53328 );
and ( n53389 , n53388 , n53339 );
and ( n53390 , n53305 , n53328 );
or ( n53391 , n53389 , n53390 );
xor ( n53392 , n52721 , n53145 );
and ( n53393 , n53392 , n53090 );
and ( n53394 , n52721 , n53145 );
or ( n53395 , n53393 , n53394 );
xor ( n53396 , n53131 , n52764 );
and ( n53397 , n53396 , n53160 );
and ( n53398 , n53131 , n52764 );
or ( n53399 , n53397 , n53398 );
xor ( n53400 , n53180 , n53194 );
and ( n53401 , n53400 , n53206 );
and ( n53402 , n53180 , n53194 );
or ( n53403 , n53401 , n53402 );
xor ( n53404 , n53237 , n53030 );
and ( n53405 , n53404 , n53034 );
and ( n53406 , n53237 , n53030 );
or ( n53407 , n53405 , n53406 );
xor ( n53408 , n53255 , n53267 );
and ( n53409 , n53408 , n53279 );
and ( n53410 , n53255 , n53267 );
or ( n53411 , n53409 , n53410 );
xor ( n53412 , n53295 , n53340 );
and ( n53413 , n53412 , n53352 );
and ( n53414 , n53295 , n53340 );
or ( n53415 , n53413 , n53414 );
not ( n53416 , n49116 );
not ( n53417 , n53085 );
or ( n53418 , n53416 , n53417 );
not ( n53419 , n52377 );
not ( n53420 , n41530 );
or ( n53421 , n53419 , n53420 );
nand ( n53422 , n41531 , n49628 );
nand ( n53423 , n53421 , n53422 );
nand ( n53424 , n53423 , n47498 );
nand ( n53425 , n53418 , n53424 );
not ( n53426 , n49737 );
not ( n53427 , n49017 );
not ( n53428 , n49245 );
or ( n53429 , n53427 , n53428 );
not ( n53430 , n47511 );
nand ( n53431 , n53430 , n48704 );
nand ( n53432 , n53429 , n53431 );
not ( n53433 , n53432 );
or ( n53434 , n53426 , n53433 );
nand ( n53435 , n50554 , n53100 );
nand ( n53436 , n53434 , n53435 );
xor ( n53437 , n53425 , n53436 );
not ( n53438 , n52723 );
buf ( n53439 , n48262 );
not ( n53440 , n53439 );
not ( n53441 , n51360 );
or ( n53442 , n53440 , n53441 );
not ( n53443 , n53439 );
nand ( n53444 , n47527 , n53443 );
nand ( n53445 , n53442 , n53444 );
not ( n53446 , n53445 );
or ( n53447 , n53438 , n53446 );
nand ( n53448 , n53116 , n50176 );
nand ( n53449 , n53447 , n53448 );
xor ( n53450 , n53437 , n53449 );
xor ( n53451 , n53425 , n53436 );
and ( n53452 , n53451 , n53449 );
and ( n53453 , n53425 , n53436 );
or ( n53454 , n53452 , n53453 );
not ( n53455 , n53128 );
not ( n53456 , n52736 );
or ( n53457 , n53455 , n53456 );
not ( n53458 , n52033 );
not ( n53459 , n50292 );
or ( n53460 , n53458 , n53459 );
not ( n53461 , n49783 );
nand ( n53462 , n53461 , n52038 );
nand ( n53463 , n53460 , n53462 );
nand ( n53464 , n53463 , n50078 );
nand ( n53465 , n53457 , n53464 );
not ( n53466 , n53221 );
not ( n53467 , n50321 );
or ( n53468 , n53466 , n53467 );
not ( n53469 , n49624 );
not ( n53470 , n50301 );
or ( n53471 , n53469 , n53470 );
nand ( n53472 , n51250 , n49630 );
nand ( n53473 , n53471 , n53472 );
nand ( n53474 , n53473 , n51452 );
nand ( n53475 , n53468 , n53474 );
xor ( n53476 , n53465 , n53475 );
not ( n53477 , n48240 );
not ( n53478 , n47855 );
not ( n53479 , n51995 );
or ( n53480 , n53478 , n53479 );
nand ( n53481 , n41576 , n52016 );
nand ( n53482 , n53480 , n53481 );
not ( n53483 , n53482 );
or ( n53484 , n53477 , n53483 );
nand ( n53485 , n53074 , n52022 );
nand ( n53486 , n53484 , n53485 );
not ( n53487 , n53066 );
not ( n53488 , n50195 );
or ( n53489 , n53487 , n53488 );
not ( n53490 , n48890 );
not ( n53491 , n48223 );
not ( n53492 , n49262 );
not ( n53493 , n53492 );
or ( n53494 , n53491 , n53493 );
nand ( n53495 , n49452 , n46880 );
nand ( n53496 , n53494 , n53495 );
nand ( n53497 , n53490 , n53496 );
nand ( n53498 , n53489 , n53497 );
and ( n53499 , n53486 , n53498 );
not ( n53500 , n53486 );
not ( n53501 , n53498 );
and ( n53502 , n53500 , n53501 );
nor ( n53503 , n53499 , n53502 );
xor ( n53504 , n53476 , n53503 );
xor ( n53505 , n53465 , n53475 );
and ( n53506 , n53505 , n53503 );
and ( n53507 , n53465 , n53475 );
or ( n53508 , n53506 , n53507 );
not ( n53509 , n47384 );
not ( n53510 , n53509 );
not ( n53511 , n53510 );
not ( n53512 , n49500 );
not ( n53513 , n41132 );
not ( n53514 , n53513 );
or ( n53515 , n53512 , n53514 );
nand ( n53516 , n52079 , n47979 );
nand ( n53517 , n53515 , n53516 );
not ( n53518 , n53517 );
or ( n53519 , n53511 , n53518 );
nand ( n53520 , n53337 , n48989 );
nand ( n53521 , n53519 , n53520 );
xor ( n53522 , n53450 , n53521 );
not ( n53523 , n53158 );
not ( n53524 , n52151 );
or ( n53525 , n53523 , n53524 );
not ( n53526 , n47765 );
not ( n53527 , n50899 );
or ( n53528 , n53526 , n53527 );
nand ( n53529 , n51461 , n48589 );
nand ( n53530 , n53528 , n53529 );
nand ( n53531 , n53530 , n51223 );
nand ( n53532 , n53525 , n53531 );
xor ( n53533 , n53522 , n53532 );
xor ( n53534 , n53403 , n53533 );
xor ( n53535 , n53534 , n53399 );
xor ( n53536 , n53403 , n53533 );
and ( n53537 , n53536 , n53399 );
and ( n53538 , n53403 , n53533 );
or ( n53539 , n53537 , n53538 );
not ( n53540 , n53178 );
buf ( n53541 , n51522 );
buf ( n53542 , n51516 );
nor ( n53543 , n53541 , n53542 );
not ( n53544 , n53543 );
or ( n53545 , n53540 , n53544 );
not ( n53546 , n49654 );
not ( n53547 , n51566 );
or ( n53548 , n53546 , n53547 );
not ( n53549 , n51504 );
buf ( n53550 , n53549 );
nand ( n53551 , n53550 , n47368 );
nand ( n53552 , n53548 , n53551 );
nand ( n53553 , n51533 , n53552 );
nand ( n53554 , n53545 , n53553 );
xor ( n53555 , n53554 , n53504 );
not ( n53556 , n53204 );
not ( n53557 , n52125 );
or ( n53558 , n53556 , n53557 );
not ( n53559 , n49734 );
not ( n53560 , n52871 );
or ( n53561 , n53559 , n53560 );
nand ( n53562 , n52490 , n47821 );
nand ( n53563 , n53561 , n53562 );
nand ( n53564 , n51766 , n53563 );
nand ( n53565 , n53558 , n53564 );
xor ( n53566 , n53555 , n53565 );
xor ( n53567 , n53407 , n53566 );
not ( n53568 , n53192 );
not ( n53569 , n53182 );
or ( n53570 , n53568 , n53569 );
buf ( n53571 , n52468 );
not ( n53572 , n46273 );
not ( n53573 , n53189 );
or ( n53574 , n53572 , n53573 );
nand ( n53575 , n52840 , n46824 );
nand ( n53576 , n53574 , n53575 );
nand ( n53577 , n53571 , n53576 );
nand ( n53578 , n53570 , n53577 );
not ( n53579 , n37671 );
not ( n53580 , n51754 );
or ( n53581 , n53579 , n53580 );
nand ( n53582 , n53581 , n37425 );
nand ( n53583 , n33535 , n33540 );
not ( n53584 , n53583 );
and ( n53585 , n53582 , n53584 );
not ( n53586 , n53582 );
and ( n53587 , n53586 , n53583 );
nor ( n53588 , n53585 , n53587 );
buf ( n53589 , n53588 );
buf ( n53590 , n53589 );
not ( n53591 , n53590 );
and ( n53592 , n46440 , n53591 );
not ( n53593 , n46440 );
not ( n53594 , n53589 );
buf ( n53595 , n53594 );
not ( n53596 , n53595 );
and ( n53597 , n53593 , n53596 );
or ( n53598 , n53592 , n53597 );
not ( n53599 , n53598 );
not ( n53600 , n53589 );
not ( n53601 , n53323 );
not ( n53602 , n53601 );
not ( n53603 , n53602 );
and ( n53604 , n53600 , n53603 );
and ( n53605 , n53589 , n53602 );
nor ( n53606 , n53604 , n53605 );
not ( n53607 , n53325 );
nand ( n53608 , n53606 , n53607 );
not ( n53609 , n53608 );
not ( n53610 , n53609 );
or ( n53611 , n53599 , n53610 );
not ( n53612 , n50914 );
not ( n53613 , n53591 );
or ( n53614 , n53612 , n53613 );
not ( n53615 , n53591 );
nand ( n53616 , n53615 , n48766 );
nand ( n53617 , n53614 , n53616 );
buf ( n53618 , n53324 );
not ( n53619 , n53618 );
buf ( n53620 , n53619 );
nand ( n53621 , n53617 , n53620 );
nand ( n53622 , n53611 , n53621 );
xor ( n53623 , n53578 , n53622 );
xor ( n53624 , n53623 , n53387 );
xor ( n53625 , n53567 , n53624 );
xor ( n53626 , n53407 , n53566 );
and ( n53627 , n53626 , n53624 );
and ( n53628 , n53407 , n53566 );
or ( n53629 , n53627 , n53628 );
xor ( n53630 , n53411 , n53415 );
not ( n53631 , n47253 );
not ( n53632 , n53631 );
not ( n53633 , n50263 );
not ( n53634 , n51602 );
or ( n53635 , n53633 , n53634 );
nand ( n53636 , n51601 , n52080 );
nand ( n53637 , n53635 , n53636 );
not ( n53638 , n53637 );
or ( n53639 , n53632 , n53638 );
nand ( n53640 , n53263 , n51157 );
nand ( n53641 , n53639 , n53640 );
xor ( n53642 , n53391 , n53641 );
and ( n53643 , n53602 , n46440 );
nor ( n53644 , n53643 , n52840 );
nor ( n53645 , n53602 , n46440 );
or ( n53646 , n53644 , n53645 );
nand ( n53647 , n53646 , n53615 );
not ( n53648 , n53647 );
xor ( n53649 , n53648 , n53094 );
xor ( n53650 , n53649 , n53135 );
xor ( n53651 , n53642 , n53650 );
xor ( n53652 , n53630 , n53651 );
xor ( n53653 , n53411 , n53415 );
and ( n53654 , n53653 , n53651 );
and ( n53655 , n53411 , n53415 );
or ( n53656 , n53654 , n53655 );
not ( n53657 , n40225 );
not ( n53658 , n46072 );
and ( n53659 , n53657 , n53658 );
not ( n53660 , n40225 );
not ( n53661 , n53660 );
and ( n53662 , n53661 , n46072 );
nor ( n53663 , n53659 , n53662 );
or ( n53664 , n53663 , n45861 );
not ( n53665 , n53292 );
nand ( n53666 , n53665 , n50659 );
nand ( n53667 , n53664 , n53666 );
xor ( n53668 , n53395 , n53667 );
not ( n53669 , n47803 );
not ( n53670 , n50958 );
or ( n53671 , n53669 , n53670 );
nand ( n53672 , n40677 , n48727 );
nand ( n53673 , n53671 , n53672 );
not ( n53674 , n53673 );
buf ( n53675 , n48929 );
not ( n53676 , n53675 );
or ( n53677 , n53674 , n53676 );
nand ( n53678 , n47407 , n53251 );
nand ( n53679 , n53677 , n53678 );
xor ( n53680 , n53668 , n53679 );
not ( n53681 , n47148 );
not ( n53682 , n51723 );
not ( n53683 , n48679 );
or ( n53684 , n53682 , n53683 );
nand ( n53685 , n49823 , n53228 );
nand ( n53686 , n53684 , n53685 );
not ( n53687 , n53686 );
or ( n53688 , n53681 , n53687 );
nand ( n53689 , n53230 , n52421 );
nand ( n53690 , n53688 , n53689 );
not ( n53691 , n51865 );
not ( n53692 , n51351 );
not ( n53693 , n52916 );
or ( n53694 , n53692 , n53693 );
nand ( n53695 , n49707 , n49809 );
nand ( n53696 , n53694 , n53695 );
not ( n53697 , n53696 );
or ( n53698 , n53691 , n53697 );
nand ( n53699 , n53143 , n49713 );
nand ( n53700 , n53698 , n53699 );
xor ( n53701 , n53690 , n53700 );
not ( n53702 , n52043 );
not ( n53703 , n50232 );
not ( n53704 , n49837 );
or ( n53705 , n53703 , n53704 );
not ( n53706 , n49837 );
nand ( n53707 , n53706 , n52048 );
nand ( n53708 , n53705 , n53707 );
not ( n53709 , n53708 );
or ( n53710 , n53702 , n53709 );
nand ( n53711 , n53301 , n50242 );
nand ( n53712 , n53710 , n53711 );
xor ( n53713 , n53701 , n53712 );
not ( n53714 , n46564 );
not ( n53715 , n53275 );
or ( n53716 , n53714 , n53715 );
not ( n53717 , n48952 );
not ( n53718 , n40635 );
not ( n53719 , n53718 );
or ( n53720 , n53717 , n53719 );
not ( n53721 , n40635 );
not ( n53722 , n53721 );
nand ( n53723 , n53722 , n52990 );
nand ( n53724 , n53720 , n53723 );
nand ( n53725 , n53724 , n49832 );
nand ( n53726 , n53716 , n53725 );
xor ( n53727 , n53713 , n53726 );
not ( n53728 , n49026 );
not ( n53729 , n46425 );
not ( n53730 , n40590 );
not ( n53731 , n53730 );
or ( n53732 , n53729 , n53731 );
nand ( n53733 , n52212 , n46422 );
nand ( n53734 , n53732 , n53733 );
not ( n53735 , n53734 );
or ( n53736 , n53728 , n53735 );
nand ( n53737 , n53349 , n46267 );
nand ( n53738 , n53736 , n53737 );
xor ( n53739 , n53727 , n53738 );
xor ( n53740 , n53680 , n53739 );
xor ( n53741 , n53740 , n53166 );
xor ( n53742 , n53680 , n53739 );
and ( n53743 , n53742 , n53166 );
and ( n53744 , n53680 , n53739 );
or ( n53745 , n53743 , n53744 );
xor ( n53746 , n53535 , n53212 );
xor ( n53747 , n53746 , n53625 );
xor ( n53748 , n53535 , n53212 );
and ( n53749 , n53748 , n53625 );
and ( n53750 , n53535 , n53212 );
or ( n53751 , n53749 , n53750 );
xor ( n53752 , n53244 , n53652 );
xor ( n53753 , n53752 , n53285 );
xor ( n53754 , n53244 , n53652 );
and ( n53755 , n53754 , n53285 );
and ( n53756 , n53244 , n53652 );
or ( n53757 , n53755 , n53756 );
xor ( n53758 , n53741 , n53359 );
xor ( n53759 , n53758 , n53747 );
xor ( n53760 , n53741 , n53359 );
and ( n53761 , n53760 , n53747 );
and ( n53762 , n53741 , n53359 );
or ( n53763 , n53761 , n53762 );
xor ( n53764 , n53365 , n53371 );
xor ( n53765 , n53764 , n53753 );
xor ( n53766 , n53365 , n53371 );
and ( n53767 , n53766 , n53753 );
and ( n53768 , n53365 , n53371 );
or ( n53769 , n53767 , n53768 );
xor ( n53770 , n53759 , n53377 );
xor ( n53771 , n53770 , n53765 );
xor ( n53772 , n53759 , n53377 );
and ( n53773 , n53772 , n53765 );
and ( n53774 , n53759 , n53377 );
or ( n53775 , n53773 , n53774 );
xor ( n53776 , n53690 , n53700 );
and ( n53777 , n53776 , n53712 );
and ( n53778 , n53690 , n53700 );
or ( n53779 , n53777 , n53778 );
xor ( n53780 , n53648 , n53094 );
and ( n53781 , n53780 , n53135 );
and ( n53782 , n53648 , n53094 );
or ( n53783 , n53781 , n53782 );
xor ( n53784 , n53450 , n53521 );
and ( n53785 , n53784 , n53532 );
and ( n53786 , n53450 , n53521 );
or ( n53787 , n53785 , n53786 );
xor ( n53788 , n53554 , n53504 );
and ( n53789 , n53788 , n53565 );
and ( n53790 , n53554 , n53504 );
or ( n53791 , n53789 , n53790 );
xor ( n53792 , n53578 , n53622 );
and ( n53793 , n53792 , n53387 );
and ( n53794 , n53578 , n53622 );
or ( n53795 , n53793 , n53794 );
xor ( n53796 , n53391 , n53641 );
and ( n53797 , n53796 , n53650 );
and ( n53798 , n53391 , n53641 );
or ( n53799 , n53797 , n53798 );
xor ( n53800 , n53713 , n53726 );
and ( n53801 , n53800 , n53738 );
and ( n53802 , n53713 , n53726 );
or ( n53803 , n53801 , n53802 );
xor ( n53804 , n53395 , n53667 );
and ( n53805 , n53804 , n53679 );
and ( n53806 , n53395 , n53667 );
or ( n53807 , n53805 , n53806 );
not ( n53808 , n50514 );
not ( n53809 , n47318 );
not ( n53810 , n53809 );
not ( n53811 , n49110 );
or ( n53812 , n53810 , n53811 );
nand ( n53813 , n47318 , n49452 );
nand ( n53814 , n53812 , n53813 );
not ( n53815 , n53814 );
or ( n53816 , n53808 , n53815 );
nand ( n53817 , n53496 , n51337 );
nand ( n53818 , n53816 , n53817 );
not ( n53819 , n48240 );
not ( n53820 , n47855 );
not ( n53821 , n49029 );
or ( n53822 , n53820 , n53821 );
not ( n53823 , n52414 );
nand ( n53824 , n53823 , n52016 );
nand ( n53825 , n53822 , n53824 );
not ( n53826 , n53825 );
or ( n53827 , n53819 , n53826 );
nand ( n53828 , n53482 , n47873 );
nand ( n53829 , n53827 , n53828 );
xor ( n53830 , n53818 , n53829 );
not ( n53831 , n49014 );
not ( n53832 , n53432 );
or ( n53833 , n53831 , n53832 );
and ( n53834 , n48758 , n48523 );
not ( n53835 , n48758 );
and ( n53836 , n53835 , n41683 );
or ( n53837 , n53834 , n53836 );
nand ( n53838 , n53837 , n49320 );
nand ( n53839 , n53833 , n53838 );
xor ( n53840 , n53830 , n53839 );
xor ( n53841 , n53818 , n53829 );
and ( n53842 , n53841 , n53839 );
and ( n53843 , n53818 , n53829 );
or ( n53844 , n53842 , n53843 );
not ( n53845 , n50176 );
not ( n53846 , n53445 );
or ( n53847 , n53845 , n53846 );
and ( n53848 , n51193 , n53439 );
not ( n53849 , n51193 );
and ( n53850 , n53849 , n48970 );
or ( n53851 , n53848 , n53850 );
nand ( n53852 , n53851 , n48277 );
nand ( n53853 , n53847 , n53852 );
not ( n53854 , n53463 );
not ( n53855 , n49779 );
or ( n53856 , n53854 , n53855 );
not ( n53857 , n51671 );
not ( n53858 , n49619 );
not ( n53859 , n53858 );
or ( n53860 , n53857 , n53859 );
nand ( n53861 , n49770 , n51670 );
nand ( n53862 , n53860 , n53861 );
nand ( n53863 , n53862 , n51809 );
nand ( n53864 , n53856 , n53863 );
xor ( n53865 , n53853 , n53864 );
not ( n53866 , n53473 );
not ( n53867 , n52749 );
or ( n53868 , n53866 , n53867 );
and ( n53869 , n50163 , n51792 );
not ( n53870 , n50163 );
and ( n53871 , n53870 , n48829 );
or ( n53872 , n53869 , n53871 );
nand ( n53873 , n53872 , n52757 );
nand ( n53874 , n53868 , n53873 );
xor ( n53875 , n53865 , n53874 );
xor ( n53876 , n53853 , n53864 );
and ( n53877 , n53876 , n53874 );
and ( n53878 , n53853 , n53864 );
or ( n53879 , n53877 , n53878 );
not ( n53880 , n50659 );
not ( n53881 , n53663 );
not ( n53882 , n53881 );
or ( n53883 , n53880 , n53882 );
not ( n53884 , n40363 );
and ( n53885 , n46072 , n53884 );
not ( n53886 , n46072 );
and ( n53887 , n53886 , n40364 );
or ( n53888 , n53885 , n53887 );
nand ( n53889 , n53888 , n47009 );
nand ( n53890 , n53883 , n53889 );
xor ( n53891 , n53454 , n53875 );
xor ( n53892 , n53891 , n53840 );
xor ( n53893 , n53890 , n53892 );
xor ( n53894 , n53893 , n53791 );
xor ( n53895 , n53890 , n53892 );
and ( n53896 , n53895 , n53791 );
and ( n53897 , n53890 , n53892 );
or ( n53898 , n53896 , n53897 );
xor ( n53899 , n53787 , n53795 );
not ( n53900 , n53530 );
not ( n53901 , n51215 );
or ( n53902 , n53900 , n53901 );
not ( n53903 , n51204 );
not ( n53904 , n50898 );
not ( n53905 , n53904 );
or ( n53906 , n53903 , n53905 );
nand ( n53907 , n51831 , n48860 );
nand ( n53908 , n53906 , n53907 );
nand ( n53909 , n53908 , n50922 );
nand ( n53910 , n53902 , n53909 );
not ( n53911 , n53563 );
not ( n53912 , n52482 );
or ( n53913 , n53911 , n53912 );
not ( n53914 , n47227 );
not ( n53915 , n52130 );
or ( n53916 , n53914 , n53915 );
buf ( n53917 , n52106 );
buf ( n53918 , n53917 );
nand ( n53919 , n53918 , n47589 );
nand ( n53920 , n53916 , n53919 );
nand ( n53921 , n51766 , n53920 );
nand ( n53922 , n53913 , n53921 );
xor ( n53923 , n53910 , n53922 );
not ( n53924 , n52139 );
not ( n53925 , n53552 );
or ( n53926 , n53924 , n53925 );
not ( n53927 , n51533 );
not ( n53928 , n53550 );
and ( n53929 , n48898 , n53928 );
not ( n53930 , n48898 );
buf ( n53931 , n51818 );
and ( n53932 , n53930 , n53931 );
nor ( n53933 , n53929 , n53932 );
or ( n53934 , n53927 , n53933 );
nand ( n53935 , n53926 , n53934 );
xor ( n53936 , n53923 , n53935 );
xor ( n53937 , n53899 , n53936 );
xor ( n53938 , n53787 , n53795 );
and ( n53939 , n53938 , n53936 );
and ( n53940 , n53787 , n53795 );
or ( n53941 , n53939 , n53940 );
not ( n53942 , n53576 );
not ( n53943 , n53182 );
or ( n53944 , n53942 , n53943 );
not ( n53945 , n47646 );
not ( n53946 , n52836 );
buf ( n53947 , n53946 );
not ( n53948 , n53947 );
or ( n53949 , n53945 , n53948 );
nand ( n53950 , n52841 , n47650 );
nand ( n53951 , n53949 , n53950 );
nand ( n53952 , n53571 , n53951 );
nand ( n53953 , n53944 , n53952 );
not ( n53954 , n53617 );
not ( n53955 , n53608 );
buf ( n53956 , n53955 );
not ( n53957 , n53956 );
or ( n53958 , n53954 , n53957 );
not ( n53959 , n46037 );
not ( n53960 , n53595 );
or ( n53961 , n53959 , n53960 );
nand ( n53962 , n53615 , n47306 );
nand ( n53963 , n53961 , n53962 );
nand ( n53964 , n53963 , n53620 );
nand ( n53965 , n53958 , n53964 );
xor ( n53966 , n53953 , n53965 );
xor ( n53967 , n53966 , n53508 );
xor ( n53968 , n53967 , n53807 );
not ( n53969 , n52004 );
not ( n53970 , n52377 );
not ( n53971 , n50084 );
or ( n53972 , n53970 , n53971 );
not ( n53973 , n52377 );
nand ( n53974 , n41407 , n53973 );
nand ( n53975 , n53972 , n53974 );
not ( n53976 , n53975 );
or ( n53977 , n53969 , n53976 );
nand ( n53978 , n53423 , n49116 );
nand ( n53979 , n53977 , n53978 );
and ( n53980 , n53486 , n53498 );
xor ( n53981 , n53979 , n53980 );
not ( n53982 , n47148 );
not ( n53983 , n51723 );
not ( n53984 , n52589 );
or ( n53985 , n53983 , n53984 );
nand ( n53986 , n49001 , n53228 );
nand ( n53987 , n53985 , n53986 );
not ( n53988 , n53987 );
or ( n53989 , n53982 , n53988 );
nand ( n53990 , n53686 , n52421 );
nand ( n53991 , n53989 , n53990 );
xor ( n53992 , n53981 , n53991 );
not ( n53993 , n47384 );
not ( n53994 , n49500 );
not ( n53995 , n51841 );
or ( n53996 , n53994 , n53995 );
not ( n53997 , n49500 );
nand ( n53998 , n40692 , n53997 );
nand ( n53999 , n53996 , n53998 );
not ( n54000 , n53999 );
or ( n54001 , n53993 , n54000 );
nand ( n54002 , n53517 , n49252 );
nand ( n54003 , n54001 , n54002 );
xor ( n54004 , n53992 , n54003 );
xor ( n54005 , n54004 , n53779 );
xor ( n54006 , n53968 , n54005 );
xor ( n54007 , n53967 , n53807 );
and ( n54008 , n54007 , n54005 );
and ( n54009 , n53967 , n53807 );
or ( n54010 , n54008 , n54009 );
xor ( n54011 , n53803 , n53799 );
xor ( n54012 , n54011 , n53539 );
xor ( n54013 , n53803 , n53799 );
and ( n54014 , n54013 , n53539 );
and ( n54015 , n53803 , n53799 );
or ( n54016 , n54014 , n54015 );
not ( n54017 , n46564 );
not ( n54018 , n53724 );
or ( n54019 , n54017 , n54018 );
not ( n54020 , n40376 );
and ( n54021 , n54020 , n48952 );
not ( n54022 , n54020 );
and ( n54023 , n54022 , n47514 );
or ( n54024 , n54021 , n54023 );
nand ( n54025 , n54024 , n49832 );
nand ( n54026 , n54019 , n54025 );
not ( n54027 , n53675 );
not ( n54028 , n50634 );
not ( n54029 , n54028 );
not ( n54030 , n40735 );
or ( n54031 , n54029 , n54030 );
not ( n54032 , n51924 );
nand ( n54033 , n54032 , n50634 );
nand ( n54034 , n54031 , n54033 );
not ( n54035 , n54034 );
or ( n54036 , n54027 , n54035 );
nand ( n54037 , n53673 , n47407 );
nand ( n54038 , n54036 , n54037 );
xor ( n54039 , n54026 , n54038 );
not ( n54040 , n46267 );
not ( n54041 , n53734 );
or ( n54042 , n54040 , n54041 );
not ( n54043 , n46425 );
not ( n54044 , n52432 );
or ( n54045 , n54043 , n54044 );
not ( n54046 , n40626 );
or ( n54047 , n54046 , n46425 );
nand ( n54048 , n54045 , n54047 );
nand ( n54049 , n54048 , n49026 );
nand ( n54050 , n54042 , n54049 );
xor ( n54051 , n54039 , n54050 );
not ( n54052 , n46776 );
not ( n54053 , n53637 );
or ( n54054 , n54052 , n54053 );
and ( n54055 , n50087 , n52570 );
not ( n54056 , n50087 );
and ( n54057 , n54056 , n51916 );
nor ( n54058 , n54055 , n54057 );
nand ( n54059 , n54058 , n47827 );
nand ( n54060 , n54054 , n54059 );
xor ( n54061 , n53783 , n54060 );
not ( n54062 , n49713 );
not ( n54063 , n53696 );
or ( n54064 , n54062 , n54063 );
and ( n54065 , n51351 , n51110 );
not ( n54066 , n51351 );
and ( n54067 , n54066 , n41036 );
nor ( n54068 , n54065 , n54067 );
nand ( n54069 , n54068 , n51865 );
nand ( n54070 , n54064 , n54069 );
and ( n54071 , n36607 , n37565 );
not ( n54072 , n36607 );
and ( n54073 , n54072 , n37564 );
nor ( n54074 , n54071 , n54073 );
xor ( n54075 , n53588 , n54074 );
not ( n54076 , n54075 );
not ( n54077 , n54076 );
and ( n54078 , n54077 , n48689 );
xor ( n54079 , n54070 , n54078 );
not ( n54080 , n50242 );
not ( n54081 , n53708 );
or ( n54082 , n54080 , n54081 );
not ( n54083 , n48645 );
not ( n54084 , n50004 );
or ( n54085 , n54083 , n54084 );
nand ( n54086 , n49549 , n52048 );
nand ( n54087 , n54085 , n54086 );
nand ( n54088 , n54087 , n52043 );
nand ( n54089 , n54082 , n54088 );
xor ( n54090 , n54079 , n54089 );
xor ( n54091 , n54061 , n54090 );
xor ( n54092 , n54051 , n54091 );
xor ( n54093 , n54092 , n53937 );
xor ( n54094 , n54051 , n54091 );
and ( n54095 , n54094 , n53937 );
and ( n54096 , n54051 , n54091 );
or ( n54097 , n54095 , n54096 );
xor ( n54098 , n53629 , n53894 );
xor ( n54099 , n54098 , n54012 );
xor ( n54100 , n53629 , n53894 );
and ( n54101 , n54100 , n54012 );
and ( n54102 , n53629 , n53894 );
or ( n54103 , n54101 , n54102 );
xor ( n54104 , n53656 , n54006 );
xor ( n54105 , n54104 , n53745 );
xor ( n54106 , n53656 , n54006 );
and ( n54107 , n54106 , n53745 );
and ( n54108 , n53656 , n54006 );
or ( n54109 , n54107 , n54108 );
xor ( n54110 , n54093 , n53751 );
xor ( n54111 , n54110 , n53757 );
xor ( n54112 , n54093 , n53751 );
and ( n54113 , n54112 , n53757 );
and ( n54114 , n54093 , n53751 );
or ( n54115 , n54113 , n54114 );
xor ( n54116 , n54099 , n54105 );
xor ( n54117 , n54116 , n53763 );
xor ( n54118 , n54099 , n54105 );
and ( n54119 , n54118 , n53763 );
and ( n54120 , n54099 , n54105 );
or ( n54121 , n54119 , n54120 );
xor ( n54122 , n54111 , n53769 );
xor ( n54123 , n54122 , n54117 );
xor ( n54124 , n54111 , n53769 );
and ( n54125 , n54124 , n54117 );
and ( n54126 , n54111 , n53769 );
or ( n54127 , n54125 , n54126 );
xor ( n54128 , n53979 , n53980 );
and ( n54129 , n54128 , n53991 );
and ( n54130 , n53979 , n53980 );
or ( n54131 , n54129 , n54130 );
xor ( n54132 , n54070 , n54078 );
and ( n54133 , n54132 , n54089 );
and ( n54134 , n54070 , n54078 );
or ( n54135 , n54133 , n54134 );
xor ( n54136 , n53454 , n53875 );
and ( n54137 , n54136 , n53840 );
and ( n54138 , n53454 , n53875 );
or ( n54139 , n54137 , n54138 );
xor ( n54140 , n53910 , n53922 );
and ( n54141 , n54140 , n53935 );
and ( n54142 , n53910 , n53922 );
or ( n54143 , n54141 , n54142 );
xor ( n54144 , n53953 , n53965 );
and ( n54145 , n54144 , n53508 );
and ( n54146 , n53953 , n53965 );
or ( n54147 , n54145 , n54146 );
xor ( n54148 , n53992 , n54003 );
and ( n54149 , n54148 , n53779 );
and ( n54150 , n53992 , n54003 );
or ( n54151 , n54149 , n54150 );
xor ( n54152 , n53783 , n54060 );
and ( n54153 , n54152 , n54090 );
and ( n54154 , n53783 , n54060 );
or ( n54155 , n54153 , n54154 );
xor ( n54156 , n54026 , n54038 );
and ( n54157 , n54156 , n54050 );
and ( n54158 , n54026 , n54038 );
or ( n54159 , n54157 , n54158 );
not ( n54160 , n49737 );
not ( n54161 , n49017 );
not ( n54162 , n47524 );
or ( n54163 , n54161 , n54162 );
nand ( n54164 , n47527 , n48704 );
nand ( n54165 , n54163 , n54164 );
not ( n54166 , n54165 );
or ( n54167 , n54160 , n54166 );
nand ( n54168 , n50554 , n53837 );
nand ( n54169 , n54167 , n54168 );
not ( n54170 , n49288 );
not ( n54171 , n49284 );
not ( n54172 , n49245 );
or ( n54173 , n54171 , n54172 );
nand ( n54174 , n47918 , n53492 );
nand ( n54175 , n54173 , n54174 );
not ( n54176 , n54175 );
or ( n54177 , n54170 , n54176 );
nand ( n54178 , n49276 , n53814 );
nand ( n54179 , n54177 , n54178 );
xor ( n54180 , n54169 , n54179 );
not ( n54181 , n53862 );
not ( n54182 , n52736 );
or ( n54183 , n54181 , n54182 );
buf ( n54184 , n46880 );
not ( n54185 , n54184 );
not ( n54186 , n54185 );
not ( n54187 , n49766 );
or ( n54188 , n54186 , n54187 );
nand ( n54189 , n49619 , n54184 );
nand ( n54190 , n54188 , n54189 );
nand ( n54191 , n54190 , n50078 );
nand ( n54192 , n54183 , n54191 );
xor ( n54193 , n54180 , n54192 );
xor ( n54194 , n54169 , n54179 );
and ( n54195 , n54194 , n54192 );
and ( n54196 , n54169 , n54179 );
or ( n54197 , n54195 , n54196 );
not ( n54198 , n52749 );
not ( n54199 , n53872 );
or ( n54200 , n54198 , n54199 );
and ( n54201 , n50301 , n52033 );
and ( n54202 , n50324 , n52038 );
nor ( n54203 , n54201 , n54202 );
or ( n54204 , n54203 , n50330 );
nand ( n54205 , n54200 , n54204 );
not ( n54206 , n48240 );
not ( n54207 , n51680 );
not ( n54208 , n48303 );
or ( n54209 , n54207 , n54208 );
not ( n54210 , n48779 );
not ( n54211 , n54210 );
nand ( n54212 , n54211 , n52016 );
nand ( n54213 , n54209 , n54212 );
not ( n54214 , n54213 );
or ( n54215 , n54206 , n54214 );
nand ( n54216 , n53825 , n47873 );
nand ( n54217 , n54215 , n54216 );
not ( n54218 , n50176 );
not ( n54219 , n53851 );
or ( n54220 , n54218 , n54219 );
not ( n54221 , n48456 );
not ( n54222 , n48736 );
or ( n54223 , n54221 , n54222 );
nand ( n54224 , n49298 , n48967 );
nand ( n54225 , n54223 , n54224 );
nand ( n54226 , n54225 , n52723 );
nand ( n54227 , n54220 , n54226 );
xor ( n54228 , n54217 , n54227 );
xor ( n54229 , n54205 , n54228 );
not ( n54230 , n52962 );
not ( n54231 , n50232 );
not ( n54232 , n49809 );
or ( n54233 , n54231 , n54232 );
nand ( n54234 , n50254 , n52048 );
nand ( n54235 , n54233 , n54234 );
not ( n54236 , n54235 );
or ( n54237 , n54230 , n54236 );
nand ( n54238 , n54087 , n52970 );
nand ( n54239 , n54237 , n54238 );
xor ( n54240 , n54229 , n54239 );
xor ( n54241 , n54205 , n54228 );
and ( n54242 , n54241 , n54239 );
and ( n54243 , n54205 , n54228 );
or ( n54244 , n54242 , n54243 );
not ( n54245 , n51865 );
not ( n54246 , n52267 );
not ( n54247 , n53513 );
or ( n54248 , n54246 , n54247 );
not ( n54249 , n52767 );
nand ( n54250 , n54249 , n52273 );
nand ( n54251 , n54248 , n54250 );
not ( n54252 , n54251 );
or ( n54253 , n54245 , n54252 );
nand ( n54254 , n54068 , n49713 );
nand ( n54255 , n54253 , n54254 );
xor ( n54256 , n53844 , n54255 );
xor ( n54257 , n54256 , n54193 );
xor ( n54258 , n54257 , n54143 );
xor ( n54259 , n54258 , n54147 );
xor ( n54260 , n54257 , n54143 );
and ( n54261 , n54260 , n54147 );
and ( n54262 , n54257 , n54143 );
or ( n54263 , n54261 , n54262 );
not ( n54264 , n53920 );
not ( n54265 , n52123 );
buf ( n54266 , n54265 );
not ( n54267 , n54266 );
or ( n54268 , n54264 , n54267 );
not ( n54269 , n49654 );
not ( n54270 , n52130 );
or ( n54271 , n54269 , n54270 );
nand ( n54272 , n52870 , n47368 );
nand ( n54273 , n54271 , n54272 );
nand ( n54274 , n54273 , n51766 );
nand ( n54275 , n54268 , n54274 );
not ( n54276 , n53951 );
not ( n54277 , n52854 );
or ( n54278 , n54276 , n54277 );
not ( n54279 , n47047 );
not ( n54280 , n53186 );
or ( n54281 , n54279 , n54280 );
not ( n54282 , n49734 );
not ( n54283 , n53947 );
nand ( n54284 , n54282 , n54283 );
nand ( n54285 , n54281 , n54284 );
nand ( n54286 , n52469 , n54285 );
nand ( n54287 , n54278 , n54286 );
xor ( n54288 , n54275 , n54287 );
buf ( n54289 , n33421 );
nand ( n54290 , n54289 , n33549 );
not ( n54291 , n54290 );
and ( n54292 , n36675 , n54291 );
not ( n54293 , n36675 );
and ( n54294 , n54293 , n54290 );
nor ( n54295 , n54292 , n54294 );
buf ( n54296 , n54295 );
buf ( n54297 , n54296 );
buf ( n54298 , n54297 );
and ( n54299 , n48689 , n54298 );
not ( n54300 , n48689 );
not ( n54301 , n54296 );
buf ( n54302 , n54301 );
and ( n54303 , n54300 , n54302 );
nor ( n54304 , n54299 , n54303 );
not ( n54305 , n54304 );
not ( n54306 , n54074 );
not ( n54307 , n54306 );
not ( n54308 , n54296 );
not ( n54309 , n54308 );
or ( n54310 , n54307 , n54309 );
nand ( n54311 , n54296 , n54074 );
nand ( n54312 , n54310 , n54311 );
nor ( n54313 , n54312 , n54075 );
not ( n54314 , n54313 );
not ( n54315 , n54314 );
buf ( n54316 , n54315 );
not ( n54317 , n54316 );
or ( n54318 , n54305 , n54317 );
not ( n54319 , n50914 );
not ( n54320 , n54302 );
or ( n54321 , n54319 , n54320 );
not ( n54322 , n54297 );
not ( n54323 , n54322 );
nand ( n54324 , n54323 , n48766 );
nand ( n54325 , n54321 , n54324 );
not ( n54326 , n54077 );
not ( n54327 , n54326 );
nand ( n54328 , n54325 , n54327 );
nand ( n54329 , n54318 , n54328 );
xor ( n54330 , n54288 , n54329 );
not ( n54331 , n53908 );
not ( n54332 , n50911 );
or ( n54333 , n54331 , n54332 );
not ( n54334 , n49624 );
not ( n54335 , n50916 );
or ( n54336 , n54334 , n54335 );
nand ( n54337 , n50898 , n49630 );
nand ( n54338 , n54336 , n54337 );
nand ( n54339 , n54338 , n50921 );
nand ( n54340 , n54333 , n54339 );
xor ( n54341 , n53879 , n54340 );
or ( n54342 , n53924 , n53933 );
not ( n54343 , n51505 );
not ( n54344 , n48589 );
and ( n54345 , n54343 , n54344 );
and ( n54346 , n53550 , n48589 );
nor ( n54347 , n54345 , n54346 );
or ( n54348 , n51146 , n54347 );
nand ( n54349 , n54342 , n54348 );
xor ( n54350 , n54341 , n54349 );
xor ( n54351 , n54330 , n54350 );
xor ( n54352 , n54351 , n54151 );
xor ( n54353 , n54330 , n54350 );
and ( n54354 , n54353 , n54151 );
and ( n54355 , n54330 , n54350 );
or ( n54356 , n54354 , n54355 );
not ( n54357 , n53963 );
not ( n54358 , n53956 );
or ( n54359 , n54357 , n54358 );
and ( n54360 , n46273 , n53591 );
not ( n54361 , n46273 );
and ( n54362 , n54361 , n53615 );
or ( n54363 , n54360 , n54362 );
not ( n54364 , n53618 );
nand ( n54365 , n54363 , n54364 );
nand ( n54366 , n54359 , n54365 );
xor ( n54367 , n54366 , n54240 );
xor ( n54368 , n54367 , n54131 );
xor ( n54369 , n54159 , n54368 );
xor ( n54370 , n54369 , n54155 );
xor ( n54371 , n54159 , n54368 );
and ( n54372 , n54371 , n54155 );
and ( n54373 , n54159 , n54368 );
or ( n54374 , n54372 , n54373 );
not ( n54375 , n47827 );
not ( n54376 , n46650 );
not ( n54377 , n40591 );
not ( n54378 , n54377 );
or ( n54379 , n54376 , n54378 );
not ( n54380 , n53730 );
nand ( n54381 , n54380 , n50087 );
nand ( n54382 , n54379 , n54381 );
not ( n54383 , n54382 );
or ( n54384 , n54375 , n54383 );
nand ( n54385 , n54058 , n48295 );
nand ( n54386 , n54384 , n54385 );
xor ( n54387 , n54135 , n54386 );
not ( n54388 , n47407 );
not ( n54389 , n54034 );
or ( n54390 , n54388 , n54389 );
not ( n54391 , n47803 );
not ( n54392 , n52894 );
or ( n54393 , n54391 , n54392 );
nand ( n54394 , n51601 , n48727 );
nand ( n54395 , n54393 , n54394 );
nand ( n54396 , n54395 , n53675 );
nand ( n54397 , n54390 , n54396 );
xor ( n54398 , n54387 , n54397 );
not ( n54399 , n47009 );
not ( n54400 , n46072 );
not ( n54401 , n40147 );
buf ( n54402 , n54401 );
not ( n54403 , n54402 );
or ( n54404 , n54400 , n54403 );
not ( n54405 , n40147 );
not ( n54406 , n54405 );
nand ( n54407 , n54406 , n50405 );
nand ( n54408 , n54404 , n54407 );
not ( n54409 , n54408 );
or ( n54410 , n54399 , n54409 );
nand ( n54411 , n53888 , n50659 );
nand ( n54412 , n54410 , n54411 );
not ( n54413 , n46188 );
not ( n54414 , n46425 );
not ( n54415 , n40635 );
not ( n54416 , n54415 );
or ( n54417 , n54414 , n54416 );
not ( n54418 , n53718 );
nand ( n54419 , n54418 , n46422 );
nand ( n54420 , n54417 , n54419 );
not ( n54421 , n54420 );
or ( n54422 , n54413 , n54421 );
nand ( n54423 , n54048 , n46267 );
nand ( n54424 , n54422 , n54423 );
xor ( n54425 , n54412 , n54424 );
xor ( n54426 , n54425 , n54139 );
xor ( n54427 , n54398 , n54426 );
not ( n54428 , n49832 );
not ( n54429 , n47508 );
not ( n54430 , n53661 );
or ( n54431 , n54429 , n54430 );
not ( n54432 , n40224 );
buf ( n54433 , n54432 );
nand ( n54434 , n54433 , n51577 );
nand ( n54435 , n54431 , n54434 );
not ( n54436 , n54435 );
or ( n54437 , n54428 , n54436 );
nand ( n54438 , n54024 , n46564 );
nand ( n54439 , n54437 , n54438 );
not ( n54440 , n52421 );
not ( n54441 , n53987 );
or ( n54442 , n54440 , n54441 );
not ( n54443 , n51723 );
not ( n54444 , n41216 );
or ( n54445 , n54443 , n54444 );
nand ( n54446 , n53706 , n53228 );
nand ( n54447 , n54445 , n54446 );
nand ( n54448 , n54447 , n47148 );
nand ( n54449 , n54442 , n54448 );
not ( n54450 , n52004 );
not ( n54451 , n52377 );
not ( n54452 , n48679 );
or ( n54453 , n54451 , n54452 );
nand ( n54454 , n52272 , n53973 );
nand ( n54455 , n54453 , n54454 );
not ( n54456 , n54455 );
or ( n54457 , n54450 , n54456 );
nand ( n54458 , n53975 , n49116 );
nand ( n54459 , n54457 , n54458 );
xor ( n54460 , n54449 , n54459 );
not ( n54461 , n53615 );
not ( n54462 , n54306 );
nand ( n54463 , n54462 , n48689 );
nand ( n54464 , n54461 , n54463 );
nand ( n54465 , n54306 , n46441 );
and ( n54466 , n54464 , n54465 );
not ( n54467 , n54297 );
buf ( n54468 , n54467 );
nor ( n54469 , n54466 , n54468 );
xor ( n54470 , n54460 , n54469 );
xor ( n54471 , n54439 , n54470 );
not ( n54472 , n53999 );
not ( n54473 , n48989 );
or ( n54474 , n54472 , n54473 );
not ( n54475 , n49500 );
not ( n54476 , n50958 );
or ( n54477 , n54475 , n54476 );
nand ( n54478 , n52284 , n47979 );
nand ( n54479 , n54477 , n54478 );
not ( n54480 , n54479 );
or ( n54481 , n54480 , n53509 );
nand ( n54482 , n54474 , n54481 );
xor ( n54483 , n54471 , n54482 );
xor ( n54484 , n54427 , n54483 );
xor ( n54485 , n54398 , n54426 );
and ( n54486 , n54485 , n54483 );
and ( n54487 , n54398 , n54426 );
or ( n54488 , n54486 , n54487 );
xor ( n54489 , n53898 , n53941 );
xor ( n54490 , n54489 , n54259 );
xor ( n54491 , n53898 , n53941 );
and ( n54492 , n54491 , n54259 );
and ( n54493 , n53898 , n53941 );
or ( n54494 , n54492 , n54493 );
xor ( n54495 , n54010 , n54352 );
xor ( n54496 , n54495 , n54370 );
xor ( n54497 , n54010 , n54352 );
and ( n54498 , n54497 , n54370 );
and ( n54499 , n54010 , n54352 );
or ( n54500 , n54498 , n54499 );
xor ( n54501 , n54016 , n54097 );
xor ( n54502 , n54501 , n54484 );
xor ( n54503 , n54016 , n54097 );
and ( n54504 , n54503 , n54484 );
and ( n54505 , n54016 , n54097 );
or ( n54506 , n54504 , n54505 );
xor ( n54507 , n54490 , n54109 );
xor ( n54508 , n54507 , n54103 );
xor ( n54509 , n54490 , n54109 );
and ( n54510 , n54509 , n54103 );
and ( n54511 , n54490 , n54109 );
or ( n54512 , n54510 , n54511 );
xor ( n54513 , n54496 , n54502 );
xor ( n54514 , n54513 , n54115 );
xor ( n54515 , n54496 , n54502 );
and ( n54516 , n54515 , n54115 );
and ( n54517 , n54496 , n54502 );
or ( n54518 , n54516 , n54517 );
xor ( n54519 , n54508 , n54121 );
xor ( n54520 , n54519 , n54514 );
xor ( n54521 , n54508 , n54121 );
and ( n54522 , n54521 , n54514 );
and ( n54523 , n54508 , n54121 );
or ( n54524 , n54522 , n54523 );
xor ( n54525 , n54449 , n54459 );
and ( n54526 , n54525 , n54469 );
and ( n54527 , n54449 , n54459 );
or ( n54528 , n54526 , n54527 );
xor ( n54529 , n53844 , n54255 );
and ( n54530 , n54529 , n54193 );
and ( n54531 , n53844 , n54255 );
or ( n54532 , n54530 , n54531 );
xor ( n54533 , n53879 , n54340 );
and ( n54534 , n54533 , n54349 );
and ( n54535 , n53879 , n54340 );
or ( n54536 , n54534 , n54535 );
xor ( n54537 , n54275 , n54287 );
and ( n54538 , n54537 , n54329 );
and ( n54539 , n54275 , n54287 );
or ( n54540 , n54538 , n54539 );
xor ( n54541 , n54366 , n54240 );
and ( n54542 , n54541 , n54131 );
and ( n54543 , n54366 , n54240 );
or ( n54544 , n54542 , n54543 );
xor ( n54545 , n54135 , n54386 );
and ( n54546 , n54545 , n54397 );
and ( n54547 , n54135 , n54386 );
or ( n54548 , n54546 , n54547 );
xor ( n54549 , n54439 , n54470 );
and ( n54550 , n54549 , n54482 );
and ( n54551 , n54439 , n54470 );
or ( n54552 , n54550 , n54551 );
xor ( n54553 , n54412 , n54424 );
and ( n54554 , n54553 , n54139 );
and ( n54555 , n54412 , n54424 );
or ( n54556 , n54554 , n54555 );
not ( n54557 , n48277 );
not ( n54558 , n53439 );
not ( n54559 , n49029 );
or ( n54560 , n54558 , n54559 );
not ( n54561 , n48510 );
nand ( n54562 , n54561 , n48967 );
nand ( n54563 , n54560 , n54562 );
not ( n54564 , n54563 );
or ( n54565 , n54557 , n54564 );
not ( n54566 , n49420 );
nand ( n54567 , n54566 , n54225 );
nand ( n54568 , n54565 , n54567 );
not ( n54569 , n49014 );
not ( n54570 , n54165 );
or ( n54571 , n54569 , n54570 );
not ( n54572 , n48758 );
not ( n54573 , n51193 );
or ( n54574 , n54572 , n54573 );
nand ( n54575 , n41415 , n48704 );
nand ( n54576 , n54574 , n54575 );
nand ( n54577 , n54576 , n49022 );
nand ( n54578 , n54571 , n54577 );
xor ( n54579 , n54568 , n54578 );
not ( n54580 , n50195 );
not ( n54581 , n54175 );
or ( n54582 , n54580 , n54581 );
not ( n54583 , n50201 );
not ( n54584 , n53114 );
not ( n54585 , n54584 );
or ( n54586 , n54583 , n54585 );
not ( n54587 , n48523 );
nand ( n54588 , n54587 , n49283 );
nand ( n54589 , n54586 , n54588 );
nand ( n54590 , n54589 , n48891 );
nand ( n54591 , n54582 , n54590 );
xor ( n54592 , n54579 , n54591 );
xor ( n54593 , n54568 , n54578 );
and ( n54594 , n54593 , n54591 );
and ( n54595 , n54568 , n54578 );
or ( n54596 , n54594 , n54595 );
not ( n54597 , n54190 );
not ( n54598 , n52058 );
or ( n54599 , n54597 , n54598 );
not ( n54600 , n30964 );
not ( n54601 , n53858 );
or ( n54602 , n54600 , n54601 );
nand ( n54603 , n49619 , n47318 );
nand ( n54604 , n54602 , n54603 );
nand ( n54605 , n54604 , n50078 );
nand ( n54606 , n54599 , n54605 );
not ( n54607 , n54203 );
not ( n54608 , n54607 );
not ( n54609 , n50321 );
or ( n54610 , n54608 , n54609 );
not ( n54611 , n51670 );
not ( n54612 , n54611 );
buf ( n54613 , n50162 );
not ( n54614 , n54613 );
not ( n54615 , n54614 );
or ( n54616 , n54612 , n54615 );
nand ( n54617 , n50304 , n51670 );
nand ( n54618 , n54616 , n54617 );
nand ( n54619 , n54618 , n51452 );
nand ( n54620 , n54610 , n54619 );
xor ( n54621 , n54606 , n54620 );
not ( n54622 , n48240 );
not ( n54623 , n54622 );
not ( n54624 , n54623 );
buf ( n54625 , n47855 );
and ( n54626 , n48951 , n54625 );
not ( n54627 , n48951 );
buf ( n54628 , n52016 );
and ( n54629 , n54627 , n54628 );
or ( n54630 , n54626 , n54629 );
not ( n54631 , n54630 );
or ( n54632 , n54624 , n54631 );
nand ( n54633 , n54213 , n52022 );
nand ( n54634 , n54632 , n54633 );
xor ( n54635 , n54621 , n54634 );
xor ( n54636 , n54606 , n54620 );
and ( n54637 , n54636 , n54634 );
and ( n54638 , n54606 , n54620 );
or ( n54639 , n54637 , n54638 );
not ( n54640 , n46267 );
not ( n54641 , n54420 );
or ( n54642 , n54640 , n54641 );
not ( n54643 , n46425 );
not ( n54644 , n53289 );
or ( n54645 , n54643 , n54644 );
not ( n54646 , n54020 );
nand ( n54647 , n54646 , n46422 );
nand ( n54648 , n54645 , n54647 );
nand ( n54649 , n54648 , n49026 );
nand ( n54650 , n54642 , n54649 );
xor ( n54651 , n54650 , n54532 );
xor ( n54652 , n54651 , n54536 );
xor ( n54653 , n54650 , n54532 );
and ( n54654 , n54653 , n54536 );
and ( n54655 , n54650 , n54532 );
or ( n54656 , n54654 , n54655 );
not ( n54657 , n54347 );
not ( n54658 , n54657 );
not ( n54659 , n52139 );
or ( n54660 , n54658 , n54659 );
not ( n54661 , n51204 );
not ( n54662 , n51566 );
or ( n54663 , n54661 , n54662 );
nand ( n54664 , n51505 , n48860 );
nand ( n54665 , n54663 , n54664 );
nand ( n54666 , n51533 , n54665 );
nand ( n54667 , n54660 , n54666 );
not ( n54668 , n54273 );
not ( n54669 , n52482 );
or ( n54670 , n54668 , n54669 );
not ( n54671 , n48898 );
not ( n54672 , n52871 );
or ( n54673 , n54671 , n54672 );
nand ( n54674 , n53918 , n48897 );
nand ( n54675 , n54673 , n54674 );
nand ( n54676 , n51766 , n54675 );
nand ( n54677 , n54670 , n54676 );
xor ( n54678 , n54667 , n54677 );
xor ( n54679 , n54678 , n54635 );
xor ( n54680 , n54540 , n54679 );
not ( n54681 , n54363 );
not ( n54682 , n53609 );
or ( n54683 , n54681 , n54682 );
not ( n54684 , n47646 );
not ( n54685 , n53591 );
or ( n54686 , n54684 , n54685 );
nand ( n54687 , n53615 , n47650 );
nand ( n54688 , n54686 , n54687 );
nand ( n54689 , n54688 , n53620 );
nand ( n54690 , n54683 , n54689 );
xor ( n54691 , n54592 , n54690 );
not ( n54692 , n52151 );
not ( n54693 , n54338 );
or ( n54694 , n54692 , n54693 );
not ( n54695 , n51792 );
not ( n54696 , n50899 );
or ( n54697 , n54695 , n54696 );
or ( n54698 , n50916 , n51792 );
nand ( n54699 , n54697 , n54698 );
not ( n54700 , n54699 );
or ( n54701 , n54700 , n50626 );
nand ( n54702 , n54694 , n54701 );
xor ( n54703 , n54691 , n54702 );
xor ( n54704 , n54680 , n54703 );
xor ( n54705 , n54540 , n54679 );
and ( n54706 , n54705 , n54703 );
and ( n54707 , n54540 , n54679 );
or ( n54708 , n54706 , n54707 );
not ( n54709 , n54285 );
not ( n54710 , n53182 );
or ( n54711 , n54709 , n54710 );
and ( n54712 , n47227 , n53189 );
not ( n54713 , n47227 );
and ( n54714 , n54713 , n52841 );
or ( n54715 , n54712 , n54714 );
nand ( n54716 , n52469 , n54715 );
nand ( n54717 , n54711 , n54716 );
not ( n54718 , n54325 );
not ( n54719 , n54316 );
or ( n54720 , n54718 , n54719 );
buf ( n54721 , n47306 );
not ( n54722 , n54721 );
and ( n54723 , n54722 , n54302 );
not ( n54724 , n54722 );
not ( n54725 , n54302 );
and ( n54726 , n54724 , n54725 );
nor ( n54727 , n54723 , n54726 );
not ( n54728 , n54727 );
nand ( n54729 , n54728 , n54327 );
nand ( n54730 , n54720 , n54729 );
xor ( n54731 , n54717 , n54730 );
not ( n54732 , n51865 );
not ( n54733 , n52267 );
not ( n54734 , n51841 );
or ( n54735 , n54733 , n54734 );
nand ( n54736 , n40692 , n51351 );
nand ( n54737 , n54735 , n54736 );
not ( n54738 , n54737 );
or ( n54739 , n54732 , n54738 );
nand ( n54740 , n54251 , n49713 );
nand ( n54741 , n54739 , n54740 );
xor ( n54742 , n54731 , n54741 );
xor ( n54743 , n54544 , n54742 );
xor ( n54744 , n54743 , n54552 );
xor ( n54745 , n54544 , n54742 );
and ( n54746 , n54745 , n54552 );
and ( n54747 , n54544 , n54742 );
or ( n54748 , n54746 , n54747 );
xor ( n54749 , n54548 , n54556 );
xor ( n54750 , n54244 , n54528 );
not ( n54751 , n48073 );
not ( n54752 , n46650 );
not ( n54753 , n53271 );
or ( n54754 , n54752 , n54753 );
nand ( n54755 , n40626 , n50087 );
nand ( n54756 , n54754 , n54755 );
not ( n54757 , n54756 );
or ( n54758 , n54751 , n54757 );
nand ( n54759 , n54382 , n46776 );
nand ( n54760 , n54758 , n54759 );
xor ( n54761 , n54750 , n54760 );
xor ( n54762 , n54749 , n54761 );
xor ( n54763 , n54548 , n54556 );
and ( n54764 , n54763 , n54761 );
and ( n54765 , n54548 , n54556 );
or ( n54766 , n54764 , n54765 );
xor ( n54767 , n54652 , n54263 );
not ( n54768 , n47407 );
not ( n54769 , n54395 );
or ( n54770 , n54768 , n54769 );
not ( n54771 , n40526 );
and ( n54772 , n54771 , n47803 );
not ( n54773 , n54771 );
and ( n54774 , n54773 , n50634 );
or ( n54775 , n54772 , n54774 );
nand ( n54776 , n54775 , n48929 );
nand ( n54777 , n54770 , n54776 );
not ( n54778 , n49252 );
not ( n54779 , n54479 );
or ( n54780 , n54778 , n54779 );
not ( n54781 , n49500 );
not ( n54782 , n53259 );
or ( n54783 , n54781 , n54782 );
nand ( n54784 , n40734 , n47979 );
nand ( n54785 , n54783 , n54784 );
nand ( n54786 , n54785 , n47384 );
nand ( n54787 , n54780 , n54786 );
xor ( n54788 , n54777 , n54787 );
not ( n54789 , n47009 );
not ( n54790 , n40388 );
not ( n54791 , n54790 );
and ( n54792 , n54791 , n50405 );
not ( n54793 , n54791 );
and ( n54794 , n54793 , n46072 );
or ( n54795 , n54792 , n54794 );
not ( n54796 , n54795 );
or ( n54797 , n54789 , n54796 );
nand ( n54798 , n54408 , n50659 );
nand ( n54799 , n54797 , n54798 );
xor ( n54800 , n54788 , n54799 );
xor ( n54801 , n54767 , n54800 );
xor ( n54802 , n54652 , n54263 );
and ( n54803 , n54802 , n54800 );
and ( n54804 , n54652 , n54263 );
or ( n54805 , n54803 , n54804 );
not ( n54806 , n46564 );
not ( n54807 , n54435 );
or ( n54808 , n54806 , n54807 );
not ( n54809 , n47508 );
not ( n54810 , n40363 );
buf ( n54811 , n54810 );
not ( n54812 , n54811 );
or ( n54813 , n54809 , n54812 );
not ( n54814 , n53884 );
nand ( n54815 , n54814 , n47514 );
nand ( n54816 , n54813 , n54815 );
nand ( n54817 , n54816 , n49832 );
nand ( n54818 , n54808 , n54817 );
not ( n54819 , n52004 );
not ( n54820 , n52377 );
not ( n54821 , n52589 );
or ( n54822 , n54820 , n54821 );
nand ( n54823 , n41286 , n53973 );
nand ( n54824 , n54822 , n54823 );
not ( n54825 , n54824 );
or ( n54826 , n54819 , n54825 );
nand ( n54827 , n54455 , n49116 );
nand ( n54828 , n54826 , n54827 );
not ( n54829 , n36640 );
nor ( n54830 , n54829 , n36560 );
not ( n54831 , n54830 );
not ( n54832 , n36286 );
or ( n54833 , n54831 , n54832 );
nand ( n54834 , n54833 , n37400 );
nand ( n54835 , n36582 , n36584 );
and ( n54836 , n54834 , n54835 );
not ( n54837 , n54834 );
not ( n54838 , n54835 );
and ( n54839 , n54837 , n54838 );
nor ( n54840 , n54836 , n54839 );
not ( n54841 , n54840 );
not ( n54842 , n54841 );
and ( n54843 , n54296 , n54842 );
not ( n54844 , n54296 );
and ( n54845 , n54844 , n54841 );
nor ( n54846 , n54843 , n54845 );
not ( n54847 , n54846 );
buf ( n54848 , n54847 );
not ( n54849 , n54848 );
nor ( n54850 , n54849 , n46441 );
xor ( n54851 , n54828 , n54850 );
xor ( n54852 , n54851 , n54197 );
xor ( n54853 , n54818 , n54852 );
and ( n54854 , n54217 , n54227 );
not ( n54855 , n50242 );
not ( n54856 , n54235 );
or ( n54857 , n54855 , n54856 );
not ( n54858 , n48645 );
not ( n54859 , n50020 );
or ( n54860 , n54858 , n54859 );
nand ( n54861 , n51891 , n52048 );
nand ( n54862 , n54860 , n54861 );
nand ( n54863 , n54862 , n52043 );
nand ( n54864 , n54857 , n54863 );
xor ( n54865 , n54854 , n54864 );
not ( n54866 , n52421 );
not ( n54867 , n54447 );
or ( n54868 , n54866 , n54867 );
not ( n54869 , n48856 );
not ( n54870 , n49549 );
not ( n54871 , n54870 );
or ( n54872 , n54869 , n54871 );
nand ( n54873 , n51740 , n53228 );
nand ( n54874 , n54872 , n54873 );
buf ( n54875 , n50767 );
nand ( n54876 , n54874 , n54875 );
nand ( n54877 , n54868 , n54876 );
xor ( n54878 , n54865 , n54877 );
xor ( n54879 , n54853 , n54878 );
xor ( n54880 , n54879 , n54356 );
xor ( n54881 , n54880 , n54374 );
xor ( n54882 , n54879 , n54356 );
and ( n54883 , n54882 , n54374 );
and ( n54884 , n54879 , n54356 );
or ( n54885 , n54883 , n54884 );
xor ( n54886 , n54744 , n54704 );
xor ( n54887 , n54886 , n54762 );
xor ( n54888 , n54744 , n54704 );
and ( n54889 , n54888 , n54762 );
and ( n54890 , n54744 , n54704 );
or ( n54891 , n54889 , n54890 );
xor ( n54892 , n54488 , n54494 );
xor ( n54893 , n54892 , n54801 );
xor ( n54894 , n54488 , n54494 );
and ( n54895 , n54894 , n54801 );
and ( n54896 , n54488 , n54494 );
or ( n54897 , n54895 , n54896 );
xor ( n54898 , n54881 , n54500 );
xor ( n54899 , n54898 , n54887 );
xor ( n54900 , n54881 , n54500 );
and ( n54901 , n54900 , n54887 );
and ( n54902 , n54881 , n54500 );
or ( n54903 , n54901 , n54902 );
xor ( n54904 , n54506 , n54893 );
xor ( n54905 , n54904 , n54512 );
xor ( n54906 , n54506 , n54893 );
and ( n54907 , n54906 , n54512 );
and ( n54908 , n54506 , n54893 );
or ( n54909 , n54907 , n54908 );
xor ( n54910 , n54854 , n54864 );
and ( n54911 , n54910 , n54877 );
and ( n54912 , n54854 , n54864 );
or ( n54913 , n54911 , n54912 );
xor ( n54914 , n54899 , n54905 );
xor ( n54915 , n54914 , n54518 );
xor ( n54916 , n54899 , n54905 );
and ( n54917 , n54916 , n54518 );
and ( n54918 , n54899 , n54905 );
or ( n54919 , n54917 , n54918 );
xor ( n54920 , n54828 , n54850 );
and ( n54921 , n54920 , n54197 );
and ( n54922 , n54828 , n54850 );
or ( n54923 , n54921 , n54922 );
xor ( n54924 , n54592 , n54690 );
and ( n54925 , n54924 , n54702 );
and ( n54926 , n54592 , n54690 );
or ( n54927 , n54925 , n54926 );
xor ( n54928 , n54667 , n54677 );
and ( n54929 , n54928 , n54635 );
and ( n54930 , n54667 , n54677 );
or ( n54931 , n54929 , n54930 );
xor ( n54932 , n54717 , n54730 );
and ( n54933 , n54932 , n54741 );
and ( n54934 , n54717 , n54730 );
or ( n54935 , n54933 , n54934 );
xor ( n54936 , n54244 , n54528 );
and ( n54937 , n54936 , n54760 );
and ( n54938 , n54244 , n54528 );
or ( n54939 , n54937 , n54938 );
xor ( n54940 , n54818 , n54852 );
and ( n54941 , n54940 , n54878 );
and ( n54942 , n54818 , n54852 );
or ( n54943 , n54941 , n54942 );
xor ( n54944 , n54777 , n54787 );
and ( n54945 , n54944 , n54799 );
and ( n54946 , n54777 , n54787 );
or ( n54947 , n54945 , n54946 );
not ( n54948 , n52191 );
not ( n54949 , n49284 );
not ( n54950 , n47524 );
or ( n54951 , n54949 , n54950 );
nand ( n54952 , n48332 , n49283 );
nand ( n54953 , n54951 , n54952 );
not ( n54954 , n54953 );
or ( n54955 , n54948 , n54954 );
nand ( n54956 , n49979 , n54589 );
nand ( n54957 , n54955 , n54956 );
not ( n54958 , n54604 );
not ( n54959 , n51234 );
not ( n54960 , n54959 );
not ( n54961 , n54960 );
or ( n54962 , n54958 , n54961 );
not ( n54963 , n41692 );
not ( n54964 , n49766 );
and ( n54965 , n54963 , n54964 );
and ( n54966 , n47918 , n49766 );
nor ( n54967 , n54965 , n54966 );
not ( n54968 , n54967 );
nand ( n54969 , n54968 , n49789 );
nand ( n54970 , n54962 , n54969 );
xor ( n54971 , n54957 , n54970 );
not ( n54972 , n54618 );
not ( n54973 , n52749 );
or ( n54974 , n54972 , n54973 );
not ( n54975 , n48223 );
not ( n54976 , n50305 );
or ( n54977 , n54975 , n54976 );
nand ( n54978 , n54613 , n52712 );
nand ( n54979 , n54977 , n54978 );
nand ( n54980 , n54979 , n52757 );
nand ( n54981 , n54974 , n54980 );
xor ( n54982 , n54971 , n54981 );
xor ( n54983 , n54957 , n54970 );
and ( n54984 , n54983 , n54981 );
and ( n54985 , n54957 , n54970 );
or ( n54986 , n54984 , n54985 );
not ( n54987 , n48277 );
and ( n54988 , n41530 , n53439 );
not ( n54989 , n41530 );
and ( n54990 , n54989 , n48967 );
or ( n54991 , n54988 , n54990 );
not ( n54992 , n54991 );
or ( n54993 , n54987 , n54992 );
nand ( n54994 , n54563 , n49421 );
nand ( n54995 , n54993 , n54994 );
not ( n54996 , n48755 );
not ( n54997 , n54576 );
or ( n54998 , n54996 , n54997 );
not ( n54999 , n49313 );
not ( n55000 , n49297 );
or ( n55001 , n54999 , n55000 );
nand ( n55002 , n41575 , n48704 );
nand ( n55003 , n55001 , n55002 );
nand ( n55004 , n55003 , n49737 );
nand ( n55005 , n54998 , n55004 );
xor ( n55006 , n54995 , n55005 );
not ( n55007 , n48894 );
not ( n55008 , n54824 );
or ( n55009 , n55007 , n55008 );
not ( n55010 , n52377 );
not ( n55011 , n41216 );
or ( n55012 , n55010 , n55011 );
not ( n55013 , n52377 );
nand ( n55014 , n49209 , n55013 );
nand ( n55015 , n55012 , n55014 );
nand ( n55016 , n55015 , n52004 );
nand ( n55017 , n55009 , n55016 );
xor ( n55018 , n55006 , n55017 );
not ( n55019 , n54623 );
not ( n55020 , n54625 );
not ( n55021 , n49190 );
or ( n55022 , n55020 , n55021 );
not ( n55023 , n54625 );
nand ( n55024 , n51476 , n55023 );
nand ( n55025 , n55022 , n55024 );
not ( n55026 , n55025 );
or ( n55027 , n55019 , n55026 );
nand ( n55028 , n54630 , n52022 );
nand ( n55029 , n55027 , n55028 );
xor ( n55030 , n55018 , n55029 );
xor ( n55031 , n55006 , n55017 );
and ( n55032 , n55031 , n55029 );
and ( n55033 , n55006 , n55017 );
or ( n55034 , n55032 , n55033 );
not ( n55035 , n52043 );
not ( n55036 , n48645 );
not ( n55037 , n52076 );
or ( n55038 , n55036 , n55037 );
nand ( n55039 , n41132 , n49679 );
nand ( n55040 , n55038 , n55039 );
not ( n55041 , n55040 );
or ( n55042 , n55035 , n55041 );
nand ( n55043 , n54862 , n52970 );
nand ( n55044 , n55042 , n55043 );
xor ( n55045 , n54982 , n55044 );
not ( n55046 , n54699 );
not ( n55047 , n50911 );
or ( n55048 , n55046 , n55047 );
not ( n55049 , n52033 );
not ( n55050 , n50916 );
or ( n55051 , n55049 , n55050 );
nand ( n55052 , n51831 , n52038 );
nand ( n55053 , n55051 , n55052 );
nand ( n55054 , n55053 , n50922 );
nand ( n55055 , n55048 , n55054 );
xor ( n55056 , n55045 , n55055 );
xor ( n55057 , n55056 , n54927 );
xor ( n55058 , n55057 , n54931 );
xor ( n55059 , n55056 , n54927 );
and ( n55060 , n55059 , n54931 );
and ( n55061 , n55056 , n54927 );
or ( n55062 , n55060 , n55061 );
not ( n55063 , n54665 );
not ( n55064 , n53543 );
or ( n55065 , n55063 , n55064 );
not ( n55066 , n51146 );
not ( n55067 , n49624 );
not ( n55068 , n51566 );
or ( n55069 , n55067 , n55068 );
nand ( n55070 , n53549 , n49630 );
nand ( n55071 , n55069 , n55070 );
nand ( n55072 , n55066 , n55071 );
nand ( n55073 , n55065 , n55072 );
not ( n55074 , n54675 );
not ( n55075 , n52482 );
or ( n55076 , n55074 , n55075 );
not ( n55077 , n47765 );
not ( n55078 , n52871 );
or ( n55079 , n55077 , n55078 );
nand ( n55080 , n53918 , n48589 );
nand ( n55081 , n55079 , n55080 );
nand ( n55082 , n51766 , n55081 );
nand ( n55083 , n55076 , n55082 );
xor ( n55084 , n55073 , n55083 );
not ( n55085 , n54688 );
not ( n55086 , n53956 );
or ( n55087 , n55085 , n55086 );
not ( n55088 , n49734 );
buf ( n55089 , n53590 );
not ( n55090 , n55089 );
not ( n55091 , n55090 );
or ( n55092 , n55088 , n55091 );
nand ( n55093 , n55089 , n47821 );
nand ( n55094 , n55092 , n55093 );
nand ( n55095 , n55094 , n53620 );
nand ( n55096 , n55087 , n55095 );
xor ( n55097 , n55084 , n55096 );
not ( n55098 , n54715 );
not ( n55099 , n53182 );
or ( n55100 , n55098 , n55099 );
not ( n55101 , n52165 );
not ( n55102 , n52835 );
not ( n55103 , n55102 );
not ( n55104 , n55103 );
not ( n55105 , n55104 );
or ( n55106 , n55101 , n55105 );
nand ( n55107 , n52840 , n47368 );
nand ( n55108 , n55106 , n55107 );
nand ( n55109 , n52469 , n55108 );
nand ( n55110 , n55100 , n55109 );
not ( n55111 , n37669 );
not ( n55112 , n55111 );
not ( n55113 , n36589 );
not ( n55114 , n55113 );
or ( n55115 , n55112 , n55114 );
nand ( n55116 , n36589 , n37669 );
nand ( n55117 , n55115 , n55116 );
buf ( n55118 , n55117 );
not ( n55119 , n55118 );
not ( n55120 , n55119 );
and ( n55121 , n48689 , n55120 );
not ( n55122 , n48689 );
buf ( n55123 , n55118 );
buf ( n55124 , n55123 );
not ( n55125 , n55124 );
and ( n55126 , n55122 , n55125 );
nor ( n55127 , n55121 , n55126 );
not ( n55128 , n55127 );
not ( n55129 , n54841 );
not ( n55130 , n55111 );
not ( n55131 , n55113 );
or ( n55132 , n55130 , n55131 );
nand ( n55133 , n55132 , n55116 );
not ( n55134 , n55133 );
and ( n55135 , n55129 , n55134 );
and ( n55136 , n55133 , n54841 );
nor ( n55137 , n55135 , n55136 );
not ( n55138 , n54296 );
or ( n55139 , n55138 , n54840 );
nand ( n55140 , n54308 , n54840 );
nand ( n55141 , n55139 , n55140 );
nand ( n55142 , n55137 , n55141 );
not ( n55143 , n55142 );
buf ( n55144 , n55143 );
not ( n55145 , n55144 );
or ( n55146 , n55128 , n55145 );
not ( n55147 , n50914 );
not ( n55148 , n55118 );
not ( n55149 , n55148 );
or ( n55150 , n55147 , n55149 );
not ( n55151 , n55123 );
not ( n55152 , n55151 );
nand ( n55153 , n55152 , n48766 );
nand ( n55154 , n55150 , n55153 );
not ( n55155 , n54846 );
not ( n55156 , n55155 );
not ( n55157 , n55156 );
nand ( n55158 , n55154 , n55157 );
nand ( n55159 , n55146 , n55158 );
xor ( n55160 , n55110 , n55159 );
not ( n55161 , n54316 );
or ( n55162 , n55161 , n54727 );
not ( n55163 , n46273 );
not ( n55164 , n54468 );
or ( n55165 , n55163 , n55164 );
nand ( n55166 , n54298 , n46824 );
nand ( n55167 , n55165 , n55166 );
not ( n55168 , n55167 );
or ( n55169 , n55168 , n54326 );
nand ( n55170 , n55162 , n55169 );
xor ( n55171 , n55160 , n55170 );
xor ( n55172 , n55097 , n55171 );
xor ( n55173 , n55172 , n54935 );
xor ( n55174 , n55097 , n55171 );
and ( n55175 , n55174 , n54935 );
and ( n55176 , n55097 , n55171 );
or ( n55177 , n55175 , n55176 );
xor ( n55178 , n54947 , n54939 );
xor ( n55179 , n54639 , n54913 );
xor ( n55180 , n55179 , n54923 );
xor ( n55181 , n55178 , n55180 );
xor ( n55182 , n54947 , n54939 );
and ( n55183 , n55182 , n55180 );
and ( n55184 , n54947 , n54939 );
or ( n55185 , n55183 , n55184 );
not ( n55186 , n48295 );
not ( n55187 , n54756 );
or ( n55188 , n55186 , n55187 );
not ( n55189 , n46650 );
not ( n55190 , n40635 );
not ( n55191 , n55190 );
or ( n55192 , n55189 , n55191 );
nand ( n55193 , n40635 , n48078 );
nand ( n55194 , n55192 , n55193 );
nand ( n55195 , n55194 , n47827 );
nand ( n55196 , n55188 , n55195 );
not ( n55197 , n44004 );
not ( n55198 , n46072 );
not ( n55199 , n40380 );
not ( n55200 , n55199 );
or ( n55201 , n55198 , n55200 );
not ( n55202 , n40380 );
not ( n55203 , n55202 );
nand ( n55204 , n55203 , n46071 );
nand ( n55205 , n55201 , n55204 );
not ( n55206 , n55205 );
or ( n55207 , n55197 , n55206 );
nand ( n55208 , n54795 , n50659 );
nand ( n55209 , n55207 , n55208 );
xor ( n55210 , n55196 , n55209 );
not ( n55211 , n46564 );
not ( n55212 , n54816 );
or ( n55213 , n55211 , n55212 );
not ( n55214 , n47508 );
not ( n55215 , n40148 );
or ( n55216 , n55214 , n55215 );
nand ( n55217 , n54406 , n47514 );
nand ( n55218 , n55216 , n55217 );
not ( n55219 , n55218 );
or ( n55220 , n55219 , n50840 );
nand ( n55221 , n55213 , n55220 );
xor ( n55222 , n55210 , n55221 );
xor ( n55223 , n54943 , n55222 );
xor ( n55224 , n55223 , n54656 );
xor ( n55225 , n54943 , n55222 );
and ( n55226 , n55225 , n54656 );
and ( n55227 , n54943 , n55222 );
or ( n55228 , n55226 , n55227 );
not ( n55229 , n53510 );
not ( n55230 , n49500 );
not ( n55231 , n52222 );
or ( n55232 , n55230 , n55231 );
not ( n55233 , n52894 );
nand ( n55234 , n55233 , n47979 );
nand ( n55235 , n55232 , n55234 );
not ( n55236 , n55235 );
or ( n55237 , n55229 , n55236 );
nand ( n55238 , n54785 , n48989 );
nand ( n55239 , n55237 , n55238 );
not ( n55240 , n49026 );
not ( n55241 , n46425 );
not ( n55242 , n54433 );
not ( n55243 , n55242 );
or ( n55244 , n55241 , n55243 );
nand ( n55245 , n53660 , n46422 );
nand ( n55246 , n55244 , n55245 );
not ( n55247 , n55246 );
or ( n55248 , n55240 , n55247 );
nand ( n55249 , n54648 , n46267 );
nand ( n55250 , n55248 , n55249 );
xor ( n55251 , n55239 , n55250 );
not ( n55252 , n51865 );
not ( n55253 , n52267 );
not ( n55254 , n51574 );
or ( n55255 , n55253 , n55254 );
nand ( n55256 , n52289 , n52273 );
nand ( n55257 , n55255 , n55256 );
not ( n55258 , n55257 );
or ( n55259 , n55252 , n55258 );
nand ( n55260 , n54737 , n49713 );
nand ( n55261 , n55259 , n55260 );
xor ( n55262 , n55251 , n55261 );
not ( n55263 , n47148 );
not ( n55264 , n48856 );
not ( n55265 , n52917 );
or ( n55266 , n55264 , n55265 );
nand ( n55267 , n53228 , n52916 );
nand ( n55268 , n55266 , n55267 );
not ( n55269 , n55268 );
or ( n55270 , n55263 , n55269 );
nand ( n55271 , n54874 , n52421 );
nand ( n55272 , n55270 , n55271 );
buf ( n55273 , n54841 );
nand ( n55274 , n55273 , n48689 );
not ( n55275 , n55274 );
not ( n55276 , n54298 );
not ( n55277 , n55276 );
or ( n55278 , n55275 , n55277 );
not ( n55279 , n55273 );
nand ( n55280 , n55279 , n46441 );
nand ( n55281 , n55278 , n55280 );
and ( n55282 , n55281 , n55152 );
xor ( n55283 , n55272 , n55282 );
xor ( n55284 , n55283 , n54596 );
not ( n55285 , n53675 );
not ( n55286 , n47803 );
not ( n55287 , n54377 );
or ( n55288 , n55286 , n55287 );
nand ( n55289 , n54380 , n48727 );
nand ( n55290 , n55288 , n55289 );
not ( n55291 , n55290 );
or ( n55292 , n55285 , n55291 );
nand ( n55293 , n54775 , n47407 );
nand ( n55294 , n55292 , n55293 );
xor ( n55295 , n55284 , n55294 );
xor ( n55296 , n55295 , n55030 );
xor ( n55297 , n55262 , n55296 );
xor ( n55298 , n55297 , n54708 );
xor ( n55299 , n55262 , n55296 );
and ( n55300 , n55299 , n54708 );
and ( n55301 , n55262 , n55296 );
or ( n55302 , n55300 , n55301 );
xor ( n55303 , n55058 , n55173 );
xor ( n55304 , n55303 , n54748 );
xor ( n55305 , n55058 , n55173 );
and ( n55306 , n55305 , n54748 );
and ( n55307 , n55058 , n55173 );
or ( n55308 , n55306 , n55307 );
xor ( n55309 , n54766 , n55181 );
xor ( n55310 , n55309 , n54805 );
xor ( n55311 , n54766 , n55181 );
and ( n55312 , n55311 , n54805 );
and ( n55313 , n54766 , n55181 );
or ( n55314 , n55312 , n55313 );
xor ( n55315 , n55298 , n55224 );
xor ( n55316 , n55315 , n54885 );
xor ( n55317 , n55298 , n55224 );
and ( n55318 , n55317 , n54885 );
and ( n55319 , n55298 , n55224 );
or ( n55320 , n55318 , n55319 );
xor ( n55321 , n55304 , n54891 );
xor ( n55322 , n55321 , n55310 );
xor ( n55323 , n55304 , n54891 );
and ( n55324 , n55323 , n55310 );
and ( n55325 , n55304 , n54891 );
or ( n55326 , n55324 , n55325 );
xor ( n55327 , n54897 , n55316 );
xor ( n55328 , n55327 , n54903 );
xor ( n55329 , n54897 , n55316 );
and ( n55330 , n55329 , n54903 );
and ( n55331 , n54897 , n55316 );
or ( n55332 , n55330 , n55331 );
xor ( n55333 , n55272 , n55282 );
and ( n55334 , n55333 , n54596 );
and ( n55335 , n55272 , n55282 );
or ( n55336 , n55334 , n55335 );
xor ( n55337 , n55322 , n55328 );
xor ( n55338 , n55337 , n54909 );
xor ( n55339 , n55322 , n55328 );
and ( n55340 , n55339 , n54909 );
and ( n55341 , n55322 , n55328 );
or ( n55342 , n55340 , n55341 );
xor ( n55343 , n54982 , n55044 );
and ( n55344 , n55343 , n55055 );
and ( n55345 , n54982 , n55044 );
or ( n55346 , n55344 , n55345 );
xor ( n55347 , n55073 , n55083 );
and ( n55348 , n55347 , n55096 );
and ( n55349 , n55073 , n55083 );
or ( n55350 , n55348 , n55349 );
xor ( n55351 , n55110 , n55159 );
and ( n55352 , n55351 , n55170 );
and ( n55353 , n55110 , n55159 );
or ( n55354 , n55352 , n55353 );
xor ( n55355 , n54639 , n54913 );
and ( n55356 , n55355 , n54923 );
and ( n55357 , n54639 , n54913 );
or ( n55358 , n55356 , n55357 );
xor ( n55359 , n55196 , n55209 );
and ( n55360 , n55359 , n55221 );
and ( n55361 , n55196 , n55209 );
or ( n55362 , n55360 , n55361 );
xor ( n55363 , n55284 , n55294 );
and ( n55364 , n55363 , n55030 );
and ( n55365 , n55284 , n55294 );
or ( n55366 , n55364 , n55365 );
xor ( n55367 , n55239 , n55250 );
and ( n55368 , n55367 , n55261 );
and ( n55369 , n55239 , n55250 );
or ( n55370 , n55368 , n55369 );
not ( n55371 , n50554 );
not ( n55372 , n55003 );
or ( n55373 , n55371 , n55372 );
not ( n55374 , n48758 );
not ( n55375 , n48510 );
or ( n55376 , n55374 , n55375 );
nand ( n55377 , n44141 , n49092 );
nand ( n55378 , n55376 , n55377 );
nand ( n55379 , n55378 , n49320 );
nand ( n55380 , n55373 , n55379 );
not ( n55381 , n49979 );
not ( n55382 , n54953 );
or ( n55383 , n55381 , n55382 );
not ( n55384 , n50201 );
not ( n55385 , n51193 );
or ( n55386 , n55384 , n55385 );
nand ( n55387 , n41415 , n49282 );
nand ( n55388 , n55386 , n55387 );
nand ( n55389 , n55388 , n49288 );
nand ( n55390 , n55383 , n55389 );
xor ( n55391 , n55380 , n55390 );
or ( n55392 , n54959 , n54967 );
not ( n55393 , n49618 );
not ( n55394 , n48523 );
or ( n55395 , n55393 , n55394 );
nand ( n55396 , n41683 , n49769 );
nand ( n55397 , n55395 , n55396 );
not ( n55398 , n55397 );
or ( n55399 , n55398 , n49788 );
nand ( n55400 , n55392 , n55399 );
xor ( n55401 , n55391 , n55400 );
xor ( n55402 , n55380 , n55390 );
and ( n55403 , n55402 , n55400 );
and ( n55404 , n55380 , n55390 );
or ( n55405 , n55403 , n55404 );
not ( n55406 , n54979 );
not ( n55407 , n50321 );
or ( n55408 , n55406 , n55407 );
not ( n55409 , n53809 );
not ( n55410 , n50163 );
or ( n55411 , n55409 , n55410 );
nand ( n55412 , n50304 , n49968 );
nand ( n55413 , n55411 , n55412 );
nand ( n55414 , n55413 , n51452 );
nand ( n55415 , n55408 , n55414 );
and ( n55416 , n54995 , n55005 );
xor ( n55417 , n55415 , n55416 );
not ( n55418 , n52723 );
not ( n55419 , n48456 );
not ( n55420 , n48483 );
or ( n55421 , n55419 , n55420 );
nand ( n55422 , n53443 , n48486 );
nand ( n55423 , n55421 , n55422 );
not ( n55424 , n55423 );
or ( n55425 , n55418 , n55424 );
nand ( n55426 , n54991 , n53104 );
nand ( n55427 , n55425 , n55426 );
xor ( n55428 , n55417 , n55427 );
xor ( n55429 , n55415 , n55416 );
and ( n55430 , n55429 , n55427 );
and ( n55431 , n55415 , n55416 );
or ( n55432 , n55430 , n55431 );
not ( n55433 , n51865 );
not ( n55434 , n52267 );
not ( n55435 , n51925 );
or ( n55436 , n55434 , n55435 );
nand ( n55437 , n53258 , n48661 );
nand ( n55438 , n55436 , n55437 );
not ( n55439 , n55438 );
or ( n55440 , n55433 , n55439 );
nand ( n55441 , n55257 , n49713 );
nand ( n55442 , n55440 , n55441 );
not ( n55443 , n55133 );
not ( n55444 , n55443 );
and ( n55445 , n36655 , n37563 );
not ( n55446 , n36655 );
and ( n55447 , n55446 , n37562 );
nor ( n55448 , n55445 , n55447 );
not ( n55449 , n55448 );
or ( n55450 , n55444 , n55449 );
and ( n55451 , n36655 , n37563 );
not ( n55452 , n36655 );
and ( n55453 , n55452 , n37562 );
nor ( n55454 , n55451 , n55453 );
not ( n55455 , n55454 );
nand ( n55456 , n55455 , n55133 );
nand ( n55457 , n55450 , n55456 );
buf ( n55458 , n55457 );
buf ( n55459 , n55458 );
and ( n55460 , n55459 , n48689 );
xor ( n55461 , n55460 , n55401 );
xor ( n55462 , n55461 , n54986 );
xor ( n55463 , n55442 , n55462 );
xor ( n55464 , n55463 , n55354 );
xor ( n55465 , n55442 , n55462 );
and ( n55466 , n55465 , n55354 );
and ( n55467 , n55442 , n55462 );
or ( n55468 , n55466 , n55467 );
xor ( n55469 , n55346 , n55350 );
xor ( n55470 , n55469 , n55358 );
xor ( n55471 , n55346 , n55350 );
and ( n55472 , n55471 , n55358 );
and ( n55473 , n55346 , n55350 );
or ( n55474 , n55472 , n55473 );
not ( n55475 , n55108 );
not ( n55476 , n52853 );
or ( n55477 , n55475 , n55476 );
not ( n55478 , n48898 );
not ( n55479 , n53946 );
or ( n55480 , n55478 , n55479 );
not ( n55481 , n52837 );
nand ( n55482 , n55481 , n48897 );
nand ( n55483 , n55480 , n55482 );
nand ( n55484 , n52469 , n55483 );
nand ( n55485 , n55477 , n55484 );
not ( n55486 , n55094 );
not ( n55487 , n53609 );
or ( n55488 , n55486 , n55487 );
not ( n55489 , n47227 );
not ( n55490 , n53595 );
or ( n55491 , n55489 , n55490 );
nand ( n55492 , n53590 , n47589 );
nand ( n55493 , n55491 , n55492 );
nand ( n55494 , n55493 , n53326 );
nand ( n55495 , n55488 , n55494 );
xor ( n55496 , n55485 , n55495 );
not ( n55497 , n55167 );
not ( n55498 , n54316 );
or ( n55499 , n55497 , n55498 );
not ( n55500 , n47646 );
not ( n55501 , n54467 );
or ( n55502 , n55500 , n55501 );
nand ( n55503 , n54297 , n47650 );
nand ( n55504 , n55502 , n55503 );
nand ( n55505 , n54077 , n55504 );
nand ( n55506 , n55499 , n55505 );
xor ( n55507 , n55496 , n55506 );
not ( n55508 , n55053 );
not ( n55509 , n51215 );
or ( n55510 , n55508 , n55509 );
not ( n55511 , n51670 );
not ( n55512 , n55511 );
not ( n55513 , n50916 );
or ( n55514 , n55512 , n55513 );
nand ( n55515 , n50898 , n51670 );
nand ( n55516 , n55514 , n55515 );
nand ( n55517 , n55516 , n51223 );
nand ( n55518 , n55510 , n55517 );
not ( n55519 , n55071 );
not ( n55520 , n52139 );
or ( n55521 , n55519 , n55520 );
and ( n55522 , n51792 , n51504 );
not ( n55523 , n51792 );
and ( n55524 , n55523 , n51818 );
or ( n55525 , n55522 , n55524 );
nand ( n55526 , n51533 , n55525 );
nand ( n55527 , n55521 , n55526 );
xor ( n55528 , n55518 , n55527 );
not ( n55529 , n55081 );
not ( n55530 , n52482 );
or ( n55531 , n55529 , n55530 );
not ( n55532 , n51204 );
not ( n55533 , n52130 );
or ( n55534 , n55532 , n55533 );
nand ( n55535 , n53918 , n48860 );
nand ( n55536 , n55534 , n55535 );
nand ( n55537 , n51766 , n55536 );
nand ( n55538 , n55531 , n55537 );
xor ( n55539 , n55528 , n55538 );
xor ( n55540 , n55507 , n55539 );
not ( n55541 , n52962 );
not ( n55542 , n50232 );
not ( n55543 , n51841 );
or ( n55544 , n55542 , n55543 );
nand ( n55545 , n40691 , n52048 );
nand ( n55546 , n55544 , n55545 );
not ( n55547 , n55546 );
or ( n55548 , n55541 , n55547 );
nand ( n55549 , n55040 , n52970 );
nand ( n55550 , n55548 , n55549 );
xor ( n55551 , n55550 , n55336 );
not ( n55552 , n46776 );
not ( n55553 , n55194 );
or ( n55554 , n55552 , n55553 );
not ( n55555 , n46650 );
not ( n55556 , n53286 );
or ( n55557 , n55555 , n55556 );
nand ( n55558 , n40377 , n50087 );
nand ( n55559 , n55557 , n55558 );
nand ( n55560 , n55559 , n53631 );
nand ( n55561 , n55554 , n55560 );
xor ( n55562 , n55551 , n55561 );
xor ( n55563 , n55540 , n55562 );
xor ( n55564 , n55507 , n55539 );
and ( n55565 , n55564 , n55562 );
and ( n55566 , n55507 , n55539 );
or ( n55567 , n55565 , n55566 );
xor ( n55568 , n55362 , n55366 );
xor ( n55569 , n55568 , n55370 );
xor ( n55570 , n55362 , n55366 );
and ( n55571 , n55570 , n55370 );
and ( n55572 , n55362 , n55366 );
or ( n55573 , n55571 , n55572 );
not ( n55574 , n55154 );
buf ( n55575 , n55142 );
not ( n55576 , n55575 );
not ( n55577 , n55576 );
or ( n55578 , n55574 , n55577 );
not ( n55579 , n54722 );
not ( n55580 , n55148 );
or ( n55581 , n55579 , n55580 );
not ( n55582 , n55148 );
nand ( n55583 , n55582 , n54721 );
nand ( n55584 , n55581 , n55583 );
nand ( n55585 , n55584 , n55157 );
nand ( n55586 , n55578 , n55585 );
xor ( n55587 , n55586 , n55428 );
xor ( n55588 , n55587 , n55034 );
not ( n55589 , n47407 );
not ( n55590 , n55290 );
or ( n55591 , n55589 , n55590 );
not ( n55592 , n47803 );
not ( n55593 , n54046 );
or ( n55594 , n55592 , n55593 );
nand ( n55595 , n40626 , n48727 );
nand ( n55596 , n55594 , n55595 );
nand ( n55597 , n55596 , n53675 );
nand ( n55598 , n55591 , n55597 );
not ( n55599 , n49252 );
not ( n55600 , n55235 );
or ( n55601 , n55599 , n55600 );
not ( n55602 , n47980 );
not ( n55603 , n40527 );
or ( n55604 , n55602 , n55603 );
nand ( n55605 , n40526 , n47979 );
nand ( n55606 , n55604 , n55605 );
nand ( n55607 , n55606 , n47384 );
nand ( n55608 , n55601 , n55607 );
xor ( n55609 , n55598 , n55608 );
not ( n55610 , n46267 );
not ( n55611 , n55246 );
or ( n55612 , n55610 , n55611 );
not ( n55613 , n46425 );
not ( n55614 , n54811 );
or ( n55615 , n55613 , n55614 );
nand ( n55616 , n40364 , n46422 );
nand ( n55617 , n55615 , n55616 );
nand ( n55618 , n55617 , n49026 );
nand ( n55619 , n55612 , n55618 );
xor ( n55620 , n55609 , n55619 );
xor ( n55621 , n55588 , n55620 );
xor ( n55622 , n55621 , n55062 );
xor ( n55623 , n55588 , n55620 );
and ( n55624 , n55623 , n55062 );
and ( n55625 , n55588 , n55620 );
or ( n55626 , n55624 , n55625 );
not ( n55627 , n50659 );
not ( n55628 , n55205 );
or ( n55629 , n55627 , n55628 );
not ( n55630 , n40451 );
and ( n55631 , n46072 , n55630 );
not ( n55632 , n46072 );
and ( n55633 , n55632 , n40452 );
or ( n55634 , n55631 , n55633 );
nand ( n55635 , n55634 , n46602 );
nand ( n55636 , n55629 , n55635 );
not ( n55637 , n46564 );
not ( n55638 , n55218 );
or ( n55639 , n55637 , n55638 );
not ( n55640 , n47514 );
not ( n55641 , n40388 );
not ( n55642 , n55641 );
not ( n55643 , n55642 );
or ( n55644 , n55640 , n55643 );
not ( n55645 , n54790 );
not ( n55646 , n55645 );
nand ( n55647 , n55646 , n48952 );
nand ( n55648 , n55644 , n55647 );
nand ( n55649 , n55648 , n49832 );
nand ( n55650 , n55639 , n55649 );
xor ( n55651 , n55636 , n55650 );
not ( n55652 , n49116 );
not ( n55653 , n55015 );
or ( n55654 , n55652 , n55653 );
not ( n55655 , n52377 );
not ( n55656 , n50546 );
or ( n55657 , n55655 , n55656 );
nand ( n55658 , n40854 , n55013 );
nand ( n55659 , n55657 , n55658 );
nand ( n55660 , n55659 , n52004 );
nand ( n55661 , n55654 , n55660 );
not ( n55662 , n52022 );
not ( n55663 , n55025 );
or ( n55664 , n55662 , n55663 );
not ( n55665 , n47855 );
not ( n55666 , n41284 );
or ( n55667 , n55665 , n55666 );
nand ( n55668 , n48996 , n52016 );
nand ( n55669 , n55667 , n55668 );
nand ( n55670 , n55669 , n54623 );
nand ( n55671 , n55664 , n55670 );
xor ( n55672 , n55661 , n55671 );
not ( n55673 , n47148 );
not ( n55674 , n51891 );
and ( n55675 , n55674 , n51723 );
not ( n55676 , n55674 );
and ( n55677 , n55676 , n51724 );
or ( n55678 , n55675 , n55677 );
not ( n55679 , n55678 );
or ( n55680 , n55673 , n55679 );
nand ( n55681 , n55268 , n52421 );
nand ( n55682 , n55680 , n55681 );
xor ( n55683 , n55672 , n55682 );
xor ( n55684 , n55651 , n55683 );
xor ( n55685 , n55684 , n55177 );
xor ( n55686 , n55685 , n55470 );
xor ( n55687 , n55684 , n55177 );
and ( n55688 , n55687 , n55470 );
and ( n55689 , n55684 , n55177 );
or ( n55690 , n55688 , n55689 );
xor ( n55691 , n55464 , n55563 );
xor ( n55692 , n55691 , n55185 );
xor ( n55693 , n55464 , n55563 );
and ( n55694 , n55693 , n55185 );
and ( n55695 , n55464 , n55563 );
or ( n55696 , n55694 , n55695 );
xor ( n55697 , n55569 , n55228 );
xor ( n55698 , n55697 , n55622 );
xor ( n55699 , n55569 , n55228 );
and ( n55700 , n55699 , n55622 );
and ( n55701 , n55569 , n55228 );
or ( n55702 , n55700 , n55701 );
xor ( n55703 , n55302 , n55686 );
xor ( n55704 , n55703 , n55308 );
xor ( n55705 , n55302 , n55686 );
and ( n55706 , n55705 , n55308 );
and ( n55707 , n55302 , n55686 );
or ( n55708 , n55706 , n55707 );
xor ( n55709 , n55314 , n55692 );
xor ( n55710 , n55709 , n55698 );
xor ( n55711 , n55314 , n55692 );
and ( n55712 , n55711 , n55698 );
and ( n55713 , n55314 , n55692 );
or ( n55714 , n55712 , n55713 );
xor ( n55715 , n55661 , n55671 );
and ( n55716 , n55715 , n55682 );
and ( n55717 , n55661 , n55671 );
or ( n55718 , n55716 , n55717 );
xor ( n55719 , n55320 , n55704 );
xor ( n55720 , n55719 , n55326 );
xor ( n55721 , n55320 , n55704 );
and ( n55722 , n55721 , n55326 );
and ( n55723 , n55320 , n55704 );
or ( n55724 , n55722 , n55723 );
xor ( n55725 , n55710 , n55332 );
xor ( n55726 , n55725 , n55720 );
xor ( n55727 , n55710 , n55332 );
and ( n55728 , n55727 , n55720 );
and ( n55729 , n55710 , n55332 );
or ( n55730 , n55728 , n55729 );
xor ( n55731 , n55460 , n55401 );
and ( n55732 , n55731 , n54986 );
and ( n55733 , n55460 , n55401 );
or ( n55734 , n55732 , n55733 );
xor ( n55735 , n55518 , n55527 );
and ( n55736 , n55735 , n55538 );
and ( n55737 , n55518 , n55527 );
or ( n55738 , n55736 , n55737 );
xor ( n55739 , n55485 , n55495 );
and ( n55740 , n55739 , n55506 );
and ( n55741 , n55485 , n55495 );
or ( n55742 , n55740 , n55741 );
xor ( n55743 , n55586 , n55428 );
and ( n55744 , n55743 , n55034 );
and ( n55745 , n55586 , n55428 );
or ( n55746 , n55744 , n55745 );
xor ( n55747 , n55550 , n55336 );
and ( n55748 , n55747 , n55561 );
and ( n55749 , n55550 , n55336 );
or ( n55750 , n55748 , n55749 );
xor ( n55751 , n55636 , n55650 );
and ( n55752 , n55751 , n55683 );
and ( n55753 , n55636 , n55650 );
or ( n55754 , n55752 , n55753 );
xor ( n55755 , n55598 , n55608 );
and ( n55756 , n55755 , n55619 );
and ( n55757 , n55598 , n55608 );
or ( n55758 , n55756 , n55757 );
not ( n55759 , n55397 );
not ( n55760 , n50565 );
or ( n55761 , n55759 , n55760 );
not ( n55762 , n49618 );
not ( n55763 , n49220 );
or ( n55764 , n55762 , n55763 );
nand ( n55765 , n30929 , n49769 );
nand ( n55766 , n55764 , n55765 );
nand ( n55767 , n55766 , n51809 );
nand ( n55768 , n55761 , n55767 );
not ( n55769 , n55413 );
not ( n55770 , n50929 );
or ( n55771 , n55769 , n55770 );
not ( n55772 , n50304 );
not ( n55773 , n47178 );
or ( n55774 , n55772 , n55773 );
nand ( n55775 , n50327 , n41692 );
nand ( n55776 , n55774 , n55775 );
nand ( n55777 , n55776 , n49920 );
nand ( n55778 , n55771 , n55777 );
xor ( n55779 , n55768 , n55778 );
not ( n55780 , n50554 );
not ( n55781 , n55378 );
or ( n55782 , n55780 , n55781 );
not ( n55783 , n49313 );
not ( n55784 , n41530 );
or ( n55785 , n55783 , n55784 );
nand ( n55786 , n49232 , n49092 );
nand ( n55787 , n55785 , n55786 );
nand ( n55788 , n55787 , n49320 );
nand ( n55789 , n55782 , n55788 );
not ( n55790 , n49452 );
not ( n55791 , n49756 );
or ( n55792 , n55790 , n55791 );
nand ( n55793 , n49110 , n41575 );
nand ( n55794 , n55792 , n55793 );
not ( n55795 , n55794 );
not ( n55796 , n49288 );
or ( n55797 , n55795 , n55796 );
nand ( n55798 , n55388 , n51337 );
nand ( n55799 , n55797 , n55798 );
xor ( n55800 , n55789 , n55799 );
xor ( n55801 , n55779 , n55800 );
xor ( n55802 , n55768 , n55778 );
and ( n55803 , n55802 , n55800 );
and ( n55804 , n55768 , n55778 );
or ( n55805 , n55803 , n55804 );
not ( n55806 , n48240 );
not ( n55807 , n51680 );
not ( n55808 , n41216 );
or ( n55809 , n55807 , n55808 );
nand ( n55810 , n50973 , n52016 );
nand ( n55811 , n55809 , n55810 );
not ( n55812 , n55811 );
or ( n55813 , n55806 , n55812 );
nand ( n55814 , n55669 , n47873 );
nand ( n55815 , n55813 , n55814 );
not ( n55816 , n52723 );
not ( n55817 , n48456 );
not ( n55818 , n48679 );
or ( n55819 , n55817 , n55818 );
nand ( n55820 , n41364 , n52728 );
nand ( n55821 , n55819 , n55820 );
not ( n55822 , n55821 );
or ( n55823 , n55816 , n55822 );
nand ( n55824 , n55423 , n50176 );
nand ( n55825 , n55823 , n55824 );
xor ( n55826 , n55815 , n55825 );
not ( n55827 , n46440 );
not ( n55828 , n55454 );
or ( n55829 , n55827 , n55828 );
nand ( n55830 , n55829 , n55151 );
not ( n55831 , n55454 );
nand ( n55832 , n55831 , n46441 );
and ( n55833 , n55830 , n55832 );
not ( n55834 , n37539 );
not ( n55835 , n36341 );
or ( n55836 , n55834 , n55835 );
nand ( n55837 , n55836 , n37443 );
nand ( n55838 , n33568 , n33393 );
not ( n55839 , n55838 );
and ( n55840 , n55837 , n55839 );
not ( n55841 , n55837 );
and ( n55842 , n55841 , n55838 );
nor ( n55843 , n55840 , n55842 );
buf ( n55844 , n55843 );
buf ( n55845 , n55844 );
not ( n55846 , n55845 );
nor ( n55847 , n55833 , n55846 );
xor ( n55848 , n55826 , n55847 );
xor ( n55849 , n55815 , n55825 );
and ( n55850 , n55849 , n55847 );
and ( n55851 , n55815 , n55825 );
or ( n55852 , n55850 , n55851 );
xor ( n55853 , n55734 , n55742 );
xor ( n55854 , n55853 , n55738 );
xor ( n55855 , n55734 , n55742 );
and ( n55856 , n55855 , n55738 );
and ( n55857 , n55734 , n55742 );
or ( n55858 , n55856 , n55857 );
not ( n55859 , n55504 );
not ( n55860 , n54315 );
or ( n55861 , n55859 , n55860 );
and ( n55862 , n49734 , n54297 );
not ( n55863 , n49734 );
and ( n55864 , n55863 , n54301 );
nor ( n55865 , n55862 , n55864 );
buf ( n55866 , n54076 );
not ( n55867 , n55866 );
nand ( n55868 , n55865 , n55867 );
nand ( n55869 , n55861 , n55868 );
xor ( n55870 , n55801 , n55869 );
not ( n55871 , n48689 );
buf ( n55872 , n55845 );
not ( n55873 , n55872 );
not ( n55874 , n55873 );
or ( n55875 , n55871 , n55874 );
not ( n55876 , n55845 );
not ( n55877 , n55876 );
nand ( n55878 , n55877 , n46441 );
nand ( n55879 , n55875 , n55878 );
not ( n55880 , n55879 );
and ( n55881 , n55117 , n55455 );
not ( n55882 , n55117 );
and ( n55883 , n55882 , n55454 );
nor ( n55884 , n55881 , n55883 );
xor ( n55885 , n55844 , n55454 );
nand ( n55886 , n55884 , n55885 );
not ( n55887 , n55886 );
not ( n55888 , n55887 );
or ( n55889 , n55880 , n55888 );
not ( n55890 , n50914 );
buf ( n55891 , n55844 );
buf ( n55892 , n55891 );
not ( n55893 , n55892 );
not ( n55894 , n55893 );
or ( n55895 , n55890 , n55894 );
nand ( n55896 , n55891 , n45767 );
nand ( n55897 , n55895 , n55896 );
nand ( n55898 , n55458 , n55897 );
nand ( n55899 , n55889 , n55898 );
xor ( n55900 , n55870 , n55899 );
xor ( n55901 , n55746 , n55900 );
not ( n55902 , n55483 );
not ( n55903 , n52853 );
or ( n55904 , n55902 , n55903 );
not ( n55905 , n47765 );
not ( n55906 , n52837 );
or ( n55907 , n55905 , n55906 );
nand ( n55908 , n55481 , n48589 );
nand ( n55909 , n55907 , n55908 );
nand ( n55910 , n55909 , n53571 );
nand ( n55911 , n55904 , n55910 );
not ( n55912 , n55493 );
and ( n55913 , n53606 , n53607 );
not ( n55914 , n55913 );
or ( n55915 , n55912 , n55914 );
not ( n55916 , n49654 );
not ( n55917 , n53590 );
buf ( n55918 , n55917 );
not ( n55919 , n55918 );
or ( n55920 , n55916 , n55919 );
nand ( n55921 , n53590 , n47368 );
nand ( n55922 , n55920 , n55921 );
nand ( n55923 , n55922 , n53326 );
nand ( n55924 , n55915 , n55923 );
xor ( n55925 , n55911 , n55924 );
not ( n55926 , n55584 );
not ( n55927 , n55576 );
or ( n55928 , n55926 , n55927 );
and ( n55929 , n46273 , n55148 );
not ( n55930 , n46273 );
and ( n55931 , n55930 , n55124 );
or ( n55932 , n55929 , n55931 );
not ( n55933 , n54846 );
buf ( n55934 , n55933 );
nand ( n55935 , n55932 , n55934 );
nand ( n55936 , n55928 , n55935 );
xor ( n55937 , n55925 , n55936 );
xor ( n55938 , n55901 , n55937 );
xor ( n55939 , n55746 , n55900 );
and ( n55940 , n55939 , n55937 );
and ( n55941 , n55746 , n55900 );
or ( n55942 , n55940 , n55941 );
not ( n55943 , n55516 );
not ( n55944 , n51215 );
or ( n55945 , n55943 , n55944 );
not ( n55946 , n48223 );
not ( n55947 , n50916 );
or ( n55948 , n55946 , n55947 );
nand ( n55949 , n50898 , n54184 );
nand ( n55950 , n55948 , n55949 );
nand ( n55951 , n55950 , n51223 );
nand ( n55952 , n55945 , n55951 );
not ( n55953 , n55525 );
not ( n55954 , n52139 );
or ( n55955 , n55953 , n55954 );
not ( n55956 , n52033 );
not ( n55957 , n51508 );
or ( n55958 , n55956 , n55957 );
not ( n55959 , n52033 );
nand ( n55960 , n51818 , n55959 );
nand ( n55961 , n55958 , n55960 );
nand ( n55962 , n55961 , n51533 );
nand ( n55963 , n55955 , n55962 );
xor ( n55964 , n55952 , n55963 );
not ( n55965 , n55536 );
not ( n55966 , n52125 );
or ( n55967 , n55965 , n55966 );
not ( n55968 , n49624 );
not ( n55969 , n52130 );
or ( n55970 , n55968 , n55969 );
nand ( n55971 , n52870 , n49630 );
nand ( n55972 , n55970 , n55971 );
nand ( n55973 , n51766 , n55972 );
nand ( n55974 , n55967 , n55973 );
xor ( n55975 , n55964 , n55974 );
xor ( n55976 , n55975 , n55750 );
xor ( n55977 , n55432 , n55718 );
not ( n55978 , n52004 );
and ( n55979 , n52377 , n49806 );
not ( n55980 , n52377 );
and ( n55981 , n55980 , n50827 );
or ( n55982 , n55979 , n55981 );
not ( n55983 , n55982 );
or ( n55984 , n55978 , n55983 );
nand ( n55985 , n55659 , n49116 );
nand ( n55986 , n55984 , n55985 );
xor ( n55987 , n55405 , n55986 );
not ( n55988 , n54875 );
not ( n55989 , n51723 );
not ( n55990 , n50400 );
or ( n55991 , n55989 , n55990 );
nand ( n55992 , n41132 , n53228 );
nand ( n55993 , n55991 , n55992 );
not ( n55994 , n55993 );
or ( n55995 , n55988 , n55994 );
nand ( n55996 , n55678 , n52421 );
nand ( n55997 , n55995 , n55996 );
xor ( n55998 , n55987 , n55997 );
xor ( n55999 , n55977 , n55998 );
xor ( n56000 , n55976 , n55999 );
xor ( n56001 , n55975 , n55750 );
and ( n56002 , n56001 , n55999 );
and ( n56003 , n55975 , n55750 );
or ( n56004 , n56002 , n56003 );
xor ( n56005 , n55758 , n55754 );
not ( n56006 , n46267 );
not ( n56007 , n55617 );
or ( n56008 , n56006 , n56007 );
not ( n56009 , n46425 );
buf ( n56010 , n40147 );
not ( n56011 , n56010 );
not ( n56012 , n56011 );
or ( n56013 , n56009 , n56012 );
nand ( n56014 , n40149 , n46422 );
nand ( n56015 , n56013 , n56014 );
nand ( n56016 , n56015 , n49026 );
nand ( n56017 , n56008 , n56016 );
not ( n56018 , n47009 );
not ( n56019 , n46072 );
not ( n56020 , n40512 );
not ( n56021 , n56020 );
or ( n56022 , n56019 , n56021 );
not ( n56023 , n56020 );
nand ( n56024 , n56023 , n50405 );
nand ( n56025 , n56022 , n56024 );
not ( n56026 , n56025 );
or ( n56027 , n56018 , n56026 );
nand ( n56028 , n55634 , n50659 );
nand ( n56029 , n56027 , n56028 );
xor ( n56030 , n56017 , n56029 );
not ( n56031 , n49713 );
not ( n56032 , n55438 );
or ( n56033 , n56031 , n56032 );
not ( n56034 , n52267 );
not ( n56035 , n52894 );
or ( n56036 , n56034 , n56035 );
nand ( n56037 , n52223 , n51351 );
nand ( n56038 , n56036 , n56037 );
nand ( n56039 , n56038 , n51865 );
nand ( n56040 , n56033 , n56039 );
xor ( n56041 , n56030 , n56040 );
xor ( n56042 , n56005 , n56041 );
xor ( n56043 , n55758 , n55754 );
and ( n56044 , n56043 , n56041 );
and ( n56045 , n55758 , n55754 );
or ( n56046 , n56044 , n56045 );
not ( n56047 , n55546 );
not ( n56048 , n52970 );
or ( n56049 , n56047 , n56048 );
and ( n56050 , n48645 , n50958 );
not ( n56051 , n48645 );
and ( n56052 , n56051 , n40677 );
nor ( n56053 , n56050 , n56052 );
or ( n56054 , n56053 , n50239 );
nand ( n56055 , n56049 , n56054 );
not ( n56056 , n49832 );
not ( n56057 , n47508 );
not ( n56058 , n40381 );
not ( n56059 , n56058 );
or ( n56060 , n56057 , n56059 );
nand ( n56061 , n55203 , n51577 );
nand ( n56062 , n56060 , n56061 );
not ( n56063 , n56062 );
or ( n56064 , n56056 , n56063 );
nand ( n56065 , n55648 , n46564 );
nand ( n56066 , n56064 , n56065 );
xor ( n56067 , n56055 , n56066 );
not ( n56068 , n55559 );
not ( n56069 , n48295 );
or ( n56070 , n56068 , n56069 );
not ( n56071 , n46650 );
not ( n56072 , n54432 );
not ( n56073 , n56072 );
not ( n56074 , n56073 );
not ( n56075 , n56074 );
or ( n56076 , n56071 , n56075 );
nand ( n56077 , n53660 , n50087 );
nand ( n56078 , n56076 , n56077 );
not ( n56079 , n56078 );
not ( n56080 , n50261 );
or ( n56081 , n56079 , n56080 );
nand ( n56082 , n56070 , n56081 );
xor ( n56083 , n56067 , n56082 );
not ( n56084 , n48929 );
not ( n56085 , n47803 );
not ( n56086 , n55190 );
or ( n56087 , n56085 , n56086 );
nand ( n56088 , n50634 , n40635 );
nand ( n56089 , n56087 , n56088 );
not ( n56090 , n56089 );
or ( n56091 , n56084 , n56090 );
nand ( n56092 , n55596 , n47407 );
nand ( n56093 , n56091 , n56092 );
xor ( n56094 , n56093 , n55848 );
not ( n56095 , n47384 );
not ( n56096 , n47980 );
not ( n56097 , n53730 );
or ( n56098 , n56096 , n56097 );
nand ( n56099 , n52212 , n47979 );
nand ( n56100 , n56098 , n56099 );
not ( n56101 , n56100 );
or ( n56102 , n56095 , n56101 );
nand ( n56103 , n55606 , n49252 );
nand ( n56104 , n56102 , n56103 );
xor ( n56105 , n56094 , n56104 );
xor ( n56106 , n56083 , n56105 );
xor ( n56107 , n56106 , n55468 );
xor ( n56108 , n56083 , n56105 );
and ( n56109 , n56108 , n55468 );
and ( n56110 , n56083 , n56105 );
or ( n56111 , n56109 , n56110 );
xor ( n56112 , n55474 , n55854 );
xor ( n56113 , n56112 , n55938 );
xor ( n56114 , n55474 , n55854 );
and ( n56115 , n56114 , n55938 );
and ( n56116 , n55474 , n55854 );
or ( n56117 , n56115 , n56116 );
xor ( n56118 , n55567 , n55573 );
xor ( n56119 , n56118 , n56042 );
xor ( n56120 , n55567 , n55573 );
and ( n56121 , n56120 , n56042 );
and ( n56122 , n55567 , n55573 );
or ( n56123 , n56121 , n56122 );
xor ( n56124 , n55626 , n56000 );
xor ( n56125 , n56124 , n55690 );
xor ( n56126 , n55626 , n56000 );
and ( n56127 , n56126 , n55690 );
and ( n56128 , n55626 , n56000 );
or ( n56129 , n56127 , n56128 );
xor ( n56130 , n56107 , n56113 );
xor ( n56131 , n56130 , n55696 );
xor ( n56132 , n56107 , n56113 );
and ( n56133 , n56132 , n55696 );
and ( n56134 , n56107 , n56113 );
or ( n56135 , n56133 , n56134 );
xor ( n56136 , n56119 , n55702 );
xor ( n56137 , n56136 , n56125 );
xor ( n56138 , n56119 , n55702 );
and ( n56139 , n56138 , n56125 );
and ( n56140 , n56119 , n55702 );
or ( n56141 , n56139 , n56140 );
xor ( n56142 , n55405 , n55986 );
and ( n56143 , n56142 , n55997 );
and ( n56144 , n55405 , n55986 );
or ( n56145 , n56143 , n56144 );
xor ( n56146 , n55708 , n56131 );
xor ( n56147 , n56146 , n55714 );
xor ( n56148 , n55708 , n56131 );
and ( n56149 , n56148 , n55714 );
and ( n56150 , n55708 , n56131 );
or ( n56151 , n56149 , n56150 );
xor ( n56152 , n56137 , n56147 );
xor ( n56153 , n56152 , n55724 );
xor ( n56154 , n56137 , n56147 );
and ( n56155 , n56154 , n55724 );
and ( n56156 , n56137 , n56147 );
or ( n56157 , n56155 , n56156 );
xor ( n56158 , n55952 , n55963 );
and ( n56159 , n56158 , n55974 );
and ( n56160 , n55952 , n55963 );
or ( n56161 , n56159 , n56160 );
xor ( n56162 , n55911 , n55924 );
and ( n56163 , n56162 , n55936 );
and ( n56164 , n55911 , n55924 );
or ( n56165 , n56163 , n56164 );
xor ( n56166 , n55801 , n55869 );
and ( n56167 , n56166 , n55899 );
and ( n56168 , n55801 , n55869 );
or ( n56169 , n56167 , n56168 );
xor ( n56170 , n55432 , n55718 );
and ( n56171 , n56170 , n55998 );
and ( n56172 , n55432 , n55718 );
or ( n56173 , n56171 , n56172 );
xor ( n56174 , n56055 , n56066 );
and ( n56175 , n56174 , n56082 );
and ( n56176 , n56055 , n56066 );
or ( n56177 , n56175 , n56176 );
xor ( n56178 , n56093 , n55848 );
and ( n56179 , n56178 , n56104 );
and ( n56180 , n56093 , n55848 );
or ( n56181 , n56179 , n56180 );
xor ( n56182 , n56017 , n56029 );
and ( n56183 , n56182 , n56040 );
and ( n56184 , n56017 , n56029 );
or ( n56185 , n56183 , n56184 );
not ( n56186 , n48891 );
not ( n56187 , n49452 );
not ( n56188 , n48510 );
or ( n56189 , n56187 , n56188 );
nand ( n56190 , n44141 , n49283 );
nand ( n56191 , n56189 , n56190 );
not ( n56192 , n56191 );
or ( n56193 , n56186 , n56192 );
nand ( n56194 , n55794 , n49979 );
nand ( n56195 , n56193 , n56194 );
not ( n56196 , n55766 );
not ( n56197 , n49779 );
or ( n56198 , n56196 , n56197 );
not ( n56199 , n49618 );
not ( n56200 , n51193 );
or ( n56201 , n56199 , n56200 );
nand ( n56202 , n52379 , n50292 );
nand ( n56203 , n56201 , n56202 );
nand ( n56204 , n56203 , n51809 );
nand ( n56205 , n56198 , n56204 );
xor ( n56206 , n56195 , n56205 );
not ( n56207 , n55776 );
not ( n56208 , n52749 );
or ( n56209 , n56207 , n56208 );
not ( n56210 , n51250 );
not ( n56211 , n48523 );
or ( n56212 , n56210 , n56211 );
nand ( n56213 , n54614 , n53114 );
nand ( n56214 , n56212 , n56213 );
nand ( n56215 , n56214 , n50331 );
nand ( n56216 , n56209 , n56215 );
xor ( n56217 , n56206 , n56216 );
xor ( n56218 , n56195 , n56205 );
and ( n56219 , n56218 , n56216 );
and ( n56220 , n56195 , n56205 );
or ( n56221 , n56219 , n56220 );
and ( n56222 , n55789 , n55799 );
not ( n56223 , n49737 );
not ( n56224 , n48705 );
not ( n56225 , n50631 );
or ( n56226 , n56224 , n56225 );
buf ( n56227 , n48749 );
nand ( n56228 , n51123 , n56227 );
nand ( n56229 , n56226 , n56228 );
not ( n56230 , n56229 );
or ( n56231 , n56223 , n56230 );
nand ( n56232 , n49309 , n55787 );
nand ( n56233 , n56231 , n56232 );
xor ( n56234 , n56222 , n56233 );
not ( n56235 , n54623 );
not ( n56236 , n47855 );
not ( n56237 , n50004 );
or ( n56238 , n56236 , n56237 );
not ( n56239 , n50546 );
nand ( n56240 , n56239 , n52016 );
nand ( n56241 , n56238 , n56240 );
not ( n56242 , n56241 );
or ( n56243 , n56235 , n56242 );
nand ( n56244 , n55811 , n47873 );
nand ( n56245 , n56243 , n56244 );
xor ( n56246 , n56234 , n56245 );
xor ( n56247 , n56222 , n56233 );
and ( n56248 , n56247 , n56245 );
and ( n56249 , n56222 , n56233 );
or ( n56250 , n56248 , n56249 );
not ( n56251 , n49713 );
not ( n56252 , n56038 );
or ( n56253 , n56251 , n56252 );
not ( n56254 , n52267 );
not ( n56255 , n54771 );
or ( n56256 , n56254 , n56255 );
nand ( n56257 , n40526 , n48661 );
nand ( n56258 , n56256 , n56257 );
nand ( n56259 , n56258 , n51865 );
nand ( n56260 , n56253 , n56259 );
xor ( n56261 , n56260 , n56145 );
xor ( n56262 , n56261 , n56165 );
xor ( n56263 , n56260 , n56145 );
and ( n56264 , n56263 , n56165 );
and ( n56265 , n56260 , n56145 );
or ( n56266 , n56264 , n56265 );
xor ( n56267 , n56169 , n56161 );
not ( n56268 , n55865 );
not ( n56269 , n54314 );
not ( n56270 , n56269 );
or ( n56271 , n56268 , n56270 );
and ( n56272 , n47589 , n54301 );
not ( n56273 , n47589 );
not ( n56274 , n54301 );
and ( n56275 , n56273 , n56274 );
nor ( n56276 , n56272 , n56275 );
not ( n56277 , n54076 );
nand ( n56278 , n56276 , n56277 );
nand ( n56279 , n56271 , n56278 );
not ( n56280 , n55897 );
not ( n56281 , n55886 );
not ( n56282 , n56281 );
or ( n56283 , n56280 , n56282 );
not ( n56284 , n54722 );
not ( n56285 , n55845 );
not ( n56286 , n56285 );
or ( n56287 , n56284 , n56286 );
nand ( n56288 , n55892 , n47306 );
nand ( n56289 , n56287 , n56288 );
nand ( n56290 , n56289 , n55459 );
nand ( n56291 , n56283 , n56290 );
xor ( n56292 , n56279 , n56291 );
not ( n56293 , n55932 );
not ( n56294 , n55576 );
or ( n56295 , n56293 , n56294 );
not ( n56296 , n47646 );
not ( n56297 , n55125 );
or ( n56298 , n56296 , n56297 );
nand ( n56299 , n55124 , n47650 );
nand ( n56300 , n56298 , n56299 );
nand ( n56301 , n56300 , n55934 );
nand ( n56302 , n56295 , n56301 );
xor ( n56303 , n56292 , n56302 );
xor ( n56304 , n56267 , n56303 );
xor ( n56305 , n56169 , n56161 );
and ( n56306 , n56305 , n56303 );
and ( n56307 , n56169 , n56161 );
or ( n56308 , n56306 , n56307 );
not ( n56309 , n55972 );
not ( n56310 , n52124 );
not ( n56311 , n56310 );
or ( n56312 , n56309 , n56311 );
not ( n56313 , n51792 );
not ( n56314 , n52130 );
or ( n56315 , n56313 , n56314 );
nand ( n56316 , n52870 , n48829 );
nand ( n56317 , n56315 , n56316 );
nand ( n56318 , n56317 , n51766 );
nand ( n56319 , n56312 , n56318 );
not ( n56320 , n55922 );
not ( n56321 , n55913 );
or ( n56322 , n56320 , n56321 );
not ( n56323 , n48898 );
not ( n56324 , n55917 );
or ( n56325 , n56323 , n56324 );
nand ( n56326 , n53590 , n48897 );
nand ( n56327 , n56325 , n56326 );
nand ( n56328 , n56327 , n54364 );
nand ( n56329 , n56322 , n56328 );
xor ( n56330 , n56319 , n56329 );
not ( n56331 , n55909 );
not ( n56332 , n52853 );
or ( n56333 , n56331 , n56332 );
not ( n56334 , n51204 );
not ( n56335 , n52837 );
or ( n56336 , n56334 , n56335 );
nand ( n56337 , n52840 , n48860 );
nand ( n56338 , n56336 , n56337 );
nand ( n56339 , n52469 , n56338 );
nand ( n56340 , n56333 , n56339 );
xor ( n56341 , n56330 , n56340 );
not ( n56342 , n55950 );
not ( n56343 , n52526 );
or ( n56344 , n56342 , n56343 );
not ( n56345 , n48983 );
not ( n56346 , n53904 );
or ( n56347 , n56345 , n56346 );
not ( n56348 , n48983 );
nand ( n56349 , n50898 , n56348 );
nand ( n56350 , n56347 , n56349 );
nand ( n56351 , n56350 , n51223 );
nand ( n56352 , n56344 , n56351 );
xor ( n56353 , n56217 , n56352 );
not ( n56354 , n55961 );
buf ( n56355 , n51525 );
not ( n56356 , n56355 );
or ( n56357 , n56354 , n56356 );
not ( n56358 , n54611 );
not ( n56359 , n51504 );
or ( n56360 , n56358 , n56359 );
buf ( n56361 , n51503 );
nand ( n56362 , n56361 , n51670 );
nand ( n56363 , n56360 , n56362 );
nand ( n56364 , n51533 , n56363 );
nand ( n56365 , n56357 , n56364 );
xor ( n56366 , n56353 , n56365 );
xor ( n56367 , n56341 , n56366 );
xor ( n56368 , n56367 , n56173 );
xor ( n56369 , n56341 , n56366 );
and ( n56370 , n56369 , n56173 );
and ( n56371 , n56341 , n56366 );
or ( n56372 , n56370 , n56371 );
xor ( n56373 , n56181 , n56177 );
not ( n56374 , n54875 );
not ( n56375 , n51723 );
not ( n56376 , n50654 );
or ( n56377 , n56375 , n56376 );
nand ( n56378 , n51724 , n40691 );
nand ( n56379 , n56377 , n56378 );
not ( n56380 , n56379 );
or ( n56381 , n56374 , n56380 );
nand ( n56382 , n55993 , n52421 );
nand ( n56383 , n56381 , n56382 );
xor ( n56384 , n55805 , n56383 );
xor ( n56385 , n56384 , n56246 );
xor ( n56386 , n56373 , n56385 );
xor ( n56387 , n56181 , n56177 );
and ( n56388 , n56387 , n56385 );
and ( n56389 , n56181 , n56177 );
or ( n56390 , n56388 , n56389 );
not ( n56391 , n52962 );
not ( n56392 , n48645 );
not ( n56393 , n51924 );
or ( n56394 , n56392 , n56393 );
nand ( n56395 , n40734 , n52048 );
nand ( n56396 , n56394 , n56395 );
not ( n56397 , n56396 );
or ( n56398 , n56391 , n56397 );
not ( n56399 , n56053 );
nand ( n56400 , n56399 , n50242 );
nand ( n56401 , n56398 , n56400 );
xor ( n56402 , n55852 , n56401 );
not ( n56403 , n46564 );
not ( n56404 , n56062 );
or ( n56405 , n56403 , n56404 );
not ( n56406 , n48952 );
not ( n56407 , n40452 );
not ( n56408 , n56407 );
or ( n56409 , n56406 , n56408 );
not ( n56410 , n47508 );
not ( n56411 , n40451 );
not ( n56412 , n56411 );
nand ( n56413 , n56410 , n56412 );
nand ( n56414 , n56409 , n56413 );
nand ( n56415 , n56414 , n49832 );
nand ( n56416 , n56405 , n56415 );
xor ( n56417 , n56402 , n56416 );
xor ( n56418 , n56185 , n56417 );
xor ( n56419 , n56418 , n55858 );
xor ( n56420 , n56185 , n56417 );
and ( n56421 , n56420 , n55858 );
and ( n56422 , n56185 , n56417 );
or ( n56423 , n56421 , n56422 );
not ( n56424 , n49252 );
not ( n56425 , n56100 );
or ( n56426 , n56424 , n56425 );
not ( n56427 , n47980 );
not ( n56428 , n54046 );
or ( n56429 , n56427 , n56428 );
nand ( n56430 , n40626 , n47979 );
nand ( n56431 , n56429 , n56430 );
nand ( n56432 , n56431 , n47384 );
nand ( n56433 , n56426 , n56432 );
not ( n56434 , n46267 );
not ( n56435 , n56015 );
or ( n56436 , n56434 , n56435 );
not ( n56437 , n46425 );
not ( n56438 , n40388 );
not ( n56439 , n56438 );
or ( n56440 , n56437 , n56439 );
not ( n56441 , n56438 );
nand ( n56442 , n56441 , n46422 );
nand ( n56443 , n56440 , n56442 );
nand ( n56444 , n49026 , n56443 );
nand ( n56445 , n56436 , n56444 );
xor ( n56446 , n56433 , n56445 );
not ( n56447 , n50659 );
not ( n56448 , n56025 );
or ( n56449 , n56447 , n56448 );
not ( n56450 , n46072 );
not ( n56451 , n40012 );
not ( n56452 , n56451 );
or ( n56453 , n56450 , n56452 );
not ( n56454 , n40011 );
not ( n56455 , n56454 );
nand ( n56456 , n56455 , n46071 );
nand ( n56457 , n56453 , n56456 );
nand ( n56458 , n56457 , n47009 );
nand ( n56459 , n56449 , n56458 );
xor ( n56460 , n56446 , n56459 );
xor ( n56461 , n56262 , n56460 );
not ( n56462 , n51157 );
not ( n56463 , n56078 );
or ( n56464 , n56462 , n56463 );
not ( n56465 , n50263 );
not ( n56466 , n53884 );
or ( n56467 , n56465 , n56466 );
nand ( n56468 , n40364 , n50087 );
nand ( n56469 , n56467 , n56468 );
nand ( n56470 , n56469 , n47827 );
nand ( n56471 , n56464 , n56470 );
not ( n56472 , n47407 );
not ( n56473 , n56089 );
or ( n56474 , n56472 , n56473 );
not ( n56475 , n47803 );
not ( n56476 , n40377 );
not ( n56477 , n56476 );
or ( n56478 , n56475 , n56477 );
nand ( n56479 , n54646 , n50634 );
nand ( n56480 , n56478 , n56479 );
nand ( n56481 , n56480 , n53675 );
nand ( n56482 , n56474 , n56481 );
xor ( n56483 , n56471 , n56482 );
not ( n56484 , n36286 );
not ( n56485 , n34094 );
or ( n56486 , n56484 , n56485 );
nand ( n56487 , n56486 , n37394 );
nand ( n56488 , n32508 , n36293 );
not ( n56489 , n56488 );
not ( n56490 , n56489 );
and ( n56491 , n56487 , n56490 );
not ( n56492 , n56487 );
and ( n56493 , n56492 , n56489 );
nor ( n56494 , n56491 , n56493 );
and ( n56495 , n55843 , n56494 );
not ( n56496 , n55843 );
not ( n56497 , n56494 );
and ( n56498 , n56496 , n56497 );
nor ( n56499 , n56495 , n56498 );
not ( n56500 , n56499 );
not ( n56501 , n56500 );
nor ( n56502 , n56501 , n46441 );
not ( n56503 , n52723 );
not ( n56504 , n53439 );
not ( n56505 , n48997 );
or ( n56506 , n56504 , n56505 );
nand ( n56507 , n41286 , n48967 );
nand ( n56508 , n56506 , n56507 );
not ( n56509 , n56508 );
or ( n56510 , n56503 , n56509 );
nand ( n56511 , n55821 , n53104 );
nand ( n56512 , n56510 , n56511 );
xor ( n56513 , n56502 , n56512 );
not ( n56514 , n55982 );
not ( n56515 , n48894 );
or ( n56516 , n56514 , n56515 );
not ( n56517 , n52377 );
not ( n56518 , n50667 );
or ( n56519 , n56517 , n56518 );
nand ( n56520 , n41036 , n53973 );
nand ( n56521 , n56519 , n56520 );
not ( n56522 , n56521 );
buf ( n56523 , n47483 );
or ( n56524 , n56522 , n56523 );
nand ( n56525 , n56516 , n56524 );
xor ( n56526 , n56513 , n56525 );
xor ( n56527 , n56483 , n56526 );
xor ( n56528 , n56461 , n56527 );
xor ( n56529 , n56262 , n56460 );
and ( n56530 , n56529 , n56527 );
and ( n56531 , n56262 , n56460 );
or ( n56532 , n56530 , n56531 );
xor ( n56533 , n56304 , n55942 );
xor ( n56534 , n56533 , n56368 );
xor ( n56535 , n56304 , n55942 );
and ( n56536 , n56535 , n56368 );
and ( n56537 , n56304 , n55942 );
or ( n56538 , n56536 , n56537 );
xor ( n56539 , n56004 , n56046 );
xor ( n56540 , n56539 , n56111 );
xor ( n56541 , n56004 , n56046 );
and ( n56542 , n56541 , n56111 );
and ( n56543 , n56004 , n56046 );
or ( n56544 , n56542 , n56543 );
xor ( n56545 , n56386 , n56528 );
xor ( n56546 , n56545 , n56419 );
xor ( n56547 , n56386 , n56528 );
and ( n56548 , n56547 , n56419 );
and ( n56549 , n56386 , n56528 );
or ( n56550 , n56548 , n56549 );
xor ( n56551 , n56534 , n56117 );
xor ( n56552 , n56551 , n56123 );
xor ( n56553 , n56534 , n56117 );
and ( n56554 , n56553 , n56123 );
and ( n56555 , n56534 , n56117 );
or ( n56556 , n56554 , n56555 );
xor ( n56557 , n56502 , n56512 );
and ( n56558 , n56557 , n56525 );
and ( n56559 , n56502 , n56512 );
or ( n56560 , n56558 , n56559 );
xor ( n56561 , n56540 , n56129 );
xor ( n56562 , n56561 , n56135 );
xor ( n56563 , n56540 , n56129 );
and ( n56564 , n56563 , n56135 );
and ( n56565 , n56540 , n56129 );
or ( n56566 , n56564 , n56565 );
xor ( n56567 , n56546 , n56552 );
xor ( n56568 , n56567 , n56141 );
xor ( n56569 , n56546 , n56552 );
and ( n56570 , n56569 , n56141 );
and ( n56571 , n56546 , n56552 );
or ( n56572 , n56570 , n56571 );
xor ( n56573 , n56562 , n56568 );
xor ( n56574 , n56573 , n56151 );
xor ( n56575 , n56562 , n56568 );
and ( n56576 , n56575 , n56151 );
and ( n56577 , n56562 , n56568 );
or ( n56578 , n56576 , n56577 );
xor ( n56579 , n56217 , n56352 );
and ( n56580 , n56579 , n56365 );
and ( n56581 , n56217 , n56352 );
or ( n56582 , n56580 , n56581 );
xor ( n56583 , n56319 , n56329 );
and ( n56584 , n56583 , n56340 );
and ( n56585 , n56319 , n56329 );
or ( n56586 , n56584 , n56585 );
xor ( n56587 , n56279 , n56291 );
and ( n56588 , n56587 , n56302 );
and ( n56589 , n56279 , n56291 );
or ( n56590 , n56588 , n56589 );
xor ( n56591 , n55805 , n56383 );
and ( n56592 , n56591 , n56246 );
and ( n56593 , n55805 , n56383 );
or ( n56594 , n56592 , n56593 );
xor ( n56595 , n55852 , n56401 );
and ( n56596 , n56595 , n56416 );
and ( n56597 , n55852 , n56401 );
or ( n56598 , n56596 , n56597 );
xor ( n56599 , n56471 , n56482 );
and ( n56600 , n56599 , n56526 );
and ( n56601 , n56471 , n56482 );
or ( n56602 , n56600 , n56601 );
xor ( n56603 , n56433 , n56445 );
and ( n56604 , n56603 , n56459 );
and ( n56605 , n56433 , n56445 );
or ( n56606 , n56604 , n56605 );
not ( n56607 , n56214 );
not ( n56608 , n52749 );
or ( n56609 , n56607 , n56608 );
and ( n56610 , n54614 , n30929 );
not ( n56611 , n54614 );
and ( n56612 , n56611 , n49220 );
or ( n56613 , n56610 , n56612 );
nand ( n56614 , n56613 , n52757 );
nand ( n56615 , n56609 , n56614 );
not ( n56616 , n49288 );
not ( n56617 , n49232 );
and ( n56618 , n50201 , n56617 );
not ( n56619 , n50201 );
and ( n56620 , n56619 , n41531 );
or ( n56621 , n56618 , n56620 );
not ( n56622 , n56621 );
or ( n56623 , n56616 , n56622 );
nand ( n56624 , n56191 , n51337 );
nand ( n56625 , n56623 , n56624 );
not ( n56626 , n56203 );
not ( n56627 , n49778 );
not ( n56628 , n56627 );
or ( n56629 , n56626 , n56628 );
not ( n56630 , n49618 );
not ( n56631 , n49297 );
or ( n56632 , n56630 , n56631 );
nand ( n56633 , n49298 , n49769 );
nand ( n56634 , n56632 , n56633 );
nand ( n56635 , n56634 , n50575 );
nand ( n56636 , n56629 , n56635 );
xor ( n56637 , n56625 , n56636 );
xor ( n56638 , n56615 , n56637 );
buf ( n56639 , n49737 );
not ( n56640 , n56639 );
not ( n56641 , n48705 );
not ( n56642 , n49190 );
or ( n56643 , n56641 , n56642 );
nand ( n56644 , n41364 , n49094 );
nand ( n56645 , n56643 , n56644 );
not ( n56646 , n56645 );
or ( n56647 , n56640 , n56646 );
nand ( n56648 , n56229 , n49309 );
nand ( n56649 , n56647 , n56648 );
xor ( n56650 , n56638 , n56649 );
xor ( n56651 , n56615 , n56637 );
and ( n56652 , n56651 , n56649 );
and ( n56653 , n56615 , n56637 );
or ( n56654 , n56652 , n56653 );
not ( n56655 , n55872 );
buf ( n56656 , n32516 );
nand ( n56657 , n56656 , n36296 );
not ( n56658 , n56657 );
not ( n56659 , n56658 );
and ( n56660 , n34067 , n32508 );
not ( n56661 , n56660 );
not ( n56662 , n53318 );
or ( n56663 , n56661 , n56662 );
not ( n56664 , n32508 );
not ( n56665 , n33571 );
or ( n56666 , n56664 , n56665 );
nand ( n56667 , n56666 , n36293 );
not ( n56668 , n56667 );
nand ( n56669 , n56663 , n56668 );
not ( n56670 , n56669 );
not ( n56671 , n56670 );
or ( n56672 , n56659 , n56671 );
not ( n56673 , n56660 );
not ( n56674 , n53318 );
or ( n56675 , n56673 , n56674 );
nand ( n56676 , n56675 , n56668 );
nand ( n56677 , n56676 , n56657 );
nand ( n56678 , n56672 , n56677 );
buf ( n56679 , n56678 );
nand ( n56680 , n56655 , n56679 );
buf ( n56681 , n56497 );
and ( n56682 , n56681 , n46440 );
or ( n56683 , n56680 , n56682 );
not ( n56684 , n46440 );
not ( n56685 , n56681 );
nand ( n56686 , n56684 , n56685 , n56679 );
nand ( n56687 , n56683 , n56686 );
not ( n56688 , n54623 );
not ( n56689 , n54625 );
not ( n56690 , n49806 );
or ( n56691 , n56689 , n56690 );
nand ( n56692 , n50827 , n51684 );
nand ( n56693 , n56691 , n56692 );
not ( n56694 , n56693 );
or ( n56695 , n56688 , n56694 );
nand ( n56696 , n56241 , n47873 );
nand ( n56697 , n56695 , n56696 );
xor ( n56698 , n56687 , n56697 );
not ( n56699 , n52723 );
not ( n56700 , n48456 );
not ( n56701 , n41216 );
or ( n56702 , n56700 , n56701 );
nand ( n56703 , n41217 , n52728 );
nand ( n56704 , n56702 , n56703 );
not ( n56705 , n56704 );
or ( n56706 , n56699 , n56705 );
nand ( n56707 , n56508 , n50176 );
nand ( n56708 , n56706 , n56707 );
xor ( n56709 , n56698 , n56708 );
xor ( n56710 , n56687 , n56697 );
and ( n56711 , n56710 , n56708 );
and ( n56712 , n56687 , n56697 );
or ( n56713 , n56711 , n56712 );
not ( n56714 , n52004 );
and ( n56715 , n52377 , n52767 );
not ( n56716 , n52377 );
and ( n56717 , n56716 , n41132 );
or ( n56718 , n56715 , n56717 );
not ( n56719 , n56718 );
or ( n56720 , n56714 , n56719 );
nand ( n56721 , n56521 , n48894 );
nand ( n56722 , n56720 , n56721 );
xor ( n56723 , n56722 , n56221 );
not ( n56724 , n56350 );
not ( n56725 , n50911 );
or ( n56726 , n56724 , n56725 );
buf ( n56727 , n47918 );
not ( n56728 , n56727 );
not ( n56729 , n53904 );
or ( n56730 , n56728 , n56729 );
not ( n56731 , n56727 );
nand ( n56732 , n50898 , n56731 );
nand ( n56733 , n56730 , n56732 );
nand ( n56734 , n56733 , n50922 );
nand ( n56735 , n56726 , n56734 );
xor ( n56736 , n56723 , n56735 );
xor ( n56737 , n56590 , n56736 );
xor ( n56738 , n56737 , n56586 );
xor ( n56739 , n56590 , n56736 );
and ( n56740 , n56739 , n56586 );
and ( n56741 , n56590 , n56736 );
or ( n56742 , n56740 , n56741 );
xor ( n56743 , n56582 , n56594 );
not ( n56744 , n56289 );
not ( n56745 , n56281 );
or ( n56746 , n56744 , n56745 );
and ( n56747 , n46273 , n55876 );
not ( n56748 , n46273 );
not ( n56749 , n55846 );
and ( n56750 , n56748 , n56749 );
or ( n56751 , n56747 , n56750 );
nand ( n56752 , n55459 , n56751 );
nand ( n56753 , n56746 , n56752 );
and ( n56754 , n56669 , n56658 );
not ( n56755 , n56669 );
and ( n56756 , n56755 , n56657 );
nor ( n56757 , n56754 , n56756 );
buf ( n56758 , n56757 );
not ( n56759 , n56758 );
and ( n56760 , n46441 , n56759 );
not ( n56761 , n46441 );
and ( n56762 , n56761 , n56679 );
nor ( n56763 , n56760 , n56762 );
not ( n56764 , n56763 );
not ( n56765 , n56658 );
not ( n56766 , n56670 );
or ( n56767 , n56765 , n56766 );
nand ( n56768 , n56767 , n56677 );
not ( n56769 , n56494 );
and ( n56770 , n56768 , n56769 );
not ( n56771 , n56768 );
not ( n56772 , n56769 );
and ( n56773 , n56771 , n56772 );
nor ( n56774 , n56770 , n56773 );
and ( n56775 , n56774 , n56499 );
buf ( n56776 , n56775 );
buf ( n56777 , n56776 );
not ( n56778 , n56777 );
or ( n56779 , n56764 , n56778 );
buf ( n56780 , n56500 );
not ( n56781 , n50914 );
not ( n56782 , n56759 );
or ( n56783 , n56781 , n56782 );
not ( n56784 , n56768 );
buf ( n56785 , n56784 );
not ( n56786 , n56785 );
nand ( n56787 , n56786 , n48766 );
nand ( n56788 , n56783 , n56787 );
nand ( n56789 , n56780 , n56788 );
nand ( n56790 , n56779 , n56789 );
xor ( n56791 , n56753 , n56790 );
xor ( n56792 , n56791 , n56650 );
xor ( n56793 , n56743 , n56792 );
xor ( n56794 , n56582 , n56594 );
and ( n56795 , n56794 , n56792 );
and ( n56796 , n56582 , n56594 );
or ( n56797 , n56795 , n56796 );
not ( n56798 , n56327 );
not ( n56799 , n53609 );
or ( n56800 , n56798 , n56799 );
not ( n56801 , n47765 );
not ( n56802 , n53590 );
not ( n56803 , n56802 );
or ( n56804 , n56801 , n56803 );
nand ( n56805 , n53590 , n48589 );
nand ( n56806 , n56804 , n56805 );
nand ( n56807 , n56806 , n54364 );
nand ( n56808 , n56800 , n56807 );
not ( n56809 , n56276 );
not ( n56810 , n54314 );
not ( n56811 , n56810 );
or ( n56812 , n56809 , n56811 );
not ( n56813 , n49654 );
not ( n56814 , n54302 );
or ( n56815 , n56813 , n56814 );
nand ( n56816 , n56274 , n47368 );
nand ( n56817 , n56815 , n56816 );
nand ( n56818 , n56817 , n55867 );
nand ( n56819 , n56812 , n56818 );
xor ( n56820 , n56808 , n56819 );
not ( n56821 , n56300 );
not ( n56822 , n55576 );
or ( n56823 , n56821 , n56822 );
not ( n56824 , n49734 );
not ( n56825 , n55119 );
or ( n56826 , n56824 , n56825 );
nand ( n56827 , n55152 , n47821 );
nand ( n56828 , n56826 , n56827 );
nand ( n56829 , n56828 , n54848 );
nand ( n56830 , n56823 , n56829 );
xor ( n56831 , n56820 , n56830 );
not ( n56832 , n56363 );
not ( n56833 , n53543 );
or ( n56834 , n56832 , n56833 );
not ( n56835 , n54185 );
not ( n56836 , n51566 );
or ( n56837 , n56835 , n56836 );
nand ( n56838 , n51505 , n54184 );
nand ( n56839 , n56837 , n56838 );
nand ( n56840 , n51533 , n56839 );
nand ( n56841 , n56834 , n56840 );
not ( n56842 , n56317 );
not ( n56843 , n52125 );
or ( n56844 , n56842 , n56843 );
not ( n56845 , n52033 );
not ( n56846 , n52110 );
or ( n56847 , n56845 , n56846 );
nand ( n56848 , n52870 , n55959 );
nand ( n56849 , n56847 , n56848 );
nand ( n56850 , n56849 , n51766 );
nand ( n56851 , n56844 , n56850 );
xor ( n56852 , n56841 , n56851 );
not ( n56853 , n53182 );
not ( n56854 , n56338 );
or ( n56855 , n56853 , n56854 );
and ( n56856 , n49630 , n52840 );
not ( n56857 , n49630 );
and ( n56858 , n56857 , n53947 );
nor ( n56859 , n56856 , n56858 );
buf ( n56860 , n52850 );
buf ( n56861 , n56860 );
or ( n56862 , n56859 , n56861 );
nand ( n56863 , n56855 , n56862 );
xor ( n56864 , n56852 , n56863 );
xor ( n56865 , n56831 , n56864 );
xor ( n56866 , n56865 , n56598 );
xor ( n56867 , n56831 , n56864 );
and ( n56868 , n56867 , n56598 );
and ( n56869 , n56831 , n56864 );
or ( n56870 , n56868 , n56869 );
xor ( n56871 , n56250 , n56560 );
not ( n56872 , n52962 );
not ( n56873 , n48645 );
not ( n56874 , n52222 );
or ( n56875 , n56873 , n56874 );
nand ( n56876 , n52893 , n52048 );
nand ( n56877 , n56875 , n56876 );
not ( n56878 , n56877 );
or ( n56879 , n56872 , n56878 );
nand ( n56880 , n56396 , n52970 );
nand ( n56881 , n56879 , n56880 );
xor ( n56882 , n56871 , n56881 );
xor ( n56883 , n56602 , n56882 );
xor ( n56884 , n56883 , n56606 );
xor ( n56885 , n56602 , n56882 );
and ( n56886 , n56885 , n56606 );
and ( n56887 , n56602 , n56882 );
or ( n56888 , n56886 , n56887 );
not ( n56889 , n47827 );
not ( n56890 , n50263 );
not ( n56891 , n40148 );
or ( n56892 , n56890 , n56891 );
nand ( n56893 , n56010 , n52080 );
nand ( n56894 , n56892 , n56893 );
not ( n56895 , n56894 );
or ( n56896 , n56889 , n56895 );
nand ( n56897 , n56469 , n48295 );
nand ( n56898 , n56896 , n56897 );
not ( n56899 , n54875 );
not ( n56900 , n51723 );
not ( n56901 , n50958 );
or ( n56902 , n56900 , n56901 );
nand ( n56903 , n52284 , n51724 );
nand ( n56904 , n56902 , n56903 );
not ( n56905 , n56904 );
or ( n56906 , n56899 , n56905 );
nand ( n56907 , n56379 , n52421 );
nand ( n56908 , n56906 , n56907 );
xor ( n56909 , n56898 , n56908 );
not ( n56910 , n53675 );
not ( n56911 , n47803 );
not ( n56912 , n40225 );
or ( n56913 , n56911 , n56912 );
nand ( n56914 , n53660 , n48727 );
nand ( n56915 , n56913 , n56914 );
not ( n56916 , n56915 );
or ( n56917 , n56910 , n56916 );
nand ( n56918 , n56480 , n47407 );
nand ( n56919 , n56917 , n56918 );
xor ( n56920 , n56909 , n56919 );
not ( n56921 , n53510 );
not ( n56922 , n49500 );
not ( n56923 , n53718 );
or ( n56924 , n56922 , n56923 );
nand ( n56925 , n40635 , n47979 );
nand ( n56926 , n56924 , n56925 );
not ( n56927 , n56926 );
or ( n56928 , n56921 , n56927 );
nand ( n56929 , n56431 , n49252 );
nand ( n56930 , n56928 , n56929 );
not ( n56931 , n49026 );
not ( n56932 , n46425 );
not ( n56933 , n56058 );
or ( n56934 , n56932 , n56933 );
nand ( n56935 , n55203 , n46422 );
nand ( n56936 , n56934 , n56935 );
not ( n56937 , n56936 );
or ( n56938 , n56931 , n56937 );
nand ( n56939 , n56443 , n46267 );
nand ( n56940 , n56938 , n56939 );
xor ( n56941 , n56930 , n56940 );
not ( n56942 , n51865 );
not ( n56943 , n52267 );
not ( n56944 , n52211 );
or ( n56945 , n56943 , n56944 );
nand ( n56946 , n40592 , n51351 );
nand ( n56947 , n56945 , n56946 );
not ( n56948 , n56947 );
or ( n56949 , n56942 , n56948 );
nand ( n56950 , n56258 , n49713 );
nand ( n56951 , n56949 , n56950 );
xor ( n56952 , n56941 , n56951 );
xor ( n56953 , n56920 , n56952 );
xor ( n56954 , n56953 , n56266 );
xor ( n56955 , n56920 , n56952 );
and ( n56956 , n56955 , n56266 );
and ( n56957 , n56920 , n56952 );
or ( n56958 , n56956 , n56957 );
not ( n56959 , n50659 );
not ( n56960 , n56457 );
or ( n56961 , n56959 , n56960 );
not ( n56962 , n39962 );
and ( n56963 , n56962 , n46071 );
not ( n56964 , n56962 );
and ( n56965 , n56964 , n46072 );
nor ( n56966 , n56963 , n56965 );
nand ( n56967 , n56966 , n46602 );
nand ( n56968 , n56961 , n56967 );
not ( n56969 , n46564 );
not ( n56970 , n56414 );
or ( n56971 , n56969 , n56970 );
not ( n56972 , n48952 );
not ( n56973 , n56020 );
or ( n56974 , n56972 , n56973 );
not ( n56975 , n40512 );
not ( n56976 , n56975 );
nand ( n56977 , n56976 , n52990 );
nand ( n56978 , n56974 , n56977 );
nand ( n56979 , n56978 , n49832 );
nand ( n56980 , n56971 , n56979 );
xor ( n56981 , n56968 , n56980 );
xor ( n56982 , n56981 , n56709 );
xor ( n56983 , n56982 , n56308 );
xor ( n56984 , n56983 , n56738 );
xor ( n56985 , n56982 , n56308 );
and ( n56986 , n56985 , n56738 );
and ( n56987 , n56982 , n56308 );
or ( n56988 , n56986 , n56987 );
xor ( n56989 , n56372 , n56390 );
xor ( n56990 , n56989 , n56866 );
xor ( n56991 , n56372 , n56390 );
and ( n56992 , n56991 , n56866 );
and ( n56993 , n56372 , n56390 );
or ( n56994 , n56992 , n56993 );
xor ( n56995 , n56793 , n56423 );
xor ( n56996 , n56995 , n56532 );
xor ( n56997 , n56793 , n56423 );
and ( n56998 , n56997 , n56532 );
and ( n56999 , n56793 , n56423 );
or ( n57000 , n56998 , n56999 );
xor ( n57001 , n56884 , n56954 );
xor ( n57002 , n57001 , n56538 );
xor ( n57003 , n56884 , n56954 );
and ( n57004 , n57003 , n56538 );
and ( n57005 , n56884 , n56954 );
or ( n57006 , n57004 , n57005 );
xor ( n57007 , n56984 , n56990 );
xor ( n57008 , n57007 , n56544 );
xor ( n57009 , n56984 , n56990 );
and ( n57010 , n57009 , n56544 );
and ( n57011 , n56984 , n56990 );
or ( n57012 , n57010 , n57011 );
xor ( n57013 , n56722 , n56221 );
and ( n57014 , n57013 , n56735 );
and ( n57015 , n56722 , n56221 );
or ( n57016 , n57014 , n57015 );
xor ( n57017 , n56550 , n56996 );
xor ( n57018 , n57017 , n57002 );
xor ( n57019 , n56550 , n56996 );
and ( n57020 , n57019 , n57002 );
and ( n57021 , n56550 , n56996 );
or ( n57022 , n57020 , n57021 );
xor ( n57023 , n56556 , n57008 );
xor ( n57024 , n57023 , n56566 );
xor ( n57025 , n56556 , n57008 );
and ( n57026 , n57025 , n56566 );
and ( n57027 , n56556 , n57008 );
or ( n57028 , n57026 , n57027 );
xor ( n57029 , n57018 , n56572 );
xor ( n57030 , n57029 , n57024 );
xor ( n57031 , n57018 , n56572 );
and ( n57032 , n57031 , n57024 );
and ( n57033 , n57018 , n56572 );
or ( n57034 , n57032 , n57033 );
xor ( n57035 , n56841 , n56851 );
and ( n57036 , n57035 , n56863 );
and ( n57037 , n56841 , n56851 );
or ( n57038 , n57036 , n57037 );
xor ( n57039 , n56808 , n56819 );
and ( n57040 , n57039 , n56830 );
and ( n57041 , n56808 , n56819 );
or ( n57042 , n57040 , n57041 );
xor ( n57043 , n56753 , n56790 );
and ( n57044 , n57043 , n56650 );
and ( n57045 , n56753 , n56790 );
or ( n57046 , n57044 , n57045 );
xor ( n57047 , n56250 , n56560 );
and ( n57048 , n57047 , n56881 );
and ( n57049 , n56250 , n56560 );
or ( n57050 , n57048 , n57049 );
xor ( n57051 , n56898 , n56908 );
and ( n57052 , n57051 , n56919 );
and ( n57053 , n56898 , n56908 );
or ( n57054 , n57052 , n57053 );
xor ( n57055 , n56968 , n56980 );
and ( n57056 , n57055 , n56709 );
and ( n57057 , n56968 , n56980 );
or ( n57058 , n57056 , n57057 );
xor ( n57059 , n56930 , n56940 );
and ( n57060 , n57059 , n56951 );
and ( n57061 , n56930 , n56940 );
or ( n57062 , n57060 , n57061 );
not ( n57063 , n56634 );
not ( n57064 , n49779 );
or ( n57065 , n57063 , n57064 );
not ( n57066 , n49770 );
not ( n57067 , n49029 );
or ( n57068 , n57066 , n57067 );
nand ( n57069 , n41668 , n50292 );
nand ( n57070 , n57068 , n57069 );
nand ( n57071 , n57070 , n51809 );
nand ( n57072 , n57065 , n57071 );
not ( n57073 , n56613 );
not ( n57074 , n50321 );
or ( n57075 , n57073 , n57074 );
not ( n57076 , n52379 );
not ( n57077 , n50301 );
or ( n57078 , n57076 , n57077 );
or ( n57079 , n52379 , n50163 );
nand ( n57080 , n57078 , n57079 );
nand ( n57081 , n57080 , n51452 );
nand ( n57082 , n57075 , n57081 );
xor ( n57083 , n57072 , n57082 );
not ( n57084 , n52191 );
not ( n57085 , n49452 );
not ( n57086 , n48951 );
or ( n57087 , n57085 , n57086 );
not ( n57088 , n49112 );
nand ( n57089 , n48486 , n57088 );
nand ( n57090 , n57087 , n57089 );
not ( n57091 , n57090 );
or ( n57092 , n57084 , n57091 );
nand ( n57093 , n56621 , n49276 );
nand ( n57094 , n57092 , n57093 );
xor ( n57095 , n57083 , n57094 );
xor ( n57096 , n57072 , n57082 );
and ( n57097 , n57096 , n57094 );
and ( n57098 , n57072 , n57082 );
or ( n57099 , n57097 , n57098 );
not ( n57100 , n56203 );
not ( n57101 , n56627 );
or ( n57102 , n57100 , n57101 );
nand ( n57103 , n57102 , n56635 );
and ( n57104 , n56625 , n57103 );
not ( n57105 , n49737 );
and ( n57106 , n48705 , n48997 );
not ( n57107 , n48705 );
and ( n57108 , n57107 , n48996 );
or ( n57109 , n57106 , n57108 );
not ( n57110 , n57109 );
or ( n57111 , n57105 , n57110 );
not ( n57112 , n48756 );
nand ( n57113 , n57112 , n56645 );
nand ( n57114 , n57111 , n57113 );
xor ( n57115 , n57104 , n57114 );
not ( n57116 , n56757 );
not ( n57117 , n36380 );
not ( n57118 , n57117 );
not ( n57119 , n34094 );
nor ( n57120 , n57119 , n37530 );
not ( n57121 , n57120 );
or ( n57122 , n57118 , n57121 );
and ( n57123 , n36347 , n37596 );
nor ( n57124 , n57123 , n36297 );
nand ( n57125 , n57122 , n57124 );
nand ( n57126 , n37548 , n32690 );
not ( n57127 , n57126 );
not ( n57128 , n57127 );
and ( n57129 , n57125 , n57128 );
not ( n57130 , n57125 );
and ( n57131 , n57130 , n57127 );
nor ( n57132 , n57129 , n57131 );
and ( n57133 , n57116 , n57132 );
not ( n57134 , n57116 );
not ( n57135 , n57132 );
and ( n57136 , n57134 , n57135 );
nor ( n57137 , n57133 , n57136 );
not ( n57138 , n57137 );
not ( n57139 , n57138 );
and ( n57140 , n57139 , n48689 );
xor ( n57141 , n57115 , n57140 );
xor ( n57142 , n57104 , n57114 );
and ( n57143 , n57142 , n57140 );
and ( n57144 , n57104 , n57114 );
or ( n57145 , n57143 , n57144 );
not ( n57146 , n44004 );
not ( n57147 , n46072 );
not ( n57148 , n39844 );
or ( n57149 , n57147 , n57148 );
nand ( n57150 , n39845 , n46071 );
nand ( n57151 , n57149 , n57150 );
not ( n57152 , n57151 );
or ( n57153 , n57146 , n57152 );
nand ( n57154 , n56966 , n50659 );
nand ( n57155 , n57153 , n57154 );
xor ( n57156 , n57155 , n57042 );
not ( n57157 , n54623 );
not ( n57158 , n54625 );
not ( n57159 , n50020 );
or ( n57160 , n57158 , n57159 );
nand ( n57161 , n41038 , n55023 );
nand ( n57162 , n57160 , n57161 );
not ( n57163 , n57162 );
or ( n57164 , n57157 , n57163 );
nand ( n57165 , n56693 , n52022 );
nand ( n57166 , n57164 , n57165 );
not ( n57167 , n53104 );
not ( n57168 , n56704 );
or ( n57169 , n57167 , n57168 );
not ( n57170 , n48456 );
not ( n57171 , n50007 );
or ( n57172 , n57170 , n57171 );
not ( n57173 , n48971 );
nand ( n57174 , n40854 , n57173 );
nand ( n57175 , n57172 , n57174 );
nand ( n57176 , n57175 , n52723 );
nand ( n57177 , n57169 , n57176 );
xor ( n57178 , n57166 , n57177 );
not ( n57179 , n56733 );
not ( n57180 , n50911 );
or ( n57181 , n57179 , n57180 );
not ( n57182 , n47332 );
not ( n57183 , n57182 );
not ( n57184 , n52781 );
or ( n57185 , n57183 , n57184 );
not ( n57186 , n57182 );
not ( n57187 , n50946 );
nand ( n57188 , n57186 , n57187 );
nand ( n57189 , n57185 , n57188 );
nand ( n57190 , n57189 , n50922 );
nand ( n57191 , n57181 , n57190 );
xor ( n57192 , n57178 , n57191 );
xor ( n57193 , n57156 , n57192 );
xor ( n57194 , n57155 , n57042 );
and ( n57195 , n57194 , n57192 );
and ( n57196 , n57155 , n57042 );
or ( n57197 , n57195 , n57196 );
xor ( n57198 , n57016 , n57038 );
xor ( n57199 , n57198 , n57046 );
xor ( n57200 , n57016 , n57038 );
and ( n57201 , n57200 , n57046 );
and ( n57202 , n57016 , n57038 );
or ( n57203 , n57201 , n57202 );
not ( n57204 , n56751 );
not ( n57205 , n56281 );
or ( n57206 , n57204 , n57205 );
not ( n57207 , n47646 );
not ( n57208 , n55893 );
or ( n57209 , n57207 , n57208 );
nand ( n57210 , n55892 , n47650 );
nand ( n57211 , n57209 , n57210 );
nand ( n57212 , n57211 , n55459 );
nand ( n57213 , n57206 , n57212 );
xor ( n57214 , n57213 , n57095 );
not ( n57215 , n56788 );
not ( n57216 , n56777 );
or ( n57217 , n57215 , n57216 );
not ( n57218 , n46037 );
not ( n57219 , n56785 );
or ( n57220 , n57218 , n57219 );
nand ( n57221 , n56758 , n47306 );
nand ( n57222 , n57220 , n57221 );
nand ( n57223 , n56780 , n57222 );
nand ( n57224 , n57217 , n57223 );
xor ( n57225 , n57214 , n57224 );
not ( n57226 , n56839 );
not ( n57227 , n53170 );
or ( n57228 , n57226 , n57227 );
not ( n57229 , n48983 );
not ( n57230 , n51504 );
or ( n57231 , n57229 , n57230 );
nand ( n57232 , n51505 , n56348 );
nand ( n57233 , n57231 , n57232 );
nand ( n57234 , n55066 , n57233 );
nand ( n57235 , n57228 , n57234 );
not ( n57236 , n56849 );
not ( n57237 , n54266 );
or ( n57238 , n57236 , n57237 );
not ( n57239 , n54611 );
not ( n57240 , n52130 );
or ( n57241 , n57239 , n57240 );
nand ( n57242 , n53918 , n51670 );
nand ( n57243 , n57241 , n57242 );
nand ( n57244 , n57243 , n51766 );
nand ( n57245 , n57238 , n57244 );
xor ( n57246 , n57235 , n57245 );
not ( n57247 , n56859 );
not ( n57248 , n57247 );
not ( n57249 , n52854 );
or ( n57250 , n57248 , n57249 );
not ( n57251 , n51792 );
not ( n57252 , n52836 );
buf ( n57253 , n57252 );
not ( n57254 , n57253 );
or ( n57255 , n57251 , n57254 );
nand ( n57256 , n55481 , n48829 );
nand ( n57257 , n57255 , n57256 );
nand ( n57258 , n52469 , n57257 );
nand ( n57259 , n57250 , n57258 );
xor ( n57260 , n57246 , n57259 );
xor ( n57261 , n57225 , n57260 );
not ( n57262 , n56806 );
not ( n57263 , n53609 );
or ( n57264 , n57262 , n57263 );
not ( n57265 , n51204 );
not ( n57266 , n55917 );
or ( n57267 , n57265 , n57266 );
nand ( n57268 , n53590 , n48860 );
nand ( n57269 , n57267 , n57268 );
nand ( n57270 , n57269 , n53326 );
nand ( n57271 , n57264 , n57270 );
not ( n57272 , n56817 );
not ( n57273 , n56810 );
or ( n57274 , n57272 , n57273 );
not ( n57275 , n48898 );
not ( n57276 , n55276 );
or ( n57277 , n57275 , n57276 );
nand ( n57278 , n54297 , n48897 );
nand ( n57279 , n57277 , n57278 );
nand ( n57280 , n57279 , n54077 );
nand ( n57281 , n57274 , n57280 );
xor ( n57282 , n57271 , n57281 );
not ( n57283 , n56828 );
not ( n57284 , n55144 );
or ( n57285 , n57283 , n57284 );
not ( n57286 , n47227 );
not ( n57287 , n55119 );
or ( n57288 , n57286 , n57287 );
nand ( n57289 , n55123 , n47589 );
nand ( n57290 , n57288 , n57289 );
nand ( n57291 , n55934 , n57290 );
nand ( n57292 , n57285 , n57291 );
xor ( n57293 , n57282 , n57292 );
xor ( n57294 , n57261 , n57293 );
xor ( n57295 , n57225 , n57260 );
and ( n57296 , n57295 , n57293 );
and ( n57297 , n57225 , n57260 );
or ( n57298 , n57296 , n57297 );
xor ( n57299 , n57050 , n57062 );
xor ( n57300 , n57299 , n57058 );
xor ( n57301 , n57050 , n57062 );
and ( n57302 , n57301 , n57058 );
and ( n57303 , n57050 , n57062 );
or ( n57304 , n57302 , n57303 );
not ( n57305 , n52004 );
not ( n57306 , n52377 );
not ( n57307 , n40691 );
not ( n57308 , n57307 );
or ( n57309 , n57306 , n57308 );
nand ( n57310 , n40691 , n53973 );
nand ( n57311 , n57309 , n57310 );
not ( n57312 , n57311 );
or ( n57313 , n57305 , n57312 );
not ( n57314 , n56515 );
nand ( n57315 , n56718 , n57314 );
nand ( n57316 , n57313 , n57315 );
xor ( n57317 , n57316 , n56654 );
xor ( n57318 , n57317 , n56713 );
xor ( n57319 , n57318 , n57054 );
not ( n57320 , n52970 );
not ( n57321 , n56877 );
or ( n57322 , n57320 , n57321 );
and ( n57323 , n48645 , n51916 );
not ( n57324 , n48645 );
and ( n57325 , n57324 , n51913 );
nor ( n57326 , n57323 , n57325 );
nand ( n57327 , n57326 , n52043 );
nand ( n57328 , n57322 , n57327 );
not ( n57329 , n54875 );
and ( n57330 , n51723 , n54032 );
not ( n57331 , n51723 );
not ( n57332 , n51928 );
not ( n57333 , n57332 );
and ( n57334 , n57331 , n57333 );
nor ( n57335 , n57330 , n57334 );
not ( n57336 , n57335 );
or ( n57337 , n57329 , n57336 );
nand ( n57338 , n56904 , n52421 );
nand ( n57339 , n57337 , n57338 );
xor ( n57340 , n57328 , n57339 );
not ( n57341 , n47407 );
not ( n57342 , n56915 );
or ( n57343 , n57341 , n57342 );
not ( n57344 , n51545 );
not ( n57345 , n54811 );
or ( n57346 , n57344 , n57345 );
nand ( n57347 , n40364 , n48727 );
nand ( n57348 , n57346 , n57347 );
nand ( n57349 , n57348 , n53675 );
nand ( n57350 , n57343 , n57349 );
xor ( n57351 , n57340 , n57350 );
xor ( n57352 , n57319 , n57351 );
xor ( n57353 , n57318 , n57054 );
and ( n57354 , n57353 , n57351 );
and ( n57355 , n57318 , n57054 );
or ( n57356 , n57354 , n57355 );
not ( n57357 , n46267 );
not ( n57358 , n56936 );
or ( n57359 , n57357 , n57358 );
not ( n57360 , n46425 );
not ( n57361 , n55630 );
or ( n57362 , n57360 , n57361 );
nand ( n57363 , n56412 , n46422 );
nand ( n57364 , n57362 , n57363 );
nand ( n57365 , n57364 , n49026 );
nand ( n57366 , n57359 , n57365 );
xor ( n57367 , n57141 , n57366 );
not ( n57368 , n49713 );
not ( n57369 , n56947 );
or ( n57370 , n57368 , n57369 );
not ( n57371 , n52267 );
not ( n57372 , n53271 );
or ( n57373 , n57371 , n57372 );
nand ( n57374 , n40626 , n51351 );
nand ( n57375 , n57373 , n57374 );
nand ( n57376 , n57375 , n51865 );
nand ( n57377 , n57370 , n57376 );
xor ( n57378 , n57367 , n57377 );
xor ( n57379 , n57378 , n56742 );
not ( n57380 , n49832 );
nand ( n57381 , n56455 , n47514 );
nand ( n57382 , n47508 , n56454 );
nand ( n57383 , n57381 , n57382 );
not ( n57384 , n57383 );
or ( n57385 , n57380 , n57384 );
nand ( n57386 , n56978 , n46564 );
nand ( n57387 , n57385 , n57386 );
not ( n57388 , n47827 );
not ( n57389 , n50263 );
not ( n57390 , n54791 );
not ( n57391 , n57390 );
or ( n57392 , n57389 , n57391 );
nand ( n57393 , n40389 , n50087 );
nand ( n57394 , n57392 , n57393 );
not ( n57395 , n57394 );
or ( n57396 , n57388 , n57395 );
nand ( n57397 , n56894 , n46776 );
nand ( n57398 , n57396 , n57397 );
xor ( n57399 , n57387 , n57398 );
not ( n57400 , n49500 );
not ( n57401 , n54020 );
or ( n57402 , n57400 , n57401 );
nand ( n57403 , n40377 , n53997 );
nand ( n57404 , n57402 , n57403 );
not ( n57405 , n57404 );
not ( n57406 , n53510 );
or ( n57407 , n57405 , n57406 );
not ( n57408 , n56926 );
or ( n57409 , n57408 , n48988 );
nand ( n57410 , n57407 , n57409 );
xor ( n57411 , n57399 , n57410 );
xor ( n57412 , n57379 , n57411 );
xor ( n57413 , n57378 , n56742 );
and ( n57414 , n57413 , n57411 );
and ( n57415 , n57378 , n56742 );
or ( n57416 , n57414 , n57415 );
xor ( n57417 , n57193 , n57199 );
xor ( n57418 , n57417 , n56797 );
xor ( n57419 , n57193 , n57199 );
and ( n57420 , n57419 , n56797 );
and ( n57421 , n57193 , n57199 );
or ( n57422 , n57420 , n57421 );
xor ( n57423 , n57294 , n56870 );
xor ( n57424 , n57423 , n56888 );
xor ( n57425 , n57294 , n56870 );
and ( n57426 , n57425 , n56888 );
and ( n57427 , n57294 , n56870 );
or ( n57428 , n57426 , n57427 );
xor ( n57429 , n57300 , n56958 );
xor ( n57430 , n57429 , n57352 );
xor ( n57431 , n57300 , n56958 );
and ( n57432 , n57431 , n57352 );
and ( n57433 , n57300 , n56958 );
or ( n57434 , n57432 , n57433 );
xor ( n57435 , n57412 , n56988 );
xor ( n57436 , n57435 , n57418 );
xor ( n57437 , n57412 , n56988 );
and ( n57438 , n57437 , n57418 );
and ( n57439 , n57412 , n56988 );
or ( n57440 , n57438 , n57439 );
xor ( n57441 , n57166 , n57177 );
and ( n57442 , n57441 , n57191 );
and ( n57443 , n57166 , n57177 );
or ( n57444 , n57442 , n57443 );
xor ( n57445 , n56994 , n57424 );
xor ( n57446 , n57445 , n57000 );
xor ( n57447 , n56994 , n57424 );
and ( n57448 , n57447 , n57000 );
and ( n57449 , n56994 , n57424 );
or ( n57450 , n57448 , n57449 );
xor ( n57451 , n57430 , n57436 );
xor ( n57452 , n57451 , n57006 );
xor ( n57453 , n57430 , n57436 );
and ( n57454 , n57453 , n57006 );
and ( n57455 , n57430 , n57436 );
or ( n57456 , n57454 , n57455 );
xor ( n57457 , n57012 , n57446 );
xor ( n57458 , n57457 , n57022 );
xor ( n57459 , n57012 , n57446 );
and ( n57460 , n57459 , n57022 );
and ( n57461 , n57012 , n57446 );
or ( n57462 , n57460 , n57461 );
xor ( n57463 , n57452 , n57458 );
xor ( n57464 , n57463 , n57028 );
xor ( n57465 , n57452 , n57458 );
and ( n57466 , n57465 , n57028 );
and ( n57467 , n57452 , n57458 );
or ( n57468 , n57466 , n57467 );
xor ( n57469 , n57235 , n57245 );
and ( n57470 , n57469 , n57259 );
and ( n57471 , n57235 , n57245 );
or ( n57472 , n57470 , n57471 );
xor ( n57473 , n57271 , n57281 );
and ( n57474 , n57473 , n57292 );
and ( n57475 , n57271 , n57281 );
or ( n57476 , n57474 , n57475 );
xor ( n57477 , n57213 , n57095 );
and ( n57478 , n57477 , n57224 );
and ( n57479 , n57213 , n57095 );
or ( n57480 , n57478 , n57479 );
xor ( n57481 , n57316 , n56654 );
and ( n57482 , n57481 , n56713 );
and ( n57483 , n57316 , n56654 );
or ( n57484 , n57482 , n57483 );
xor ( n57485 , n57328 , n57339 );
and ( n57486 , n57485 , n57350 );
and ( n57487 , n57328 , n57339 );
or ( n57488 , n57486 , n57487 );
xor ( n57489 , n57387 , n57398 );
and ( n57490 , n57489 , n57410 );
and ( n57491 , n57387 , n57398 );
or ( n57492 , n57490 , n57491 );
xor ( n57493 , n57141 , n57366 );
and ( n57494 , n57493 , n57377 );
and ( n57495 , n57141 , n57366 );
or ( n57496 , n57494 , n57495 );
not ( n57497 , n52723 );
not ( n57498 , n48456 );
not ( n57499 , n49809 );
or ( n57500 , n57498 , n57499 );
nand ( n57501 , n52916 , n57173 );
nand ( n57502 , n57500 , n57501 );
not ( n57503 , n57502 );
or ( n57504 , n57497 , n57503 );
nand ( n57505 , n57175 , n50176 );
nand ( n57506 , n57504 , n57505 );
and ( n57507 , n57125 , n57127 );
not ( n57508 , n57125 );
and ( n57509 , n57508 , n57126 );
nor ( n57510 , n57507 , n57509 );
not ( n57511 , n57510 );
nand ( n57512 , n57511 , n46441 );
not ( n57513 , n46440 );
not ( n57514 , n57510 );
or ( n57515 , n57513 , n57514 );
nand ( n57516 , n57515 , n56785 );
and ( n57517 , n57512 , n57516 );
not ( n57518 , n37531 );
not ( n57519 , n34069 );
or ( n57520 , n57518 , n57519 );
and ( n57521 , n37532 , n51754 );
nor ( n57522 , n57521 , n37549 );
nand ( n57523 , n57520 , n57522 );
not ( n57524 , n36303 );
nand ( n57525 , n57524 , n32772 );
not ( n57526 , n57525 );
and ( n57527 , n57523 , n57526 );
not ( n57528 , n57523 );
and ( n57529 , n57528 , n57525 );
nor ( n57530 , n57527 , n57529 );
not ( n57531 , n57530 );
not ( n57532 , n57531 );
buf ( n57533 , n57532 );
not ( n57534 , n57533 );
nor ( n57535 , n57517 , n57534 );
xor ( n57536 , n57506 , n57535 );
not ( n57537 , n57080 );
not ( n57538 , n50321 );
or ( n57539 , n57537 , n57538 );
not ( n57540 , n50163 );
not ( n57541 , n57540 );
not ( n57542 , n49297 );
or ( n57543 , n57541 , n57542 );
nand ( n57544 , n49298 , n50163 );
nand ( n57545 , n57543 , n57544 );
nand ( n57546 , n57545 , n50331 );
nand ( n57547 , n57539 , n57546 );
not ( n57548 , n57070 );
not ( n57549 , n52057 );
or ( n57550 , n57548 , n57549 );
not ( n57551 , n48306 );
not ( n57552 , n50292 );
and ( n57553 , n57551 , n57552 );
not ( n57554 , n54210 );
and ( n57555 , n57554 , n49769 );
nor ( n57556 , n57553 , n57555 );
not ( n57557 , n57556 );
nand ( n57558 , n57557 , n50575 );
nand ( n57559 , n57550 , n57558 );
xor ( n57560 , n57547 , n57559 );
xor ( n57561 , n57536 , n57560 );
xor ( n57562 , n57506 , n57535 );
and ( n57563 , n57562 , n57560 );
and ( n57564 , n57506 , n57535 );
or ( n57565 , n57563 , n57564 );
not ( n57566 , n49309 );
not ( n57567 , n57109 );
or ( n57568 , n57566 , n57567 );
and ( n57569 , n56227 , n41216 );
not ( n57570 , n56227 );
not ( n57571 , n41216 );
and ( n57572 , n57570 , n57571 );
or ( n57573 , n57569 , n57572 );
not ( n57574 , n57573 );
nand ( n57575 , n57574 , n56639 );
nand ( n57576 , n57568 , n57575 );
not ( n57577 , n49288 );
not ( n57578 , n49112 );
not ( n57579 , n49820 );
or ( n57580 , n57578 , n57579 );
nand ( n57581 , n52272 , n57088 );
nand ( n57582 , n57580 , n57581 );
not ( n57583 , n57582 );
or ( n57584 , n57577 , n57583 );
buf ( n57585 , n49275 );
not ( n57586 , n57585 );
nand ( n57587 , n57090 , n57586 );
nand ( n57588 , n57584 , n57587 );
xor ( n57589 , n57576 , n57588 );
not ( n57590 , n54623 );
not ( n57591 , n54625 );
not ( n57592 , n50400 );
or ( n57593 , n57591 , n57592 );
nand ( n57594 , n50404 , n51684 );
nand ( n57595 , n57593 , n57594 );
not ( n57596 , n57595 );
or ( n57597 , n57590 , n57596 );
nand ( n57598 , n57162 , n47873 );
nand ( n57599 , n57597 , n57598 );
xor ( n57600 , n57589 , n57599 );
xor ( n57601 , n57576 , n57588 );
and ( n57602 , n57601 , n57599 );
and ( n57603 , n57576 , n57588 );
or ( n57604 , n57602 , n57603 );
xor ( n57605 , n57476 , n57480 );
xor ( n57606 , n57605 , n57444 );
xor ( n57607 , n57476 , n57480 );
and ( n57608 , n57607 , n57444 );
and ( n57609 , n57476 , n57480 );
or ( n57610 , n57608 , n57609 );
xor ( n57611 , n57472 , n57484 );
not ( n57612 , n46440 );
buf ( n57613 , n57530 );
buf ( n57614 , n57613 );
not ( n57615 , n57614 );
not ( n57616 , n57615 );
or ( n57617 , n57612 , n57616 );
not ( n57618 , n48689 );
buf ( n57619 , n57613 );
nand ( n57620 , n57618 , n57619 );
nand ( n57621 , n57617 , n57620 );
not ( n57622 , n57621 );
and ( n57623 , n57613 , n57510 );
not ( n57624 , n57613 );
and ( n57625 , n57624 , n57511 );
nor ( n57626 , n57623 , n57625 );
nand ( n57627 , n57138 , n57626 );
not ( n57628 , n57627 );
not ( n57629 , n57628 );
or ( n57630 , n57622 , n57629 );
buf ( n57631 , n57139 );
not ( n57632 , n45767 );
buf ( n57633 , n57531 );
not ( n57634 , n57633 );
not ( n57635 , n57634 );
or ( n57636 , n57632 , n57635 );
not ( n57637 , n57619 );
nand ( n57638 , n57637 , n50914 );
nand ( n57639 , n57636 , n57638 );
nand ( n57640 , n57631 , n57639 );
nand ( n57641 , n57630 , n57640 );
xor ( n57642 , n57641 , n57099 );
xor ( n57643 , n57642 , n57145 );
xor ( n57644 , n57611 , n57643 );
xor ( n57645 , n57472 , n57484 );
and ( n57646 , n57645 , n57643 );
and ( n57647 , n57472 , n57484 );
or ( n57648 , n57646 , n57647 );
not ( n57649 , n57290 );
not ( n57650 , n55143 );
or ( n57651 , n57649 , n57650 );
not ( n57652 , n52165 );
not ( n57653 , n55148 );
or ( n57654 , n57652 , n57653 );
not ( n57655 , n55119 );
nand ( n57656 , n57655 , n47368 );
nand ( n57657 , n57654 , n57656 );
nand ( n57658 , n57657 , n55155 );
nand ( n57659 , n57651 , n57658 );
not ( n57660 , n57222 );
not ( n57661 , n56776 );
or ( n57662 , n57660 , n57661 );
not ( n57663 , n46273 );
not ( n57664 , n56784 );
not ( n57665 , n57664 );
not ( n57666 , n57665 );
or ( n57667 , n57663 , n57666 );
nand ( n57668 , n56758 , n46824 );
nand ( n57669 , n57667 , n57668 );
nand ( n57670 , n56780 , n57669 );
nand ( n57671 , n57662 , n57670 );
xor ( n57672 , n57659 , n57671 );
not ( n57673 , n57211 );
not ( n57674 , n55887 );
or ( n57675 , n57673 , n57674 );
not ( n57676 , n55845 );
and ( n57677 , n47821 , n57676 );
not ( n57678 , n47821 );
and ( n57679 , n57678 , n55845 );
or ( n57680 , n57677 , n57679 );
not ( n57681 , n57680 );
nand ( n57682 , n57681 , n55459 );
nand ( n57683 , n57675 , n57682 );
xor ( n57684 , n57672 , n57683 );
not ( n57685 , n57257 );
not ( n57686 , n52853 );
or ( n57687 , n57685 , n57686 );
not ( n57688 , n52033 );
not ( n57689 , n57253 );
or ( n57690 , n57688 , n57689 );
nand ( n57691 , n55481 , n52038 );
nand ( n57692 , n57690 , n57691 );
nand ( n57693 , n57692 , n53571 );
nand ( n57694 , n57687 , n57693 );
not ( n57695 , n57269 );
not ( n57696 , n55913 );
or ( n57697 , n57695 , n57696 );
not ( n57698 , n49624 );
not ( n57699 , n55918 );
or ( n57700 , n57698 , n57699 );
nand ( n57701 , n53590 , n49630 );
nand ( n57702 , n57700 , n57701 );
nand ( n57703 , n57702 , n53619 );
nand ( n57704 , n57697 , n57703 );
xor ( n57705 , n57694 , n57704 );
not ( n57706 , n57279 );
not ( n57707 , n56810 );
or ( n57708 , n57706 , n57707 );
and ( n57709 , n54297 , n48589 );
not ( n57710 , n54297 );
and ( n57711 , n57710 , n47765 );
nor ( n57712 , n57709 , n57711 );
not ( n57713 , n57712 );
nand ( n57714 , n57713 , n54077 );
nand ( n57715 , n57708 , n57714 );
xor ( n57716 , n57705 , n57715 );
xor ( n57717 , n57684 , n57716 );
not ( n57718 , n57189 );
not ( n57719 , n50911 );
or ( n57720 , n57718 , n57719 );
and ( n57721 , n47527 , n51461 );
not ( n57722 , n47527 );
and ( n57723 , n57722 , n53904 );
nor ( n57724 , n57721 , n57723 );
nand ( n57725 , n57724 , n50921 );
nand ( n57726 , n57720 , n57725 );
not ( n57727 , n57233 );
not ( n57728 , n51525 );
or ( n57729 , n57727 , n57728 );
not ( n57730 , n56727 );
not ( n57731 , n51504 );
or ( n57732 , n57730 , n57731 );
nand ( n57733 , n51818 , n56731 );
nand ( n57734 , n57732 , n57733 );
nand ( n57735 , n57734 , n51533 );
nand ( n57736 , n57729 , n57735 );
xor ( n57737 , n57726 , n57736 );
not ( n57738 , n57243 );
not ( n57739 , n54266 );
or ( n57740 , n57738 , n57739 );
not ( n57741 , n54185 );
not ( n57742 , n52130 );
or ( n57743 , n57741 , n57742 );
nand ( n57744 , n53918 , n54184 );
nand ( n57745 , n57743 , n57744 );
nand ( n57746 , n51766 , n57745 );
nand ( n57747 , n57740 , n57746 );
xor ( n57748 , n57737 , n57747 );
xor ( n57749 , n57717 , n57748 );
xor ( n57750 , n57684 , n57716 );
and ( n57751 , n57750 , n57748 );
and ( n57752 , n57684 , n57716 );
or ( n57753 , n57751 , n57752 );
xor ( n57754 , n57496 , n57492 );
xor ( n57755 , n57754 , n57488 );
xor ( n57756 , n57496 , n57492 );
and ( n57757 , n57756 , n57488 );
and ( n57758 , n57496 , n57492 );
or ( n57759 , n57757 , n57758 );
not ( n57760 , n46267 );
not ( n57761 , n57364 );
or ( n57762 , n57760 , n57761 );
not ( n57763 , n46425 );
not ( n57764 , n56020 );
or ( n57765 , n57763 , n57764 );
nand ( n57766 , n56976 , n46422 );
nand ( n57767 , n57765 , n57766 );
nand ( n57768 , n57767 , n49026 );
nand ( n57769 , n57762 , n57768 );
not ( n57770 , n51865 );
not ( n57771 , n52267 );
not ( n57772 , n53718 );
or ( n57773 , n57771 , n57772 );
nand ( n57774 , n40635 , n51351 );
nand ( n57775 , n57773 , n57774 );
not ( n57776 , n57775 );
or ( n57777 , n57770 , n57776 );
nand ( n57778 , n57375 , n49713 );
nand ( n57779 , n57777 , n57778 );
xor ( n57780 , n57769 , n57779 );
not ( n57781 , n50659 );
not ( n57782 , n57151 );
or ( n57783 , n57781 , n57782 );
not ( n57784 , n46072 );
not ( n57785 , n39893 );
or ( n57786 , n57784 , n57785 );
not ( n57787 , n39893 );
nand ( n57788 , n57787 , n50405 );
nand ( n57789 , n57786 , n57788 );
nand ( n57790 , n57789 , n44004 );
nand ( n57791 , n57783 , n57790 );
xor ( n57792 , n57780 , n57791 );
xor ( n57793 , n57792 , n57197 );
not ( n57794 , n46564 );
not ( n57795 , n57383 );
or ( n57796 , n57794 , n57795 );
not ( n57797 , n47508 );
not ( n57798 , n39962 );
not ( n57799 , n57798 );
or ( n57800 , n57797 , n57799 );
not ( n57801 , n57798 );
nand ( n57802 , n57801 , n51577 );
nand ( n57803 , n57800 , n57802 );
nand ( n57804 , n57803 , n49832 );
nand ( n57805 , n57796 , n57804 );
xor ( n57806 , n57600 , n57805 );
not ( n57807 , n52970 );
not ( n57808 , n57326 );
or ( n57809 , n57807 , n57808 );
not ( n57810 , n52048 );
not ( n57811 , n57810 );
not ( n57812 , n53730 );
or ( n57813 , n57811 , n57812 );
nand ( n57814 , n40591 , n49679 );
nand ( n57815 , n57813 , n57814 );
nand ( n57816 , n57815 , n52043 );
nand ( n57817 , n57809 , n57816 );
xor ( n57818 , n57806 , n57817 );
xor ( n57819 , n57793 , n57818 );
xor ( n57820 , n57792 , n57197 );
and ( n57821 , n57820 , n57818 );
and ( n57822 , n57792 , n57197 );
or ( n57823 , n57821 , n57822 );
not ( n57824 , n52421 );
not ( n57825 , n57335 );
or ( n57826 , n57824 , n57825 );
not ( n57827 , n48856 );
not ( n57828 , n52894 );
or ( n57829 , n57827 , n57828 );
not ( n57830 , n52222 );
nand ( n57831 , n57830 , n53228 );
nand ( n57832 , n57829 , n57831 );
nand ( n57833 , n57832 , n54875 );
nand ( n57834 , n57826 , n57833 );
not ( n57835 , n52004 );
not ( n57836 , n52377 );
not ( n57837 , n52285 );
or ( n57838 , n57836 , n57837 );
nand ( n57839 , n52289 , n53973 );
nand ( n57840 , n57838 , n57839 );
not ( n57841 , n57840 );
or ( n57842 , n57835 , n57841 );
nand ( n57843 , n57311 , n57314 );
nand ( n57844 , n57842 , n57843 );
xor ( n57845 , n57834 , n57844 );
not ( n57846 , n46776 );
not ( n57847 , n57394 );
or ( n57848 , n57846 , n57847 );
not ( n57849 , n50263 );
not ( n57850 , n55202 );
or ( n57851 , n57849 , n57850 );
nand ( n57852 , n40380 , n50087 );
nand ( n57853 , n57851 , n57852 );
nand ( n57854 , n57853 , n53631 );
nand ( n57855 , n57848 , n57854 );
xor ( n57856 , n57845 , n57855 );
not ( n57857 , n47407 );
not ( n57858 , n57348 );
or ( n57859 , n57857 , n57858 );
not ( n57860 , n54028 );
not ( n57861 , n40148 );
or ( n57862 , n57860 , n57861 );
not ( n57863 , n47803 );
nand ( n57864 , n57863 , n54406 );
nand ( n57865 , n57862 , n57864 );
nand ( n57866 , n57865 , n53675 );
nand ( n57867 , n57859 , n57866 );
not ( n57868 , n53510 );
not ( n57869 , n49500 );
not ( n57870 , n40225 );
or ( n57871 , n57869 , n57870 );
not ( n57872 , n47980 );
nand ( n57873 , n57872 , n56073 );
nand ( n57874 , n57871 , n57873 );
not ( n57875 , n57874 );
or ( n57876 , n57868 , n57875 );
nand ( n57877 , n57404 , n48989 );
nand ( n57878 , n57876 , n57877 );
xor ( n57879 , n57867 , n57878 );
xor ( n57880 , n57879 , n57561 );
xor ( n57881 , n57856 , n57880 );
xor ( n57882 , n57881 , n57606 );
xor ( n57883 , n57856 , n57880 );
and ( n57884 , n57883 , n57606 );
and ( n57885 , n57856 , n57880 );
or ( n57886 , n57884 , n57885 );
xor ( n57887 , n57203 , n57298 );
xor ( n57888 , n57887 , n57749 );
xor ( n57889 , n57203 , n57298 );
and ( n57890 , n57889 , n57749 );
and ( n57891 , n57203 , n57298 );
or ( n57892 , n57890 , n57891 );
xor ( n57893 , n57304 , n57644 );
xor ( n57894 , n57893 , n57416 );
xor ( n57895 , n57304 , n57644 );
and ( n57896 , n57895 , n57416 );
and ( n57897 , n57304 , n57644 );
or ( n57898 , n57896 , n57897 );
xor ( n57899 , n57356 , n57755 );
xor ( n57900 , n57899 , n57422 );
xor ( n57901 , n57356 , n57755 );
and ( n57902 , n57901 , n57422 );
and ( n57903 , n57356 , n57755 );
or ( n57904 , n57902 , n57903 );
xor ( n57905 , n57819 , n57882 );
xor ( n57906 , n57905 , n57888 );
xor ( n57907 , n57819 , n57882 );
and ( n57908 , n57907 , n57888 );
and ( n57909 , n57819 , n57882 );
or ( n57910 , n57908 , n57909 );
xor ( n57911 , n57726 , n57736 );
and ( n57912 , n57911 , n57747 );
and ( n57913 , n57726 , n57736 );
or ( n57914 , n57912 , n57913 );
xor ( n57915 , n57428 , n57894 );
xor ( n57916 , n57915 , n57434 );
xor ( n57917 , n57428 , n57894 );
and ( n57918 , n57917 , n57434 );
and ( n57919 , n57428 , n57894 );
or ( n57920 , n57918 , n57919 );
xor ( n57921 , n57900 , n57906 );
xor ( n57922 , n57921 , n57440 );
xor ( n57923 , n57900 , n57906 );
and ( n57924 , n57923 , n57440 );
and ( n57925 , n57900 , n57906 );
or ( n57926 , n57924 , n57925 );
xor ( n57927 , n57450 , n57916 );
xor ( n57928 , n57927 , n57456 );
xor ( n57929 , n57450 , n57916 );
and ( n57930 , n57929 , n57456 );
and ( n57931 , n57450 , n57916 );
or ( n57932 , n57930 , n57931 );
xor ( n57933 , n57922 , n57928 );
xor ( n57934 , n57933 , n57462 );
xor ( n57935 , n57922 , n57928 );
and ( n57936 , n57935 , n57462 );
and ( n57937 , n57922 , n57928 );
or ( n57938 , n57936 , n57937 );
xor ( n57939 , n57694 , n57704 );
and ( n57940 , n57939 , n57715 );
and ( n57941 , n57694 , n57704 );
or ( n57942 , n57940 , n57941 );
xor ( n57943 , n57659 , n57671 );
and ( n57944 , n57943 , n57683 );
and ( n57945 , n57659 , n57671 );
or ( n57946 , n57944 , n57945 );
xor ( n57947 , n57641 , n57099 );
and ( n57948 , n57947 , n57145 );
and ( n57949 , n57641 , n57099 );
or ( n57950 , n57948 , n57949 );
xor ( n57951 , n57600 , n57805 );
and ( n57952 , n57951 , n57817 );
and ( n57953 , n57600 , n57805 );
or ( n57954 , n57952 , n57953 );
xor ( n57955 , n57834 , n57844 );
and ( n57956 , n57955 , n57855 );
and ( n57957 , n57834 , n57844 );
or ( n57958 , n57956 , n57957 );
xor ( n57959 , n57867 , n57878 );
and ( n57960 , n57959 , n57561 );
and ( n57961 , n57867 , n57878 );
or ( n57962 , n57960 , n57961 );
xor ( n57963 , n57769 , n57779 );
and ( n57964 , n57963 , n57791 );
and ( n57965 , n57769 , n57779 );
or ( n57966 , n57964 , n57965 );
not ( n57967 , n57545 );
not ( n57968 , n50929 );
or ( n57969 , n57967 , n57968 );
and ( n57970 , n41668 , n50163 );
not ( n57971 , n41668 );
and ( n57972 , n57971 , n54613 );
or ( n57973 , n57970 , n57972 );
nand ( n57974 , n57973 , n49920 );
nand ( n57975 , n57969 , n57974 );
and ( n57976 , n41407 , n50292 );
not ( n57977 , n41407 );
and ( n57978 , n57977 , n49618 );
or ( n57979 , n57976 , n57978 );
not ( n57980 , n57979 );
or ( n57981 , n57980 , n49788 );
or ( n57982 , n50566 , n57556 );
nand ( n57983 , n57981 , n57982 );
xor ( n57984 , n57975 , n57983 );
not ( n57985 , n53104 );
not ( n57986 , n57502 );
or ( n57987 , n57985 , n57986 );
not ( n57988 , n48456 );
not ( n57989 , n41037 );
or ( n57990 , n57988 , n57989 );
nand ( n57991 , n41036 , n48967 );
nand ( n57992 , n57990 , n57991 );
nand ( n57993 , n57992 , n52723 );
nand ( n57994 , n57987 , n57993 );
xor ( n57995 , n57984 , n57994 );
xor ( n57996 , n57975 , n57983 );
and ( n57997 , n57996 , n57994 );
and ( n57998 , n57975 , n57983 );
or ( n57999 , n57997 , n57998 );
not ( n58000 , n57532 );
not ( n58001 , n36356 );
not ( n58002 , n58001 );
or ( n58003 , n58000 , n58002 );
nand ( n58004 , n57531 , n36356 );
nand ( n58005 , n58003 , n58004 );
not ( n58006 , n58005 );
nor ( n58007 , n58006 , n46441 );
not ( n58008 , n49309 );
not ( n58009 , n57573 );
not ( n58010 , n58009 );
or ( n58011 , n58008 , n58010 );
not ( n58012 , n56227 );
not ( n58013 , n40853 );
not ( n58014 , n58013 );
or ( n58015 , n58012 , n58014 );
or ( n58016 , n56227 , n58013 );
nand ( n58017 , n58015 , n58016 );
not ( n58018 , n49737 );
or ( n58019 , n58017 , n58018 );
nand ( n58020 , n58011 , n58019 );
xor ( n58021 , n58007 , n58020 );
and ( n58022 , n57547 , n57559 );
xor ( n58023 , n58021 , n58022 );
xor ( n58024 , n58007 , n58020 );
and ( n58025 , n58024 , n58022 );
and ( n58026 , n58007 , n58020 );
or ( n58027 , n58025 , n58026 );
not ( n58028 , n46564 );
not ( n58029 , n57803 );
or ( n58030 , n58028 , n58029 );
not ( n58031 , n48952 );
not ( n58032 , n39844 );
or ( n58033 , n58031 , n58032 );
not ( n58034 , n39844 );
nand ( n58035 , n58034 , n47514 );
nand ( n58036 , n58033 , n58035 );
nand ( n58037 , n58036 , n49832 );
nand ( n58038 , n58030 , n58037 );
xor ( n58039 , n58038 , n57942 );
xor ( n58040 , n58039 , n57946 );
xor ( n58041 , n58038 , n57942 );
and ( n58042 , n58041 , n57946 );
and ( n58043 , n58038 , n57942 );
or ( n58044 , n58042 , n58043 );
not ( n58045 , n46602 );
not ( n58046 , n46072 );
not ( n58047 , n39779 );
not ( n58048 , n58047 );
or ( n58049 , n58046 , n58048 );
nand ( n58050 , n39779 , n50405 );
nand ( n58051 , n58049 , n58050 );
not ( n58052 , n58051 );
or ( n58053 , n58045 , n58052 );
nand ( n58054 , n57789 , n50659 );
nand ( n58055 , n58053 , n58054 );
xor ( n58056 , n58055 , n57914 );
xor ( n58057 , n58056 , n57950 );
xor ( n58058 , n58055 , n57914 );
and ( n58059 , n58058 , n57950 );
and ( n58060 , n58055 , n57914 );
or ( n58061 , n58059 , n58060 );
and ( n58062 , n47589 , n56285 );
not ( n58063 , n47589 );
and ( n58064 , n58063 , n55891 );
or ( n58065 , n58062 , n58064 );
not ( n58066 , n55458 );
or ( n58067 , n58065 , n58066 );
not ( n58068 , n57680 );
nand ( n58069 , n55885 , n55884 );
not ( n58070 , n58069 );
nand ( n58071 , n58068 , n58070 );
nand ( n58072 , n58067 , n58071 );
not ( n58073 , n57639 );
not ( n58074 , n57628 );
or ( n58075 , n58073 , n58074 );
not ( n58076 , n54721 );
not ( n58077 , n57533 );
or ( n58078 , n58076 , n58077 );
not ( n58079 , n57619 );
nand ( n58080 , n58079 , n46037 );
nand ( n58081 , n58078 , n58080 );
nand ( n58082 , n58081 , n57139 );
nand ( n58083 , n58075 , n58082 );
xor ( n58084 , n58072 , n58083 );
not ( n58085 , n57595 );
not ( n58086 , n47873 );
or ( n58087 , n58085 , n58086 );
not ( n58088 , n40691 );
not ( n58089 , n54628 );
and ( n58090 , n58088 , n58089 );
and ( n58091 , n40691 , n51684 );
nor ( n58092 , n58090 , n58091 );
or ( n58093 , n58092 , n54622 );
nand ( n58094 , n58087 , n58093 );
xor ( n58095 , n58084 , n58094 );
or ( n58096 , n54314 , n57712 );
and ( n58097 , n51204 , n54297 );
not ( n58098 , n51204 );
and ( n58099 , n58098 , n54301 );
nor ( n58100 , n58097 , n58099 );
not ( n58101 , n58100 );
or ( n58102 , n58101 , n54076 );
nand ( n58103 , n58096 , n58102 );
not ( n58104 , n57657 );
not ( n58105 , n55143 );
or ( n58106 , n58104 , n58105 );
not ( n58107 , n48898 );
not ( n58108 , n55118 );
not ( n58109 , n58108 );
or ( n58110 , n58107 , n58109 );
nand ( n58111 , n55118 , n48897 );
nand ( n58112 , n58110 , n58111 );
nand ( n58113 , n58112 , n54848 );
nand ( n58114 , n58106 , n58113 );
xor ( n58115 , n58103 , n58114 );
not ( n58116 , n57669 );
not ( n58117 , n56776 );
or ( n58118 , n58116 , n58117 );
not ( n58119 , n47646 );
not ( n58120 , n56784 );
or ( n58121 , n58119 , n58120 );
nand ( n58122 , n56758 , n47650 );
nand ( n58123 , n58121 , n58122 );
nand ( n58124 , n56780 , n58123 );
nand ( n58125 , n58118 , n58124 );
xor ( n58126 , n58115 , n58125 );
xor ( n58127 , n58095 , n58126 );
not ( n58128 , n57745 );
not ( n58129 , n54266 );
or ( n58130 , n58128 , n58129 );
not ( n58131 , n48983 );
not ( n58132 , n52129 );
or ( n58133 , n58131 , n58132 );
nand ( n58134 , n52108 , n48980 );
nand ( n58135 , n58133 , n58134 );
nand ( n58136 , n51766 , n58135 );
nand ( n58137 , n58130 , n58136 );
not ( n58138 , n57692 );
not ( n58139 , n52853 );
or ( n58140 , n58138 , n58139 );
not ( n58141 , n54611 );
not ( n58142 , n52837 );
or ( n58143 , n58141 , n58142 );
not ( n58144 , n53946 );
nand ( n58145 , n58144 , n51670 );
nand ( n58146 , n58143 , n58145 );
nand ( n58147 , n53571 , n58146 );
nand ( n58148 , n58140 , n58147 );
xor ( n58149 , n58137 , n58148 );
not ( n58150 , n57702 );
not ( n58151 , n53956 );
or ( n58152 , n58150 , n58151 );
not ( n58153 , n51792 );
not ( n58154 , n53594 );
or ( n58155 , n58153 , n58154 );
nand ( n58156 , n53590 , n48829 );
nand ( n58157 , n58155 , n58156 );
not ( n58158 , n58157 );
or ( n58159 , n58158 , n53618 );
nand ( n58160 , n58152 , n58159 );
xor ( n58161 , n58149 , n58160 );
xor ( n58162 , n58127 , n58161 );
xor ( n58163 , n58095 , n58126 );
and ( n58164 , n58163 , n58161 );
and ( n58165 , n58095 , n58126 );
or ( n58166 , n58164 , n58165 );
not ( n58167 , n50195 );
not ( n58168 , n58167 );
not ( n58169 , n58168 );
not ( n58170 , n57582 );
or ( n58171 , n58169 , n58170 );
not ( n58172 , n41284 );
xor ( n58173 , n49109 , n58172 );
nand ( n58174 , n58173 , n52191 );
nand ( n58175 , n58171 , n58174 );
not ( n58176 , n57724 );
not ( n58177 , n52151 );
or ( n58178 , n58176 , n58177 );
buf ( n58179 , n51193 );
not ( n58180 , n58179 );
not ( n58181 , n58180 );
not ( n58182 , n50916 );
or ( n58183 , n58181 , n58182 );
nand ( n58184 , n51461 , n41416 );
nand ( n58185 , n58183 , n58184 );
nand ( n58186 , n58185 , n50921 );
nand ( n58187 , n58178 , n58186 );
xor ( n58188 , n58175 , n58187 );
not ( n58189 , n53543 );
not ( n58190 , n57734 );
or ( n58191 , n58189 , n58190 );
not ( n58192 , n57182 );
not ( n58193 , n51508 );
or ( n58194 , n58192 , n58193 );
buf ( n58195 , n47332 );
nand ( n58196 , n53549 , n58195 );
nand ( n58197 , n58194 , n58196 );
not ( n58198 , n58197 );
or ( n58199 , n53927 , n58198 );
nand ( n58200 , n58191 , n58199 );
xor ( n58201 , n58188 , n58200 );
xor ( n58202 , n58201 , n57958 );
xor ( n58203 , n57995 , n57565 );
not ( n58204 , n46267 );
not ( n58205 , n57767 );
or ( n58206 , n58204 , n58205 );
and ( n58207 , n40011 , n46422 );
not ( n58208 , n40011 );
and ( n58209 , n58208 , n46425 );
or ( n58210 , n58207 , n58209 );
nand ( n58211 , n58210 , n49026 );
nand ( n58212 , n58206 , n58211 );
xor ( n58213 , n58203 , n58212 );
xor ( n58214 , n58202 , n58213 );
xor ( n58215 , n58201 , n57958 );
and ( n58216 , n58215 , n58213 );
and ( n58217 , n58201 , n57958 );
or ( n58218 , n58216 , n58217 );
xor ( n58219 , n57962 , n57954 );
not ( n58220 , n52043 );
not ( n58221 , n48645 );
not ( n58222 , n54046 );
or ( n58223 , n58221 , n58222 );
nand ( n58224 , n40626 , n49679 );
nand ( n58225 , n58223 , n58224 );
not ( n58226 , n58225 );
or ( n58227 , n58220 , n58226 );
nand ( n58228 , n57815 , n50242 );
nand ( n58229 , n58227 , n58228 );
not ( n58230 , n52421 );
not ( n58231 , n57832 );
or ( n58232 , n58230 , n58231 );
not ( n58233 , n48856 );
not ( n58234 , n52570 );
or ( n58235 , n58233 , n58234 );
not ( n58236 , n54771 );
nand ( n58237 , n58236 , n51724 );
nand ( n58238 , n58235 , n58237 );
nand ( n58239 , n58238 , n54875 );
nand ( n58240 , n58232 , n58239 );
xor ( n58241 , n58229 , n58240 );
not ( n58242 , n52004 );
not ( n58243 , n52377 );
not ( n58244 , n51928 );
or ( n58245 , n58243 , n58244 );
not ( n58246 , n40732 );
nand ( n58247 , n58246 , n53973 );
nand ( n58248 , n58245 , n58247 );
not ( n58249 , n58248 );
or ( n58250 , n58242 , n58249 );
not ( n58251 , n57840 );
or ( n58252 , n58251 , n56515 );
nand ( n58253 , n58250 , n58252 );
xor ( n58254 , n58241 , n58253 );
xor ( n58255 , n58219 , n58254 );
xor ( n58256 , n57962 , n57954 );
and ( n58257 , n58256 , n58254 );
and ( n58258 , n57962 , n57954 );
or ( n58259 , n58257 , n58258 );
not ( n58260 , n49252 );
not ( n58261 , n57874 );
or ( n58262 , n58260 , n58261 );
not ( n58263 , n49500 );
not ( n58264 , n54810 );
or ( n58265 , n58263 , n58264 );
nand ( n58266 , n40363 , n47979 );
nand ( n58267 , n58265 , n58266 );
nand ( n58268 , n58267 , n53510 );
nand ( n58269 , n58262 , n58268 );
not ( n58270 , n49713 );
not ( n58271 , n57775 );
or ( n58272 , n58270 , n58271 );
not ( n58273 , n52267 );
not ( n58274 , n53289 );
or ( n58275 , n58273 , n58274 );
nand ( n58276 , n40377 , n52273 );
nand ( n58277 , n58275 , n58276 );
nand ( n58278 , n58277 , n51865 );
nand ( n58279 , n58272 , n58278 );
xor ( n58280 , n58269 , n58279 );
xor ( n58281 , n58280 , n57604 );
xor ( n58282 , n58281 , n57966 );
xor ( n58283 , n58282 , n57610 );
xor ( n58284 , n58281 , n57966 );
and ( n58285 , n58284 , n57610 );
and ( n58286 , n58281 , n57966 );
or ( n58287 , n58285 , n58286 );
not ( n58288 , n47827 );
and ( n58289 , n40451 , n50087 );
not ( n58290 , n40451 );
and ( n58291 , n58290 , n50263 );
or ( n58292 , n58289 , n58291 );
not ( n58293 , n58292 );
or ( n58294 , n58288 , n58293 );
nand ( n58295 , n57853 , n46776 );
nand ( n58296 , n58294 , n58295 );
not ( n58297 , n47407 );
not ( n58298 , n57865 );
or ( n58299 , n58297 , n58298 );
not ( n58300 , n54028 );
not ( n58301 , n54790 );
or ( n58302 , n58300 , n58301 );
nand ( n58303 , n40388 , n48727 );
nand ( n58304 , n58302 , n58303 );
nand ( n58305 , n58304 , n53675 );
nand ( n58306 , n58299 , n58305 );
xor ( n58307 , n58296 , n58306 );
xor ( n58308 , n58307 , n58023 );
xor ( n58309 , n58308 , n57753 );
xor ( n58310 , n58309 , n57648 );
xor ( n58311 , n58308 , n57753 );
and ( n58312 , n58311 , n57648 );
and ( n58313 , n58308 , n57753 );
or ( n58314 , n58312 , n58313 );
xor ( n58315 , n58057 , n58040 );
xor ( n58316 , n58315 , n58162 );
xor ( n58317 , n58057 , n58040 );
and ( n58318 , n58317 , n58162 );
and ( n58319 , n58057 , n58040 );
or ( n58320 , n58318 , n58319 );
xor ( n58321 , n57759 , n57823 );
xor ( n58322 , n58321 , n58255 );
xor ( n58323 , n57759 , n57823 );
and ( n58324 , n58323 , n58255 );
and ( n58325 , n57759 , n57823 );
or ( n58326 , n58324 , n58325 );
xor ( n58327 , n58214 , n57886 );
xor ( n58328 , n58327 , n58283 );
xor ( n58329 , n58214 , n57886 );
and ( n58330 , n58329 , n58283 );
and ( n58331 , n58214 , n57886 );
or ( n58332 , n58330 , n58331 );
xor ( n58333 , n58175 , n58187 );
and ( n58334 , n58333 , n58200 );
and ( n58335 , n58175 , n58187 );
or ( n58336 , n58334 , n58335 );
xor ( n58337 , n58316 , n58310 );
xor ( n58338 , n58337 , n57892 );
xor ( n58339 , n58316 , n58310 );
and ( n58340 , n58339 , n57892 );
and ( n58341 , n58316 , n58310 );
or ( n58342 , n58340 , n58341 );
xor ( n58343 , n57898 , n57904 );
xor ( n58344 , n58343 , n58322 );
xor ( n58345 , n57898 , n57904 );
and ( n58346 , n58345 , n58322 );
and ( n58347 , n57898 , n57904 );
or ( n58348 , n58346 , n58347 );
xor ( n58349 , n58328 , n57910 );
xor ( n58350 , n58349 , n57920 );
xor ( n58351 , n58328 , n57910 );
and ( n58352 , n58351 , n57920 );
and ( n58353 , n58328 , n57910 );
or ( n58354 , n58352 , n58353 );
xor ( n58355 , n58338 , n58344 );
xor ( n58356 , n58355 , n57926 );
xor ( n58357 , n58338 , n58344 );
and ( n58358 , n58357 , n57926 );
and ( n58359 , n58338 , n58344 );
or ( n58360 , n58358 , n58359 );
xor ( n58361 , n58350 , n57932 );
xor ( n58362 , n58361 , n58356 );
xor ( n58363 , n58350 , n57932 );
and ( n58364 , n58363 , n58356 );
and ( n58365 , n58350 , n57932 );
or ( n58366 , n58364 , n58365 );
xor ( n58367 , n58137 , n58148 );
and ( n58368 , n58367 , n58160 );
and ( n58369 , n58137 , n58148 );
or ( n58370 , n58368 , n58369 );
xor ( n58371 , n58103 , n58114 );
and ( n58372 , n58371 , n58125 );
and ( n58373 , n58103 , n58114 );
or ( n58374 , n58372 , n58373 );
xor ( n58375 , n58072 , n58083 );
and ( n58376 , n58375 , n58094 );
and ( n58377 , n58072 , n58083 );
or ( n58378 , n58376 , n58377 );
xor ( n58379 , n57995 , n57565 );
and ( n58380 , n58379 , n58212 );
and ( n58381 , n57995 , n57565 );
or ( n58382 , n58380 , n58381 );
xor ( n58383 , n58229 , n58240 );
and ( n58384 , n58383 , n58253 );
and ( n58385 , n58229 , n58240 );
or ( n58386 , n58384 , n58385 );
xor ( n58387 , n58296 , n58306 );
and ( n58388 , n58387 , n58023 );
and ( n58389 , n58296 , n58306 );
or ( n58390 , n58388 , n58389 );
xor ( n58391 , n58269 , n58279 );
and ( n58392 , n58391 , n57604 );
and ( n58393 , n58269 , n58279 );
or ( n58394 , n58392 , n58393 );
not ( n58395 , n49979 );
not ( n58396 , n58173 );
or ( n58397 , n58395 , n58396 );
not ( n58398 , n49283 );
and ( n58399 , n831 , n41213 );
not ( n58400 , n831 );
and ( n58401 , n58400 , n41174 );
nor ( n58402 , n58399 , n58401 );
or ( n58403 , n58398 , n58402 );
nand ( n58404 , n58402 , n50201 );
nand ( n58405 , n58403 , n58404 );
nand ( n58406 , n58405 , n50514 );
nand ( n58407 , n58397 , n58406 );
not ( n58408 , n49789 );
not ( n58409 , n49619 );
not ( n58410 , n50980 );
or ( n58411 , n58409 , n58410 );
nand ( n58412 , n41363 , n49766 );
nand ( n58413 , n58411 , n58412 );
not ( n58414 , n58413 );
or ( n58415 , n58408 , n58414 );
nand ( n58416 , n57979 , n51234 );
nand ( n58417 , n58415 , n58416 );
xor ( n58418 , n58407 , n58417 );
not ( n58419 , n46440 );
not ( n58420 , n36356 );
not ( n58421 , n58420 );
not ( n58422 , n58421 );
or ( n58423 , n58419 , n58422 );
nand ( n58424 , n58423 , n57633 );
nand ( n58425 , n58420 , n46441 );
and ( n58426 , n58424 , n58425 );
and ( n58427 , n36389 , n37572 );
not ( n58428 , n36389 );
not ( n58429 , n37572 );
and ( n58430 , n58428 , n58429 );
nor ( n58431 , n58427 , n58430 );
not ( n58432 , n58431 );
not ( n58433 , n58432 );
nor ( n58434 , n58426 , n58433 );
xor ( n58435 , n58418 , n58434 );
xor ( n58436 , n58407 , n58417 );
and ( n58437 , n58436 , n58434 );
and ( n58438 , n58407 , n58417 );
or ( n58439 , n58437 , n58438 );
not ( n58440 , n57992 );
not ( n58441 , n50176 );
or ( n58442 , n58440 , n58441 );
not ( n58443 , n52722 );
and ( n58444 , n41132 , n48456 );
not ( n58445 , n41132 );
and ( n58446 , n58445 , n52728 );
nor ( n58447 , n58444 , n58446 );
nand ( n58448 , n58443 , n58447 );
nand ( n58449 , n58442 , n58448 );
not ( n58450 , n58185 );
not ( n58451 , n50911 );
or ( n58452 , n58450 , n58451 );
not ( n58453 , n52954 );
not ( n58454 , n58453 );
not ( n58455 , n58454 );
not ( n58456 , n53904 );
or ( n58457 , n58455 , n58456 );
not ( n58458 , n49297 );
not ( n58459 , n58458 );
nand ( n58460 , n50898 , n58459 );
nand ( n58461 , n58457 , n58460 );
nand ( n58462 , n58461 , n50921 );
nand ( n58463 , n58452 , n58462 );
xor ( n58464 , n58449 , n58463 );
not ( n58465 , n58197 );
not ( n58466 , n51525 );
or ( n58467 , n58465 , n58466 );
not ( n58468 , n47527 );
not ( n58469 , n51504 );
or ( n58470 , n58468 , n58469 );
nand ( n58471 , n56361 , n51360 );
nand ( n58472 , n58470 , n58471 );
nand ( n58473 , n51533 , n58472 );
nand ( n58474 , n58467 , n58473 );
xor ( n58475 , n58464 , n58474 );
xor ( n58476 , n58449 , n58463 );
and ( n58477 , n58476 , n58474 );
and ( n58478 , n58449 , n58463 );
or ( n58479 , n58477 , n58478 );
not ( n58480 , n47009 );
not ( n58481 , n46072 );
not ( n58482 , n39678 );
not ( n58483 , n58482 );
or ( n58484 , n58481 , n58483 );
not ( n58485 , n39679 );
nand ( n58486 , n58485 , n46071 );
nand ( n58487 , n58484 , n58486 );
not ( n58488 , n58487 );
or ( n58489 , n58480 , n58488 );
nand ( n58490 , n58051 , n50659 );
nand ( n58491 , n58489 , n58490 );
xor ( n58492 , n58374 , n58491 );
xor ( n58493 , n58492 , n58336 );
xor ( n58494 , n58374 , n58491 );
and ( n58495 , n58494 , n58336 );
and ( n58496 , n58374 , n58491 );
or ( n58497 , n58495 , n58496 );
not ( n58498 , n58135 );
not ( n58499 , n54265 );
or ( n58500 , n58498 , n58499 );
xor ( n58501 , n47510 , n52129 );
nand ( n58502 , n58501 , n51765 );
nand ( n58503 , n58500 , n58502 );
not ( n58504 , n58146 );
not ( n58505 , n52852 );
or ( n58506 , n58504 , n58505 );
not ( n58507 , n54185 );
not ( n58508 , n57252 );
or ( n58509 , n58507 , n58508 );
nand ( n58510 , n58144 , n52712 );
nand ( n58511 , n58509 , n58510 );
nand ( n58512 , n58511 , n52468 );
nand ( n58513 , n58506 , n58512 );
xor ( n58514 , n58503 , n58513 );
not ( n58515 , n58157 );
not ( n58516 , n55913 );
or ( n58517 , n58515 , n58516 );
not ( n58518 , n52033 );
not ( n58519 , n56802 );
or ( n58520 , n58518 , n58519 );
nand ( n58521 , n53590 , n55959 );
nand ( n58522 , n58520 , n58521 );
nand ( n58523 , n58522 , n53619 );
nand ( n58524 , n58517 , n58523 );
xor ( n58525 , n58514 , n58524 );
xor ( n58526 , n58525 , n58378 );
not ( n58527 , n58123 );
not ( n58528 , n56774 );
nor ( n58529 , n58528 , n56500 );
not ( n58530 , n58529 );
or ( n58531 , n58527 , n58530 );
and ( n58532 , n49734 , n57664 );
not ( n58533 , n49734 );
not ( n58534 , n57664 );
and ( n58535 , n58533 , n58534 );
nor ( n58536 , n58532 , n58535 );
nand ( n58537 , n58536 , n56500 );
nand ( n58538 , n58531 , n58537 );
not ( n58539 , n58081 );
nand ( n58540 , n57138 , n57626 );
not ( n58541 , n58540 );
not ( n58542 , n58541 );
or ( n58543 , n58539 , n58542 );
not ( n58544 , n46273 );
not ( n58545 , n57633 );
or ( n58546 , n58544 , n58545 );
nand ( n58547 , n57619 , n46824 );
nand ( n58548 , n58546 , n58547 );
nand ( n58549 , n58548 , n57139 );
nand ( n58550 , n58543 , n58549 );
xor ( n58551 , n58538 , n58550 );
not ( n58552 , n57973 );
not ( n58553 , n50321 );
or ( n58554 , n58552 , n58553 );
not ( n58555 , n50304 );
buf ( n58556 , n41530 );
not ( n58557 , n58556 );
or ( n58558 , n58555 , n58557 );
nand ( n58559 , n50301 , n41531 );
nand ( n58560 , n58558 , n58559 );
nand ( n58561 , n58560 , n50331 );
nand ( n58562 , n58554 , n58561 );
not ( n58563 , n49320 );
and ( n58564 , n49809 , n48764 );
not ( n58565 , n49809 );
and ( n58566 , n58565 , n49314 );
or ( n58567 , n58564 , n58566 );
not ( n58568 , n58567 );
or ( n58569 , n58563 , n58568 );
not ( n58570 , n58017 );
nand ( n58571 , n58570 , n49309 );
nand ( n58572 , n58569 , n58571 );
xor ( n58573 , n58562 , n58572 );
xor ( n58574 , n58551 , n58573 );
xor ( n58575 , n58526 , n58574 );
xor ( n58576 , n58525 , n58378 );
and ( n58577 , n58576 , n58574 );
and ( n58578 , n58525 , n58378 );
or ( n58579 , n58577 , n58578 );
not ( n58580 , n56277 );
not ( n58581 , n49624 );
not ( n58582 , n54301 );
or ( n58583 , n58581 , n58582 );
nand ( n58584 , n54297 , n49630 );
nand ( n58585 , n58583 , n58584 );
not ( n58586 , n58585 );
or ( n58587 , n58580 , n58586 );
nand ( n58588 , n58100 , n54313 );
nand ( n58589 , n58587 , n58588 );
not ( n58590 , n58112 );
nand ( n58591 , n55137 , n55141 );
not ( n58592 , n58591 );
not ( n58593 , n58592 );
or ( n58594 , n58590 , n58593 );
not ( n58595 , n47765 );
not ( n58596 , n58108 );
or ( n58597 , n58595 , n58596 );
nand ( n58598 , n55118 , n48589 );
nand ( n58599 , n58597 , n58598 );
nand ( n58600 , n54847 , n58599 );
nand ( n58601 , n58594 , n58600 );
xor ( n58602 , n58589 , n58601 );
not ( n58603 , n49654 );
not ( n58604 , n55891 );
not ( n58605 , n58604 );
or ( n58606 , n58603 , n58605 );
nand ( n58607 , n55891 , n47368 );
nand ( n58608 , n58606 , n58607 );
not ( n58609 , n58608 );
not ( n58610 , n55458 );
or ( n58611 , n58609 , n58610 );
not ( n58612 , n58065 );
nand ( n58613 , n58612 , n55887 );
nand ( n58614 , n58611 , n58613 );
xor ( n58615 , n58602 , n58614 );
xor ( n58616 , n58615 , n58475 );
xor ( n58617 , n58616 , n58386 );
xor ( n58618 , n58615 , n58475 );
and ( n58619 , n58618 , n58386 );
and ( n58620 , n58615 , n58475 );
or ( n58621 , n58619 , n58620 );
xor ( n58622 , n58390 , n58394 );
not ( n58623 , n48689 );
not ( n58624 , n58433 );
or ( n58625 , n58623 , n58624 );
not ( n58626 , n58433 );
nand ( n58627 , n58626 , n46441 );
nand ( n58628 , n58625 , n58627 );
not ( n58629 , n58628 );
buf ( n58630 , n58431 );
and ( n58631 , n58630 , n58420 );
not ( n58632 , n58630 );
and ( n58633 , n58632 , n36356 );
nor ( n58634 , n58631 , n58633 );
and ( n58635 , n58006 , n58634 );
not ( n58636 , n58635 );
or ( n58637 , n58629 , n58636 );
not ( n58638 , n58006 );
not ( n58639 , n45816 );
not ( n58640 , n58630 );
or ( n58641 , n58639 , n58640 );
buf ( n58642 , n58432 );
nand ( n58643 , n58642 , n48766 );
nand ( n58644 , n58641 , n58643 );
nand ( n58645 , n58638 , n58644 );
nand ( n58646 , n58637 , n58645 );
xor ( n58647 , n58646 , n57999 );
xor ( n58648 , n58647 , n58027 );
xor ( n58649 , n58622 , n58648 );
xor ( n58650 , n58390 , n58394 );
and ( n58651 , n58650 , n58648 );
and ( n58652 , n58390 , n58394 );
or ( n58653 , n58651 , n58652 );
not ( n58654 , n46188 );
xnor ( n58655 , n46422 , n39962 );
not ( n58656 , n58655 );
or ( n58657 , n58654 , n58656 );
nand ( n58658 , n58210 , n46267 );
nand ( n58659 , n58657 , n58658 );
xor ( n58660 , n58659 , n58435 );
not ( n58661 , n51865 );
not ( n58662 , n49707 );
not ( n58663 , n56074 );
or ( n58664 , n58662 , n58663 );
nand ( n58665 , n54433 , n51351 );
nand ( n58666 , n58664 , n58665 );
not ( n58667 , n58666 );
or ( n58668 , n58661 , n58667 );
nand ( n58669 , n58277 , n49713 );
nand ( n58670 , n58668 , n58669 );
xor ( n58671 , n58660 , n58670 );
xor ( n58672 , n58382 , n58671 );
not ( n58673 , n58292 );
or ( n58674 , n58673 , n46775 );
not ( n58675 , n40512 );
not ( n58676 , n48078 );
and ( n58677 , n58675 , n58676 );
and ( n58678 , n40512 , n50087 );
nor ( n58679 , n58677 , n58678 );
or ( n58680 , n56080 , n58679 );
nand ( n58681 , n58674 , n58680 );
not ( n58682 , n58225 );
or ( n58683 , n58682 , n50241 );
and ( n58684 , n40635 , n48645 );
not ( n58685 , n40635 );
and ( n58686 , n58685 , n52048 );
or ( n58687 , n58684 , n58686 );
or ( n58688 , n50239 , n58687 );
nand ( n58689 , n58683 , n58688 );
xor ( n58690 , n58681 , n58689 );
not ( n58691 , n54875 );
not ( n58692 , n48856 );
and ( n58693 , n40590 , n58692 );
not ( n58694 , n40590 );
and ( n58695 , n58694 , n51723 );
or ( n58696 , n58693 , n58695 );
not ( n58697 , n58696 );
or ( n58698 , n58691 , n58697 );
not ( n58699 , n58238 );
not ( n58700 , n52421 );
or ( n58701 , n58699 , n58700 );
nand ( n58702 , n58698 , n58701 );
xor ( n58703 , n58690 , n58702 );
xor ( n58704 , n58672 , n58703 );
xor ( n58705 , n58382 , n58671 );
and ( n58706 , n58705 , n58703 );
and ( n58707 , n58382 , n58671 );
or ( n58708 , n58706 , n58707 );
not ( n58709 , n48894 );
not ( n58710 , n58248 );
or ( n58711 , n58709 , n58710 );
and ( n58712 , n53973 , n52222 );
not ( n58713 , n53973 );
and ( n58714 , n58713 , n40769 );
nor ( n58715 , n58712 , n58714 );
nand ( n58716 , n58715 , n52004 );
nand ( n58717 , n58711 , n58716 );
not ( n58718 , n47407 );
not ( n58719 , n58304 );
or ( n58720 , n58718 , n58719 );
and ( n58721 , n40380 , n48727 );
not ( n58722 , n40380 );
and ( n58723 , n58722 , n47803 );
or ( n58724 , n58721 , n58723 );
nand ( n58725 , n58724 , n53675 );
nand ( n58726 , n58720 , n58725 );
xor ( n58727 , n58717 , n58726 );
not ( n58728 , n51680 );
not ( n58729 , n51573 );
or ( n58730 , n58728 , n58729 );
nand ( n58731 , n40677 , n51684 );
nand ( n58732 , n58730 , n58731 );
not ( n58733 , n58732 );
or ( n58734 , n58733 , n54622 );
not ( n58735 , n58092 );
nand ( n58736 , n58735 , n52022 );
nand ( n58737 , n58734 , n58736 );
xor ( n58738 , n58727 , n58737 );
xor ( n58739 , n58044 , n58738 );
not ( n58740 , n53510 );
not ( n58741 , n49500 );
not ( n58742 , n40148 );
or ( n58743 , n58741 , n58742 );
nand ( n58744 , n56010 , n47979 );
nand ( n58745 , n58743 , n58744 );
not ( n58746 , n58745 );
or ( n58747 , n58740 , n58746 );
nand ( n58748 , n58267 , n48989 );
nand ( n58749 , n58747 , n58748 );
not ( n58750 , n46564 );
not ( n58751 , n58036 );
or ( n58752 , n58750 , n58751 );
not ( n58753 , n52990 );
not ( n58754 , n57787 );
or ( n58755 , n58753 , n58754 );
nand ( n58756 , n39893 , n48952 );
nand ( n58757 , n58755 , n58756 );
nand ( n58758 , n58757 , n49832 );
nand ( n58759 , n58752 , n58758 );
xor ( n58760 , n58749 , n58759 );
xor ( n58761 , n58760 , n58370 );
xor ( n58762 , n58739 , n58761 );
xor ( n58763 , n58044 , n58738 );
and ( n58764 , n58763 , n58761 );
and ( n58765 , n58044 , n58738 );
or ( n58766 , n58764 , n58765 );
xor ( n58767 , n58061 , n58166 );
xor ( n58768 , n58767 , n58493 );
xor ( n58769 , n58061 , n58166 );
and ( n58770 , n58769 , n58493 );
and ( n58771 , n58061 , n58166 );
or ( n58772 , n58770 , n58771 );
xor ( n58773 , n58575 , n58617 );
xor ( n58774 , n58773 , n58218 );
xor ( n58775 , n58575 , n58617 );
and ( n58776 , n58775 , n58218 );
and ( n58777 , n58575 , n58617 );
or ( n58778 , n58776 , n58777 );
xor ( n58779 , n58649 , n58287 );
xor ( n58780 , n58779 , n58259 );
xor ( n58781 , n58649 , n58287 );
and ( n58782 , n58781 , n58259 );
and ( n58783 , n58649 , n58287 );
or ( n58784 , n58782 , n58783 );
xor ( n58785 , n58314 , n58704 );
xor ( n58786 , n58785 , n58762 );
xor ( n58787 , n58314 , n58704 );
and ( n58788 , n58787 , n58762 );
and ( n58789 , n58314 , n58704 );
or ( n58790 , n58788 , n58789 );
xor ( n58791 , n58503 , n58513 );
and ( n58792 , n58791 , n58524 );
and ( n58793 , n58503 , n58513 );
or ( n58794 , n58792 , n58793 );
xor ( n58795 , n58768 , n58320 );
xor ( n58796 , n58795 , n58774 );
xor ( n58797 , n58768 , n58320 );
and ( n58798 , n58797 , n58774 );
and ( n58799 , n58768 , n58320 );
or ( n58800 , n58798 , n58799 );
xor ( n58801 , n58326 , n58780 );
xor ( n58802 , n58801 , n58332 );
xor ( n58803 , n58326 , n58780 );
and ( n58804 , n58803 , n58332 );
and ( n58805 , n58326 , n58780 );
or ( n58806 , n58804 , n58805 );
xor ( n58807 , n58342 , n58786 );
xor ( n58808 , n58807 , n58796 );
xor ( n58809 , n58342 , n58786 );
and ( n58810 , n58809 , n58796 );
and ( n58811 , n58342 , n58786 );
or ( n58812 , n58810 , n58811 );
xor ( n58813 , n58348 , n58802 );
xor ( n58814 , n58813 , n58354 );
xor ( n58815 , n58348 , n58802 );
and ( n58816 , n58815 , n58354 );
and ( n58817 , n58348 , n58802 );
or ( n58818 , n58816 , n58817 );
xor ( n58819 , n58808 , n58360 );
xor ( n58820 , n58819 , n58814 );
xor ( n58821 , n58808 , n58360 );
and ( n58822 , n58821 , n58814 );
and ( n58823 , n58808 , n58360 );
or ( n58824 , n58822 , n58823 );
xor ( n58825 , n58589 , n58601 );
and ( n58826 , n58825 , n58614 );
and ( n58827 , n58589 , n58601 );
or ( n58828 , n58826 , n58827 );
xor ( n58829 , n58538 , n58550 );
and ( n58830 , n58829 , n58573 );
and ( n58831 , n58538 , n58550 );
or ( n58832 , n58830 , n58831 );
xor ( n58833 , n58646 , n57999 );
and ( n58834 , n58833 , n58027 );
and ( n58835 , n58646 , n57999 );
or ( n58836 , n58834 , n58835 );
xor ( n58837 , n58681 , n58689 );
and ( n58838 , n58837 , n58702 );
and ( n58839 , n58681 , n58689 );
or ( n58840 , n58838 , n58839 );
xor ( n58841 , n58717 , n58726 );
and ( n58842 , n58841 , n58737 );
and ( n58843 , n58717 , n58726 );
or ( n58844 , n58842 , n58843 );
xor ( n58845 , n58659 , n58435 );
and ( n58846 , n58845 , n58670 );
and ( n58847 , n58659 , n58435 );
or ( n58848 , n58846 , n58847 );
xor ( n58849 , n58749 , n58759 );
and ( n58850 , n58849 , n58370 );
and ( n58851 , n58749 , n58759 );
or ( n58852 , n58850 , n58851 );
not ( n58853 , n51452 );
not ( n58854 , n51250 );
not ( n58855 , n48483 );
or ( n58856 , n58854 , n58855 );
not ( n58857 , n54613 );
nand ( n58858 , n58857 , n41407 );
nand ( n58859 , n58856 , n58858 );
not ( n58860 , n58859 );
or ( n58861 , n58853 , n58860 );
not ( n58862 , n50319 );
nand ( n58863 , n58862 , n58560 );
nand ( n58864 , n58861 , n58863 );
not ( n58865 , n49309 );
not ( n58866 , n58567 );
or ( n58867 , n58865 , n58866 );
not ( n58868 , n48705 );
not ( n58869 , n51110 );
or ( n58870 , n58868 , n58869 );
nand ( n58871 , n41036 , n49094 );
nand ( n58872 , n58870 , n58871 );
nand ( n58873 , n58872 , n56639 );
nand ( n58874 , n58867 , n58873 );
xor ( n58875 , n58864 , n58874 );
not ( n58876 , n49288 );
not ( n58877 , n49452 );
not ( n58878 , n51741 );
or ( n58879 , n58877 , n58878 );
nand ( n58880 , n51740 , n57088 );
nand ( n58881 , n58879 , n58880 );
not ( n58882 , n58881 );
or ( n58883 , n58876 , n58882 );
buf ( n58884 , n58405 );
nand ( n58885 , n50195 , n58884 );
nand ( n58886 , n58883 , n58885 );
xor ( n58887 , n58875 , n58886 );
xor ( n58888 , n58864 , n58874 );
and ( n58889 , n58888 , n58886 );
and ( n58890 , n58864 , n58874 );
or ( n58891 , n58889 , n58890 );
not ( n58892 , n50078 );
not ( n58893 , n49619 );
not ( n58894 , n41285 );
or ( n58895 , n58893 , n58894 );
nand ( n58896 , n49001 , n52740 );
nand ( n58897 , n58895 , n58896 );
not ( n58898 , n58897 );
or ( n58899 , n58892 , n58898 );
nand ( n58900 , n58413 , n52058 );
nand ( n58901 , n58899 , n58900 );
not ( n58902 , n36337 );
and ( n58903 , n58432 , n58902 );
not ( n58904 , n58432 );
and ( n58905 , n58904 , n36337 );
nor ( n58906 , n58903 , n58905 );
buf ( n58907 , n58906 );
not ( n58908 , n58907 );
and ( n58909 , n58908 , n46440 );
xor ( n58910 , n58901 , n58909 );
not ( n58911 , n58461 );
not ( n58912 , n50911 );
or ( n58913 , n58911 , n58912 );
buf ( n58914 , n49029 );
not ( n58915 , n58914 );
not ( n58916 , n58915 );
not ( n58917 , n51462 );
or ( n58918 , n58916 , n58917 );
nand ( n58919 , n50898 , n58914 );
nand ( n58920 , n58918 , n58919 );
nand ( n58921 , n58920 , n50921 );
nand ( n58922 , n58913 , n58921 );
xor ( n58923 , n58910 , n58922 );
xor ( n58924 , n58901 , n58909 );
and ( n58925 , n58924 , n58922 );
and ( n58926 , n58901 , n58909 );
or ( n58927 , n58925 , n58926 );
xor ( n58928 , n58828 , n58832 );
not ( n58929 , n50659 );
not ( n58930 , n58487 );
or ( n58931 , n58929 , n58930 );
not ( n58932 , n46072 );
not ( n58933 , n39714 );
not ( n58934 , n58933 );
or ( n58935 , n58932 , n58934 );
nand ( n58936 , n39714 , n50405 );
nand ( n58937 , n58935 , n58936 );
nand ( n58938 , n58937 , n44004 );
nand ( n58939 , n58931 , n58938 );
xor ( n58940 , n58928 , n58939 );
xor ( n58941 , n58828 , n58832 );
and ( n58942 , n58941 , n58939 );
and ( n58943 , n58828 , n58832 );
or ( n58944 , n58942 , n58943 );
not ( n58945 , n58655 );
not ( n58946 , n46267 );
or ( n58947 , n58945 , n58946 );
and ( n58948 , n46425 , n39844 );
not ( n58949 , n46425 );
and ( n58950 , n58949 , n39845 );
nor ( n58951 , n58948 , n58950 );
or ( n58952 , n58951 , n49025 );
nand ( n58953 , n58947 , n58952 );
xor ( n58954 , n58923 , n58953 );
xor ( n58955 , n58954 , n58479 );
xor ( n58956 , n58923 , n58953 );
and ( n58957 , n58956 , n58479 );
and ( n58958 , n58923 , n58953 );
or ( n58959 , n58957 , n58958 );
not ( n58960 , n58644 );
nand ( n58961 , n58006 , n58634 );
not ( n58962 , n58961 );
not ( n58963 , n58962 );
or ( n58964 , n58960 , n58963 );
not ( n58965 , n54722 );
not ( n58966 , n58642 );
not ( n58967 , n58966 );
or ( n58968 , n58965 , n58967 );
not ( n58969 , n46037 );
nand ( n58970 , n58969 , n58642 );
nand ( n58971 , n58968 , n58970 );
nand ( n58972 , n58971 , n58638 );
nand ( n58973 , n58964 , n58972 );
and ( n58974 , n58572 , n58562 );
xor ( n58975 , n58973 , n58974 );
not ( n58976 , n52723 );
not ( n58977 , n58976 );
not ( n58978 , n58977 );
not ( n58979 , n52728 );
not ( n58980 , n40691 );
or ( n58981 , n58979 , n58980 );
buf ( n58982 , n53439 );
nand ( n58983 , n57307 , n58982 );
nand ( n58984 , n58981 , n58983 );
not ( n58985 , n58984 );
or ( n58986 , n58978 , n58985 );
nand ( n58987 , n58447 , n53104 );
nand ( n58988 , n58986 , n58987 );
xor ( n58989 , n58975 , n58988 );
xor ( n58990 , n58836 , n58989 );
not ( n58991 , n58472 );
not ( n58992 , n53169 );
or ( n58993 , n58991 , n58992 );
buf ( n58994 , n52379 );
not ( n58995 , n58994 );
not ( n58996 , n51504 );
or ( n58997 , n58995 , n58996 );
nand ( n58998 , n52816 , n58179 );
nand ( n58999 , n58997 , n58998 );
nand ( n59000 , n58999 , n51145 );
nand ( n59001 , n58993 , n59000 );
not ( n59002 , n58501 );
not ( n59003 , n56310 );
or ( n59004 , n59002 , n59003 );
not ( n59005 , n57182 );
not ( n59006 , n52113 );
or ( n59007 , n59005 , n59006 );
nand ( n59008 , n52133 , n47332 );
nand ( n59009 , n59007 , n59008 );
nand ( n59010 , n59009 , n51766 );
nand ( n59011 , n59004 , n59010 );
xor ( n59012 , n59001 , n59011 );
not ( n59013 , n58511 );
not ( n59014 , n53182 );
or ( n59015 , n59013 , n59014 );
not ( n59016 , n48983 );
not ( n59017 , n55102 );
or ( n59018 , n59016 , n59017 );
nand ( n59019 , n58144 , n56348 );
nand ( n59020 , n59018 , n59019 );
nand ( n59021 , n52469 , n59020 );
nand ( n59022 , n59015 , n59021 );
xor ( n59023 , n59012 , n59022 );
xor ( n59024 , n58990 , n59023 );
xor ( n59025 , n58836 , n58989 );
and ( n59026 , n59025 , n59023 );
and ( n59027 , n58836 , n58989 );
or ( n59028 , n59026 , n59027 );
not ( n59029 , n58070 );
not ( n59030 , n58608 );
or ( n59031 , n59029 , n59030 );
not ( n59032 , n48898 );
not ( n59033 , n56285 );
or ( n59034 , n59032 , n59033 );
nand ( n59035 , n55845 , n48897 );
nand ( n59036 , n59034 , n59035 );
nand ( n59037 , n59036 , n55458 );
nand ( n59038 , n59031 , n59037 );
not ( n59039 , n58536 );
not ( n59040 , n56776 );
or ( n59041 , n59039 , n59040 );
not ( n59042 , n47227 );
not ( n59043 , n56759 );
or ( n59044 , n59042 , n59043 );
not ( n59045 , n56759 );
nand ( n59046 , n59045 , n47589 );
nand ( n59047 , n59044 , n59046 );
nand ( n59048 , n56780 , n59047 );
nand ( n59049 , n59041 , n59048 );
xor ( n59050 , n59038 , n59049 );
not ( n59051 , n58548 );
not ( n59052 , n57628 );
or ( n59053 , n59051 , n59052 );
and ( n59054 , n57533 , n47650 );
not ( n59055 , n57533 );
and ( n59056 , n59055 , n47646 );
or ( n59057 , n59054 , n59056 );
nand ( n59058 , n59057 , n57631 );
nand ( n59059 , n59053 , n59058 );
xor ( n59060 , n59050 , n59059 );
not ( n59061 , n58522 );
not ( n59062 , n55913 );
or ( n59063 , n59061 , n59062 );
not ( n59064 , n55511 );
not ( n59065 , n55917 );
or ( n59066 , n59064 , n59065 );
not ( n59067 , n53594 );
nand ( n59068 , n59067 , n51670 );
nand ( n59069 , n59066 , n59068 );
nand ( n59070 , n59069 , n54364 );
nand ( n59071 , n59063 , n59070 );
not ( n59072 , n58585 );
not ( n59073 , n56810 );
or ( n59074 , n59072 , n59073 );
not ( n59075 , n51792 );
not ( n59076 , n54467 );
or ( n59077 , n59075 , n59076 );
not ( n59078 , n54302 );
nand ( n59079 , n59078 , n48829 );
nand ( n59080 , n59077 , n59079 );
nand ( n59081 , n59080 , n54077 );
nand ( n59082 , n59074 , n59081 );
xor ( n59083 , n59071 , n59082 );
not ( n59084 , n58599 );
not ( n59085 , n55144 );
or ( n59086 , n59084 , n59085 );
not ( n59087 , n51204 );
not ( n59088 , n55119 );
or ( n59089 , n59087 , n59088 );
nand ( n59090 , n55118 , n48860 );
nand ( n59091 , n59089 , n59090 );
nand ( n59092 , n55157 , n59091 );
nand ( n59093 , n59086 , n59092 );
xor ( n59094 , n59083 , n59093 );
xor ( n59095 , n59060 , n59094 );
xor ( n59096 , n59095 , n58840 );
xor ( n59097 , n59060 , n59094 );
and ( n59098 , n59097 , n58840 );
and ( n59099 , n59060 , n59094 );
or ( n59100 , n59098 , n59099 );
xor ( n59101 , n58848 , n58844 );
xor ( n59102 , n59101 , n58852 );
xor ( n59103 , n58848 , n58844 );
and ( n59104 , n59103 , n58852 );
and ( n59105 , n58848 , n58844 );
or ( n59106 , n59104 , n59105 );
not ( n59107 , n47827 );
not ( n59108 , n50263 );
not ( n59109 , n56451 );
or ( n59110 , n59108 , n59109 );
nand ( n59111 , n40012 , n50087 );
nand ( n59112 , n59110 , n59111 );
not ( n59113 , n59112 );
or ( n59114 , n59107 , n59113 );
not ( n59115 , n58679 );
nand ( n59116 , n59115 , n48295 );
nand ( n59117 , n59114 , n59116 );
xor ( n59118 , n58887 , n59117 );
not ( n59119 , n47384 );
not ( n59120 , n49500 );
not ( n59121 , n56438 );
or ( n59122 , n59120 , n59121 );
nand ( n59123 , n40389 , n47979 );
nand ( n59124 , n59122 , n59123 );
not ( n59125 , n59124 );
or ( n59126 , n59119 , n59125 );
nand ( n59127 , n58745 , n49252 );
nand ( n59128 , n59126 , n59127 );
xor ( n59129 , n59118 , n59128 );
not ( n59130 , n47407 );
not ( n59131 , n58724 );
or ( n59132 , n59130 , n59131 );
not ( n59133 , n47803 );
not ( n59134 , n40451 );
not ( n59135 , n59134 );
or ( n59136 , n59133 , n59135 );
nand ( n59137 , n40451 , n50634 );
nand ( n59138 , n59136 , n59137 );
nand ( n59139 , n59138 , n48929 );
nand ( n59140 , n59132 , n59139 );
xor ( n59141 , n58439 , n59140 );
or ( n59142 , n58687 , n50241 );
xor ( n59143 , n52048 , n40376 );
or ( n59144 , n59143 , n50239 );
nand ( n59145 , n59142 , n59144 );
xor ( n59146 , n59141 , n59145 );
xor ( n59147 , n59129 , n59146 );
xor ( n59148 , n59147 , n58497 );
xor ( n59149 , n59129 , n59146 );
and ( n59150 , n59149 , n58497 );
and ( n59151 , n59129 , n59146 );
or ( n59152 , n59150 , n59151 );
not ( n59153 , n52421 );
not ( n59154 , n58696 );
or ( n59155 , n59153 , n59154 );
and ( n59156 , n40625 , n53228 );
not ( n59157 , n40625 );
and ( n59158 , n59157 , n51723 );
or ( n59159 , n59156 , n59158 );
nand ( n59160 , n59159 , n47148 );
nand ( n59161 , n59155 , n59160 );
not ( n59162 , n57314 );
not ( n59163 , n58715 );
or ( n59164 , n59162 , n59163 );
not ( n59165 , n52377 );
not ( n59166 , n54771 );
or ( n59167 , n59165 , n59166 );
nand ( n59168 , n40526 , n53973 );
nand ( n59169 , n59167 , n59168 );
nand ( n59170 , n59169 , n52004 );
nand ( n59171 , n59164 , n59170 );
xor ( n59172 , n59161 , n59171 );
not ( n59173 , n54623 );
not ( n59174 , n54628 );
not ( n59175 , n59174 );
buf ( n59176 , n51928 );
not ( n59177 , n59176 );
or ( n59178 , n59175 , n59177 );
buf ( n59179 , n58246 );
nand ( n59180 , n59179 , n51684 );
nand ( n59181 , n59178 , n59180 );
not ( n59182 , n59181 );
or ( n59183 , n59173 , n59182 );
nand ( n59184 , n58732 , n47873 );
nand ( n59185 , n59183 , n59184 );
xor ( n59186 , n59172 , n59185 );
xor ( n59187 , n59186 , n58579 );
not ( n59188 , n49713 );
not ( n59189 , n58666 );
or ( n59190 , n59188 , n59189 );
not ( n59191 , n52267 );
not ( n59192 , n54811 );
or ( n59193 , n59191 , n59192 );
not ( n59194 , n40363 );
not ( n59195 , n59194 );
nand ( n59196 , n59195 , n51351 );
nand ( n59197 , n59193 , n59196 );
nand ( n59198 , n59197 , n51865 );
nand ( n59199 , n59190 , n59198 );
not ( n59200 , n46564 );
not ( n59201 , n58757 );
or ( n59202 , n59200 , n59201 );
not ( n59203 , n47508 );
not ( n59204 , n58047 );
or ( n59205 , n59203 , n59204 );
nand ( n59206 , n39779 , n48955 );
nand ( n59207 , n59205 , n59206 );
nand ( n59208 , n59207 , n49832 );
nand ( n59209 , n59202 , n59208 );
xor ( n59210 , n59199 , n59209 );
xor ( n59211 , n59210 , n58794 );
xor ( n59212 , n59187 , n59211 );
xor ( n59213 , n59186 , n58579 );
and ( n59214 , n59213 , n59211 );
and ( n59215 , n59186 , n58579 );
or ( n59216 , n59214 , n59215 );
xor ( n59217 , n58940 , n58955 );
xor ( n59218 , n59217 , n59024 );
xor ( n59219 , n58940 , n58955 );
and ( n59220 , n59219 , n59024 );
and ( n59221 , n58940 , n58955 );
or ( n59222 , n59220 , n59221 );
xor ( n59223 , n58621 , n59096 );
xor ( n59224 , n59223 , n58653 );
xor ( n59225 , n58621 , n59096 );
and ( n59226 , n59225 , n58653 );
and ( n59227 , n58621 , n59096 );
or ( n59228 , n59226 , n59227 );
xor ( n59229 , n58708 , n59102 );
xor ( n59230 , n59229 , n58766 );
xor ( n59231 , n58708 , n59102 );
and ( n59232 , n59231 , n58766 );
and ( n59233 , n58708 , n59102 );
or ( n59234 , n59232 , n59233 );
xor ( n59235 , n59001 , n59011 );
and ( n59236 , n59235 , n59022 );
and ( n59237 , n59001 , n59011 );
or ( n59238 , n59236 , n59237 );
xor ( n59239 , n58772 , n59148 );
xor ( n59240 , n59239 , n58778 );
xor ( n59241 , n58772 , n59148 );
and ( n59242 , n59241 , n58778 );
and ( n59243 , n58772 , n59148 );
or ( n59244 , n59242 , n59243 );
xor ( n59245 , n59212 , n59218 );
xor ( n59246 , n59245 , n59224 );
xor ( n59247 , n59212 , n59218 );
and ( n59248 , n59247 , n59224 );
and ( n59249 , n59212 , n59218 );
or ( n59250 , n59248 , n59249 );
xor ( n59251 , n58784 , n59230 );
xor ( n59252 , n59251 , n58790 );
xor ( n59253 , n58784 , n59230 );
and ( n59254 , n59253 , n58790 );
and ( n59255 , n58784 , n59230 );
or ( n59256 , n59254 , n59255 );
xor ( n59257 , n59240 , n58800 );
xor ( n59258 , n59257 , n59246 );
xor ( n59259 , n59240 , n58800 );
and ( n59260 , n59259 , n59246 );
and ( n59261 , n59240 , n58800 );
or ( n59262 , n59260 , n59261 );
xor ( n59263 , n58806 , n59252 );
xor ( n59264 , n59263 , n58812 );
xor ( n59265 , n58806 , n59252 );
and ( n59266 , n59265 , n58812 );
and ( n59267 , n58806 , n59252 );
or ( n59268 , n59266 , n59267 );
xor ( n59269 , n59258 , n59264 );
xor ( n59270 , n59269 , n58818 );
xor ( n59271 , n59258 , n59264 );
and ( n59272 , n59271 , n58818 );
and ( n59273 , n59258 , n59264 );
or ( n59274 , n59272 , n59273 );
xor ( n59275 , n59071 , n59082 );
and ( n59276 , n59275 , n59093 );
and ( n59277 , n59071 , n59082 );
or ( n59278 , n59276 , n59277 );
xor ( n59279 , n59038 , n59049 );
and ( n59280 , n59279 , n59059 );
and ( n59281 , n59038 , n59049 );
or ( n59282 , n59280 , n59281 );
xor ( n59283 , n58973 , n58974 );
and ( n59284 , n59283 , n58988 );
and ( n59285 , n58973 , n58974 );
or ( n59286 , n59284 , n59285 );
xor ( n59287 , n58439 , n59140 );
and ( n59288 , n59287 , n59145 );
and ( n59289 , n58439 , n59140 );
or ( n59290 , n59288 , n59289 );
xor ( n59291 , n59161 , n59171 );
and ( n59292 , n59291 , n59185 );
and ( n59293 , n59161 , n59171 );
or ( n59294 , n59292 , n59293 );
xor ( n59295 , n58887 , n59117 );
and ( n59296 , n59295 , n59128 );
and ( n59297 , n58887 , n59117 );
or ( n59298 , n59296 , n59297 );
xor ( n59299 , n59199 , n59209 );
and ( n59300 , n59299 , n58794 );
and ( n59301 , n59199 , n59209 );
or ( n59302 , n59300 , n59301 );
not ( n59303 , n52736 );
not ( n59304 , n58897 );
or ( n59305 , n59303 , n59304 );
not ( n59306 , n49619 );
not ( n59307 , n49837 );
or ( n59308 , n59306 , n59307 );
nand ( n59309 , n57571 , n49766 );
nand ( n59310 , n59308 , n59309 );
nand ( n59311 , n59310 , n50078 );
nand ( n59312 , n59305 , n59311 );
not ( n59313 , n58433 );
not ( n59314 , n58902 );
nand ( n59315 , n59314 , n46440 );
not ( n59316 , n59315 );
or ( n59317 , n59313 , n59316 );
nand ( n59318 , n58902 , n46441 );
nand ( n59319 , n59317 , n59318 );
not ( n59320 , n36542 );
nand ( n59321 , n59320 , n36524 );
not ( n59322 , n59321 );
nand ( n59323 , n37528 , n36287 );
and ( n59324 , n37526 , n36307 );
not ( n59325 , n36328 );
not ( n59326 , n36316 );
or ( n59327 , n59325 , n59326 );
nand ( n59328 , n59327 , n36331 );
nor ( n59329 , n59324 , n59328 );
nand ( n59330 , n37662 , n59323 , n59329 );
not ( n59331 , n59330 );
or ( n59332 , n59322 , n59331 );
not ( n59333 , n59321 );
and ( n59334 , n59329 , n59333 );
nand ( n59335 , n59334 , n37662 , n59323 );
nand ( n59336 , n59332 , n59335 );
buf ( n59337 , n59336 );
buf ( n59338 , n59337 );
not ( n59339 , n59338 );
buf ( n59340 , n59339 );
not ( n59341 , n59340 );
and ( n59342 , n59319 , n59341 );
xor ( n59343 , n59312 , n59342 );
not ( n59344 , n56639 );
buf ( n59345 , n48705 );
not ( n59346 , n59345 );
not ( n59347 , n52076 );
or ( n59348 , n59346 , n59347 );
nand ( n59349 , n41132 , n51426 );
nand ( n59350 , n59348 , n59349 );
not ( n59351 , n59350 );
or ( n59352 , n59344 , n59351 );
nand ( n59353 , n58872 , n49309 );
nand ( n59354 , n59352 , n59353 );
xor ( n59355 , n59343 , n59354 );
xor ( n59356 , n59312 , n59342 );
and ( n59357 , n59356 , n59354 );
and ( n59358 , n59312 , n59342 );
or ( n59359 , n59357 , n59358 );
not ( n59360 , n58920 );
not ( n59361 , n50911 );
or ( n59362 , n59360 , n59361 );
not ( n59363 , n41532 );
not ( n59364 , n53904 );
or ( n59365 , n59363 , n59364 );
nand ( n59366 , n51461 , n49233 );
nand ( n59367 , n59365 , n59366 );
nand ( n59368 , n59367 , n50921 );
nand ( n59369 , n59362 , n59368 );
not ( n59370 , n58999 );
not ( n59371 , n52139 );
or ( n59372 , n59370 , n59371 );
not ( n59373 , n58454 );
not ( n59374 , n51566 );
or ( n59375 , n59373 , n59374 );
nand ( n59376 , n53549 , n58459 );
nand ( n59377 , n59375 , n59376 );
nand ( n59378 , n59377 , n51145 );
nand ( n59379 , n59372 , n59378 );
xor ( n59380 , n59369 , n59379 );
not ( n59381 , n59009 );
not ( n59382 , n52125 );
or ( n59383 , n59381 , n59382 );
not ( n59384 , n47527 );
not ( n59385 , n52109 );
or ( n59386 , n59384 , n59385 );
not ( n59387 , n52129 );
not ( n59388 , n47527 );
nand ( n59389 , n59387 , n59388 );
nand ( n59390 , n59386 , n59389 );
nand ( n59391 , n51766 , n59390 );
nand ( n59392 , n59383 , n59391 );
xor ( n59393 , n59380 , n59392 );
xor ( n59394 , n59369 , n59379 );
and ( n59395 , n59394 , n59392 );
and ( n59396 , n59369 , n59379 );
or ( n59397 , n59395 , n59396 );
not ( n59398 , n46602 );
not ( n59399 , n39574 );
and ( n59400 , n46072 , n59399 );
not ( n59401 , n46072 );
not ( n59402 , n39573 );
not ( n59403 , n59402 );
and ( n59404 , n59401 , n59403 );
or ( n59405 , n59400 , n59404 );
not ( n59406 , n59405 );
or ( n59407 , n59398 , n59406 );
nand ( n59408 , n58937 , n50659 );
nand ( n59409 , n59407 , n59408 );
xor ( n59410 , n59282 , n59409 );
not ( n59411 , n49026 );
not ( n59412 , n46425 );
not ( n59413 , n39893 );
not ( n59414 , n59413 );
not ( n59415 , n59414 );
or ( n59416 , n59412 , n59415 );
not ( n59417 , n39894 );
nand ( n59418 , n59417 , n46422 );
nand ( n59419 , n59416 , n59418 );
not ( n59420 , n59419 );
or ( n59421 , n59411 , n59420 );
not ( n59422 , n58951 );
nand ( n59423 , n59422 , n46267 );
nand ( n59424 , n59421 , n59423 );
xor ( n59425 , n59410 , n59424 );
xor ( n59426 , n59282 , n59409 );
and ( n59427 , n59426 , n59424 );
and ( n59428 , n59282 , n59409 );
or ( n59429 , n59427 , n59428 );
xor ( n59430 , n58927 , n59286 );
not ( n59431 , n59057 );
not ( n59432 , n57627 );
not ( n59433 , n59432 );
or ( n59434 , n59431 , n59433 );
not ( n59435 , n57138 );
not ( n59436 , n49734 );
not ( n59437 , n57613 );
not ( n59438 , n59437 );
or ( n59439 , n59436 , n59438 );
nand ( n59440 , n57614 , n47821 );
nand ( n59441 , n59439 , n59440 );
nand ( n59442 , n59435 , n59441 );
nand ( n59443 , n59434 , n59442 );
not ( n59444 , n58971 );
not ( n59445 , n58961 );
not ( n59446 , n59445 );
or ( n59447 , n59444 , n59446 );
and ( n59448 , n58642 , n46824 );
not ( n59449 , n58642 );
and ( n59450 , n59449 , n46273 );
or ( n59451 , n59448 , n59450 );
nand ( n59452 , n58638 , n59451 );
nand ( n59453 , n59447 , n59452 );
xor ( n59454 , n59443 , n59453 );
not ( n59455 , n51452 );
not ( n59456 , n50304 );
not ( n59457 , n48679 );
or ( n59458 , n59456 , n59457 );
nand ( n59459 , n41364 , n54614 );
nand ( n59460 , n59458 , n59459 );
not ( n59461 , n59460 );
or ( n59462 , n59455 , n59461 );
nand ( n59463 , n58859 , n50580 );
nand ( n59464 , n59462 , n59463 );
not ( n59465 , n52191 );
not ( n59466 , n49284 );
not ( n59467 , n49805 );
or ( n59468 , n59466 , n59467 );
nand ( n59469 , n57088 , n52916 );
nand ( n59470 , n59468 , n59469 );
not ( n59471 , n59470 );
or ( n59472 , n59465 , n59471 );
nand ( n59473 , n58881 , n51337 );
nand ( n59474 , n59472 , n59473 );
xor ( n59475 , n59464 , n59474 );
xor ( n59476 , n59454 , n59475 );
xor ( n59477 , n59430 , n59476 );
xor ( n59478 , n58927 , n59286 );
and ( n59479 , n59478 , n59476 );
and ( n59480 , n58927 , n59286 );
or ( n59481 , n59479 , n59480 );
not ( n59482 , n59091 );
not ( n59483 , n55143 );
or ( n59484 , n59482 , n59483 );
not ( n59485 , n49624 );
not ( n59486 , n58108 );
or ( n59487 , n59485 , n59486 );
nand ( n59488 , n55118 , n49630 );
nand ( n59489 , n59487 , n59488 );
nand ( n59490 , n54847 , n59489 );
nand ( n59491 , n59484 , n59490 );
not ( n59492 , n59036 );
not ( n59493 , n58070 );
or ( n59494 , n59492 , n59493 );
not ( n59495 , n47765 );
not ( n59496 , n55872 );
not ( n59497 , n59496 );
or ( n59498 , n59495 , n59497 );
not ( n59499 , n57676 );
nand ( n59500 , n59499 , n48589 );
nand ( n59501 , n59498 , n59500 );
nand ( n59502 , n59501 , n55458 );
nand ( n59503 , n59494 , n59502 );
xor ( n59504 , n59491 , n59503 );
not ( n59505 , n59047 );
not ( n59506 , n56776 );
or ( n59507 , n59505 , n59506 );
and ( n59508 , n56758 , n47368 );
not ( n59509 , n56758 );
and ( n59510 , n59509 , n52165 );
or ( n59511 , n59508 , n59510 );
nand ( n59512 , n56780 , n59511 );
nand ( n59513 , n59507 , n59512 );
xor ( n59514 , n59504 , n59513 );
xor ( n59515 , n59514 , n59393 );
not ( n59516 , n59020 );
not ( n59517 , n52852 );
or ( n59518 , n59516 , n59517 );
not ( n59519 , n47918 );
not ( n59520 , n52837 );
or ( n59521 , n59519 , n59520 );
nand ( n59522 , n58144 , n47510 );
nand ( n59523 , n59521 , n59522 );
nand ( n59524 , n59523 , n52468 );
nand ( n59525 , n59518 , n59524 );
not ( n59526 , n59069 );
not ( n59527 , n55913 );
or ( n59528 , n59526 , n59527 );
not ( n59529 , n41802 );
not ( n59530 , n55917 );
or ( n59531 , n59529 , n59530 );
nand ( n59532 , n53590 , n54184 );
nand ( n59533 , n59531 , n59532 );
nand ( n59534 , n59533 , n53619 );
nand ( n59535 , n59528 , n59534 );
xor ( n59536 , n59525 , n59535 );
not ( n59537 , n59080 );
not ( n59538 , n54315 );
or ( n59539 , n59537 , n59538 );
not ( n59540 , n52033 );
not ( n59541 , n54467 );
or ( n59542 , n59540 , n59541 );
nand ( n59543 , n54298 , n52038 );
nand ( n59544 , n59542 , n59543 );
nand ( n59545 , n59544 , n56277 );
nand ( n59546 , n59539 , n59545 );
xor ( n59547 , n59536 , n59546 );
xor ( n59548 , n59515 , n59547 );
xor ( n59549 , n59514 , n59393 );
and ( n59550 , n59549 , n59547 );
and ( n59551 , n59514 , n59393 );
or ( n59552 , n59550 , n59551 );
xor ( n59553 , n59290 , n59294 );
xor ( n59554 , n59553 , n59298 );
xor ( n59555 , n59290 , n59294 );
and ( n59556 , n59555 , n59298 );
and ( n59557 , n59290 , n59294 );
or ( n59558 , n59556 , n59557 );
not ( n59559 , n48689 );
not ( n59560 , n59339 );
or ( n59561 , n59559 , n59560 );
nand ( n59562 , n59338 , n46441 );
nand ( n59563 , n59561 , n59562 );
not ( n59564 , n59563 );
and ( n59565 , n59337 , n36337 );
not ( n59566 , n59337 );
and ( n59567 , n59566 , n58902 );
nor ( n59568 , n59565 , n59567 );
nand ( n59569 , n58906 , n59568 );
not ( n59570 , n59569 );
buf ( n59571 , n59570 );
not ( n59572 , n59571 );
or ( n59573 , n59564 , n59572 );
buf ( n59574 , n58907 );
not ( n59575 , n59574 );
not ( n59576 , n50914 );
not ( n59577 , n59336 );
buf ( n59578 , n59577 );
not ( n59579 , n59578 );
or ( n59580 , n59576 , n59579 );
nand ( n59581 , n59338 , n48766 );
nand ( n59582 , n59580 , n59581 );
nand ( n59583 , n59575 , n59582 );
nand ( n59584 , n59573 , n59583 );
xor ( n59585 , n59584 , n58891 );
xor ( n59586 , n59585 , n59355 );
not ( n59587 , n48929 );
not ( n59588 , n47803 );
not ( n59589 , n56975 );
or ( n59590 , n59588 , n59589 );
nand ( n59591 , n40512 , n50634 );
nand ( n59592 , n59590 , n59591 );
not ( n59593 , n59592 );
or ( n59594 , n59587 , n59593 );
nand ( n59595 , n59138 , n47407 );
nand ( n59596 , n59594 , n59595 );
not ( n59597 , n52043 );
not ( n59598 , n48645 );
not ( n59599 , n56074 );
or ( n59600 , n59598 , n59599 );
not ( n59601 , n40225 );
nand ( n59602 , n59601 , n49679 );
nand ( n59603 , n59600 , n59602 );
not ( n59604 , n59603 );
or ( n59605 , n59597 , n59604 );
not ( n59606 , n59143 );
nand ( n59607 , n59606 , n50242 );
nand ( n59608 , n59605 , n59607 );
xor ( n59609 , n59596 , n59608 );
not ( n59610 , n54875 );
not ( n59611 , n40635 );
not ( n59612 , n59611 );
not ( n59613 , n59612 );
not ( n59614 , n53228 );
or ( n59615 , n59613 , n59614 );
nand ( n59616 , n54415 , n51723 );
nand ( n59617 , n59615 , n59616 );
not ( n59618 , n59617 );
or ( n59619 , n59610 , n59618 );
nand ( n59620 , n59159 , n52421 );
nand ( n59621 , n59619 , n59620 );
xor ( n59622 , n59609 , n59621 );
xor ( n59623 , n59586 , n59622 );
not ( n59624 , n58982 );
not ( n59625 , n51573 );
or ( n59626 , n59624 , n59625 );
nand ( n59627 , n40677 , n52728 );
nand ( n59628 , n59626 , n59627 );
not ( n59629 , n59628 );
buf ( n59630 , n52722 );
or ( n59631 , n59629 , n59630 );
not ( n59632 , n50176 );
not ( n59633 , n59632 );
nand ( n59634 , n58984 , n59633 );
nand ( n59635 , n59631 , n59634 );
not ( n59636 , n49713 );
not ( n59637 , n59197 );
or ( n59638 , n59636 , n59637 );
not ( n59639 , n52267 );
not ( n59640 , n56011 );
or ( n59641 , n59639 , n59640 );
nand ( n59642 , n54406 , n51351 );
nand ( n59643 , n59641 , n59642 );
nand ( n59644 , n59643 , n51865 );
nand ( n59645 , n59638 , n59644 );
xor ( n59646 , n59635 , n59645 );
not ( n59647 , n51157 );
not ( n59648 , n59112 );
or ( n59649 , n59647 , n59648 );
not ( n59650 , n50263 );
buf ( n59651 , n56962 );
not ( n59652 , n59651 );
or ( n59653 , n59650 , n59652 );
buf ( n59654 , n57801 );
nand ( n59655 , n59654 , n52080 );
nand ( n59656 , n59653 , n59655 );
nand ( n59657 , n59656 , n47827 );
nand ( n59658 , n59649 , n59657 );
xor ( n59659 , n59646 , n59658 );
xor ( n59660 , n59623 , n59659 );
xor ( n59661 , n59586 , n59622 );
and ( n59662 , n59661 , n59659 );
and ( n59663 , n59586 , n59622 );
or ( n59664 , n59662 , n59663 );
xor ( n59665 , n58944 , n58959 );
xor ( n59666 , n59665 , n59302 );
xor ( n59667 , n58944 , n58959 );
and ( n59668 , n59667 , n59302 );
and ( n59669 , n58944 , n58959 );
or ( n59670 , n59668 , n59669 );
not ( n59671 , n48894 );
not ( n59672 , n59169 );
or ( n59673 , n59671 , n59672 );
not ( n59674 , n40591 );
not ( n59675 , n53973 );
and ( n59676 , n59674 , n59675 );
and ( n59677 , n52212 , n53973 );
nor ( n59678 , n59676 , n59677 );
or ( n59679 , n59678 , n56523 );
nand ( n59680 , n59673 , n59679 );
not ( n59681 , n54623 );
not ( n59682 , n54625 );
not ( n59683 , n52894 );
or ( n59684 , n59682 , n59683 );
nand ( n59685 , n51601 , n54628 );
nand ( n59686 , n59684 , n59685 );
not ( n59687 , n59686 );
or ( n59688 , n59681 , n59687 );
nand ( n59689 , n59181 , n47873 );
nand ( n59690 , n59688 , n59689 );
xor ( n59691 , n59680 , n59690 );
not ( n59692 , n47384 );
not ( n59693 , n49500 );
buf ( n59694 , n55202 );
not ( n59695 , n59694 );
or ( n59696 , n59693 , n59695 );
not ( n59697 , n55199 );
nand ( n59698 , n59697 , n53997 );
nand ( n59699 , n59696 , n59698 );
not ( n59700 , n59699 );
or ( n59701 , n59692 , n59700 );
nand ( n59702 , n59124 , n48989 );
nand ( n59703 , n59701 , n59702 );
xor ( n59704 , n59691 , n59703 );
xor ( n59705 , n59704 , n59028 );
not ( n59706 , n49832 );
not ( n59707 , n48952 );
not ( n59708 , n58482 );
or ( n59709 , n59707 , n59708 );
nand ( n59710 , n39680 , n47514 );
nand ( n59711 , n59709 , n59710 );
not ( n59712 , n59711 );
or ( n59713 , n59706 , n59712 );
nand ( n59714 , n59207 , n46564 );
nand ( n59715 , n59713 , n59714 );
xor ( n59716 , n59715 , n59238 );
xor ( n59717 , n59716 , n59278 );
xor ( n59718 , n59705 , n59717 );
xor ( n59719 , n59704 , n59028 );
and ( n59720 , n59719 , n59717 );
and ( n59721 , n59704 , n59028 );
or ( n59722 , n59720 , n59721 );
xor ( n59723 , n59425 , n59100 );
xor ( n59724 , n59723 , n59548 );
xor ( n59725 , n59425 , n59100 );
and ( n59726 , n59725 , n59548 );
and ( n59727 , n59425 , n59100 );
or ( n59728 , n59726 , n59727 );
xor ( n59729 , n59477 , n59554 );
xor ( n59730 , n59729 , n59152 );
xor ( n59731 , n59477 , n59554 );
and ( n59732 , n59731 , n59152 );
and ( n59733 , n59477 , n59554 );
or ( n59734 , n59732 , n59733 );
xor ( n59735 , n59106 , n59216 );
xor ( n59736 , n59735 , n59660 );
xor ( n59737 , n59106 , n59216 );
and ( n59738 , n59737 , n59660 );
and ( n59739 , n59106 , n59216 );
or ( n59740 , n59738 , n59739 );
xor ( n59741 , n59525 , n59535 );
and ( n59742 , n59741 , n59546 );
and ( n59743 , n59525 , n59535 );
or ( n59744 , n59742 , n59743 );
xor ( n59745 , n59666 , n59222 );
xor ( n59746 , n59745 , n59718 );
xor ( n59747 , n59666 , n59222 );
and ( n59748 , n59747 , n59718 );
and ( n59749 , n59666 , n59222 );
or ( n59750 , n59748 , n59749 );
xor ( n59751 , n59228 , n59724 );
xor ( n59752 , n59751 , n59730 );
xor ( n59753 , n59228 , n59724 );
and ( n59754 , n59753 , n59730 );
and ( n59755 , n59228 , n59724 );
or ( n59756 , n59754 , n59755 );
xor ( n59757 , n59234 , n59736 );
xor ( n59758 , n59757 , n59244 );
xor ( n59759 , n59234 , n59736 );
and ( n59760 , n59759 , n59244 );
and ( n59761 , n59234 , n59736 );
or ( n59762 , n59760 , n59761 );
xor ( n59763 , n59746 , n59250 );
xor ( n59764 , n59763 , n59752 );
xor ( n59765 , n59746 , n59250 );
and ( n59766 , n59765 , n59752 );
and ( n59767 , n59746 , n59250 );
or ( n59768 , n59766 , n59767 );
xor ( n59769 , n59256 , n59758 );
xor ( n59770 , n59769 , n59262 );
xor ( n59771 , n59256 , n59758 );
and ( n59772 , n59771 , n59262 );
and ( n59773 , n59256 , n59758 );
or ( n59774 , n59772 , n59773 );
xor ( n59775 , n59764 , n59268 );
xor ( n59776 , n59775 , n59770 );
xor ( n59777 , n59764 , n59268 );
and ( n59778 , n59777 , n59770 );
and ( n59779 , n59764 , n59268 );
or ( n59780 , n59778 , n59779 );
xor ( n59781 , n59491 , n59503 );
and ( n59782 , n59781 , n59513 );
and ( n59783 , n59491 , n59503 );
or ( n59784 , n59782 , n59783 );
xor ( n59785 , n59443 , n59453 );
and ( n59786 , n59785 , n59475 );
and ( n59787 , n59443 , n59453 );
or ( n59788 , n59786 , n59787 );
xor ( n59789 , n59584 , n58891 );
and ( n59790 , n59789 , n59355 );
and ( n59791 , n59584 , n58891 );
or ( n59792 , n59790 , n59791 );
xor ( n59793 , n59596 , n59608 );
and ( n59794 , n59793 , n59621 );
and ( n59795 , n59596 , n59608 );
or ( n59796 , n59794 , n59795 );
xor ( n59797 , n59680 , n59690 );
and ( n59798 , n59797 , n59703 );
and ( n59799 , n59680 , n59690 );
or ( n59800 , n59798 , n59799 );
xor ( n59801 , n59635 , n59645 );
and ( n59802 , n59801 , n59658 );
and ( n59803 , n59635 , n59645 );
or ( n59804 , n59802 , n59803 );
xor ( n59805 , n59715 , n59238 );
and ( n59806 , n59805 , n59278 );
and ( n59807 , n59715 , n59238 );
or ( n59808 , n59806 , n59807 );
not ( n59809 , n59470 );
or ( n59810 , n59809 , n57585 );
not ( n59811 , n52191 );
not ( n59812 , n41036 );
not ( n59813 , n49259 );
and ( n59814 , n59812 , n59813 );
and ( n59815 , n51891 , n49283 );
nor ( n59816 , n59814 , n59815 );
or ( n59817 , n59811 , n59816 );
nand ( n59818 , n59810 , n59817 );
not ( n59819 , n59460 );
not ( n59820 , n52749 );
or ( n59821 , n59819 , n59820 );
not ( n59822 , n51250 );
not ( n59823 , n41285 );
or ( n59824 , n59822 , n59823 );
nand ( n59825 , n50327 , n48996 );
nand ( n59826 , n59824 , n59825 );
not ( n59827 , n59826 );
not ( n59828 , n52757 );
or ( n59829 , n59827 , n59828 );
nand ( n59830 , n59821 , n59829 );
xor ( n59831 , n59818 , n59830 );
not ( n59832 , n50078 );
not ( n59833 , n49619 );
not ( n59834 , n54870 );
or ( n59835 , n59833 , n59834 );
nand ( n59836 , n40854 , n49766 );
nand ( n59837 , n59835 , n59836 );
not ( n59838 , n59837 );
or ( n59839 , n59832 , n59838 );
nand ( n59840 , n59310 , n52058 );
nand ( n59841 , n59839 , n59840 );
xor ( n59842 , n59831 , n59841 );
xor ( n59843 , n59818 , n59830 );
and ( n59844 , n59843 , n59841 );
and ( n59845 , n59818 , n59830 );
or ( n59846 , n59844 , n59845 );
not ( n59847 , n37569 );
not ( n59848 , n59847 );
not ( n59849 , n36549 );
not ( n59850 , n59849 );
or ( n59851 , n59848 , n59850 );
nand ( n59852 , n36549 , n37569 );
nand ( n59853 , n59851 , n59852 );
xor ( n59854 , n59577 , n59853 );
not ( n59855 , n59854 );
and ( n59856 , n59855 , n48689 );
not ( n59857 , n59367 );
not ( n59858 , n52526 );
or ( n59859 , n59857 , n59858 );
not ( n59860 , n48486 );
not ( n59861 , n50916 );
or ( n59862 , n59860 , n59861 );
nand ( n59863 , n51461 , n48951 );
nand ( n59864 , n59862 , n59863 );
nand ( n59865 , n59864 , n50921 );
nand ( n59866 , n59859 , n59865 );
xor ( n59867 , n59856 , n59866 );
not ( n59868 , n59377 );
not ( n59869 , n52139 );
or ( n59870 , n59868 , n59869 );
not ( n59871 , n41668 );
not ( n59872 , n51566 );
or ( n59873 , n59871 , n59872 );
nand ( n59874 , n56361 , n58914 );
nand ( n59875 , n59873 , n59874 );
nand ( n59876 , n51145 , n59875 );
nand ( n59877 , n59870 , n59876 );
xor ( n59878 , n59867 , n59877 );
xor ( n59879 , n59856 , n59866 );
and ( n59880 , n59879 , n59877 );
and ( n59881 , n59856 , n59866 );
or ( n59882 , n59880 , n59881 );
xor ( n59883 , n59744 , n59784 );
xor ( n59884 , n59883 , n59788 );
xor ( n59885 , n59744 , n59784 );
and ( n59886 , n59885 , n59788 );
and ( n59887 , n59744 , n59784 );
or ( n59888 , n59886 , n59887 );
not ( n59889 , n44004 );
not ( n59890 , n46072 );
not ( n59891 , n39055 );
not ( n59892 , n59891 );
or ( n59893 , n59890 , n59892 );
nand ( n59894 , n39055 , n50405 );
nand ( n59895 , n59893 , n59894 );
not ( n59896 , n59895 );
or ( n59897 , n59889 , n59896 );
nand ( n59898 , n59405 , n50659 );
nand ( n59899 , n59897 , n59898 );
not ( n59900 , n49832 );
not ( n59901 , n48952 );
not ( n59902 , n39715 );
or ( n59903 , n59901 , n59902 );
nand ( n59904 , n39714 , n47514 );
nand ( n59905 , n59903 , n59904 );
not ( n59906 , n59905 );
or ( n59907 , n59900 , n59906 );
nand ( n59908 , n59711 , n46564 );
nand ( n59909 , n59907 , n59908 );
xor ( n59910 , n59899 , n59909 );
not ( n59911 , n49026 );
not ( n59912 , n46425 );
buf ( n59913 , n39779 );
not ( n59914 , n59913 );
not ( n59915 , n59914 );
or ( n59916 , n59912 , n59915 );
nand ( n59917 , n59913 , n46422 );
nand ( n59918 , n59916 , n59917 );
not ( n59919 , n59918 );
or ( n59920 , n59911 , n59919 );
nand ( n59921 , n59419 , n46267 );
nand ( n59922 , n59920 , n59921 );
xor ( n59923 , n59910 , n59922 );
xor ( n59924 , n59899 , n59909 );
and ( n59925 , n59924 , n59922 );
and ( n59926 , n59899 , n59909 );
or ( n59927 , n59925 , n59926 );
not ( n59928 , n59582 );
not ( n59929 , n59570 );
or ( n59930 , n59928 , n59929 );
not ( n59931 , n58907 );
not ( n59932 , n46037 );
not ( n59933 , n59339 );
or ( n59934 , n59932 , n59933 );
not ( n59935 , n59578 );
nand ( n59936 , n59935 , n54721 );
nand ( n59937 , n59934 , n59936 );
nand ( n59938 , n59931 , n59937 );
nand ( n59939 , n59930 , n59938 );
and ( n59940 , n59474 , n59464 );
xor ( n59941 , n59939 , n59940 );
not ( n59942 , n56639 );
not ( n59943 , n59345 );
not ( n59944 , n57307 );
or ( n59945 , n59943 , n59944 );
nand ( n59946 , n40691 , n51426 );
nand ( n59947 , n59945 , n59946 );
not ( n59948 , n59947 );
or ( n59949 , n59942 , n59948 );
buf ( n59950 , n49309 );
nand ( n59951 , n59350 , n59950 );
nand ( n59952 , n59949 , n59951 );
xor ( n59953 , n59941 , n59952 );
xor ( n59954 , n59953 , n59878 );
not ( n59955 , n59544 );
not ( n59956 , n54315 );
or ( n59957 , n59955 , n59956 );
not ( n59958 , n54611 );
not ( n59959 , n54467 );
or ( n59960 , n59958 , n59959 );
nand ( n59961 , n54298 , n51670 );
nand ( n59962 , n59960 , n59961 );
nand ( n59963 , n59962 , n54077 );
nand ( n59964 , n59957 , n59963 );
not ( n59965 , n59489 );
not ( n59966 , n55143 );
or ( n59967 , n59965 , n59966 );
not ( n59968 , n51792 );
not ( n59969 , n55148 );
or ( n59970 , n59968 , n59969 );
nand ( n59971 , n55152 , n48829 );
nand ( n59972 , n59970 , n59971 );
nand ( n59973 , n59972 , n54848 );
nand ( n59974 , n59967 , n59973 );
xor ( n59975 , n59964 , n59974 );
not ( n59976 , n55887 );
not ( n59977 , n59501 );
or ( n59978 , n59976 , n59977 );
not ( n59979 , n51204 );
not ( n59980 , n55876 );
or ( n59981 , n59979 , n59980 );
nand ( n59982 , n55872 , n48860 );
nand ( n59983 , n59981 , n59982 );
buf ( n59984 , n55457 );
nand ( n59985 , n59983 , n59984 );
nand ( n59986 , n59978 , n59985 );
xor ( n59987 , n59975 , n59986 );
xor ( n59988 , n59954 , n59987 );
xor ( n59989 , n59953 , n59878 );
and ( n59990 , n59989 , n59987 );
and ( n59991 , n59953 , n59878 );
or ( n59992 , n59990 , n59991 );
not ( n59993 , n59390 );
not ( n59994 , n54265 );
or ( n59995 , n59993 , n59994 );
not ( n59996 , n52379 );
not ( n59997 , n52113 );
or ( n59998 , n59996 , n59997 );
not ( n59999 , n52113 );
nand ( n60000 , n59999 , n41416 );
nand ( n60001 , n59998 , n60000 );
nand ( n60002 , n60001 , n51765 );
nand ( n60003 , n59995 , n60002 );
not ( n60004 , n59523 );
not ( n60005 , n52853 );
or ( n60006 , n60004 , n60005 );
not ( n60007 , n57182 );
not ( n60008 , n55102 );
or ( n60009 , n60007 , n60008 );
not ( n60010 , n52837 );
nand ( n60011 , n60010 , n47332 );
nand ( n60012 , n60009 , n60011 );
nand ( n60013 , n60012 , n53571 );
nand ( n60014 , n60006 , n60013 );
xor ( n60015 , n60003 , n60014 );
not ( n60016 , n55913 );
not ( n60017 , n59533 );
or ( n60018 , n60016 , n60017 );
xor ( n60019 , n53590 , n56348 );
or ( n60020 , n60019 , n53618 );
nand ( n60021 , n60018 , n60020 );
xor ( n60022 , n60015 , n60021 );
not ( n60023 , n59511 );
not ( n60024 , n58529 );
or ( n60025 , n60023 , n60024 );
not ( n60026 , n48898 );
not ( n60027 , n56784 );
or ( n60028 , n60026 , n60027 );
nand ( n60029 , n56757 , n48897 );
nand ( n60030 , n60028 , n60029 );
nand ( n60031 , n56500 , n60030 );
nand ( n60032 , n60025 , n60031 );
not ( n60033 , n59441 );
not ( n60034 , n58541 );
or ( n60035 , n60033 , n60034 );
not ( n60036 , n47227 );
not ( n60037 , n57633 );
or ( n60038 , n60036 , n60037 );
nand ( n60039 , n57614 , n47589 );
nand ( n60040 , n60038 , n60039 );
nand ( n60041 , n60040 , n57139 );
nand ( n60042 , n60035 , n60041 );
xor ( n60043 , n60032 , n60042 );
not ( n60044 , n59451 );
not ( n60045 , n59445 );
or ( n60046 , n60044 , n60045 );
and ( n60047 , n58642 , n47650 );
not ( n60048 , n58642 );
and ( n60049 , n60048 , n47646 );
or ( n60050 , n60047 , n60049 );
nand ( n60051 , n58638 , n60050 );
nand ( n60052 , n60046 , n60051 );
xor ( n60053 , n60043 , n60052 );
xor ( n60054 , n60022 , n60053 );
xor ( n60055 , n60054 , n59796 );
xor ( n60056 , n60022 , n60053 );
and ( n60057 , n60056 , n59796 );
and ( n60058 , n60022 , n60053 );
or ( n60059 , n60057 , n60058 );
xor ( n60060 , n59792 , n59800 );
xor ( n60061 , n60060 , n59804 );
xor ( n60062 , n59792 , n59800 );
and ( n60063 , n60062 , n59804 );
and ( n60064 , n59792 , n59800 );
or ( n60065 , n60063 , n60064 );
not ( n60066 , n53104 );
not ( n60067 , n59628 );
or ( n60068 , n60066 , n60067 );
not ( n60069 , n58982 );
not ( n60070 , n40733 );
or ( n60071 , n60069 , n60070 );
nand ( n60072 , n51929 , n52728 );
nand ( n60073 , n60071 , n60072 );
nand ( n60074 , n60073 , n52723 );
nand ( n60075 , n60068 , n60074 );
not ( n60076 , n49713 );
not ( n60077 , n59643 );
or ( n60078 , n60076 , n60077 );
not ( n60079 , n52267 );
not ( n60080 , n55641 );
or ( n60081 , n60079 , n60080 );
nand ( n60082 , n55645 , n51351 );
nand ( n60083 , n60081 , n60082 );
nand ( n60084 , n60083 , n51865 );
nand ( n60085 , n60078 , n60084 );
xor ( n60086 , n60075 , n60085 );
not ( n60087 , n53675 );
and ( n60088 , n56454 , n54028 );
not ( n60089 , n56454 );
and ( n60090 , n60089 , n48727 );
or ( n60091 , n60088 , n60090 );
not ( n60092 , n60091 );
or ( n60093 , n60087 , n60092 );
nand ( n60094 , n59592 , n47407 );
nand ( n60095 , n60093 , n60094 );
xor ( n60096 , n60086 , n60095 );
xor ( n60097 , n60096 , n59808 );
xor ( n60098 , n60097 , n59429 );
xor ( n60099 , n60096 , n59808 );
and ( n60100 , n60099 , n59429 );
and ( n60101 , n60096 , n59808 );
or ( n60102 , n60100 , n60101 );
not ( n60103 , n52962 );
not ( n60104 , n50232 );
not ( n60105 , n54811 );
or ( n60106 , n60104 , n60105 );
nand ( n60107 , n40364 , n52048 );
nand ( n60108 , n60106 , n60107 );
not ( n60109 , n60108 );
or ( n60110 , n60103 , n60109 );
nand ( n60111 , n59603 , n52970 );
nand ( n60112 , n60110 , n60111 );
not ( n60113 , n51368 );
not ( n60114 , n59617 );
or ( n60115 , n60113 , n60114 );
not ( n60116 , n48856 );
not ( n60117 , n53289 );
or ( n60118 , n60116 , n60117 );
nand ( n60119 , n40376 , n53228 );
nand ( n60120 , n60118 , n60119 );
nand ( n60121 , n60120 , n54875 );
nand ( n60122 , n60115 , n60121 );
xor ( n60123 , n60112 , n60122 );
xor ( n60124 , n60123 , n59842 );
not ( n60125 , n52004 );
not ( n60126 , n52377 );
not ( n60127 , n53271 );
or ( n60128 , n60126 , n60127 );
nand ( n60129 , n40626 , n55013 );
nand ( n60130 , n60128 , n60129 );
not ( n60131 , n60130 );
or ( n60132 , n60125 , n60131 );
not ( n60133 , n59678 );
nand ( n60134 , n60133 , n57314 );
nand ( n60135 , n60132 , n60134 );
not ( n60136 , n54623 );
not ( n60137 , n54625 );
not ( n60138 , n51916 );
not ( n60139 , n60138 );
or ( n60140 , n60137 , n60139 );
nand ( n60141 , n51912 , n54628 );
nand ( n60142 , n60140 , n60141 );
not ( n60143 , n60142 );
or ( n60144 , n60136 , n60143 );
nand ( n60145 , n59686 , n47873 );
nand ( n60146 , n60144 , n60145 );
xor ( n60147 , n60135 , n60146 );
not ( n60148 , n49252 );
not ( n60149 , n59699 );
or ( n60150 , n60148 , n60149 );
not ( n60151 , n49500 );
not ( n60152 , n55630 );
or ( n60153 , n60151 , n60152 );
nand ( n60154 , n40452 , n47979 );
nand ( n60155 , n60153 , n60154 );
nand ( n60156 , n60155 , n47384 );
nand ( n60157 , n60150 , n60156 );
xor ( n60158 , n60147 , n60157 );
xor ( n60159 , n60124 , n60158 );
xor ( n60160 , n60159 , n59481 );
xor ( n60161 , n60124 , n60158 );
and ( n60162 , n60161 , n59481 );
and ( n60163 , n60124 , n60158 );
or ( n60164 , n60162 , n60163 );
not ( n60165 , n47827 );
not ( n60166 , n46650 );
not ( n60167 , n39845 );
not ( n60168 , n60167 );
or ( n60169 , n60166 , n60168 );
nand ( n60170 , n58034 , n48078 );
nand ( n60171 , n60169 , n60170 );
not ( n60172 , n60171 );
or ( n60173 , n60165 , n60172 );
nand ( n60174 , n59656 , n46776 );
nand ( n60175 , n60173 , n60174 );
xor ( n60176 , n59359 , n60175 );
xor ( n60177 , n60176 , n59397 );
xor ( n60178 , n59884 , n60177 );
xor ( n60179 , n60178 , n59923 );
xor ( n60180 , n59884 , n60177 );
and ( n60181 , n60180 , n59923 );
and ( n60182 , n59884 , n60177 );
or ( n60183 , n60181 , n60182 );
xor ( n60184 , n59552 , n59558 );
xor ( n60185 , n60184 , n60055 );
xor ( n60186 , n59552 , n59558 );
and ( n60187 , n60186 , n60055 );
and ( n60188 , n59552 , n59558 );
or ( n60189 , n60187 , n60188 );
xor ( n60190 , n59988 , n59670 );
xor ( n60191 , n60190 , n60061 );
xor ( n60192 , n59988 , n59670 );
and ( n60193 , n60192 , n60061 );
and ( n60194 , n59988 , n59670 );
or ( n60195 , n60193 , n60194 );
xor ( n60196 , n60003 , n60014 );
and ( n60197 , n60196 , n60021 );
and ( n60198 , n60003 , n60014 );
or ( n60199 , n60197 , n60198 );
xor ( n60200 , n59664 , n59722 );
xor ( n60201 , n60200 , n60160 );
xor ( n60202 , n59664 , n59722 );
and ( n60203 , n60202 , n60160 );
and ( n60204 , n59664 , n59722 );
or ( n60205 , n60203 , n60204 );
xor ( n60206 , n60098 , n59728 );
xor ( n60207 , n60206 , n60179 );
xor ( n60208 , n60098 , n59728 );
and ( n60209 , n60208 , n60179 );
and ( n60210 , n60098 , n59728 );
or ( n60211 , n60209 , n60210 );
xor ( n60212 , n60185 , n59734 );
xor ( n60213 , n60212 , n59740 );
xor ( n60214 , n60185 , n59734 );
and ( n60215 , n60214 , n59740 );
and ( n60216 , n60185 , n59734 );
or ( n60217 , n60215 , n60216 );
xor ( n60218 , n60191 , n60201 );
xor ( n60219 , n60218 , n59750 );
xor ( n60220 , n60191 , n60201 );
and ( n60221 , n60220 , n59750 );
and ( n60222 , n60191 , n60201 );
or ( n60223 , n60221 , n60222 );
xor ( n60224 , n60207 , n60213 );
xor ( n60225 , n60224 , n59756 );
xor ( n60226 , n60207 , n60213 );
and ( n60227 , n60226 , n59756 );
and ( n60228 , n60207 , n60213 );
or ( n60229 , n60227 , n60228 );
xor ( n60230 , n59762 , n60219 );
xor ( n60231 , n60230 , n59768 );
xor ( n60232 , n59762 , n60219 );
and ( n60233 , n60232 , n59768 );
and ( n60234 , n59762 , n60219 );
or ( n60235 , n60233 , n60234 );
xor ( n60236 , n60225 , n59774 );
xor ( n60237 , n60236 , n60231 );
xor ( n60238 , n60225 , n59774 );
and ( n60239 , n60238 , n60231 );
and ( n60240 , n60225 , n59774 );
or ( n60241 , n60239 , n60240 );
xor ( n60242 , n59964 , n59974 );
and ( n60243 , n60242 , n59986 );
and ( n60244 , n59964 , n59974 );
or ( n60245 , n60243 , n60244 );
xor ( n60246 , n60032 , n60042 );
and ( n60247 , n60246 , n60052 );
and ( n60248 , n60032 , n60042 );
or ( n60249 , n60247 , n60248 );
xor ( n60250 , n59939 , n59940 );
and ( n60251 , n60250 , n59952 );
and ( n60252 , n59939 , n59940 );
or ( n60253 , n60251 , n60252 );
xor ( n60254 , n60112 , n60122 );
and ( n60255 , n60254 , n59842 );
and ( n60256 , n60112 , n60122 );
or ( n60257 , n60255 , n60256 );
xor ( n60258 , n60135 , n60146 );
and ( n60259 , n60258 , n60157 );
and ( n60260 , n60135 , n60146 );
or ( n60261 , n60259 , n60260 );
xor ( n60262 , n60075 , n60085 );
and ( n60263 , n60262 , n60095 );
and ( n60264 , n60075 , n60085 );
or ( n60265 , n60263 , n60264 );
xor ( n60266 , n59359 , n60175 );
and ( n60267 , n60266 , n59397 );
and ( n60268 , n59359 , n60175 );
or ( n60269 , n60267 , n60268 );
not ( n60270 , n59338 );
not ( n60271 , n59847 );
not ( n60272 , n59849 );
or ( n60273 , n60271 , n60272 );
nand ( n60274 , n60273 , n59852 );
buf ( n60275 , n60274 );
nand ( n60276 , n60275 , n46440 );
nand ( n60277 , n60270 , n60276 );
not ( n60278 , n60275 );
nand ( n60279 , n60278 , n46441 );
and ( n60280 , n60277 , n60279 );
and ( n60281 , n36913 , n37408 );
nand ( n60282 , n37524 , n57117 );
nand ( n60283 , n60282 , n37066 , n37418 );
xor ( n60284 , n60281 , n60283 );
buf ( n60285 , n60284 );
not ( n60286 , n60285 );
nor ( n60287 , n60280 , n60286 );
not ( n60288 , n54249 );
not ( n60289 , n49112 );
not ( n60290 , n60289 );
and ( n60291 , n60288 , n60290 );
not ( n60292 , n49112 );
and ( n60293 , n41132 , n60292 );
nor ( n60294 , n60291 , n60293 );
not ( n60295 , n49288 );
or ( n60296 , n60294 , n60295 );
not ( n60297 , n59816 );
nand ( n60298 , n60297 , n57586 );
nand ( n60299 , n60296 , n60298 );
xor ( n60300 , n60287 , n60299 );
not ( n60301 , n59864 );
or ( n60302 , n50910 , n60301 );
and ( n60303 , n41363 , n50894 );
not ( n60304 , n41363 );
and ( n60305 , n60304 , n50907 );
or ( n60306 , n60303 , n60305 );
not ( n60307 , n60306 );
or ( n60308 , n60307 , n50626 );
nand ( n60309 , n60302 , n60308 );
xor ( n60310 , n60300 , n60309 );
xor ( n60311 , n60287 , n60299 );
and ( n60312 , n60311 , n60309 );
and ( n60313 , n60287 , n60299 );
or ( n60314 , n60312 , n60313 );
not ( n60315 , n59875 );
not ( n60316 , n51525 );
or ( n60317 , n60315 , n60316 );
not ( n60318 , n41531 );
not ( n60319 , n51504 );
or ( n60320 , n60318 , n60319 );
not ( n60321 , n51565 );
nand ( n60322 , n60321 , n49233 );
nand ( n60323 , n60320 , n60322 );
nand ( n60324 , n51145 , n60323 );
nand ( n60325 , n60317 , n60324 );
not ( n60326 , n60001 );
not ( n60327 , n56310 );
or ( n60328 , n60326 , n60327 );
not ( n60329 , n49756 );
not ( n60330 , n60329 );
not ( n60331 , n52130 );
or ( n60332 , n60330 , n60331 );
nand ( n60333 , n53917 , n58453 );
nand ( n60334 , n60332 , n60333 );
nand ( n60335 , n51766 , n60334 );
nand ( n60336 , n60328 , n60335 );
xor ( n60337 , n60325 , n60336 );
not ( n60338 , n60012 );
not ( n60339 , n52853 );
or ( n60340 , n60338 , n60339 );
and ( n60341 , n47524 , n57252 );
not ( n60342 , n47524 );
and ( n60343 , n60342 , n52836 );
or ( n60344 , n60341 , n60343 );
not ( n60345 , n60344 );
nand ( n60346 , n60345 , n52469 );
nand ( n60347 , n60340 , n60346 );
xor ( n60348 , n60337 , n60347 );
xor ( n60349 , n60325 , n60336 );
and ( n60350 , n60349 , n60347 );
and ( n60351 , n60325 , n60336 );
or ( n60352 , n60350 , n60351 );
not ( n60353 , n46474 );
not ( n60354 , n59895 );
or ( n60355 , n60353 , n60354 );
not ( n60356 , n46072 );
not ( n60357 , n38498 );
not ( n60358 , n60357 );
or ( n60359 , n60356 , n60358 );
nand ( n60360 , n38498 , n50405 );
nand ( n60361 , n60359 , n60360 );
nand ( n60362 , n60361 , n46602 );
nand ( n60363 , n60355 , n60362 );
xor ( n60364 , n60249 , n60363 );
not ( n60365 , n46564 );
not ( n60366 , n59905 );
or ( n60367 , n60365 , n60366 );
and ( n60368 , n39573 , n47514 );
not ( n60369 , n39573 );
and ( n60370 , n60369 , n48952 );
or ( n60371 , n60368 , n60370 );
nand ( n60372 , n60371 , n49832 );
nand ( n60373 , n60367 , n60372 );
xor ( n60374 , n60364 , n60373 );
xor ( n60375 , n60249 , n60363 );
and ( n60376 , n60375 , n60373 );
and ( n60377 , n60249 , n60363 );
or ( n60378 , n60376 , n60377 );
not ( n60379 , n46267 );
not ( n60380 , n59918 );
or ( n60381 , n60379 , n60380 );
not ( n60382 , n46425 );
not ( n60383 , n39680 );
not ( n60384 , n60383 );
or ( n60385 , n60382 , n60384 );
not ( n60386 , n58482 );
nand ( n60387 , n60386 , n46422 );
nand ( n60388 , n60385 , n60387 );
nand ( n60389 , n60388 , n49026 );
nand ( n60390 , n60381 , n60389 );
xor ( n60391 , n60310 , n60390 );
xor ( n60392 , n60391 , n60253 );
xor ( n60393 , n60310 , n60390 );
and ( n60394 , n60393 , n60253 );
and ( n60395 , n60310 , n60390 );
or ( n60396 , n60394 , n60395 );
not ( n60397 , n60050 );
not ( n60398 , n58635 );
or ( n60399 , n60397 , n60398 );
not ( n60400 , n58006 );
and ( n60401 , n58642 , n47821 );
not ( n60402 , n58642 );
and ( n60403 , n60402 , n49734 );
or ( n60404 , n60401 , n60403 );
nand ( n60405 , n60400 , n60404 );
nand ( n60406 , n60399 , n60405 );
not ( n60407 , n46441 );
not ( n60408 , n60285 );
or ( n60409 , n60407 , n60408 );
nand ( n60410 , n60286 , n46440 );
nand ( n60411 , n60409 , n60410 );
not ( n60412 , n60411 );
not ( n60413 , n60284 );
not ( n60414 , n60274 );
and ( n60415 , n60413 , n60414 );
not ( n60416 , n60413 );
and ( n60417 , n60416 , n60274 );
nor ( n60418 , n60415 , n60417 );
and ( n60419 , n59337 , n60414 );
not ( n60420 , n59337 );
and ( n60421 , n60420 , n59853 );
nor ( n60422 , n60419 , n60421 );
nand ( n60423 , n60418 , n60422 );
not ( n60424 , n60423 );
not ( n60425 , n60424 );
or ( n60426 , n60412 , n60425 );
not ( n60427 , n59854 );
and ( n60428 , n60285 , n45767 );
not ( n60429 , n60285 );
and ( n60430 , n60429 , n50914 );
or ( n60431 , n60428 , n60430 );
nand ( n60432 , n60427 , n60431 );
nand ( n60433 , n60426 , n60432 );
xor ( n60434 , n60406 , n60433 );
not ( n60435 , n50078 );
not ( n60436 , n49770 );
not ( n60437 , n40949 );
not ( n60438 , n60437 );
or ( n60439 , n60436 , n60438 );
nand ( n60440 , n40949 , n50292 );
nand ( n60441 , n60439 , n60440 );
not ( n60442 , n60441 );
or ( n60443 , n60435 , n60442 );
nand ( n60444 , n59837 , n52058 );
nand ( n60445 , n60443 , n60444 );
not ( n60446 , n50580 );
not ( n60447 , n59826 );
or ( n60448 , n60446 , n60447 );
not ( n60449 , n54613 );
not ( n60450 , n41216 );
or ( n60451 , n60449 , n60450 );
nand ( n60452 , n50973 , n50301 );
nand ( n60453 , n60451 , n60452 );
nand ( n60454 , n60453 , n50331 );
nand ( n60455 , n60448 , n60454 );
xor ( n60456 , n60445 , n60455 );
xor ( n60457 , n60434 , n60456 );
xor ( n60458 , n60348 , n60457 );
not ( n60459 , n59983 );
not ( n60460 , n55887 );
or ( n60461 , n60459 , n60460 );
not ( n60462 , n49624 );
not ( n60463 , n58604 );
or ( n60464 , n60462 , n60463 );
nand ( n60465 , n55872 , n49630 );
nand ( n60466 , n60464 , n60465 );
nand ( n60467 , n55459 , n60466 );
nand ( n60468 , n60461 , n60467 );
not ( n60469 , n60030 );
not ( n60470 , n56777 );
or ( n60471 , n60469 , n60470 );
buf ( n60472 , n56780 );
not ( n60473 , n47765 );
not ( n60474 , n56759 );
or ( n60475 , n60473 , n60474 );
nand ( n60476 , n57664 , n48589 );
nand ( n60477 , n60475 , n60476 );
nand ( n60478 , n60472 , n60477 );
nand ( n60479 , n60471 , n60478 );
xor ( n60480 , n60468 , n60479 );
not ( n60481 , n60040 );
buf ( n60482 , n59432 );
not ( n60483 , n60482 );
or ( n60484 , n60481 , n60483 );
not ( n60485 , n52165 );
not ( n60486 , n57534 );
or ( n60487 , n60485 , n60486 );
nand ( n60488 , n57533 , n47368 );
nand ( n60489 , n60487 , n60488 );
nand ( n60490 , n57631 , n60489 );
nand ( n60491 , n60484 , n60490 );
xor ( n60492 , n60480 , n60491 );
xor ( n60493 , n60458 , n60492 );
xor ( n60494 , n60348 , n60457 );
and ( n60495 , n60494 , n60492 );
and ( n60496 , n60348 , n60457 );
or ( n60497 , n60495 , n60496 );
not ( n60498 , n53619 );
not ( n60499 , n47918 );
not ( n60500 , n53594 );
or ( n60501 , n60499 , n60500 );
nand ( n60502 , n59067 , n47510 );
nand ( n60503 , n60501 , n60502 );
not ( n60504 , n60503 );
or ( n60505 , n60498 , n60504 );
not ( n60506 , n60019 );
nand ( n60507 , n60506 , n55913 );
nand ( n60508 , n60505 , n60507 );
not ( n60509 , n54316 );
not ( n60510 , n59962 );
or ( n60511 , n60509 , n60510 );
not ( n60512 , n54185 );
not ( n60513 , n54467 );
or ( n60514 , n60512 , n60513 );
nand ( n60515 , n54298 , n52712 );
nand ( n60516 , n60514 , n60515 );
nand ( n60517 , n54077 , n60516 );
nand ( n60518 , n60511 , n60517 );
xor ( n60519 , n60508 , n60518 );
not ( n60520 , n59972 );
not ( n60521 , n55144 );
or ( n60522 , n60520 , n60521 );
not ( n60523 , n52033 );
not ( n60524 , n55119 );
or ( n60525 , n60523 , n60524 );
nand ( n60526 , n55118 , n55959 );
nand ( n60527 , n60525 , n60526 );
nand ( n60528 , n55157 , n60527 );
nand ( n60529 , n60522 , n60528 );
xor ( n60530 , n60519 , n60529 );
xor ( n60531 , n60530 , n60265 );
xor ( n60532 , n60531 , n60257 );
xor ( n60533 , n60530 , n60265 );
and ( n60534 , n60533 , n60257 );
and ( n60535 , n60530 , n60265 );
or ( n60536 , n60534 , n60535 );
not ( n60537 , n59937 );
buf ( n60538 , n59569 );
not ( n60539 , n60538 );
not ( n60540 , n60539 );
or ( n60541 , n60537 , n60540 );
buf ( n60542 , n58908 );
not ( n60543 , n46273 );
not ( n60544 , n59340 );
or ( n60545 , n60543 , n60544 );
nand ( n60546 , n59338 , n46824 );
nand ( n60547 , n60545 , n60546 );
nand ( n60548 , n60542 , n60547 );
nand ( n60549 , n60541 , n60548 );
xor ( n60550 , n60549 , n59846 );
not ( n60551 , n60108 );
or ( n60552 , n60551 , n50241 );
not ( n60553 , n50232 );
not ( n60554 , n54401 );
or ( n60555 , n60553 , n60554 );
nand ( n60556 , n40147 , n52048 );
nand ( n60557 , n60555 , n60556 );
not ( n60558 , n60557 );
or ( n60559 , n60558 , n50239 );
nand ( n60560 , n60552 , n60559 );
xor ( n60561 , n60550 , n60560 );
xor ( n60562 , n60261 , n60561 );
not ( n60563 , n47407 );
not ( n60564 , n60091 );
or ( n60565 , n60563 , n60564 );
not ( n60566 , n54028 );
not ( n60567 , n56962 );
or ( n60568 , n60566 , n60567 );
nand ( n60569 , n39962 , n48727 );
nand ( n60570 , n60568 , n60569 );
nand ( n60571 , n60570 , n48929 );
nand ( n60572 , n60565 , n60571 );
not ( n60573 , n48989 );
not ( n60574 , n60155 );
or ( n60575 , n60573 , n60574 );
not ( n60576 , n47980 );
not ( n60577 , n40513 );
or ( n60578 , n60576 , n60577 );
nand ( n60579 , n40512 , n47979 );
nand ( n60580 , n60578 , n60579 );
nand ( n60581 , n60580 , n53510 );
nand ( n60582 , n60575 , n60581 );
xor ( n60583 , n60572 , n60582 );
not ( n60584 , n51157 );
not ( n60585 , n60171 );
or ( n60586 , n60584 , n60585 );
not ( n60587 , n50263 );
not ( n60588 , n39894 );
or ( n60589 , n60587 , n60588 );
not ( n60590 , n39893 );
nand ( n60591 , n60590 , n50087 );
nand ( n60592 , n60589 , n60591 );
nand ( n60593 , n60592 , n48073 );
nand ( n60594 , n60586 , n60593 );
xor ( n60595 , n60583 , n60594 );
xor ( n60596 , n60562 , n60595 );
xor ( n60597 , n60261 , n60561 );
and ( n60598 , n60597 , n60595 );
and ( n60599 , n60261 , n60561 );
or ( n60600 , n60598 , n60599 );
not ( n60601 , n58977 );
not ( n60602 , n52728 );
not ( n60603 , n60602 );
not ( n60604 , n52222 );
or ( n60605 , n60603 , n60604 );
buf ( n60606 , n40768 );
nand ( n60607 , n60606 , n52728 );
nand ( n60608 , n60605 , n60607 );
not ( n60609 , n60608 );
or ( n60610 , n60601 , n60609 );
nand ( n60611 , n60073 , n59633 );
nand ( n60612 , n60610 , n60611 );
not ( n60613 , n56639 );
not ( n60614 , n59345 );
not ( n60615 , n50958 );
or ( n60616 , n60614 , n60615 );
not ( n60617 , n59345 );
nand ( n60618 , n51572 , n60617 );
nand ( n60619 , n60616 , n60618 );
not ( n60620 , n60619 );
or ( n60621 , n60613 , n60620 );
nand ( n60622 , n59947 , n59950 );
nand ( n60623 , n60621 , n60622 );
xor ( n60624 , n60612 , n60623 );
not ( n60625 , n60083 );
or ( n60626 , n60625 , n50057 );
not ( n60627 , n49707 );
not ( n60628 , n55202 );
or ( n60629 , n60627 , n60628 );
nand ( n60630 , n40381 , n48661 );
nand ( n60631 , n60629 , n60630 );
not ( n60632 , n60631 );
not ( n60633 , n51865 );
or ( n60634 , n60632 , n60633 );
nand ( n60635 , n60626 , n60634 );
xor ( n60636 , n60624 , n60635 );
xor ( n60637 , n59927 , n60636 );
xor ( n60638 , n60637 , n60269 );
xor ( n60639 , n59927 , n60636 );
and ( n60640 , n60639 , n60269 );
and ( n60641 , n59927 , n60636 );
or ( n60642 , n60640 , n60641 );
not ( n60643 , n54875 );
and ( n60644 , n40225 , n51723 );
not ( n60645 , n40225 );
and ( n60646 , n60645 , n53228 );
or ( n60647 , n60644 , n60646 );
not ( n60648 , n60647 );
or ( n60649 , n60643 , n60648 );
nand ( n60650 , n60120 , n52421 );
nand ( n60651 , n60649 , n60650 );
not ( n60652 , n48894 );
not ( n60653 , n60130 );
or ( n60654 , n60652 , n60653 );
not ( n60655 , n52377 );
not ( n60656 , n55190 );
or ( n60657 , n60655 , n60656 );
nand ( n60658 , n40635 , n55013 );
nand ( n60659 , n60657 , n60658 );
nand ( n60660 , n60659 , n52004 );
nand ( n60661 , n60654 , n60660 );
xor ( n60662 , n60651 , n60661 );
not ( n60663 , n54623 );
not ( n60664 , n54625 );
not ( n60665 , n52211 );
or ( n60666 , n60664 , n60665 );
nand ( n60667 , n40591 , n55023 );
nand ( n60668 , n60666 , n60667 );
not ( n60669 , n60668 );
or ( n60670 , n60663 , n60669 );
nand ( n60671 , n60142 , n47873 );
nand ( n60672 , n60670 , n60671 );
xor ( n60673 , n60662 , n60672 );
xor ( n60674 , n60673 , n59888 );
xor ( n60675 , n60674 , n59992 );
xor ( n60676 , n60673 , n59888 );
and ( n60677 , n60676 , n59992 );
and ( n60678 , n60673 , n59888 );
or ( n60679 , n60677 , n60678 );
xor ( n60680 , n59882 , n60199 );
xor ( n60681 , n60680 , n60245 );
xor ( n60682 , n60374 , n60681 );
xor ( n60683 , n60682 , n60392 );
xor ( n60684 , n60374 , n60681 );
and ( n60685 , n60684 , n60392 );
and ( n60686 , n60374 , n60681 );
or ( n60687 , n60685 , n60686 );
xor ( n60688 , n60493 , n60065 );
xor ( n60689 , n60688 , n60059 );
xor ( n60690 , n60493 , n60065 );
and ( n60691 , n60690 , n60059 );
and ( n60692 , n60493 , n60065 );
or ( n60693 , n60691 , n60692 );
xor ( n60694 , n60532 , n60102 );
xor ( n60695 , n60694 , n60596 );
xor ( n60696 , n60532 , n60102 );
and ( n60697 , n60696 , n60596 );
and ( n60698 , n60532 , n60102 );
or ( n60699 , n60697 , n60698 );
xor ( n60700 , n60508 , n60518 );
and ( n60701 , n60700 , n60529 );
and ( n60702 , n60508 , n60518 );
or ( n60703 , n60701 , n60702 );
xor ( n60704 , n60675 , n60164 );
xor ( n60705 , n60704 , n60638 );
xor ( n60706 , n60675 , n60164 );
and ( n60707 , n60706 , n60638 );
and ( n60708 , n60675 , n60164 );
or ( n60709 , n60707 , n60708 );
xor ( n60710 , n60183 , n60683 );
xor ( n60711 , n60710 , n60189 );
xor ( n60712 , n60183 , n60683 );
and ( n60713 , n60712 , n60189 );
and ( n60714 , n60183 , n60683 );
or ( n60715 , n60713 , n60714 );
xor ( n60716 , n60195 , n60689 );
xor ( n60717 , n60716 , n60695 );
xor ( n60718 , n60195 , n60689 );
and ( n60719 , n60718 , n60695 );
and ( n60720 , n60195 , n60689 );
or ( n60721 , n60719 , n60720 );
xor ( n60722 , n60205 , n60211 );
xor ( n60723 , n60722 , n60705 );
xor ( n60724 , n60205 , n60211 );
and ( n60725 , n60724 , n60705 );
and ( n60726 , n60205 , n60211 );
or ( n60727 , n60725 , n60726 );
xor ( n60728 , n60711 , n60217 );
xor ( n60729 , n60728 , n60717 );
xor ( n60730 , n60711 , n60217 );
and ( n60731 , n60730 , n60717 );
and ( n60732 , n60711 , n60217 );
or ( n60733 , n60731 , n60732 );
xor ( n60734 , n60223 , n60723 );
xor ( n60735 , n60734 , n60229 );
xor ( n60736 , n60223 , n60723 );
and ( n60737 , n60736 , n60229 );
and ( n60738 , n60223 , n60723 );
or ( n60739 , n60737 , n60738 );
xor ( n60740 , n60729 , n60735 );
xor ( n60741 , n60740 , n60235 );
xor ( n60742 , n60729 , n60735 );
and ( n60743 , n60742 , n60235 );
and ( n60744 , n60729 , n60735 );
or ( n60745 , n60743 , n60744 );
xor ( n60746 , n60468 , n60479 );
and ( n60747 , n60746 , n60491 );
and ( n60748 , n60468 , n60479 );
or ( n60749 , n60747 , n60748 );
xor ( n60750 , n60406 , n60433 );
and ( n60751 , n60750 , n60456 );
and ( n60752 , n60406 , n60433 );
or ( n60753 , n60751 , n60752 );
xor ( n60754 , n60549 , n59846 );
and ( n60755 , n60754 , n60560 );
and ( n60756 , n60549 , n59846 );
or ( n60757 , n60755 , n60756 );
xor ( n60758 , n60651 , n60661 );
and ( n60759 , n60758 , n60672 );
and ( n60760 , n60651 , n60661 );
or ( n60761 , n60759 , n60760 );
xor ( n60762 , n60612 , n60623 );
and ( n60763 , n60762 , n60635 );
and ( n60764 , n60612 , n60623 );
or ( n60765 , n60763 , n60764 );
xor ( n60766 , n60572 , n60582 );
and ( n60767 , n60766 , n60594 );
and ( n60768 , n60572 , n60582 );
or ( n60769 , n60767 , n60768 );
xor ( n60770 , n59882 , n60199 );
and ( n60771 , n60770 , n60245 );
and ( n60772 , n59882 , n60199 );
or ( n60773 , n60771 , n60772 );
not ( n60774 , n51234 );
not ( n60775 , n60441 );
or ( n60776 , n60774 , n60775 );
and ( n60777 , n41035 , n50292 );
not ( n60778 , n41035 );
and ( n60779 , n60778 , n49619 );
or ( n60780 , n60777 , n60779 );
nand ( n60781 , n60780 , n49789 );
nand ( n60782 , n60776 , n60781 );
not ( n60783 , n50580 );
not ( n60784 , n60453 );
or ( n60785 , n60783 , n60784 );
not ( n60786 , n54613 );
not ( n60787 , n49548 );
or ( n60788 , n60786 , n60787 );
or ( n60789 , n58013 , n57540 );
nand ( n60790 , n60788 , n60789 );
nand ( n60791 , n60790 , n51452 );
nand ( n60792 , n60785 , n60791 );
xor ( n60793 , n60782 , n60792 );
not ( n60794 , n37570 );
nand ( n60795 , n36927 , n37658 , n37412 );
not ( n60796 , n60795 );
or ( n60797 , n60794 , n60796 );
not ( n60798 , n37570 );
nand ( n60799 , n60798 , n36927 , n37658 , n37412 );
nand ( n60800 , n60797 , n60799 );
not ( n60801 , n60800 );
and ( n60802 , n60284 , n60801 );
not ( n60803 , n60284 );
and ( n60804 , n60803 , n60800 );
nor ( n60805 , n60802 , n60804 );
buf ( n60806 , n60805 );
nor ( n60807 , n60806 , n46441 );
xor ( n60808 , n60793 , n60807 );
xor ( n60809 , n60782 , n60792 );
and ( n60810 , n60809 , n60807 );
and ( n60811 , n60782 , n60792 );
or ( n60812 , n60810 , n60811 );
not ( n60813 , n60306 );
not ( n60814 , n50909 );
not ( n60815 , n60814 );
or ( n60816 , n60813 , n60815 );
not ( n60817 , n50625 );
not ( n60818 , n49000 );
not ( n60819 , n50894 );
or ( n60820 , n60818 , n60819 );
nand ( n60821 , n41284 , n50907 );
nand ( n60822 , n60820 , n60821 );
nand ( n60823 , n60817 , n60822 );
nand ( n60824 , n60816 , n60823 );
not ( n60825 , n60323 );
nor ( n60826 , n51522 , n51516 );
not ( n60827 , n60826 );
or ( n60828 , n60825 , n60827 );
not ( n60829 , n41407 );
not ( n60830 , n51504 );
or ( n60831 , n60829 , n60830 );
nand ( n60832 , n56361 , n50631 );
nand ( n60833 , n60831 , n60832 );
nand ( n60834 , n60833 , n51144 );
nand ( n60835 , n60828 , n60834 );
xor ( n60836 , n60824 , n60835 );
not ( n60837 , n60334 );
not ( n60838 , n54265 );
or ( n60839 , n60837 , n60838 );
not ( n60840 , n41668 );
not ( n60841 , n52109 );
or ( n60842 , n60840 , n60841 );
nand ( n60843 , n53917 , n58914 );
nand ( n60844 , n60842 , n60843 );
nand ( n60845 , n60844 , n51765 );
nand ( n60846 , n60839 , n60845 );
xor ( n60847 , n60836 , n60846 );
xor ( n60848 , n60824 , n60835 );
and ( n60849 , n60848 , n60846 );
and ( n60850 , n60824 , n60835 );
or ( n60851 , n60849 , n60850 );
not ( n60852 , n47009 );
not ( n60853 , n46072 );
buf ( n60854 , n39330 );
not ( n60855 , n60854 );
not ( n60856 , n60855 );
or ( n60857 , n60853 , n60856 );
nand ( n60858 , n39332 , n46071 );
nand ( n60859 , n60857 , n60858 );
not ( n60860 , n60859 );
or ( n60861 , n60852 , n60860 );
nand ( n60862 , n60361 , n50659 );
nand ( n60863 , n60861 , n60862 );
xor ( n60864 , n60863 , n60703 );
xor ( n60865 , n60864 , n60749 );
xor ( n60866 , n60863 , n60703 );
and ( n60867 , n60866 , n60749 );
and ( n60868 , n60863 , n60703 );
or ( n60869 , n60867 , n60868 );
not ( n60870 , n46564 );
not ( n60871 , n60371 );
or ( n60872 , n60870 , n60871 );
not ( n60873 , n48952 );
not ( n60874 , n39055 );
not ( n60875 , n60874 );
or ( n60876 , n60873 , n60875 );
nand ( n60877 , n39055 , n48955 );
nand ( n60878 , n60876 , n60877 );
nand ( n60879 , n60878 , n49832 );
nand ( n60880 , n60872 , n60879 );
xor ( n60881 , n60880 , n60753 );
not ( n60882 , n60570 );
not ( n60883 , n47407 );
or ( n60884 , n60882 , n60883 );
buf ( n60885 , n39845 );
and ( n60886 , n50634 , n60885 );
not ( n60887 , n50634 );
and ( n60888 , n60887 , n39846 );
nor ( n60889 , n60886 , n60888 );
or ( n60890 , n60889 , n53676 );
nand ( n60891 , n60884 , n60890 );
xor ( n60892 , n60881 , n60891 );
xor ( n60893 , n60880 , n60753 );
and ( n60894 , n60893 , n60891 );
and ( n60895 , n60880 , n60753 );
or ( n60896 , n60894 , n60895 );
not ( n60897 , n46267 );
not ( n60898 , n60388 );
or ( n60899 , n60897 , n60898 );
not ( n60900 , n46425 );
and ( n60901 , n831 , n18376 );
not ( n60902 , n831 );
and ( n60903 , n60902 , n39710 );
nor ( n60904 , n60901 , n60903 );
not ( n60905 , n60904 );
not ( n60906 , n60905 );
not ( n60907 , n60906 );
or ( n60908 , n60900 , n60907 );
nand ( n60909 , n39714 , n46422 );
nand ( n60910 , n60908 , n60909 );
nand ( n60911 , n60910 , n49026 );
nand ( n60912 , n60899 , n60911 );
not ( n60913 , n60547 );
not ( n60914 , n60539 );
or ( n60915 , n60913 , n60914 );
and ( n60916 , n47650 , n59338 );
not ( n60917 , n47650 );
and ( n60918 , n60917 , n59339 );
nor ( n60919 , n60916 , n60918 );
not ( n60920 , n60919 );
nand ( n60921 , n60920 , n59931 );
nand ( n60922 , n60915 , n60921 );
and ( n60923 , n60445 , n60455 );
xor ( n60924 , n60922 , n60923 );
not ( n60925 , n60294 );
nand ( n60926 , n60925 , n58168 );
not ( n60927 , n59811 );
not ( n60928 , n49112 );
not ( n60929 , n57307 );
or ( n60930 , n60928 , n60929 );
nand ( n60931 , n40691 , n60292 );
nand ( n60932 , n60930 , n60931 );
nand ( n60933 , n60927 , n60932 );
nand ( n60934 , n60926 , n60933 );
xor ( n60935 , n60924 , n60934 );
xor ( n60936 , n60912 , n60935 );
not ( n60937 , n60404 );
not ( n60938 , n58635 );
or ( n60939 , n60937 , n60938 );
not ( n60940 , n47589 );
not ( n60941 , n58642 );
or ( n60942 , n60940 , n60941 );
not ( n60943 , n58626 );
nand ( n60944 , n60943 , n47227 );
nand ( n60945 , n60942 , n60944 );
nand ( n60946 , n60400 , n60945 );
nand ( n60947 , n60939 , n60946 );
not ( n60948 , n60466 );
not ( n60949 , n56281 );
or ( n60950 , n60948 , n60949 );
not ( n60951 , n55845 );
not ( n60952 , n53126 );
and ( n60953 , n60951 , n60952 );
and ( n60954 , n55891 , n53126 );
nor ( n60955 , n60953 , n60954 );
not ( n60956 , n60955 );
nand ( n60957 , n60956 , n55459 );
nand ( n60958 , n60950 , n60957 );
xor ( n60959 , n60947 , n60958 );
buf ( n60960 , n60423 );
not ( n60961 , n60431 );
or ( n60962 , n60960 , n60961 );
not ( n60963 , n60427 );
not ( n60964 , n60413 );
not ( n60965 , n60964 );
not ( n60966 , n47306 );
and ( n60967 , n60965 , n60966 );
not ( n60968 , n60285 );
not ( n60969 , n60968 );
and ( n60970 , n60969 , n54721 );
nor ( n60971 , n60967 , n60970 );
or ( n60972 , n60963 , n60971 );
nand ( n60973 , n60962 , n60972 );
xor ( n60974 , n60959 , n60973 );
xor ( n60975 , n60936 , n60974 );
xor ( n60976 , n60912 , n60935 );
and ( n60977 , n60976 , n60974 );
and ( n60978 , n60912 , n60935 );
or ( n60979 , n60977 , n60978 );
not ( n60980 , n60527 );
not ( n60981 , n58592 );
or ( n60982 , n60980 , n60981 );
and ( n60983 , n55511 , n55118 );
not ( n60984 , n55511 );
not ( n60985 , n55118 );
and ( n60986 , n60984 , n60985 );
nor ( n60987 , n60983 , n60986 );
nand ( n60988 , n60987 , n54847 );
nand ( n60989 , n60982 , n60988 );
not ( n60990 , n60477 );
not ( n60991 , n56776 );
or ( n60992 , n60990 , n60991 );
not ( n60993 , n51204 );
not ( n60994 , n56759 );
or ( n60995 , n60993 , n60994 );
not ( n60996 , n56784 );
nand ( n60997 , n60996 , n48860 );
nand ( n60998 , n60995 , n60997 );
nand ( n60999 , n56780 , n60998 );
nand ( n61000 , n60992 , n60999 );
xor ( n61001 , n60989 , n61000 );
not ( n61002 , n60489 );
not ( n61003 , n59432 );
or ( n61004 , n61002 , n61003 );
not ( n61005 , n48898 );
not ( n61006 , n57534 );
or ( n61007 , n61005 , n61006 );
nand ( n61008 , n57634 , n48897 );
nand ( n61009 , n61007 , n61008 );
nand ( n61010 , n59435 , n61009 );
nand ( n61011 , n61004 , n61010 );
xor ( n61012 , n61001 , n61011 );
not ( n61013 , n60344 );
not ( n61014 , n61013 );
nand ( n61015 , n52846 , n52847 );
nor ( n61016 , n52467 , n61015 );
not ( n61017 , n61016 );
or ( n61018 , n61014 , n61017 );
not ( n61019 , n56860 );
not ( n61020 , n53946 );
not ( n61021 , n41415 );
or ( n61022 , n61020 , n61021 );
not ( n61023 , n52836 );
or ( n61024 , n61023 , n41417 );
nand ( n61025 , n61022 , n61024 );
nand ( n61026 , n61019 , n61025 );
nand ( n61027 , n61018 , n61026 );
not ( n61028 , n60503 );
not ( n61029 , n53589 );
nand ( n61030 , n61029 , n53601 );
nand ( n61031 , n53589 , n53602 );
and ( n61032 , n61030 , n53324 , n61031 );
not ( n61033 , n61032 );
or ( n61034 , n61028 , n61033 );
not ( n61035 , n57182 );
not ( n61036 , n53594 );
or ( n61037 , n61035 , n61036 );
nand ( n61038 , n59067 , n48523 );
nand ( n61039 , n61037 , n61038 );
nand ( n61040 , n61039 , n53619 );
nand ( n61041 , n61034 , n61040 );
xor ( n61042 , n61027 , n61041 );
not ( n61043 , n60516 );
not ( n61044 , n54315 );
or ( n61045 , n61043 , n61044 );
not ( n61046 , n48983 );
not ( n61047 , n54467 );
or ( n61048 , n61046 , n61047 );
nand ( n61049 , n54298 , n56348 );
nand ( n61050 , n61048 , n61049 );
nand ( n61051 , n61050 , n54077 );
nand ( n61052 , n61045 , n61051 );
xor ( n61053 , n61042 , n61052 );
xor ( n61054 , n61012 , n61053 );
xor ( n61055 , n61054 , n60847 );
xor ( n61056 , n61012 , n61053 );
and ( n61057 , n61056 , n60847 );
and ( n61058 , n61012 , n61053 );
or ( n61059 , n61057 , n61058 );
xor ( n61060 , n60765 , n60757 );
xor ( n61061 , n61060 , n60761 );
xor ( n61062 , n60765 , n60757 );
and ( n61063 , n61062 , n60761 );
and ( n61064 , n60765 , n60757 );
or ( n61065 , n61063 , n61064 );
not ( n61066 , n49252 );
not ( n61067 , n60580 );
or ( n61068 , n61066 , n61067 );
not ( n61069 , n47980 );
not ( n61070 , n56454 );
or ( n61071 , n61069 , n61070 );
nand ( n61072 , n40012 , n47979 );
nand ( n61073 , n61071 , n61072 );
nand ( n61074 , n61073 , n47384 );
nand ( n61075 , n61068 , n61074 );
xor ( n61076 , n60808 , n61075 );
not ( n61077 , n49713 );
not ( n61078 , n60631 );
or ( n61079 , n61077 , n61078 );
and ( n61080 , n40451 , n51351 );
not ( n61081 , n40451 );
and ( n61082 , n61081 , n52267 );
or ( n61083 , n61080 , n61082 );
nand ( n61084 , n61083 , n51865 );
nand ( n61085 , n61079 , n61084 );
xor ( n61086 , n61076 , n61085 );
xor ( n61087 , n61086 , n60769 );
xor ( n61088 , n61087 , n60773 );
xor ( n61089 , n61086 , n60769 );
and ( n61090 , n61089 , n60773 );
and ( n61091 , n61086 , n60769 );
or ( n61092 , n61090 , n61091 );
not ( n61093 , n52970 );
not ( n61094 , n60557 );
or ( n61095 , n61093 , n61094 );
not ( n61096 , n50232 );
not ( n61097 , n56438 );
or ( n61098 , n61096 , n61097 );
nand ( n61099 , n40388 , n49679 );
nand ( n61100 , n61098 , n61099 );
nand ( n61101 , n61100 , n52962 );
nand ( n61102 , n61095 , n61101 );
not ( n61103 , n52421 );
not ( n61104 , n60647 );
or ( n61105 , n61103 , n61104 );
and ( n61106 , n40363 , n51724 );
not ( n61107 , n40363 );
and ( n61108 , n61107 , n51723 );
or ( n61109 , n61106 , n61108 );
nand ( n61110 , n61109 , n54875 );
nand ( n61111 , n61105 , n61110 );
xor ( n61112 , n61102 , n61111 );
not ( n61113 , n57314 );
not ( n61114 , n60659 );
or ( n61115 , n61113 , n61114 );
not ( n61116 , n52377 );
not ( n61117 , n53289 );
or ( n61118 , n61116 , n61117 );
nand ( n61119 , n40377 , n55013 );
nand ( n61120 , n61118 , n61119 );
nand ( n61121 , n61120 , n52004 );
nand ( n61122 , n61115 , n61121 );
xor ( n61123 , n61112 , n61122 );
xor ( n61124 , n60378 , n61123 );
not ( n61125 , n52022 );
not ( n61126 , n60668 );
or ( n61127 , n61125 , n61126 );
not ( n61128 , n59174 );
not ( n61129 , n54046 );
or ( n61130 , n61128 , n61129 );
nand ( n61131 , n40626 , n54628 );
nand ( n61132 , n61130 , n61131 );
nand ( n61133 , n61132 , n54623 );
nand ( n61134 , n61127 , n61133 );
not ( n61135 , n59633 );
not ( n61136 , n60608 );
or ( n61137 , n61135 , n61136 );
not ( n61138 , n60602 );
not ( n61139 , n51916 );
not ( n61140 , n61139 );
or ( n61141 , n61138 , n61140 );
not ( n61142 , n51916 );
or ( n61143 , n61142 , n60602 );
nand ( n61144 , n61141 , n61143 );
nand ( n61145 , n61144 , n58977 );
nand ( n61146 , n61137 , n61145 );
xor ( n61147 , n61134 , n61146 );
not ( n61148 , n59950 );
not ( n61149 , n60619 );
or ( n61150 , n61148 , n61149 );
and ( n61151 , n58246 , n51426 );
not ( n61152 , n58246 );
and ( n61153 , n61152 , n59345 );
or ( n61154 , n61151 , n61153 );
nand ( n61155 , n61154 , n56639 );
nand ( n61156 , n61150 , n61155 );
xor ( n61157 , n61147 , n61156 );
xor ( n61158 , n61124 , n61157 );
xor ( n61159 , n60378 , n61123 );
and ( n61160 , n61159 , n61157 );
and ( n61161 , n60378 , n61123 );
or ( n61162 , n61160 , n61161 );
not ( n61163 , n46776 );
not ( n61164 , n60592 );
or ( n61165 , n61163 , n61164 );
and ( n61166 , n39779 , n52080 );
not ( n61167 , n39779 );
and ( n61168 , n61167 , n50263 );
or ( n61169 , n61166 , n61168 );
nand ( n61170 , n61169 , n48073 );
nand ( n61171 , n61165 , n61170 );
xor ( n61172 , n61171 , n60314 );
xor ( n61173 , n61172 , n60352 );
xor ( n61174 , n60892 , n61173 );
xor ( n61175 , n61174 , n60865 );
xor ( n61176 , n60892 , n61173 );
and ( n61177 , n61176 , n60865 );
and ( n61178 , n60892 , n61173 );
or ( n61179 , n61177 , n61178 );
xor ( n61180 , n60497 , n60396 );
xor ( n61181 , n61180 , n60975 );
xor ( n61182 , n60497 , n60396 );
and ( n61183 , n61182 , n60975 );
and ( n61184 , n60497 , n60396 );
or ( n61185 , n61183 , n61184 );
xor ( n61186 , n60536 , n61055 );
xor ( n61187 , n61186 , n60600 );
xor ( n61188 , n60536 , n61055 );
and ( n61189 , n61188 , n60600 );
and ( n61190 , n60536 , n61055 );
or ( n61191 , n61189 , n61190 );
xor ( n61192 , n61027 , n61041 );
and ( n61193 , n61192 , n61052 );
and ( n61194 , n61027 , n61041 );
or ( n61195 , n61193 , n61194 );
xor ( n61196 , n60642 , n61061 );
xor ( n61197 , n61196 , n60687 );
xor ( n61198 , n60642 , n61061 );
and ( n61199 , n61198 , n60687 );
and ( n61200 , n60642 , n61061 );
or ( n61201 , n61199 , n61200 );
xor ( n61202 , n61088 , n60679 );
xor ( n61203 , n61202 , n61158 );
xor ( n61204 , n61088 , n60679 );
and ( n61205 , n61204 , n61158 );
and ( n61206 , n61088 , n60679 );
or ( n61207 , n61205 , n61206 );
xor ( n61208 , n60693 , n61181 );
xor ( n61209 , n61208 , n61175 );
xor ( n61210 , n60693 , n61181 );
and ( n61211 , n61210 , n61175 );
and ( n61212 , n60693 , n61181 );
or ( n61213 , n61211 , n61212 );
xor ( n61214 , n61187 , n60699 );
xor ( n61215 , n61214 , n61197 );
xor ( n61216 , n61187 , n60699 );
and ( n61217 , n61216 , n61197 );
and ( n61218 , n61187 , n60699 );
or ( n61219 , n61217 , n61218 );
xor ( n61220 , n60709 , n60715 );
xor ( n61221 , n61220 , n61203 );
xor ( n61222 , n60709 , n60715 );
and ( n61223 , n61222 , n61203 );
and ( n61224 , n60709 , n60715 );
or ( n61225 , n61223 , n61224 );
xor ( n61226 , n61209 , n60721 );
xor ( n61227 , n61226 , n61215 );
xor ( n61228 , n61209 , n60721 );
and ( n61229 , n61228 , n61215 );
and ( n61230 , n61209 , n60721 );
or ( n61231 , n61229 , n61230 );
xor ( n61232 , n60727 , n61221 );
xor ( n61233 , n61232 , n60733 );
xor ( n61234 , n60727 , n61221 );
and ( n61235 , n61234 , n60733 );
and ( n61236 , n60727 , n61221 );
or ( n61237 , n61235 , n61236 );
xor ( n61238 , n61227 , n61233 );
xor ( n61239 , n61238 , n60739 );
xor ( n61240 , n61227 , n61233 );
and ( n61241 , n61240 , n60739 );
and ( n61242 , n61227 , n61233 );
or ( n61243 , n61241 , n61242 );
xor ( n61244 , n60989 , n61000 );
and ( n61245 , n61244 , n61011 );
and ( n61246 , n60989 , n61000 );
or ( n61247 , n61245 , n61246 );
xor ( n61248 , n60947 , n60958 );
and ( n61249 , n61248 , n60973 );
and ( n61250 , n60947 , n60958 );
or ( n61251 , n61249 , n61250 );
xor ( n61252 , n60922 , n60923 );
and ( n61253 , n61252 , n60934 );
and ( n61254 , n60922 , n60923 );
or ( n61255 , n61253 , n61254 );
xor ( n61256 , n61102 , n61111 );
and ( n61257 , n61256 , n61122 );
and ( n61258 , n61102 , n61111 );
or ( n61259 , n61257 , n61258 );
xor ( n61260 , n61134 , n61146 );
and ( n61261 , n61260 , n61156 );
and ( n61262 , n61134 , n61146 );
or ( n61263 , n61261 , n61262 );
xor ( n61264 , n60808 , n61075 );
and ( n61265 , n61264 , n61085 );
and ( n61266 , n60808 , n61075 );
or ( n61267 , n61265 , n61266 );
xor ( n61268 , n61171 , n60314 );
and ( n61269 , n61268 , n60352 );
and ( n61270 , n61171 , n60314 );
or ( n61271 , n61269 , n61270 );
not ( n61272 , n50078 );
not ( n61273 , n49619 );
not ( n61274 , n52767 );
or ( n61275 , n61273 , n61274 );
nand ( n61276 , n41131 , n49766 );
nand ( n61277 , n61275 , n61276 );
not ( n61278 , n61277 );
or ( n61279 , n61272 , n61278 );
nand ( n61280 , n60780 , n54960 );
nand ( n61281 , n61279 , n61280 );
not ( n61282 , n60822 );
not ( n61283 , n50911 );
or ( n61284 , n61282 , n61283 );
not ( n61285 , n57571 );
not ( n61286 , n50916 );
or ( n61287 , n61285 , n61286 );
nand ( n61288 , n51461 , n41216 );
nand ( n61289 , n61287 , n61288 );
nand ( n61290 , n61289 , n50921 );
nand ( n61291 , n61284 , n61290 );
xor ( n61292 , n61281 , n61291 );
not ( n61293 , n60833 );
not ( n61294 , n51525 );
or ( n61295 , n61293 , n61294 );
not ( n61296 , n41363 );
not ( n61297 , n51504 );
or ( n61298 , n61296 , n61297 );
nand ( n61299 , n60321 , n52271 );
nand ( n61300 , n61298 , n61299 );
nand ( n61301 , n51145 , n61300 );
nand ( n61302 , n61295 , n61301 );
xor ( n61303 , n61292 , n61302 );
xor ( n61304 , n61281 , n61291 );
and ( n61305 , n61304 , n61302 );
and ( n61306 , n61281 , n61291 );
or ( n61307 , n61305 , n61306 );
not ( n61308 , n60844 );
not ( n61309 , n54265 );
or ( n61310 , n61308 , n61309 );
and ( n61311 , n41532 , n53917 );
not ( n61312 , n41532 );
and ( n61313 , n61312 , n52113 );
nor ( n61314 , n61311 , n61313 );
nand ( n61315 , n51765 , n61314 );
nand ( n61316 , n61310 , n61315 );
not ( n61317 , n61025 );
not ( n61318 , n52853 );
or ( n61319 , n61317 , n61318 );
not ( n61320 , n58458 );
not ( n61321 , n55102 );
or ( n61322 , n61320 , n61321 );
not ( n61323 , n57252 );
nand ( n61324 , n61323 , n58453 );
nand ( n61325 , n61322 , n61324 );
nand ( n61326 , n52469 , n61325 );
nand ( n61327 , n61319 , n61326 );
xor ( n61328 , n61316 , n61327 );
not ( n61329 , n53955 );
not ( n61330 , n61039 );
or ( n61331 , n61329 , n61330 );
not ( n61332 , n47527 );
not ( n61333 , n56802 );
or ( n61334 , n61332 , n61333 );
nand ( n61335 , n59067 , n51360 );
nand ( n61336 , n61334 , n61335 );
not ( n61337 , n61336 );
not ( n61338 , n53326 );
or ( n61339 , n61337 , n61338 );
nand ( n61340 , n61331 , n61339 );
xor ( n61341 , n61328 , n61340 );
xor ( n61342 , n61316 , n61327 );
and ( n61343 , n61342 , n61340 );
and ( n61344 , n61316 , n61327 );
or ( n61345 , n61343 , n61344 );
not ( n61346 , n49832 );
not ( n61347 , n38498 );
and ( n61348 , n48952 , n61347 );
not ( n61349 , n48952 );
and ( n61350 , n61349 , n38498 );
nor ( n61351 , n61348 , n61350 );
not ( n61352 , n61351 );
not ( n61353 , n61352 );
or ( n61354 , n61346 , n61353 );
nand ( n61355 , n60878 , n45842 );
nand ( n61356 , n61354 , n61355 );
xor ( n61357 , n61356 , n61251 );
not ( n61358 , n51545 );
not ( n61359 , n39893 );
or ( n61360 , n61358 , n61359 );
nand ( n61361 , n57787 , n50634 );
nand ( n61362 , n61360 , n61361 );
not ( n61363 , n61362 );
not ( n61364 , n53675 );
or ( n61365 , n61363 , n61364 );
not ( n61366 , n47407 );
or ( n61367 , n60889 , n61366 );
nand ( n61368 , n61365 , n61367 );
xor ( n61369 , n61357 , n61368 );
xor ( n61370 , n61356 , n61251 );
and ( n61371 , n61370 , n61368 );
and ( n61372 , n61356 , n61251 );
or ( n61373 , n61371 , n61372 );
not ( n61374 , n46267 );
not ( n61375 , n60910 );
or ( n61376 , n61374 , n61375 );
and ( n61377 , n39573 , n46422 );
not ( n61378 , n39573 );
and ( n61379 , n61378 , n46425 );
or ( n61380 , n61377 , n61379 );
nand ( n61381 , n61380 , n49026 );
nand ( n61382 , n61376 , n61381 );
not ( n61383 , n50659 );
not ( n61384 , n60859 );
or ( n61385 , n61383 , n61384 );
or ( n61386 , n46071 , n39253 );
nand ( n61387 , n46071 , n39253 );
nand ( n61388 , n61386 , n61387 );
nand ( n61389 , n61388 , n47009 );
nand ( n61390 , n61385 , n61389 );
xor ( n61391 , n61382 , n61390 );
xor ( n61392 , n61391 , n61255 );
xor ( n61393 , n61382 , n61390 );
and ( n61394 , n61393 , n61255 );
and ( n61395 , n61382 , n61390 );
or ( n61396 , n61394 , n61395 );
nand ( n61397 , n60422 , n60418 );
or ( n61398 , n60971 , n61397 );
and ( n61399 , n60968 , n46273 );
and ( n61400 , n60285 , n46824 );
nor ( n61401 , n61399 , n61400 );
or ( n61402 , n61401 , n59854 );
nand ( n61403 , n61398 , n61402 );
not ( n61404 , n60801 );
and ( n61405 , n61404 , n48689 );
not ( n61406 , n37585 );
not ( n61407 , n37455 );
nor ( n61408 , n36697 , n37654 );
nand ( n61409 , n61408 , n51754 );
nand ( n61410 , n61407 , n61409 , n37656 );
not ( n61411 , n61410 );
not ( n61412 , n61411 );
or ( n61413 , n61406 , n61412 );
nand ( n61414 , n61410 , n37586 );
nand ( n61415 , n61413 , n61414 );
buf ( n61416 , n61415 );
not ( n61417 , n61416 );
nor ( n61418 , n61405 , n61417 );
or ( n61419 , n61404 , n48689 );
nand ( n61420 , n61419 , n60964 );
nand ( n61421 , n61418 , n61420 );
not ( n61422 , n61421 );
not ( n61423 , n61422 );
not ( n61424 , n49920 );
not ( n61425 , n50304 );
not ( n61426 , n60437 );
or ( n61427 , n61425 , n61426 );
nand ( n61428 , n40949 , n50163 );
nand ( n61429 , n61427 , n61428 );
not ( n61430 , n61429 );
or ( n61431 , n61424 , n61430 );
not ( n61432 , n50319 );
nand ( n61433 , n61432 , n60790 );
nand ( n61434 , n61431 , n61433 );
not ( n61435 , n61434 );
not ( n61436 , n61435 );
or ( n61437 , n61423 , n61436 );
or ( n61438 , n61435 , n61422 );
nand ( n61439 , n61437 , n61438 );
xor ( n61440 , n61403 , n61439 );
not ( n61441 , n59931 );
and ( n61442 , n49734 , n59578 );
not ( n61443 , n49734 );
and ( n61444 , n61443 , n59935 );
or ( n61445 , n61442 , n61444 );
not ( n61446 , n61445 );
or ( n61447 , n61441 , n61446 );
or ( n61448 , n60538 , n60919 );
nand ( n61449 , n61447 , n61448 );
xor ( n61450 , n61440 , n61449 );
xor ( n61451 , n61303 , n61450 );
not ( n61452 , n61009 );
not ( n61453 , n59432 );
or ( n61454 , n61452 , n61453 );
not ( n61455 , n47765 );
not ( n61456 , n57534 );
or ( n61457 , n61455 , n61456 );
nand ( n61458 , n57619 , n48589 );
nand ( n61459 , n61457 , n61458 );
nand ( n61460 , n57139 , n61459 );
nand ( n61461 , n61454 , n61460 );
not ( n61462 , n60945 );
not ( n61463 , n59445 );
or ( n61464 , n61462 , n61463 );
not ( n61465 , n58006 );
not ( n61466 , n49654 );
not ( n61467 , n58433 );
or ( n61468 , n61466 , n61467 );
nand ( n61469 , n58642 , n47368 );
nand ( n61470 , n61468 , n61469 );
nand ( n61471 , n61465 , n61470 );
nand ( n61472 , n61464 , n61471 );
xor ( n61473 , n61461 , n61472 );
not ( n61474 , n60955 );
not ( n61475 , n61474 );
not ( n61476 , n55887 );
or ( n61477 , n61475 , n61476 );
not ( n61478 , n52033 );
not ( n61479 , n55846 );
or ( n61480 , n61478 , n61479 );
nand ( n61481 , n55872 , n52038 );
nand ( n61482 , n61480 , n61481 );
nand ( n61483 , n59984 , n61482 );
nand ( n61484 , n61477 , n61483 );
xor ( n61485 , n61473 , n61484 );
xor ( n61486 , n61451 , n61485 );
xor ( n61487 , n61303 , n61450 );
and ( n61488 , n61487 , n61485 );
and ( n61489 , n61303 , n61450 );
or ( n61490 , n61488 , n61489 );
not ( n61491 , n61050 );
not ( n61492 , n56810 );
or ( n61493 , n61491 , n61492 );
not ( n61494 , n56727 );
not ( n61495 , n54322 );
or ( n61496 , n61494 , n61495 );
nand ( n61497 , n54297 , n47511 );
nand ( n61498 , n61496 , n61497 );
nand ( n61499 , n61498 , n56277 );
nand ( n61500 , n61493 , n61499 );
not ( n61501 , n60987 );
not ( n61502 , n55143 );
or ( n61503 , n61501 , n61502 );
not ( n61504 , n48223 );
not ( n61505 , n58108 );
or ( n61506 , n61504 , n61505 );
not ( n61507 , n60985 );
nand ( n61508 , n61507 , n52712 );
nand ( n61509 , n61506 , n61508 );
nand ( n61510 , n61509 , n55155 );
nand ( n61511 , n61503 , n61510 );
xor ( n61512 , n61500 , n61511 );
not ( n61513 , n60998 );
not ( n61514 , n56776 );
or ( n61515 , n61513 , n61514 );
and ( n61516 , n49624 , n56759 );
not ( n61517 , n49624 );
not ( n61518 , n57665 );
and ( n61519 , n61517 , n61518 );
or ( n61520 , n61516 , n61519 );
nand ( n61521 , n60472 , n61520 );
nand ( n61522 , n61515 , n61521 );
xor ( n61523 , n61512 , n61522 );
xor ( n61524 , n61523 , n61341 );
xor ( n61525 , n61524 , n61263 );
xor ( n61526 , n61523 , n61341 );
and ( n61527 , n61526 , n61263 );
and ( n61528 , n61523 , n61341 );
or ( n61529 , n61527 , n61528 );
xor ( n61530 , n61259 , n61267 );
not ( n61531 , n46440 );
not ( n61532 , n37585 );
not ( n61533 , n61411 );
or ( n61534 , n61532 , n61533 );
nand ( n61535 , n61534 , n61414 );
not ( n61536 , n61535 );
buf ( n61537 , n61536 );
not ( n61538 , n61537 );
or ( n61539 , n61531 , n61538 );
not ( n61540 , n61537 );
nand ( n61541 , n61540 , n46441 );
nand ( n61542 , n61539 , n61541 );
not ( n61543 , n61542 );
and ( n61544 , n60801 , n61536 );
and ( n61545 , n60800 , n61535 );
nor ( n61546 , n61544 , n61545 );
nand ( n61547 , n60805 , n61546 );
not ( n61548 , n61547 );
not ( n61549 , n61548 );
not ( n61550 , n61549 );
not ( n61551 , n61550 );
or ( n61552 , n61543 , n61551 );
and ( n61553 , n61536 , n50914 );
and ( n61554 , n61416 , n48766 );
nor ( n61555 , n61553 , n61554 );
not ( n61556 , n61555 );
not ( n61557 , n60806 );
buf ( n61558 , n61557 );
nand ( n61559 , n61556 , n61558 );
nand ( n61560 , n61552 , n61559 );
xor ( n61561 , n61560 , n60812 );
not ( n61562 , n50242 );
not ( n61563 , n61100 );
or ( n61564 , n61562 , n61563 );
and ( n61565 , n40380 , n52048 );
not ( n61566 , n40380 );
and ( n61567 , n61566 , n48645 );
or ( n61568 , n61565 , n61567 );
nand ( n61569 , n61568 , n52962 );
nand ( n61570 , n61564 , n61569 );
xor ( n61571 , n61561 , n61570 );
xor ( n61572 , n61530 , n61571 );
xor ( n61573 , n61259 , n61267 );
and ( n61574 , n61573 , n61571 );
and ( n61575 , n61259 , n61267 );
or ( n61576 , n61574 , n61575 );
not ( n61577 , n59950 );
not ( n61578 , n61154 );
or ( n61579 , n61577 , n61578 );
and ( n61580 , n40768 , n51426 );
not ( n61581 , n40768 );
and ( n61582 , n61581 , n59345 );
or ( n61583 , n61580 , n61582 );
nand ( n61584 , n61583 , n56639 );
nand ( n61585 , n61579 , n61584 );
not ( n61586 , n52191 );
not ( n61587 , n49112 );
not ( n61588 , n51573 );
or ( n61589 , n61587 , n61588 );
nand ( n61590 , n51572 , n60289 );
nand ( n61591 , n61589 , n61590 );
not ( n61592 , n61591 );
or ( n61593 , n61586 , n61592 );
nand ( n61594 , n60932 , n58168 );
nand ( n61595 , n61593 , n61594 );
xor ( n61596 , n61585 , n61595 );
not ( n61597 , n50261 );
and ( n61598 , n39680 , n52080 );
not ( n61599 , n39680 );
and ( n61600 , n61599 , n46650 );
or ( n61601 , n61598 , n61600 );
not ( n61602 , n61601 );
or ( n61603 , n61597 , n61602 );
nand ( n61604 , n61169 , n51157 );
nand ( n61605 , n61603 , n61604 );
xor ( n61606 , n61596 , n61605 );
xor ( n61607 , n61606 , n61271 );
xor ( n61608 , n61607 , n60869 );
xor ( n61609 , n61606 , n61271 );
and ( n61610 , n61609 , n60869 );
and ( n61611 , n61606 , n61271 );
or ( n61612 , n61610 , n61611 );
not ( n61613 , n52421 );
not ( n61614 , n61109 );
or ( n61615 , n61613 , n61614 );
and ( n61616 , n40147 , n58692 );
not ( n61617 , n40147 );
and ( n61618 , n61617 , n51723 );
or ( n61619 , n61616 , n61618 );
nand ( n61620 , n61619 , n47148 );
nand ( n61621 , n61615 , n61620 );
not ( n61622 , n49713 );
not ( n61623 , n61083 );
or ( n61624 , n61622 , n61623 );
not ( n61625 , n49707 );
not ( n61626 , n56975 );
or ( n61627 , n61625 , n61626 );
nand ( n61628 , n40512 , n51351 );
nand ( n61629 , n61627 , n61628 );
nand ( n61630 , n61629 , n51865 );
nand ( n61631 , n61624 , n61630 );
xor ( n61632 , n61621 , n61631 );
not ( n61633 , n52004 );
not ( n61634 , n52377 );
not ( n61635 , n40225 );
or ( n61636 , n61634 , n61635 );
nand ( n61637 , n56073 , n53973 );
nand ( n61638 , n61636 , n61637 );
not ( n61639 , n61638 );
or ( n61640 , n61633 , n61639 );
nand ( n61641 , n61120 , n57314 );
nand ( n61642 , n61640 , n61641 );
xor ( n61643 , n61632 , n61642 );
xor ( n61644 , n61643 , n60896 );
not ( n61645 , n47873 );
not ( n61646 , n61132 );
or ( n61647 , n61645 , n61646 );
not ( n61648 , n54625 );
not ( n61649 , n55190 );
or ( n61650 , n61648 , n61649 );
nand ( n61651 , n40635 , n51684 );
nand ( n61652 , n61650 , n61651 );
nand ( n61653 , n61652 , n54623 );
nand ( n61654 , n61647 , n61653 );
not ( n61655 , n48989 );
not ( n61656 , n61073 );
or ( n61657 , n61655 , n61656 );
not ( n61658 , n47980 );
not ( n61659 , n39963 );
or ( n61660 , n61658 , n61659 );
nand ( n61661 , n39962 , n47979 );
nand ( n61662 , n61660 , n61661 );
nand ( n61663 , n61662 , n47384 );
nand ( n61664 , n61657 , n61663 );
xor ( n61665 , n61654 , n61664 );
not ( n61666 , n61144 );
or ( n61667 , n61666 , n59632 );
not ( n61668 , n60602 );
not ( n61669 , n53730 );
or ( n61670 , n61668 , n61669 );
nand ( n61671 , n54380 , n52728 );
nand ( n61672 , n61670 , n61671 );
not ( n61673 , n61672 );
or ( n61674 , n61673 , n59630 );
nand ( n61675 , n61667 , n61674 );
xor ( n61676 , n61665 , n61675 );
xor ( n61677 , n61644 , n61676 );
xor ( n61678 , n61643 , n60896 );
and ( n61679 , n61678 , n61676 );
and ( n61680 , n61643 , n60896 );
or ( n61681 , n61679 , n61680 );
xor ( n61682 , n61059 , n61392 );
xor ( n61683 , n60851 , n61195 );
xor ( n61684 , n61683 , n61247 );
xor ( n61685 , n61682 , n61684 );
xor ( n61686 , n61059 , n61392 );
and ( n61687 , n61686 , n61684 );
and ( n61688 , n61059 , n61392 );
or ( n61689 , n61687 , n61688 );
xor ( n61690 , n61369 , n60979 );
xor ( n61691 , n61690 , n61065 );
xor ( n61692 , n61369 , n60979 );
and ( n61693 , n61692 , n61065 );
and ( n61694 , n61369 , n60979 );
or ( n61695 , n61693 , n61694 );
xor ( n61696 , n61486 , n61525 );
xor ( n61697 , n61696 , n61162 );
xor ( n61698 , n61486 , n61525 );
and ( n61699 , n61698 , n61162 );
and ( n61700 , n61486 , n61525 );
or ( n61701 , n61699 , n61700 );
xor ( n61702 , n61500 , n61511 );
and ( n61703 , n61702 , n61522 );
and ( n61704 , n61500 , n61511 );
or ( n61705 , n61703 , n61704 );
xor ( n61706 , n61572 , n61092 );
xor ( n61707 , n61706 , n61608 );
xor ( n61708 , n61572 , n61092 );
and ( n61709 , n61708 , n61608 );
and ( n61710 , n61572 , n61092 );
or ( n61711 , n61709 , n61710 );
xor ( n61712 , n61677 , n61179 );
xor ( n61713 , n61712 , n61185 );
xor ( n61714 , n61677 , n61179 );
and ( n61715 , n61714 , n61185 );
and ( n61716 , n61677 , n61179 );
or ( n61717 , n61715 , n61716 );
xor ( n61718 , n61685 , n61691 );
xor ( n61719 , n61718 , n61191 );
xor ( n61720 , n61685 , n61691 );
and ( n61721 , n61720 , n61191 );
and ( n61722 , n61685 , n61691 );
or ( n61723 , n61721 , n61722 );
xor ( n61724 , n61697 , n61207 );
xor ( n61725 , n61724 , n61707 );
xor ( n61726 , n61697 , n61207 );
and ( n61727 , n61726 , n61707 );
and ( n61728 , n61697 , n61207 );
or ( n61729 , n61727 , n61728 );
xor ( n61730 , n61201 , n61213 );
xor ( n61731 , n61730 , n61713 );
xor ( n61732 , n61201 , n61213 );
and ( n61733 , n61732 , n61713 );
and ( n61734 , n61201 , n61213 );
or ( n61735 , n61733 , n61734 );
xor ( n61736 , n61719 , n61219 );
xor ( n61737 , n61736 , n61225 );
xor ( n61738 , n61719 , n61219 );
and ( n61739 , n61738 , n61225 );
and ( n61740 , n61719 , n61219 );
or ( n61741 , n61739 , n61740 );
xor ( n61742 , n61725 , n61731 );
xor ( n61743 , n61742 , n61231 );
xor ( n61744 , n61725 , n61731 );
and ( n61745 , n61744 , n61231 );
and ( n61746 , n61725 , n61731 );
or ( n61747 , n61745 , n61746 );
xor ( n61748 , n61737 , n61743 );
xor ( n61749 , n61748 , n61237 );
xor ( n61750 , n61737 , n61743 );
and ( n61751 , n61750 , n61237 );
and ( n61752 , n61737 , n61743 );
or ( n61753 , n61751 , n61752 );
xor ( n61754 , n61461 , n61472 );
and ( n61755 , n61754 , n61484 );
and ( n61756 , n61461 , n61472 );
or ( n61757 , n61755 , n61756 );
xor ( n61758 , n61403 , n61439 );
and ( n61759 , n61758 , n61449 );
and ( n61760 , n61403 , n61439 );
or ( n61761 , n61759 , n61760 );
xor ( n61762 , n61560 , n60812 );
and ( n61763 , n61762 , n61570 );
and ( n61764 , n61560 , n60812 );
or ( n61765 , n61763 , n61764 );
xor ( n61766 , n61621 , n61631 );
and ( n61767 , n61766 , n61642 );
and ( n61768 , n61621 , n61631 );
or ( n61769 , n61767 , n61768 );
xor ( n61770 , n61654 , n61664 );
and ( n61771 , n61770 , n61675 );
and ( n61772 , n61654 , n61664 );
or ( n61773 , n61771 , n61772 );
xor ( n61774 , n61585 , n61595 );
and ( n61775 , n61774 , n61605 );
and ( n61776 , n61585 , n61595 );
or ( n61777 , n61775 , n61776 );
xor ( n61778 , n60851 , n61195 );
and ( n61779 , n61778 , n61247 );
and ( n61780 , n60851 , n61195 );
or ( n61781 , n61779 , n61780 );
not ( n61782 , n52757 );
not ( n61783 , n50304 );
not ( n61784 , n51110 );
or ( n61785 , n61783 , n61784 );
nand ( n61786 , n41036 , n54614 );
nand ( n61787 , n61785 , n61786 );
not ( n61788 , n61787 );
or ( n61789 , n61782 , n61788 );
nand ( n61790 , n61429 , n52749 );
nand ( n61791 , n61789 , n61790 );
not ( n61792 , n61416 );
buf ( n61793 , n51754 );
not ( n61794 , n37523 );
not ( n61795 , n61794 );
nor ( n61796 , n61795 , n37542 );
nand ( n61797 , n61793 , n61796 );
nand ( n61798 , n61797 , n37660 , n37645 );
nand ( n61799 , n37496 , n37490 );
not ( n61800 , n61799 );
and ( n61801 , n61798 , n61800 );
not ( n61802 , n61798 );
and ( n61803 , n61802 , n61799 );
nor ( n61804 , n61801 , n61803 );
not ( n61805 , n61804 );
not ( n61806 , n61805 );
or ( n61807 , n61792 , n61806 );
and ( n61808 , n61798 , n61800 );
not ( n61809 , n61798 );
and ( n61810 , n61809 , n61799 );
nor ( n61811 , n61808 , n61810 );
nand ( n61812 , n61536 , n61811 );
nand ( n61813 , n61807 , n61812 );
and ( n61814 , n61813 , n48689 );
xor ( n61815 , n61791 , n61814 );
not ( n61816 , n61289 );
not ( n61817 , n51215 );
or ( n61818 , n61816 , n61817 );
not ( n61819 , n56239 );
not ( n61820 , n51462 );
or ( n61821 , n61819 , n61820 );
nand ( n61822 , n51461 , n50004 );
nand ( n61823 , n61821 , n61822 );
nand ( n61824 , n61823 , n50921 );
nand ( n61825 , n61818 , n61824 );
xor ( n61826 , n61815 , n61825 );
xor ( n61827 , n61791 , n61814 );
and ( n61828 , n61827 , n61825 );
and ( n61829 , n61791 , n61814 );
or ( n61830 , n61828 , n61829 );
not ( n61831 , n61300 );
not ( n61832 , n60826 );
or ( n61833 , n61831 , n61832 );
and ( n61834 , n48996 , n51504 );
not ( n61835 , n48996 );
and ( n61836 , n61835 , n53549 );
or ( n61837 , n61834 , n61836 );
nand ( n61838 , n61837 , n51144 );
nand ( n61839 , n61833 , n61838 );
and ( n61840 , n61434 , n61422 );
xor ( n61841 , n61839 , n61840 );
not ( n61842 , n61314 );
not ( n61843 , n52125 );
or ( n61844 , n61842 , n61843 );
not ( n61845 , n41407 );
not ( n61846 , n52109 );
or ( n61847 , n61845 , n61846 );
nand ( n61848 , n48951 , n52870 );
nand ( n61849 , n61847 , n61848 );
nand ( n61850 , n61849 , n51766 );
nand ( n61851 , n61844 , n61850 );
xor ( n61852 , n61841 , n61851 );
xor ( n61853 , n61839 , n61840 );
and ( n61854 , n61853 , n61851 );
and ( n61855 , n61839 , n61840 );
or ( n61856 , n61854 , n61855 );
not ( n61857 , n49832 );
and ( n61858 , n39331 , n48952 );
not ( n61859 , n39331 );
and ( n61860 , n61859 , n47514 );
or ( n61861 , n61858 , n61860 );
not ( n61862 , n61861 );
or ( n61863 , n61857 , n61862 );
not ( n61864 , n61351 );
nand ( n61865 , n61864 , n46564 );
nand ( n61866 , n61863 , n61865 );
xor ( n61867 , n61826 , n61866 );
xor ( n61868 , n61867 , n61757 );
xor ( n61869 , n61826 , n61866 );
and ( n61870 , n61869 , n61757 );
and ( n61871 , n61826 , n61866 );
or ( n61872 , n61870 , n61871 );
not ( n61873 , n47407 );
not ( n61874 , n61362 );
or ( n61875 , n61873 , n61874 );
not ( n61876 , n47803 );
not ( n61877 , n58047 );
or ( n61878 , n61876 , n61877 );
nand ( n61879 , n39779 , n50634 );
nand ( n61880 , n61878 , n61879 );
nand ( n61881 , n61880 , n53675 );
nand ( n61882 , n61875 , n61881 );
xor ( n61883 , n61761 , n61882 );
not ( n61884 , n47384 );
not ( n61885 , n47980 );
not ( n61886 , n39844 );
or ( n61887 , n61885 , n61886 );
not ( n61888 , n39843 );
nand ( n61889 , n61888 , n47979 );
nand ( n61890 , n61887 , n61889 );
not ( n61891 , n61890 );
or ( n61892 , n61884 , n61891 );
nand ( n61893 , n61662 , n49252 );
nand ( n61894 , n61892 , n61893 );
xor ( n61895 , n61883 , n61894 );
xor ( n61896 , n61761 , n61882 );
and ( n61897 , n61896 , n61894 );
and ( n61898 , n61761 , n61882 );
or ( n61899 , n61897 , n61898 );
not ( n61900 , n46474 );
not ( n61901 , n61388 );
or ( n61902 , n61900 , n61901 );
nand ( n61903 , n42458 , n42451 );
not ( n61904 , n61903 );
and ( n61905 , n50405 , n61904 );
not ( n61906 , n50405 );
not ( n61907 , n61904 );
and ( n61908 , n61906 , n61907 );
nor ( n61909 , n61905 , n61908 );
nand ( n61910 , n61909 , n47009 );
nand ( n61911 , n61902 , n61910 );
not ( n61912 , n46267 );
not ( n61913 , n61380 );
or ( n61914 , n61912 , n61913 );
not ( n61915 , n46425 );
not ( n61916 , n60874 );
or ( n61917 , n61915 , n61916 );
nand ( n61918 , n46422 , n39055 );
nand ( n61919 , n61917 , n61918 );
nand ( n61920 , n61919 , n49026 );
nand ( n61921 , n61914 , n61920 );
xor ( n61922 , n61911 , n61921 );
xor ( n61923 , n61922 , n61852 );
xor ( n61924 , n61911 , n61921 );
and ( n61925 , n61924 , n61852 );
and ( n61926 , n61911 , n61921 );
or ( n61927 , n61925 , n61926 );
not ( n61928 , n61445 );
not ( n61929 , n59570 );
or ( n61930 , n61928 , n61929 );
not ( n61931 , n47227 );
not ( n61932 , n59578 );
or ( n61933 , n61931 , n61932 );
nand ( n61934 , n59935 , n47589 );
nand ( n61935 , n61933 , n61934 );
nand ( n61936 , n61935 , n58908 );
nand ( n61937 , n61930 , n61936 );
or ( n61938 , n61547 , n61555 );
not ( n61939 , n61416 );
and ( n61940 , n61939 , n46037 );
and ( n61941 , n61416 , n54721 );
nor ( n61942 , n61940 , n61941 );
or ( n61943 , n61942 , n60806 );
nand ( n61944 , n61938 , n61943 );
xor ( n61945 , n61937 , n61944 );
not ( n61946 , n50078 );
buf ( n61947 , n49766 );
not ( n61948 , n61947 );
not ( n61949 , n40691 );
or ( n61950 , n61948 , n61949 );
buf ( n61951 , n49618 );
not ( n61952 , n61951 );
or ( n61953 , n40691 , n61952 );
nand ( n61954 , n61950 , n61953 );
not ( n61955 , n61954 );
or ( n61956 , n61946 , n61955 );
nand ( n61957 , n61277 , n52736 );
nand ( n61958 , n61956 , n61957 );
xor ( n61959 , n61945 , n61958 );
not ( n61960 , n61470 );
not ( n61961 , n58961 );
not ( n61962 , n61961 );
or ( n61963 , n61960 , n61962 );
not ( n61964 , n48898 );
not ( n61965 , n58433 );
or ( n61966 , n61964 , n61965 );
nand ( n61967 , n58642 , n48897 );
nand ( n61968 , n61966 , n61967 );
nand ( n61969 , n61968 , n58638 );
nand ( n61970 , n61963 , n61969 );
not ( n61971 , n61482 );
not ( n61972 , n55887 );
or ( n61973 , n61971 , n61972 );
not ( n61974 , n54611 );
not ( n61975 , n59496 );
or ( n61976 , n61974 , n61975 );
nand ( n61977 , n55892 , n51670 );
nand ( n61978 , n61976 , n61977 );
nand ( n61979 , n61978 , n55459 );
nand ( n61980 , n61973 , n61979 );
xor ( n61981 , n61970 , n61980 );
or ( n61982 , n60960 , n61401 );
and ( n61983 , n60285 , n47650 );
not ( n61984 , n60285 );
and ( n61985 , n61984 , n47646 );
or ( n61986 , n61983 , n61985 );
not ( n61987 , n61986 );
or ( n61988 , n61987 , n60963 );
nand ( n61989 , n61982 , n61988 );
xor ( n61990 , n61981 , n61989 );
xor ( n61991 , n61959 , n61990 );
not ( n61992 , n61509 );
not ( n61993 , n55143 );
or ( n61994 , n61992 , n61993 );
and ( n61995 , n48983 , n58108 );
not ( n61996 , n48983 );
and ( n61997 , n61996 , n61507 );
or ( n61998 , n61995 , n61997 );
nand ( n61999 , n61998 , n55933 );
nand ( n62000 , n61994 , n61999 );
not ( n62001 , n61520 );
not ( n62002 , n56776 );
or ( n62003 , n62001 , n62002 );
not ( n62004 , n51792 );
not ( n62005 , n56785 );
or ( n62006 , n62004 , n62005 );
nand ( n62007 , n61518 , n53126 );
nand ( n62008 , n62006 , n62007 );
nand ( n62009 , n56780 , n62008 );
nand ( n62010 , n62003 , n62009 );
xor ( n62011 , n62000 , n62010 );
not ( n62012 , n61459 );
not ( n62013 , n59432 );
or ( n62014 , n62012 , n62013 );
not ( n62015 , n51204 );
not ( n62016 , n57534 );
or ( n62017 , n62015 , n62016 );
nand ( n62018 , n57619 , n48860 );
nand ( n62019 , n62017 , n62018 );
nand ( n62020 , n62019 , n57631 );
nand ( n62021 , n62014 , n62020 );
xor ( n62022 , n62011 , n62021 );
xor ( n62023 , n61991 , n62022 );
xor ( n62024 , n61959 , n61990 );
and ( n62025 , n62024 , n62022 );
and ( n62026 , n61959 , n61990 );
or ( n62027 , n62025 , n62026 );
not ( n62028 , n61325 );
not ( n62029 , n52852 );
or ( n62030 , n62028 , n62029 );
not ( n62031 , n41668 );
not ( n62032 , n53946 );
or ( n62033 , n62031 , n62032 );
nand ( n62034 , n58144 , n48118 );
nand ( n62035 , n62033 , n62034 );
nand ( n62036 , n62035 , n52468 );
nand ( n62037 , n62030 , n62036 );
not ( n62038 , n61336 );
not ( n62039 , n55913 );
or ( n62040 , n62038 , n62039 );
not ( n62041 , n58180 );
not ( n62042 , n55917 );
or ( n62043 , n62041 , n62042 );
nand ( n62044 , n53590 , n41416 );
nand ( n62045 , n62043 , n62044 );
nand ( n62046 , n62045 , n53619 );
nand ( n62047 , n62040 , n62046 );
xor ( n62048 , n62037 , n62047 );
not ( n62049 , n61498 );
not ( n62050 , n54315 );
or ( n62051 , n62049 , n62050 );
not ( n62052 , n57182 );
not ( n62053 , n54467 );
or ( n62054 , n62052 , n62053 );
nand ( n62055 , n54298 , n47332 );
nand ( n62056 , n62054 , n62055 );
nand ( n62057 , n62056 , n54077 );
nand ( n62058 , n62051 , n62057 );
xor ( n62059 , n62048 , n62058 );
xor ( n62060 , n62059 , n61765 );
xor ( n62061 , n62060 , n61769 );
xor ( n62062 , n62059 , n61765 );
and ( n62063 , n62062 , n61769 );
and ( n62064 , n62059 , n61765 );
or ( n62065 , n62063 , n62064 );
xor ( n62066 , n61773 , n61373 );
not ( n62067 , n59633 );
not ( n62068 , n61672 );
or ( n62069 , n62067 , n62068 );
and ( n62070 , n40626 , n52728 );
not ( n62071 , n40626 );
and ( n62072 , n62071 , n60602 );
or ( n62073 , n62070 , n62072 );
nand ( n62074 , n62073 , n52723 );
nand ( n62075 , n62069 , n62074 );
not ( n62076 , n60927 );
not ( n62077 , n60289 );
not ( n62078 , n62077 );
not ( n62079 , n53259 );
or ( n62080 , n62078 , n62079 );
nand ( n62081 , n57332 , n60289 );
nand ( n62082 , n62080 , n62081 );
not ( n62083 , n62082 );
or ( n62084 , n62076 , n62083 );
buf ( n62085 , n58168 );
nand ( n62086 , n61591 , n62085 );
nand ( n62087 , n62084 , n62086 );
xor ( n62088 , n62075 , n62087 );
not ( n62089 , n51157 );
not ( n62090 , n61601 );
or ( n62091 , n62089 , n62090 );
not ( n62092 , n50263 );
not ( n62093 , n58933 );
or ( n62094 , n62092 , n62093 );
nand ( n62095 , n60905 , n52080 );
nand ( n62096 , n62094 , n62095 );
nand ( n62097 , n62096 , n47827 );
nand ( n62098 , n62091 , n62097 );
xor ( n62099 , n62088 , n62098 );
xor ( n62100 , n62066 , n62099 );
xor ( n62101 , n61773 , n61373 );
and ( n62102 , n62101 , n62099 );
and ( n62103 , n61773 , n61373 );
or ( n62104 , n62102 , n62103 );
xor ( n62105 , n61777 , n61781 );
not ( n62106 , n47873 );
not ( n62107 , n61652 );
or ( n62108 , n62106 , n62107 );
and ( n62109 , n40376 , n51684 );
not ( n62110 , n40376 );
and ( n62111 , n62110 , n51680 );
or ( n62112 , n62109 , n62111 );
nand ( n62113 , n62112 , n54623 );
nand ( n62114 , n62108 , n62113 );
not ( n62115 , n51865 );
not ( n62116 , n49707 );
not ( n62117 , n56451 );
or ( n62118 , n62116 , n62117 );
nand ( n62119 , n40012 , n52273 );
nand ( n62120 , n62118 , n62119 );
not ( n62121 , n62120 );
or ( n62122 , n62115 , n62121 );
nand ( n62123 , n61629 , n49713 );
nand ( n62124 , n62122 , n62123 );
xor ( n62125 , n62114 , n62124 );
not ( n62126 , n56639 );
not ( n62127 , n59345 );
not ( n62128 , n61139 );
or ( n62129 , n62127 , n62128 );
nand ( n62130 , n51912 , n60617 );
nand ( n62131 , n62129 , n62130 );
not ( n62132 , n62131 );
or ( n62133 , n62126 , n62132 );
nand ( n62134 , n61583 , n59950 );
nand ( n62135 , n62133 , n62134 );
xor ( n62136 , n62125 , n62135 );
xor ( n62137 , n62105 , n62136 );
xor ( n62138 , n61777 , n61781 );
and ( n62139 , n62138 , n62136 );
and ( n62140 , n61777 , n61781 );
or ( n62141 , n62139 , n62140 );
not ( n62142 , n52970 );
not ( n62143 , n61568 );
or ( n62144 , n62142 , n62143 );
not ( n62145 , n48645 );
not ( n62146 , n59134 );
or ( n62147 , n62145 , n62146 );
nand ( n62148 , n40451 , n52048 );
nand ( n62149 , n62147 , n62148 );
nand ( n62150 , n62149 , n52043 );
nand ( n62151 , n62144 , n62150 );
not ( n62152 , n52421 );
not ( n62153 , n61619 );
or ( n62154 , n62152 , n62153 );
and ( n62155 , n40388 , n53228 );
not ( n62156 , n40388 );
and ( n62157 , n62156 , n51723 );
or ( n62158 , n62155 , n62157 );
nand ( n62159 , n62158 , n47148 );
nand ( n62160 , n62154 , n62159 );
xor ( n62161 , n62151 , n62160 );
not ( n62162 , n57314 );
not ( n62163 , n61638 );
or ( n62164 , n62162 , n62163 );
not ( n62165 , n52377 );
not ( n62166 , n54810 );
or ( n62167 , n62165 , n62166 );
nand ( n62168 , n40363 , n53973 );
nand ( n62169 , n62167 , n62168 );
nand ( n62170 , n62169 , n52004 );
nand ( n62171 , n62164 , n62170 );
xor ( n62172 , n62161 , n62171 );
xor ( n62173 , n62172 , n61923 );
xor ( n62174 , n61307 , n61345 );
xor ( n62175 , n62174 , n61705 );
xor ( n62176 , n62173 , n62175 );
xor ( n62177 , n62172 , n61923 );
and ( n62178 , n62177 , n62175 );
and ( n62179 , n62172 , n61923 );
or ( n62180 , n62178 , n62179 );
xor ( n62181 , n61868 , n61895 );
xor ( n62182 , n62181 , n61396 );
xor ( n62183 , n61868 , n61895 );
and ( n62184 , n62183 , n61396 );
and ( n62185 , n61868 , n61895 );
or ( n62186 , n62184 , n62185 );
xor ( n62187 , n61490 , n62023 );
xor ( n62188 , n62187 , n61576 );
xor ( n62189 , n61490 , n62023 );
and ( n62190 , n62189 , n61576 );
and ( n62191 , n61490 , n62023 );
or ( n62192 , n62190 , n62191 );
xor ( n62193 , n62037 , n62047 );
and ( n62194 , n62193 , n62058 );
and ( n62195 , n62037 , n62047 );
or ( n62196 , n62194 , n62195 );
xor ( n62197 , n61529 , n61681 );
xor ( n62198 , n62197 , n61612 );
xor ( n62199 , n61529 , n61681 );
and ( n62200 , n62199 , n61612 );
and ( n62201 , n61529 , n61681 );
or ( n62202 , n62200 , n62201 );
xor ( n62203 , n62061 , n61689 );
xor ( n62204 , n62203 , n62100 );
xor ( n62205 , n62061 , n61689 );
and ( n62206 , n62205 , n62100 );
and ( n62207 , n62061 , n61689 );
or ( n62208 , n62206 , n62207 );
xor ( n62209 , n62137 , n61695 );
xor ( n62210 , n62209 , n62182 );
xor ( n62211 , n62137 , n61695 );
and ( n62212 , n62211 , n62182 );
and ( n62213 , n62137 , n61695 );
or ( n62214 , n62212 , n62213 );
xor ( n62215 , n62176 , n62188 );
xor ( n62216 , n62215 , n61701 );
xor ( n62217 , n62176 , n62188 );
and ( n62218 , n62217 , n61701 );
and ( n62219 , n62176 , n62188 );
or ( n62220 , n62218 , n62219 );
xor ( n62221 , n62198 , n61711 );
xor ( n62222 , n62221 , n62204 );
xor ( n62223 , n62198 , n61711 );
and ( n62224 , n62223 , n62204 );
and ( n62225 , n62198 , n61711 );
or ( n62226 , n62224 , n62225 );
xor ( n62227 , n61717 , n61723 );
xor ( n62228 , n62227 , n62210 );
xor ( n62229 , n61717 , n61723 );
and ( n62230 , n62229 , n62210 );
and ( n62231 , n61717 , n61723 );
or ( n62232 , n62230 , n62231 );
xor ( n62233 , n61729 , n62216 );
xor ( n62234 , n62233 , n62222 );
xor ( n62235 , n61729 , n62216 );
and ( n62236 , n62235 , n62222 );
and ( n62237 , n61729 , n62216 );
or ( n62238 , n62236 , n62237 );
xor ( n62239 , n61735 , n62228 );
xor ( n62240 , n62239 , n61741 );
xor ( n62241 , n61735 , n62228 );
and ( n62242 , n62241 , n61741 );
and ( n62243 , n61735 , n62228 );
or ( n62244 , n62242 , n62243 );
xor ( n62245 , n62234 , n61747 );
xor ( n62246 , n62245 , n62240 );
xor ( n62247 , n62234 , n61747 );
and ( n62248 , n62247 , n62240 );
and ( n62249 , n62234 , n61747 );
or ( n62250 , n62248 , n62249 );
xor ( n62251 , n62000 , n62010 );
and ( n62252 , n62251 , n62021 );
and ( n62253 , n62000 , n62010 );
or ( n62254 , n62252 , n62253 );
xor ( n62255 , n61970 , n61980 );
and ( n62256 , n62255 , n61989 );
and ( n62257 , n61970 , n61980 );
or ( n62258 , n62256 , n62257 );
xor ( n62259 , n61937 , n61944 );
and ( n62260 , n62259 , n61958 );
and ( n62261 , n61937 , n61944 );
or ( n62262 , n62260 , n62261 );
xor ( n62263 , n62151 , n62160 );
and ( n62264 , n62263 , n62171 );
and ( n62265 , n62151 , n62160 );
or ( n62266 , n62264 , n62265 );
xor ( n62267 , n62114 , n62124 );
and ( n62268 , n62267 , n62135 );
and ( n62269 , n62114 , n62124 );
or ( n62270 , n62268 , n62269 );
xor ( n62271 , n62075 , n62087 );
and ( n62272 , n62271 , n62098 );
and ( n62273 , n62075 , n62087 );
or ( n62274 , n62272 , n62273 );
xor ( n62275 , n61307 , n61345 );
and ( n62276 , n62275 , n61705 );
and ( n62277 , n61307 , n61345 );
or ( n62278 , n62276 , n62277 );
not ( n62279 , n61823 );
not ( n62280 , n50911 );
or ( n62281 , n62279 , n62280 );
not ( n62282 , n50827 );
not ( n62283 , n50916 );
or ( n62284 , n62282 , n62283 );
nand ( n62285 , n51465 , n49806 );
nand ( n62286 , n62284 , n62285 );
nand ( n62287 , n62286 , n51223 );
nand ( n62288 , n62281 , n62287 );
not ( n62289 , n61837 );
not ( n62290 , n53170 );
or ( n62291 , n62289 , n62290 );
not ( n62292 , n51566 );
not ( n62293 , n53706 );
or ( n62294 , n62292 , n62293 );
nand ( n62295 , n53549 , n41216 );
nand ( n62296 , n62294 , n62295 );
nand ( n62297 , n62296 , n55066 );
nand ( n62298 , n62291 , n62297 );
xor ( n62299 , n62288 , n62298 );
not ( n62300 , n61849 );
or ( n62301 , n52481 , n62300 );
not ( n62302 , n51766 );
not ( n62303 , n51476 );
not ( n62304 , n52130 );
or ( n62305 , n62303 , n62304 );
nand ( n62306 , n53917 , n48679 );
nand ( n62307 , n62305 , n62306 );
not ( n62308 , n62307 );
or ( n62309 , n62302 , n62308 );
nand ( n62310 , n62301 , n62309 );
xor ( n62311 , n62299 , n62310 );
xor ( n62312 , n62288 , n62298 );
and ( n62313 , n62312 , n62310 );
and ( n62314 , n62288 , n62298 );
or ( n62315 , n62313 , n62314 );
not ( n62316 , n62035 );
not ( n62317 , n52853 );
or ( n62318 , n62316 , n62317 );
not ( n62319 , n49233 );
not ( n62320 , n62319 );
not ( n62321 , n52837 );
or ( n62322 , n62320 , n62321 );
nand ( n62323 , n52840 , n49233 );
nand ( n62324 , n62322 , n62323 );
nand ( n62325 , n53571 , n62324 );
nand ( n62326 , n62318 , n62325 );
not ( n62327 , n62045 );
not ( n62328 , n53609 );
or ( n62329 , n62327 , n62328 );
not ( n62330 , n58458 );
not ( n62331 , n53591 );
or ( n62332 , n62330 , n62331 );
nand ( n62333 , n55089 , n58459 );
nand ( n62334 , n62332 , n62333 );
nand ( n62335 , n62334 , n53326 );
nand ( n62336 , n62329 , n62335 );
xor ( n62337 , n62326 , n62336 );
not ( n62338 , n56810 );
not ( n62339 , n62056 );
or ( n62340 , n62338 , n62339 );
not ( n62341 , n47527 );
not ( n62342 , n54467 );
or ( n62343 , n62341 , n62342 );
nand ( n62344 , n54297 , n59388 );
nand ( n62345 , n62343 , n62344 );
not ( n62346 , n62345 );
or ( n62347 , n55866 , n62346 );
nand ( n62348 , n62340 , n62347 );
xor ( n62349 , n62337 , n62348 );
xor ( n62350 , n62326 , n62336 );
and ( n62351 , n62350 , n62348 );
and ( n62352 , n62326 , n62336 );
or ( n62353 , n62351 , n62352 );
xor ( n62354 , n62254 , n62258 );
not ( n62355 , n53675 );
not ( n62356 , n47803 );
not ( n62357 , n58485 );
not ( n62358 , n62357 );
or ( n62359 , n62356 , n62358 );
nand ( n62360 , n39680 , n50634 );
nand ( n62361 , n62359 , n62360 );
not ( n62362 , n62361 );
or ( n62363 , n62355 , n62362 );
nand ( n62364 , n61880 , n47407 );
nand ( n62365 , n62363 , n62364 );
xor ( n62366 , n62354 , n62365 );
xor ( n62367 , n62254 , n62258 );
and ( n62368 , n62367 , n62365 );
and ( n62369 , n62254 , n62258 );
or ( n62370 , n62368 , n62369 );
not ( n62371 , n48989 );
not ( n62372 , n61890 );
or ( n62373 , n62371 , n62372 );
or ( n62374 , n49500 , n39893 );
nand ( n62375 , n39893 , n49500 );
nand ( n62376 , n62374 , n62375 );
nand ( n62377 , n62376 , n53510 );
nand ( n62378 , n62373 , n62377 );
not ( n62379 , n46602 );
not ( n62380 , n46072 );
not ( n62381 , n42397 );
not ( n62382 , n62381 );
or ( n62383 , n62380 , n62382 );
not ( n62384 , n42398 );
nand ( n62385 , n62384 , n50405 );
nand ( n62386 , n62383 , n62385 );
not ( n62387 , n62386 );
or ( n62388 , n62379 , n62387 );
nand ( n62389 , n61909 , n50659 );
nand ( n62390 , n62388 , n62389 );
xor ( n62391 , n62378 , n62390 );
not ( n62392 , n49026 );
not ( n62393 , n46425 );
buf ( n62394 , n61347 );
not ( n62395 , n62394 );
or ( n62396 , n62393 , n62395 );
or ( n62397 , n60357 , n46425 );
nand ( n62398 , n62396 , n62397 );
not ( n62399 , n62398 );
or ( n62400 , n62392 , n62399 );
nand ( n62401 , n61919 , n46267 );
nand ( n62402 , n62400 , n62401 );
xor ( n62403 , n62391 , n62402 );
xor ( n62404 , n62378 , n62390 );
and ( n62405 , n62404 , n62402 );
and ( n62406 , n62378 , n62390 );
or ( n62407 , n62405 , n62406 );
xor ( n62408 , n62262 , n62311 );
not ( n62409 , n61986 );
not ( n62410 , n60424 );
or ( n62411 , n62409 , n62410 );
not ( n62412 , n49734 );
not ( n62413 , n60968 );
or ( n62414 , n62412 , n62413 );
nand ( n62415 , n60285 , n47821 );
nand ( n62416 , n62414 , n62415 );
nand ( n62417 , n60427 , n62416 );
nand ( n62418 , n62411 , n62417 );
not ( n62419 , n61942 );
not ( n62420 , n62419 );
not ( n62421 , n61548 );
or ( n62422 , n62420 , n62421 );
not ( n62423 , n46273 );
not ( n62424 , n61939 );
or ( n62425 , n62423 , n62424 );
nand ( n62426 , n61416 , n46824 );
nand ( n62427 , n62425 , n62426 );
not ( n62428 , n60806 );
nand ( n62429 , n62427 , n62428 );
nand ( n62430 , n62422 , n62429 );
xor ( n62431 , n62418 , n62430 );
not ( n62432 , n37639 );
not ( n62433 , n37544 );
nand ( n62434 , n62433 , n37067 );
nor ( n62435 , n36697 , n37544 );
nand ( n62436 , n62435 , n36287 );
not ( n62437 , n36547 );
not ( n62438 , n37543 );
or ( n62439 , n62437 , n62438 );
nand ( n62440 , n62439 , n37501 );
not ( n62441 , n62440 );
nand ( n62442 , n62434 , n62436 , n62441 );
not ( n62443 , n62442 );
or ( n62444 , n62432 , n62443 );
not ( n62445 , n37639 );
nand ( n62446 , n62434 , n62441 , n62436 , n62445 );
nand ( n62447 , n62444 , n62446 );
buf ( n62448 , n62447 );
buf ( n62449 , n62448 );
or ( n62450 , n62449 , n46441 );
buf ( n62451 , n62448 );
not ( n62452 , n62451 );
or ( n62453 , n62452 , n48689 );
nand ( n62454 , n62450 , n62453 );
not ( n62455 , n62454 );
not ( n62456 , n62447 );
not ( n62457 , n62456 );
not ( n62458 , n61805 );
or ( n62459 , n62457 , n62458 );
nand ( n62460 , n62448 , n61811 );
nand ( n62461 , n62459 , n62460 );
nor ( n62462 , n61813 , n62461 );
buf ( n62463 , n62462 );
not ( n62464 , n62463 );
or ( n62465 , n62455 , n62464 );
not ( n62466 , n61813 );
not ( n62467 , n62466 );
not ( n62468 , n50914 );
not ( n62469 , n62452 );
or ( n62470 , n62468 , n62469 );
nand ( n62471 , n62451 , n48766 );
nand ( n62472 , n62470 , n62471 );
nand ( n62473 , n62467 , n62472 );
nand ( n62474 , n62465 , n62473 );
xor ( n62475 , n62431 , n62474 );
xor ( n62476 , n62408 , n62475 );
xor ( n62477 , n62262 , n62311 );
and ( n62478 , n62477 , n62475 );
and ( n62479 , n62262 , n62311 );
or ( n62480 , n62478 , n62479 );
not ( n62481 , n62019 );
not ( n62482 , n59432 );
or ( n62483 , n62481 , n62482 );
not ( n62484 , n49624 );
not ( n62485 , n57619 );
not ( n62486 , n62485 );
or ( n62487 , n62484 , n62486 );
nand ( n62488 , n57619 , n49630 );
nand ( n62489 , n62487 , n62488 );
nand ( n62490 , n62489 , n59435 );
nand ( n62491 , n62483 , n62490 );
not ( n62492 , n61968 );
not ( n62493 , n61961 );
or ( n62494 , n62492 , n62493 );
not ( n62495 , n47765 );
not ( n62496 , n58630 );
not ( n62497 , n62496 );
not ( n62498 , n62497 );
or ( n62499 , n62495 , n62498 );
nand ( n62500 , n58642 , n48589 );
nand ( n62501 , n62499 , n62500 );
nand ( n62502 , n61465 , n62501 );
nand ( n62503 , n62494 , n62502 );
xor ( n62504 , n62491 , n62503 );
not ( n62505 , n61935 );
not ( n62506 , n60538 );
not ( n62507 , n62506 );
or ( n62508 , n62505 , n62507 );
not ( n62509 , n49654 );
not ( n62510 , n59338 );
not ( n62511 , n62510 );
or ( n62512 , n62509 , n62511 );
buf ( n62513 , n59337 );
nand ( n62514 , n62513 , n47368 );
nand ( n62515 , n62512 , n62514 );
nand ( n62516 , n59575 , n62515 );
nand ( n62517 , n62508 , n62516 );
xor ( n62518 , n62504 , n62517 );
xor ( n62519 , n62518 , n62349 );
not ( n62520 , n61998 );
not ( n62521 , n55143 );
or ( n62522 , n62520 , n62521 );
not ( n62523 , n56727 );
not ( n62524 , n55148 );
or ( n62525 , n62523 , n62524 );
not ( n62526 , n58108 );
nand ( n62527 , n62526 , n47511 );
nand ( n62528 , n62525 , n62527 );
nand ( n62529 , n62528 , n54848 );
nand ( n62530 , n62522 , n62529 );
not ( n62531 , n61978 );
not ( n62532 , n56281 );
or ( n62533 , n62531 , n62532 );
not ( n62534 , n47158 );
not ( n62535 , n58604 );
or ( n62536 , n62534 , n62535 );
nand ( n62537 , n55872 , n54184 );
nand ( n62538 , n62536 , n62537 );
nand ( n62539 , n62538 , n55459 );
nand ( n62540 , n62533 , n62539 );
xor ( n62541 , n62530 , n62540 );
not ( n62542 , n62008 );
not ( n62543 , n56777 );
or ( n62544 , n62542 , n62543 );
not ( n62545 , n52033 );
not ( n62546 , n57665 );
or ( n62547 , n62545 , n62546 );
nand ( n62548 , n57664 , n52038 );
nand ( n62549 , n62547 , n62548 );
nand ( n62550 , n60472 , n62549 );
nand ( n62551 , n62544 , n62550 );
xor ( n62552 , n62541 , n62551 );
xor ( n62553 , n62519 , n62552 );
xor ( n62554 , n62518 , n62349 );
and ( n62555 , n62554 , n62552 );
and ( n62556 , n62518 , n62349 );
or ( n62557 , n62555 , n62556 );
xor ( n62558 , n62266 , n62270 );
xor ( n62559 , n62558 , n61872 );
xor ( n62560 , n62266 , n62270 );
and ( n62561 , n62560 , n61872 );
and ( n62562 , n62266 , n62270 );
or ( n62563 , n62561 , n62562 );
not ( n62564 , n54623 );
and ( n62565 , n54432 , n51684 );
not ( n62566 , n54432 );
and ( n62567 , n62566 , n51680 );
or ( n62568 , n62565 , n62567 );
not ( n62569 , n62568 );
or ( n62570 , n62564 , n62569 );
nand ( n62571 , n52022 , n62112 );
nand ( n62572 , n62570 , n62571 );
not ( n62573 , n52723 );
not ( n62574 , n58982 );
not ( n62575 , n55190 );
or ( n62576 , n62574 , n62575 );
not ( n62577 , n58982 );
nand ( n62578 , n40635 , n62577 );
nand ( n62579 , n62576 , n62578 );
not ( n62580 , n62579 );
or ( n62581 , n62573 , n62580 );
nand ( n62582 , n62073 , n59633 );
nand ( n62583 , n62581 , n62582 );
xor ( n62584 , n62572 , n62583 );
not ( n62585 , n56639 );
not ( n62586 , n59345 );
not ( n62587 , n54377 );
or ( n62588 , n62586 , n62587 );
nand ( n62589 , n52212 , n60617 );
nand ( n62590 , n62588 , n62589 );
not ( n62591 , n62590 );
or ( n62592 , n62585 , n62591 );
nand ( n62593 , n62131 , n59950 );
nand ( n62594 , n62592 , n62593 );
xor ( n62595 , n62584 , n62594 );
xor ( n62596 , n62595 , n62274 );
xor ( n62597 , n62596 , n62278 );
xor ( n62598 , n62595 , n62274 );
and ( n62599 , n62598 , n62278 );
and ( n62600 , n62595 , n62274 );
or ( n62601 , n62599 , n62600 );
not ( n62602 , n54875 );
not ( n62603 , n51723 );
not ( n62604 , n56058 );
or ( n62605 , n62603 , n62604 );
nand ( n62606 , n55203 , n51724 );
nand ( n62607 , n62605 , n62606 );
not ( n62608 , n62607 );
or ( n62609 , n62602 , n62608 );
nand ( n62610 , n62158 , n52421 );
nand ( n62611 , n62609 , n62610 );
not ( n62612 , n49713 );
not ( n62613 , n62120 );
or ( n62614 , n62612 , n62613 );
not ( n62615 , n49707 );
not ( n62616 , n59651 );
or ( n62617 , n62615 , n62616 );
not ( n62618 , n59651 );
nand ( n62619 , n62618 , n51351 );
nand ( n62620 , n62617 , n62619 );
nand ( n62621 , n62620 , n51865 );
nand ( n62622 , n62614 , n62621 );
xor ( n62623 , n62611 , n62622 );
not ( n62624 , n52004 );
not ( n62625 , n52377 );
buf ( n62626 , n40148 );
not ( n62627 , n62626 );
or ( n62628 , n62625 , n62627 );
nand ( n62629 , n40149 , n53973 );
nand ( n62630 , n62628 , n62629 );
not ( n62631 , n62630 );
or ( n62632 , n62624 , n62631 );
nand ( n62633 , n62169 , n48894 );
nand ( n62634 , n62632 , n62633 );
xor ( n62635 , n62623 , n62634 );
xor ( n62636 , n61899 , n62635 );
nand ( n62637 , n61811 , n46440 );
not ( n62638 , n46441 );
not ( n62639 , n61805 );
or ( n62640 , n62638 , n62639 );
nand ( n62641 , n62640 , n61416 );
and ( n62642 , n62637 , n62451 , n62641 );
not ( n62643 , n52757 );
not ( n62644 , n50306 );
not ( n62645 , n53513 );
or ( n62646 , n62644 , n62645 );
nand ( n62647 , n50404 , n50943 );
nand ( n62648 , n62646 , n62647 );
not ( n62649 , n62648 );
or ( n62650 , n62643 , n62649 );
nand ( n62651 , n61787 , n50321 );
nand ( n62652 , n62650 , n62651 );
xor ( n62653 , n62642 , n62652 );
buf ( n62654 , n50078 );
not ( n62655 , n62654 );
not ( n62656 , n61951 );
not ( n62657 , n50958 );
or ( n62658 , n62656 , n62657 );
nand ( n62659 , n52284 , n61952 );
nand ( n62660 , n62658 , n62659 );
not ( n62661 , n62660 );
or ( n62662 , n62655 , n62661 );
not ( n62663 , n52058 );
not ( n62664 , n62663 );
nand ( n62665 , n61954 , n62664 );
nand ( n62666 , n62662 , n62665 );
xor ( n62667 , n62653 , n62666 );
not ( n62668 , n52962 );
not ( n62669 , n50232 );
not ( n62670 , n56020 );
or ( n62671 , n62669 , n62670 );
nand ( n62672 , n56023 , n49679 );
nand ( n62673 , n62671 , n62672 );
not ( n62674 , n62673 );
or ( n62675 , n62668 , n62674 );
nand ( n62676 , n62149 , n52970 );
nand ( n62677 , n62675 , n62676 );
xor ( n62678 , n62667 , n62677 );
xor ( n62679 , n62636 , n62678 );
xor ( n62680 , n61899 , n62635 );
and ( n62681 , n62680 , n62678 );
and ( n62682 , n61899 , n62635 );
or ( n62683 , n62681 , n62682 );
not ( n62684 , n58168 );
not ( n62685 , n62082 );
or ( n62686 , n62684 , n62685 );
not ( n62687 , n49112 );
not ( n62688 , n52894 );
or ( n62689 , n62687 , n62688 );
nand ( n62690 , n51601 , n60292 );
nand ( n62691 , n62689 , n62690 );
nand ( n62692 , n62691 , n52191 );
nand ( n62693 , n62686 , n62692 );
not ( n62694 , n47827 );
not ( n62695 , n50263 );
not ( n62696 , n59402 );
or ( n62697 , n62695 , n62696 );
nand ( n62698 , n39574 , n48078 );
nand ( n62699 , n62697 , n62698 );
not ( n62700 , n62699 );
or ( n62701 , n62694 , n62700 );
nand ( n62702 , n62096 , n51157 );
nand ( n62703 , n62701 , n62702 );
xor ( n62704 , n62693 , n62703 );
xor ( n62705 , n62704 , n61830 );
xor ( n62706 , n62705 , n62403 );
xor ( n62707 , n62706 , n62366 );
xor ( n62708 , n62705 , n62403 );
and ( n62709 , n62708 , n62366 );
and ( n62710 , n62705 , n62403 );
or ( n62711 , n62709 , n62710 );
xor ( n62712 , n61856 , n62196 );
not ( n62713 , n49832 );
not ( n62714 , n47508 );
not ( n62715 , n39253 );
not ( n62716 , n62715 );
or ( n62717 , n62714 , n62716 );
nand ( n62718 , n39253 , n47514 );
nand ( n62719 , n62717 , n62718 );
not ( n62720 , n62719 );
or ( n62721 , n62713 , n62720 );
nand ( n62722 , n61861 , n46564 );
nand ( n62723 , n62721 , n62722 );
xor ( n62724 , n62712 , n62723 );
xor ( n62725 , n62724 , n62027 );
xor ( n62726 , n62725 , n61927 );
xor ( n62727 , n62724 , n62027 );
and ( n62728 , n62727 , n61927 );
and ( n62729 , n62724 , n62027 );
or ( n62730 , n62728 , n62729 );
xor ( n62731 , n62553 , n62476 );
xor ( n62732 , n62731 , n62065 );
xor ( n62733 , n62553 , n62476 );
and ( n62734 , n62733 , n62065 );
and ( n62735 , n62553 , n62476 );
or ( n62736 , n62734 , n62735 );
xor ( n62737 , n62530 , n62540 );
and ( n62738 , n62737 , n62551 );
and ( n62739 , n62530 , n62540 );
or ( n62740 , n62738 , n62739 );
xor ( n62741 , n62141 , n62104 );
xor ( n62742 , n62741 , n62559 );
xor ( n62743 , n62141 , n62104 );
and ( n62744 , n62743 , n62559 );
and ( n62745 , n62141 , n62104 );
or ( n62746 , n62744 , n62745 );
xor ( n62747 , n62180 , n62597 );
xor ( n62748 , n62747 , n62186 );
xor ( n62749 , n62180 , n62597 );
and ( n62750 , n62749 , n62186 );
and ( n62751 , n62180 , n62597 );
or ( n62752 , n62750 , n62751 );
xor ( n62753 , n62679 , n62726 );
xor ( n62754 , n62753 , n62707 );
xor ( n62755 , n62679 , n62726 );
and ( n62756 , n62755 , n62707 );
and ( n62757 , n62679 , n62726 );
or ( n62758 , n62756 , n62757 );
xor ( n62759 , n62192 , n62202 );
xor ( n62760 , n62759 , n62732 );
xor ( n62761 , n62192 , n62202 );
and ( n62762 , n62761 , n62732 );
and ( n62763 , n62192 , n62202 );
or ( n62764 , n62762 , n62763 );
xor ( n62765 , n62742 , n62208 );
xor ( n62766 , n62765 , n62748 );
xor ( n62767 , n62742 , n62208 );
and ( n62768 , n62767 , n62748 );
and ( n62769 , n62742 , n62208 );
or ( n62770 , n62768 , n62769 );
xor ( n62771 , n62214 , n62220 );
xor ( n62772 , n62771 , n62754 );
xor ( n62773 , n62214 , n62220 );
and ( n62774 , n62773 , n62754 );
and ( n62775 , n62214 , n62220 );
or ( n62776 , n62774 , n62775 );
xor ( n62777 , n62760 , n62226 );
xor ( n62778 , n62777 , n62766 );
xor ( n62779 , n62760 , n62226 );
and ( n62780 , n62779 , n62766 );
and ( n62781 , n62760 , n62226 );
or ( n62782 , n62780 , n62781 );
xor ( n62783 , n62232 , n62772 );
xor ( n62784 , n62783 , n62238 );
xor ( n62785 , n62232 , n62772 );
and ( n62786 , n62785 , n62238 );
and ( n62787 , n62232 , n62772 );
or ( n62788 , n62786 , n62787 );
xor ( n62789 , n62778 , n62784 );
xor ( n62790 , n62789 , n62244 );
xor ( n62791 , n62778 , n62784 );
and ( n62792 , n62791 , n62244 );
and ( n62793 , n62778 , n62784 );
or ( n62794 , n62792 , n62793 );
xor ( n62795 , n62491 , n62503 );
and ( n62796 , n62795 , n62517 );
and ( n62797 , n62491 , n62503 );
or ( n62798 , n62796 , n62797 );
xor ( n62799 , n62418 , n62430 );
and ( n62800 , n62799 , n62474 );
and ( n62801 , n62418 , n62430 );
or ( n62802 , n62800 , n62801 );
xor ( n62803 , n62653 , n62666 );
and ( n62804 , n62803 , n62677 );
and ( n62805 , n62653 , n62666 );
or ( n62806 , n62804 , n62805 );
xor ( n62807 , n62611 , n62622 );
and ( n62808 , n62807 , n62634 );
and ( n62809 , n62611 , n62622 );
or ( n62810 , n62808 , n62809 );
xor ( n62811 , n62572 , n62583 );
and ( n62812 , n62811 , n62594 );
and ( n62813 , n62572 , n62583 );
or ( n62814 , n62812 , n62813 );
xor ( n62815 , n62693 , n62703 );
and ( n62816 , n62815 , n61830 );
and ( n62817 , n62693 , n62703 );
or ( n62818 , n62816 , n62817 );
xor ( n62819 , n61856 , n62196 );
and ( n62820 , n62819 , n62723 );
and ( n62821 , n61856 , n62196 );
or ( n62822 , n62820 , n62821 );
not ( n62823 , n37541 );
nand ( n62824 , n37067 , n62823 );
nor ( n62825 , n61795 , n37541 );
nand ( n62826 , n61793 , n62825 );
and ( n62827 , n37540 , n36547 );
nor ( n62828 , n62827 , n37495 );
nand ( n62829 , n62824 , n62826 , n62828 );
not ( n62830 , n37507 );
nand ( n62831 , n62830 , n37379 );
not ( n62832 , n62831 );
and ( n62833 , n62829 , n62832 );
not ( n62834 , n62829 );
and ( n62835 , n62834 , n62831 );
nor ( n62836 , n62833 , n62835 );
not ( n62837 , n62836 );
or ( n62838 , n62456 , n62837 );
not ( n62839 , n62836 );
not ( n62840 , n62447 );
nand ( n62841 , n62839 , n62840 );
nand ( n62842 , n62838 , n62841 );
not ( n62843 , n62842 );
and ( n62844 , n62843 , n48689 );
not ( n62845 , n62286 );
not ( n62846 , n52526 );
or ( n62847 , n62845 , n62846 );
and ( n62848 , n41036 , n57187 );
not ( n62849 , n41036 );
and ( n62850 , n62849 , n50946 );
nor ( n62851 , n62848 , n62850 );
nand ( n62852 , n62851 , n51223 );
nand ( n62853 , n62847 , n62852 );
xor ( n62854 , n62844 , n62853 );
not ( n62855 , n62296 );
or ( n62856 , n58189 , n62855 );
not ( n62857 , n49549 );
not ( n62858 , n56361 );
not ( n62859 , n62858 );
or ( n62860 , n62857 , n62859 );
not ( n62861 , n51740 );
nand ( n62862 , n62861 , n52816 );
nand ( n62863 , n62860 , n62862 );
not ( n62864 , n62863 );
or ( n62865 , n51146 , n62864 );
nand ( n62866 , n62856 , n62865 );
xor ( n62867 , n62854 , n62866 );
xor ( n62868 , n62844 , n62853 );
and ( n62869 , n62868 , n62866 );
and ( n62870 , n62844 , n62853 );
or ( n62871 , n62869 , n62870 );
not ( n62872 , n62307 );
not ( n62873 , n52125 );
or ( n62874 , n62872 , n62873 );
not ( n62875 , n52592 );
not ( n62876 , n52109 );
or ( n62877 , n62875 , n62876 );
nand ( n62878 , n52870 , n52589 );
nand ( n62879 , n62877 , n62878 );
nand ( n62880 , n51766 , n62879 );
nand ( n62881 , n62874 , n62880 );
not ( n62882 , n62324 );
not ( n62883 , n52853 );
or ( n62884 , n62882 , n62883 );
not ( n62885 , n41407 );
not ( n62886 , n55102 );
or ( n62887 , n62885 , n62886 );
nand ( n62888 , n52835 , n48483 );
nand ( n62889 , n62887 , n62888 );
nand ( n62890 , n52469 , n62889 );
nand ( n62891 , n62884 , n62890 );
xor ( n62892 , n62881 , n62891 );
not ( n62893 , n62334 );
or ( n62894 , n61329 , n62893 );
not ( n62895 , n41668 );
not ( n62896 , n53594 );
or ( n62897 , n62895 , n62896 );
nand ( n62898 , n53589 , n49029 );
nand ( n62899 , n62897 , n62898 );
not ( n62900 , n62899 );
or ( n62901 , n53618 , n62900 );
nand ( n62902 , n62894 , n62901 );
xor ( n62903 , n62892 , n62902 );
xor ( n62904 , n62881 , n62891 );
and ( n62905 , n62904 , n62902 );
and ( n62906 , n62881 , n62891 );
or ( n62907 , n62905 , n62906 );
not ( n62908 , n47508 );
not ( n62909 , n61907 );
not ( n62910 , n62909 );
or ( n62911 , n62908 , n62910 );
not ( n62912 , n61904 );
buf ( n62913 , n62912 );
nand ( n62914 , n62913 , n52990 );
nand ( n62915 , n62911 , n62914 );
not ( n62916 , n62915 );
not ( n62917 , n49832 );
or ( n62918 , n62916 , n62917 );
nand ( n62919 , n62719 , n46564 );
nand ( n62920 , n62918 , n62919 );
xor ( n62921 , n62920 , n62740 );
xor ( n62922 , n62921 , n62798 );
xor ( n62923 , n62920 , n62740 );
and ( n62924 , n62923 , n62798 );
and ( n62925 , n62920 , n62740 );
or ( n62926 , n62924 , n62925 );
not ( n62927 , n47407 );
not ( n62928 , n62361 );
or ( n62929 , n62927 , n62928 );
not ( n62930 , n51545 );
not ( n62931 , n39714 );
not ( n62932 , n62931 );
or ( n62933 , n62930 , n62932 );
nand ( n62934 , n60905 , n48727 );
nand ( n62935 , n62933 , n62934 );
nand ( n62936 , n62935 , n53675 );
nand ( n62937 , n62929 , n62936 );
xor ( n62938 , n62802 , n62937 );
not ( n62939 , n62376 );
not ( n62940 , n48989 );
or ( n62941 , n62939 , n62940 );
not ( n62942 , n49500 );
not ( n62943 , n59914 );
or ( n62944 , n62942 , n62943 );
nand ( n62945 , n59913 , n53997 );
nand ( n62946 , n62944 , n62945 );
not ( n62947 , n62946 );
or ( n62948 , n62947 , n53509 );
nand ( n62949 , n62941 , n62948 );
xor ( n62950 , n62938 , n62949 );
xor ( n62951 , n62802 , n62937 );
and ( n62952 , n62951 , n62949 );
and ( n62953 , n62802 , n62937 );
or ( n62954 , n62952 , n62953 );
not ( n62955 , n46267 );
not ( n62956 , n62398 );
or ( n62957 , n62955 , n62956 );
not ( n62958 , n46425 );
not ( n62959 , n60854 );
buf ( n62960 , n62959 );
not ( n62961 , n62960 );
or ( n62962 , n62958 , n62961 );
not ( n62963 , n62959 );
nand ( n62964 , n62963 , n46422 );
nand ( n62965 , n62962 , n62964 );
nand ( n62966 , n62965 , n49026 );
nand ( n62967 , n62957 , n62966 );
not ( n62968 , n51865 );
not ( n62969 , n52267 );
not ( n62970 , n58034 );
not ( n62971 , n62970 );
or ( n62972 , n62969 , n62971 );
nand ( n62973 , n60885 , n51351 );
nand ( n62974 , n62972 , n62973 );
not ( n62975 , n62974 );
or ( n62976 , n62968 , n62975 );
nand ( n62977 , n62620 , n49713 );
nand ( n62978 , n62976 , n62977 );
xor ( n62979 , n62967 , n62978 );
xor ( n62980 , n62979 , n62903 );
xor ( n62981 , n62967 , n62978 );
and ( n62982 , n62981 , n62903 );
and ( n62983 , n62967 , n62978 );
or ( n62984 , n62982 , n62983 );
not ( n62985 , n62345 );
not ( n62986 , n56269 );
or ( n62987 , n62985 , n62986 );
not ( n62988 , n58180 );
not ( n62989 , n54467 );
or ( n62990 , n62988 , n62989 );
nand ( n62991 , n52380 , n56274 );
nand ( n62992 , n62990 , n62991 );
nand ( n62993 , n56277 , n62992 );
nand ( n62994 , n62987 , n62993 );
not ( n62995 , n62528 );
not ( n62996 , n55143 );
or ( n62997 , n62995 , n62996 );
not ( n62998 , n55118 );
not ( n62999 , n54584 );
or ( n63000 , n62998 , n62999 );
or ( n63001 , n61507 , n57186 );
nand ( n63002 , n63000 , n63001 );
nand ( n63003 , n54848 , n63002 );
nand ( n63004 , n62997 , n63003 );
xor ( n63005 , n62994 , n63004 );
not ( n63006 , n62538 );
not ( n63007 , n56281 );
or ( n63008 , n63006 , n63007 );
not ( n63009 , n48983 );
not ( n63010 , n56285 );
or ( n63011 , n63009 , n63010 );
nand ( n63012 , n55891 , n48980 );
nand ( n63013 , n63011 , n63012 );
nand ( n63014 , n55459 , n63013 );
nand ( n63015 , n63008 , n63014 );
xor ( n63016 , n63005 , n63015 );
xor ( n63017 , n62867 , n63016 );
not ( n63018 , n62515 );
not ( n63019 , n60539 );
or ( n63020 , n63018 , n63019 );
not ( n63021 , n48898 );
not ( n63022 , n62510 );
or ( n63023 , n63021 , n63022 );
nand ( n63024 , n62513 , n48897 );
nand ( n63025 , n63023 , n63024 );
nand ( n63026 , n63025 , n59931 );
nand ( n63027 , n63020 , n63026 );
not ( n63028 , n62416 );
not ( n63029 , n60960 );
not ( n63030 , n63029 );
or ( n63031 , n63028 , n63030 );
not ( n63032 , n47227 );
not ( n63033 , n60968 );
or ( n63034 , n63032 , n63033 );
nand ( n63035 , n60964 , n47589 );
nand ( n63036 , n63034 , n63035 );
nand ( n63037 , n60427 , n63036 );
nand ( n63038 , n63031 , n63037 );
xor ( n63039 , n63027 , n63038 );
not ( n63040 , n62427 );
not ( n63041 , n61550 );
or ( n63042 , n63040 , n63041 );
not ( n63043 , n47646 );
not ( n63044 , n61537 );
or ( n63045 , n63043 , n63044 );
nand ( n63046 , n61416 , n47650 );
nand ( n63047 , n63045 , n63046 );
nand ( n63048 , n62428 , n63047 );
nand ( n63049 , n63042 , n63048 );
xor ( n63050 , n63039 , n63049 );
xor ( n63051 , n63017 , n63050 );
xor ( n63052 , n62867 , n63016 );
and ( n63053 , n63052 , n63050 );
and ( n63054 , n62867 , n63016 );
or ( n63055 , n63053 , n63054 );
not ( n63056 , n62549 );
not ( n63057 , n56776 );
or ( n63058 , n63056 , n63057 );
not ( n63059 , n56679 );
not ( n63060 , n63059 );
not ( n63061 , n54611 );
or ( n63062 , n63060 , n63061 );
nand ( n63063 , n57664 , n51670 );
nand ( n63064 , n63062 , n63063 );
nand ( n63065 , n56780 , n63064 );
nand ( n63066 , n63058 , n63065 );
not ( n63067 , n62489 );
not ( n63068 , n59432 );
or ( n63069 , n63067 , n63068 );
not ( n63070 , n51792 );
not ( n63071 , n59437 );
or ( n63072 , n63070 , n63071 );
nand ( n63073 , n57619 , n53126 );
nand ( n63074 , n63072 , n63073 );
nand ( n63075 , n63074 , n59435 );
nand ( n63076 , n63069 , n63075 );
xor ( n63077 , n63066 , n63076 );
not ( n63078 , n62501 );
not ( n63079 , n58962 );
not ( n63080 , n63079 );
not ( n63081 , n63080 );
or ( n63082 , n63078 , n63081 );
not ( n63083 , n51204 );
not ( n63084 , n58966 );
or ( n63085 , n63083 , n63084 );
nand ( n63086 , n62496 , n48860 );
nand ( n63087 , n63085 , n63086 );
nand ( n63088 , n61465 , n63087 );
nand ( n63089 , n63082 , n63088 );
xor ( n63090 , n63077 , n63089 );
xor ( n63091 , n63090 , n62806 );
xor ( n63092 , n63091 , n62810 );
xor ( n63093 , n63090 , n62806 );
and ( n63094 , n63093 , n62810 );
and ( n63095 , n63090 , n62806 );
or ( n63096 , n63094 , n63095 );
not ( n63097 , n62472 );
not ( n63098 , n62463 );
or ( n63099 , n63097 , n63098 );
and ( n63100 , n46037 , n62456 );
not ( n63101 , n46037 );
and ( n63102 , n63101 , n62448 );
nor ( n63103 , n63100 , n63102 );
not ( n63104 , n63103 );
nand ( n63105 , n63104 , n62467 );
nand ( n63106 , n63099 , n63105 );
and ( n63107 , n62642 , n62652 );
xor ( n63108 , n63106 , n63107 );
not ( n63109 , n52757 );
not ( n63110 , n50304 );
not ( n63111 , n50654 );
or ( n63112 , n63110 , n63111 );
nand ( n63113 , n40692 , n50943 );
nand ( n63114 , n63112 , n63113 );
not ( n63115 , n63114 );
or ( n63116 , n63109 , n63115 );
nand ( n63117 , n62648 , n52749 );
nand ( n63118 , n63116 , n63117 );
xor ( n63119 , n63108 , n63118 );
xor ( n63120 , n62814 , n63119 );
xor ( n63121 , n63120 , n62407 );
xor ( n63122 , n62814 , n63119 );
and ( n63123 , n63122 , n62407 );
and ( n63124 , n62814 , n63119 );
or ( n63125 , n63123 , n63124 );
not ( n63126 , n60927 );
not ( n63127 , n62077 );
not ( n63128 , n52570 );
or ( n63129 , n63127 , n63128 );
not ( n63130 , n54771 );
nand ( n63131 , n63130 , n60289 );
nand ( n63132 , n63129 , n63131 );
not ( n63133 , n63132 );
or ( n63134 , n63126 , n63133 );
nand ( n63135 , n62691 , n62085 );
nand ( n63136 , n63134 , n63135 );
not ( n63137 , n62654 );
not ( n63138 , n61951 );
not ( n63139 , n51928 );
or ( n63140 , n63138 , n63139 );
nand ( n63141 , n53258 , n61947 );
nand ( n63142 , n63140 , n63141 );
not ( n63143 , n63142 );
or ( n63144 , n63137 , n63143 );
nand ( n63145 , n62660 , n52058 );
nand ( n63146 , n63144 , n63145 );
xor ( n63147 , n63136 , n63146 );
not ( n63148 , n48073 );
not ( n63149 , n50263 );
not ( n63150 , n59891 );
or ( n63151 , n63149 , n63150 );
not ( n63152 , n60874 );
nand ( n63153 , n63152 , n50087 );
nand ( n63154 , n63151 , n63153 );
not ( n63155 , n63154 );
or ( n63156 , n63148 , n63155 );
nand ( n63157 , n62699 , n51157 );
nand ( n63158 , n63156 , n63157 );
xor ( n63159 , n63147 , n63158 );
xor ( n63160 , n62822 , n63159 );
xor ( n63161 , n63160 , n62818 );
xor ( n63162 , n62822 , n63159 );
and ( n63163 , n63162 , n62818 );
and ( n63164 , n62822 , n63159 );
or ( n63165 , n63163 , n63164 );
not ( n63166 , n54875 );
not ( n63167 , n51723 );
not ( n63168 , n56411 );
or ( n63169 , n63167 , n63168 );
nand ( n63170 , n56412 , n58692 );
nand ( n63171 , n63169 , n63170 );
not ( n63172 , n63171 );
or ( n63173 , n63166 , n63172 );
nand ( n63174 , n62607 , n52421 );
nand ( n63175 , n63173 , n63174 );
not ( n63176 , n50242 );
not ( n63177 , n62673 );
or ( n63178 , n63176 , n63177 );
not ( n63179 , n48645 );
not ( n63180 , n56455 );
not ( n63181 , n63180 );
or ( n63182 , n63179 , n63181 );
nand ( n63183 , n56455 , n52048 );
nand ( n63184 , n63182 , n63183 );
nand ( n63185 , n63184 , n52962 );
nand ( n63186 , n63178 , n63185 );
xor ( n63187 , n63175 , n63186 );
not ( n63188 , n52004 );
and ( n63189 , n56438 , n52377 );
not ( n63190 , n56438 );
and ( n63191 , n63190 , n53973 );
or ( n63192 , n63189 , n63191 );
not ( n63193 , n63192 );
or ( n63194 , n63188 , n63193 );
nand ( n63195 , n62630 , n57314 );
nand ( n63196 , n63194 , n63195 );
xor ( n63197 , n63187 , n63196 );
xor ( n63198 , n62370 , n63197 );
not ( n63199 , n54623 );
not ( n63200 , n59174 );
not ( n63201 , n40364 );
not ( n63202 , n63201 );
or ( n63203 , n63200 , n63202 );
not ( n63204 , n54811 );
nand ( n63205 , n63204 , n54628 );
nand ( n63206 , n63203 , n63205 );
not ( n63207 , n63206 );
or ( n63208 , n63199 , n63207 );
nand ( n63209 , n62568 , n47873 );
nand ( n63210 , n63208 , n63209 );
not ( n63211 , n59633 );
not ( n63212 , n62579 );
or ( n63213 , n63211 , n63212 );
not ( n63214 , n58982 );
not ( n63215 , n53289 );
or ( n63216 , n63214 , n63215 );
not ( n63217 , n54020 );
nand ( n63218 , n63217 , n62577 );
nand ( n63219 , n63216 , n63218 );
nand ( n63220 , n63219 , n58977 );
nand ( n63221 , n63213 , n63220 );
xor ( n63222 , n63210 , n63221 );
not ( n63223 , n56639 );
not ( n63224 , n59345 );
not ( n63225 , n53271 );
or ( n63226 , n63224 , n63225 );
nand ( n63227 , n40628 , n60617 );
nand ( n63228 , n63226 , n63227 );
not ( n63229 , n63228 );
or ( n63230 , n63223 , n63229 );
nand ( n63231 , n62590 , n59950 );
nand ( n63232 , n63230 , n63231 );
xor ( n63233 , n63222 , n63232 );
xor ( n63234 , n63198 , n63233 );
xor ( n63235 , n62370 , n63197 );
and ( n63236 , n63235 , n63233 );
and ( n63237 , n62370 , n63197 );
or ( n63238 , n63236 , n63237 );
not ( n63239 , n50659 );
not ( n63240 , n62386 );
or ( n63241 , n63239 , n63240 );
not ( n63242 , n46072 );
and ( n63243 , n831 , n38980 );
not ( n63244 , n831 );
and ( n63245 , n63244 , n42551 );
nor ( n63246 , n63243 , n63245 );
not ( n63247 , n63246 );
or ( n63248 , n63242 , n63247 );
nand ( n63249 , n42554 , n50405 );
nand ( n63250 , n63248 , n63249 );
nand ( n63251 , n63250 , n46602 );
nand ( n63252 , n63241 , n63251 );
xor ( n63253 , n63252 , n62315 );
xor ( n63254 , n63253 , n62353 );
xor ( n63255 , n63254 , n62922 );
xor ( n63256 , n63255 , n62980 );
xor ( n63257 , n63254 , n62922 );
and ( n63258 , n63257 , n62980 );
and ( n63259 , n63254 , n62922 );
or ( n63260 , n63258 , n63259 );
xor ( n63261 , n62950 , n62480 );
xor ( n63262 , n63261 , n62557 );
xor ( n63263 , n62950 , n62480 );
and ( n63264 , n63263 , n62557 );
and ( n63265 , n62950 , n62480 );
or ( n63266 , n63264 , n63265 );
xor ( n63267 , n62994 , n63004 );
and ( n63268 , n63267 , n63015 );
and ( n63269 , n62994 , n63004 );
or ( n63270 , n63268 , n63269 );
xor ( n63271 , n63051 , n63092 );
xor ( n63272 , n63271 , n62683 );
xor ( n63273 , n63051 , n63092 );
and ( n63274 , n63273 , n62683 );
and ( n63275 , n63051 , n63092 );
or ( n63276 , n63274 , n63275 );
xor ( n63277 , n63121 , n62563 );
xor ( n63278 , n63277 , n62601 );
xor ( n63279 , n63121 , n62563 );
and ( n63280 , n63279 , n62601 );
and ( n63281 , n63121 , n62563 );
or ( n63282 , n63280 , n63281 );
xor ( n63283 , n62730 , n62711 );
xor ( n63284 , n63283 , n63234 );
xor ( n63285 , n62730 , n62711 );
and ( n63286 , n63285 , n63234 );
and ( n63287 , n62730 , n62711 );
or ( n63288 , n63286 , n63287 );
xor ( n63289 , n63161 , n62736 );
xor ( n63290 , n63289 , n63262 );
xor ( n63291 , n63161 , n62736 );
and ( n63292 , n63291 , n63262 );
and ( n63293 , n63161 , n62736 );
or ( n63294 , n63292 , n63293 );
xor ( n63295 , n63256 , n62746 );
xor ( n63296 , n63295 , n63278 );
xor ( n63297 , n63256 , n62746 );
and ( n63298 , n63297 , n63278 );
and ( n63299 , n63256 , n62746 );
or ( n63300 , n63298 , n63299 );
xor ( n63301 , n62752 , n63272 );
xor ( n63302 , n63301 , n63284 );
xor ( n63303 , n62752 , n63272 );
and ( n63304 , n63303 , n63284 );
and ( n63305 , n62752 , n63272 );
or ( n63306 , n63304 , n63305 );
xor ( n63307 , n62758 , n63290 );
xor ( n63308 , n63307 , n62764 );
xor ( n63309 , n62758 , n63290 );
and ( n63310 , n63309 , n62764 );
and ( n63311 , n62758 , n63290 );
or ( n63312 , n63310 , n63311 );
xor ( n63313 , n63296 , n63302 );
xor ( n63314 , n63313 , n62770 );
xor ( n63315 , n63296 , n63302 );
and ( n63316 , n63315 , n62770 );
and ( n63317 , n63296 , n63302 );
or ( n63318 , n63316 , n63317 );
xor ( n63319 , n62776 , n63308 );
xor ( n63320 , n63319 , n62782 );
xor ( n63321 , n62776 , n63308 );
and ( n63322 , n63321 , n62782 );
and ( n63323 , n62776 , n63308 );
or ( n63324 , n63322 , n63323 );
xor ( n63325 , n63314 , n63320 );
xor ( n63326 , n63325 , n62788 );
xor ( n63327 , n63314 , n63320 );
and ( n63328 , n63327 , n62788 );
and ( n63329 , n63314 , n63320 );
or ( n63330 , n63328 , n63329 );
xor ( n63331 , n63066 , n63076 );
and ( n63332 , n63331 , n63089 );
and ( n63333 , n63066 , n63076 );
or ( n63334 , n63332 , n63333 );
xor ( n63335 , n63027 , n63038 );
and ( n63336 , n63335 , n63049 );
and ( n63337 , n63027 , n63038 );
or ( n63338 , n63336 , n63337 );
xor ( n63339 , n63106 , n63107 );
and ( n63340 , n63339 , n63118 );
and ( n63341 , n63106 , n63107 );
or ( n63342 , n63340 , n63341 );
xor ( n63343 , n63175 , n63186 );
and ( n63344 , n63343 , n63196 );
and ( n63345 , n63175 , n63186 );
or ( n63346 , n63344 , n63345 );
xor ( n63347 , n63210 , n63221 );
and ( n63348 , n63347 , n63232 );
and ( n63349 , n63210 , n63221 );
or ( n63350 , n63348 , n63349 );
xor ( n63351 , n63136 , n63146 );
and ( n63352 , n63351 , n63158 );
and ( n63353 , n63136 , n63146 );
or ( n63354 , n63352 , n63353 );
xor ( n63355 , n63252 , n62315 );
and ( n63356 , n63355 , n62353 );
and ( n63357 , n63252 , n62315 );
or ( n63358 , n63356 , n63357 );
not ( n63359 , n62863 );
not ( n63360 , n53169 );
or ( n63361 , n63359 , n63360 );
not ( n63362 , n50827 );
not ( n63363 , n62858 );
or ( n63364 , n63362 , n63363 );
nand ( n63365 , n49809 , n51505 );
nand ( n63366 , n63364 , n63365 );
nand ( n63367 , n63366 , n51145 );
nand ( n63368 , n63361 , n63367 );
not ( n63369 , n62879 );
not ( n63370 , n56310 );
or ( n63371 , n63369 , n63370 );
not ( n63372 , n49838 );
not ( n63373 , n52130 );
or ( n63374 , n63372 , n63373 );
nand ( n63375 , n52108 , n49837 );
nand ( n63376 , n63374 , n63375 );
nand ( n63377 , n51766 , n63376 );
nand ( n63378 , n63371 , n63377 );
xor ( n63379 , n63368 , n63378 );
not ( n63380 , n45816 );
not ( n63381 , n37637 );
not ( n63382 , n37523 );
nand ( n63383 , n63382 , n36287 , n37382 );
nand ( n63384 , n37383 , n37647 , n63383 );
not ( n63385 , n63384 );
or ( n63386 , n63381 , n63385 );
not ( n63387 , n37637 );
nand ( n63388 , n37383 , n37647 , n63383 , n63387 );
nand ( n63389 , n63386 , n63388 );
not ( n63390 , n63389 );
not ( n63391 , n63390 );
or ( n63392 , n63380 , n63391 );
not ( n63393 , n63389 );
not ( n63394 , n63393 );
nand ( n63395 , n63394 , n48766 );
nand ( n63396 , n63392 , n63395 );
not ( n63397 , n63396 );
buf ( n63398 , n62843 );
not ( n63399 , n63398 );
or ( n63400 , n63397 , n63399 );
not ( n63401 , n63393 );
not ( n63402 , n62837 );
not ( n63403 , n63402 );
or ( n63404 , n63401 , n63403 );
not ( n63405 , n63389 );
not ( n63406 , n62837 );
or ( n63407 , n63405 , n63406 );
nand ( n63408 , n63404 , n63407 );
nand ( n63409 , n62842 , n63408 );
not ( n63410 , n63409 );
not ( n63411 , n63410 );
buf ( n63412 , n63405 );
and ( n63413 , n46440 , n63412 );
not ( n63414 , n46440 );
buf ( n63415 , n63390 );
not ( n63416 , n63415 );
and ( n63417 , n63414 , n63416 );
nor ( n63418 , n63413 , n63417 );
or ( n63419 , n63411 , n63418 );
nand ( n63420 , n63400 , n63419 );
xor ( n63421 , n63379 , n63420 );
xor ( n63422 , n63368 , n63378 );
and ( n63423 , n63422 , n63420 );
and ( n63424 , n63368 , n63378 );
or ( n63425 , n63423 , n63424 );
not ( n63426 , n62889 );
not ( n63427 , n61016 );
or ( n63428 , n63426 , n63427 );
not ( n63429 , n57252 );
not ( n63430 , n41363 );
or ( n63431 , n63429 , n63430 );
not ( n63432 , n41363 );
nand ( n63433 , n63432 , n52836 );
nand ( n63434 , n63431 , n63433 );
nand ( n63435 , n63434 , n52467 );
nand ( n63436 , n63428 , n63435 );
not ( n63437 , n62899 );
not ( n63438 , n61032 );
or ( n63439 , n63437 , n63438 );
not ( n63440 , n58556 );
not ( n63441 , n63440 );
not ( n63442 , n53594 );
or ( n63443 , n63441 , n63442 );
nand ( n63444 , n53589 , n41530 );
nand ( n63445 , n63443 , n63444 );
nand ( n63446 , n63445 , n53325 );
nand ( n63447 , n63439 , n63446 );
xor ( n63448 , n63436 , n63447 );
not ( n63449 , n62992 );
not ( n63450 , n54313 );
or ( n63451 , n63449 , n63450 );
not ( n63452 , n60329 );
not ( n63453 , n54301 );
or ( n63454 , n63452 , n63453 );
nand ( n63455 , n56274 , n58459 );
nand ( n63456 , n63454 , n63455 );
nand ( n63457 , n63456 , n54077 );
nand ( n63458 , n63451 , n63457 );
xor ( n63459 , n63448 , n63458 );
xor ( n63460 , n63436 , n63447 );
and ( n63461 , n63460 , n63458 );
and ( n63462 , n63436 , n63447 );
or ( n63463 , n63461 , n63462 );
xor ( n63464 , n63270 , n63334 );
xor ( n63465 , n63464 , n63338 );
xor ( n63466 , n63270 , n63334 );
and ( n63467 , n63466 , n63338 );
and ( n63468 , n63270 , n63334 );
or ( n63469 , n63467 , n63468 );
not ( n63470 , n47407 );
not ( n63471 , n62935 );
or ( n63472 , n63470 , n63471 );
not ( n63473 , n51545 );
not ( n63474 , n59402 );
or ( n63475 , n63473 , n63474 );
nand ( n63476 , n39574 , n50634 );
nand ( n63477 , n63475 , n63476 );
nand ( n63478 , n63477 , n53675 );
nand ( n63479 , n63472 , n63478 );
not ( n63480 , n49252 );
not ( n63481 , n62946 );
or ( n63482 , n63480 , n63481 );
not ( n63483 , n47980 );
not ( n63484 , n39679 );
or ( n63485 , n63483 , n63484 );
or ( n63486 , n39679 , n47980 );
nand ( n63487 , n63485 , n63486 );
nand ( n63488 , n63487 , n53510 );
nand ( n63489 , n63482 , n63488 );
xor ( n63490 , n63479 , n63489 );
not ( n63491 , n46267 );
not ( n63492 , n62965 );
or ( n63493 , n63491 , n63492 );
not ( n63494 , n46425 );
not ( n63495 , n62715 );
or ( n63496 , n63494 , n63495 );
nand ( n63497 , n39253 , n46422 );
nand ( n63498 , n63496 , n63497 );
nand ( n63499 , n63498 , n49026 );
nand ( n63500 , n63493 , n63499 );
xor ( n63501 , n63490 , n63500 );
xor ( n63502 , n63479 , n63489 );
and ( n63503 , n63502 , n63500 );
and ( n63504 , n63479 , n63489 );
or ( n63505 , n63503 , n63504 );
not ( n63506 , n49713 );
not ( n63507 , n62974 );
or ( n63508 , n63506 , n63507 );
not ( n63509 , n57787 );
not ( n63510 , n63509 );
and ( n63511 , n51351 , n63510 );
not ( n63512 , n51351 );
and ( n63513 , n63512 , n39894 );
nor ( n63514 , n63511 , n63513 );
not ( n63515 , n63514 );
nand ( n63516 , n63515 , n51865 );
nand ( n63517 , n63508 , n63516 );
xor ( n63518 , n63517 , n63342 );
xor ( n63519 , n63518 , n63421 );
xor ( n63520 , n63517 , n63342 );
and ( n63521 , n63520 , n63421 );
and ( n63522 , n63517 , n63342 );
or ( n63523 , n63521 , n63522 );
not ( n63524 , n63036 );
not ( n63525 , n61397 );
not ( n63526 , n63525 );
or ( n63527 , n63524 , n63526 );
not ( n63528 , n49654 );
not ( n63529 , n60968 );
or ( n63530 , n63528 , n63529 );
nand ( n63531 , n60285 , n47368 );
nand ( n63532 , n63530 , n63531 );
nand ( n63533 , n59855 , n63532 );
nand ( n63534 , n63527 , n63533 );
not ( n63535 , n63047 );
not ( n63536 , n61548 );
or ( n63537 , n63535 , n63536 );
not ( n63538 , n47047 );
not ( n63539 , n61537 );
or ( n63540 , n63538 , n63539 );
not ( n63541 , n61536 );
nand ( n63542 , n63541 , n47821 );
nand ( n63543 , n63540 , n63542 );
nand ( n63544 , n61557 , n63543 );
nand ( n63545 , n63537 , n63544 );
xor ( n63546 , n63534 , n63545 );
not ( n63547 , n62461 );
and ( n63548 , n61416 , n61805 );
not ( n63549 , n61416 );
and ( n63550 , n63549 , n61804 );
nor ( n63551 , n63548 , n63550 );
nand ( n63552 , n63547 , n63551 );
or ( n63553 , n63552 , n63103 );
and ( n63554 , n62448 , n46824 );
not ( n63555 , n62448 );
and ( n63556 , n63555 , n46273 );
nor ( n63557 , n63554 , n63556 );
or ( n63558 , n63557 , n63551 );
nand ( n63559 , n63553 , n63558 );
xor ( n63560 , n63546 , n63559 );
xor ( n63561 , n63560 , n63459 );
not ( n63562 , n63074 );
not ( n63563 , n58541 );
or ( n63564 , n63562 , n63563 );
not ( n63565 , n52033 );
not ( n63566 , n57534 );
or ( n63567 , n63565 , n63566 );
nand ( n63568 , n57634 , n55959 );
nand ( n63569 , n63567 , n63568 );
nand ( n63570 , n63569 , n57139 );
nand ( n63571 , n63564 , n63570 );
not ( n63572 , n63087 );
not ( n63573 , n58962 );
or ( n63574 , n63572 , n63573 );
not ( n63575 , n58630 );
not ( n63576 , n49624 );
or ( n63577 , n63575 , n63576 );
nand ( n63578 , n58626 , n49630 );
nand ( n63579 , n63577 , n63578 );
nand ( n63580 , n63579 , n60400 );
nand ( n63581 , n63574 , n63580 );
xor ( n63582 , n63571 , n63581 );
not ( n63583 , n63025 );
not ( n63584 , n60539 );
or ( n63585 , n63583 , n63584 );
not ( n63586 , n47765 );
buf ( n63587 , n59578 );
not ( n63588 , n63587 );
or ( n63589 , n63586 , n63588 );
nand ( n63590 , n62513 , n48589 );
nand ( n63591 , n63589 , n63590 );
nand ( n63592 , n63591 , n59931 );
nand ( n63593 , n63585 , n63592 );
xor ( n63594 , n63582 , n63593 );
xor ( n63595 , n63561 , n63594 );
xor ( n63596 , n63560 , n63459 );
and ( n63597 , n63596 , n63594 );
and ( n63598 , n63560 , n63459 );
or ( n63599 , n63597 , n63598 );
not ( n63600 , n63002 );
not ( n63601 , n58592 );
or ( n63602 , n63600 , n63601 );
not ( n63603 , n47527 );
not ( n63604 , n60985 );
or ( n63605 , n63603 , n63604 );
nand ( n63606 , n55118 , n51360 );
nand ( n63607 , n63605 , n63606 );
nand ( n63608 , n63607 , n54847 );
nand ( n63609 , n63602 , n63608 );
not ( n63610 , n63013 );
not ( n63611 , n58070 );
or ( n63612 , n63610 , n63611 );
not ( n63613 , n47918 );
not ( n63614 , n57676 );
or ( n63615 , n63613 , n63614 );
nand ( n63616 , n55845 , n49245 );
nand ( n63617 , n63615 , n63616 );
nand ( n63618 , n55458 , n63617 );
nand ( n63619 , n63612 , n63618 );
xor ( n63620 , n63609 , n63619 );
not ( n63621 , n63064 );
not ( n63622 , n56776 );
or ( n63623 , n63621 , n63622 );
not ( n63624 , n54185 );
not ( n63625 , n57665 );
or ( n63626 , n63624 , n63625 );
nand ( n63627 , n56679 , n52712 );
nand ( n63628 , n63626 , n63627 );
nand ( n63629 , n56780 , n63628 );
nand ( n63630 , n63623 , n63629 );
xor ( n63631 , n63620 , n63630 );
xor ( n63632 , n63631 , n63346 );
xor ( n63633 , n63632 , n63350 );
xor ( n63634 , n63631 , n63346 );
and ( n63635 , n63634 , n63350 );
and ( n63636 , n63631 , n63346 );
or ( n63637 , n63635 , n63636 );
xor ( n63638 , n62954 , n63358 );
xor ( n63639 , n63638 , n63354 );
xor ( n63640 , n62954 , n63358 );
and ( n63641 , n63640 , n63354 );
and ( n63642 , n62954 , n63358 );
or ( n63643 , n63641 , n63642 );
not ( n63644 , n58977 );
not ( n63645 , n58982 );
not ( n63646 , n40225 );
or ( n63647 , n63645 , n63646 );
nand ( n63648 , n56073 , n62577 );
nand ( n63649 , n63647 , n63648 );
not ( n63650 , n63649 );
or ( n63651 , n63644 , n63650 );
nand ( n63652 , n63219 , n53104 );
nand ( n63653 , n63651 , n63652 );
not ( n63654 , n56639 );
not ( n63655 , n59345 );
buf ( n63656 , n52906 );
not ( n63657 , n63656 );
or ( n63658 , n63655 , n63657 );
nand ( n63659 , n59612 , n60617 );
nand ( n63660 , n63658 , n63659 );
not ( n63661 , n63660 );
or ( n63662 , n63654 , n63661 );
nand ( n63663 , n63228 , n59950 );
nand ( n63664 , n63662 , n63663 );
xor ( n63665 , n63653 , n63664 );
not ( n63666 , n62085 );
not ( n63667 , n63132 );
or ( n63668 , n63666 , n63667 );
not ( n63669 , n62077 );
not ( n63670 , n54377 );
or ( n63671 , n63669 , n63670 );
nand ( n63672 , n52212 , n60289 );
nand ( n63673 , n63671 , n63672 );
nand ( n63674 , n63673 , n60927 );
nand ( n63675 , n63668 , n63674 );
xor ( n63676 , n63665 , n63675 );
xor ( n63677 , n62926 , n63676 );
not ( n63678 , n62837 );
or ( n63679 , n63678 , n46440 );
nand ( n63680 , n63679 , n62451 );
not ( n63681 , n63412 );
nand ( n63682 , n63678 , n48689 );
and ( n63683 , n63680 , n63681 , n63682 );
not ( n63684 , n63683 );
not ( n63685 , n62851 );
not ( n63686 , n51215 );
or ( n63687 , n63685 , n63686 );
not ( n63688 , n51461 );
not ( n63689 , n52767 );
or ( n63690 , n63688 , n63689 );
nand ( n63691 , n51462 , n54249 );
nand ( n63692 , n63690 , n63691 );
nand ( n63693 , n63692 , n50921 );
nand ( n63694 , n63687 , n63693 );
not ( n63695 , n63694 );
not ( n63696 , n63695 );
or ( n63697 , n63684 , n63696 );
or ( n63698 , n63695 , n63683 );
nand ( n63699 , n63697 , n63698 );
not ( n63700 , n50304 );
not ( n63701 , n50958 );
or ( n63702 , n63700 , n63701 );
nand ( n63703 , n52284 , n50943 );
nand ( n63704 , n63702 , n63703 );
not ( n63705 , n63704 );
not ( n63706 , n52757 );
or ( n63707 , n63705 , n63706 );
not ( n63708 , n59820 );
nand ( n63709 , n63114 , n63708 );
nand ( n63710 , n63707 , n63709 );
xor ( n63711 , n63699 , n63710 );
not ( n63712 , n63184 );
or ( n63713 , n63712 , n50241 );
not ( n63714 , n57810 );
not ( n63715 , n39963 );
or ( n63716 , n63714 , n63715 );
nand ( n63717 , n57801 , n49679 );
nand ( n63718 , n63716 , n63717 );
not ( n63719 , n63718 );
or ( n63720 , n63719 , n50239 );
nand ( n63721 , n63713 , n63720 );
xor ( n63722 , n63711 , n63721 );
xor ( n63723 , n63677 , n63722 );
xor ( n63724 , n62926 , n63676 );
and ( n63725 , n63724 , n63722 );
and ( n63726 , n62926 , n63676 );
or ( n63727 , n63725 , n63726 );
not ( n63728 , n54875 );
not ( n63729 , n48856 );
not ( n63730 , n56020 );
or ( n63731 , n63729 , n63730 );
not ( n63732 , n40513 );
nand ( n63733 , n63732 , n58692 );
nand ( n63734 , n63731 , n63733 );
not ( n63735 , n63734 );
or ( n63736 , n63728 , n63735 );
nand ( n63737 , n63171 , n52421 );
nand ( n63738 , n63736 , n63737 );
not ( n63739 , n52004 );
not ( n63740 , n52377 );
not ( n63741 , n55199 );
or ( n63742 , n63740 , n63741 );
nand ( n63743 , n55203 , n53973 );
nand ( n63744 , n63742 , n63743 );
not ( n63745 , n63744 );
or ( n63746 , n63739 , n63745 );
nand ( n63747 , n63192 , n48894 );
nand ( n63748 , n63746 , n63747 );
xor ( n63749 , n63738 , n63748 );
not ( n63750 , n47873 );
not ( n63751 , n63206 );
or ( n63752 , n63750 , n63751 );
not ( n63753 , n59174 );
not ( n63754 , n54405 );
or ( n63755 , n63753 , n63754 );
nand ( n63756 , n54406 , n54628 );
nand ( n63757 , n63755 , n63756 );
nand ( n63758 , n63757 , n54623 );
nand ( n63759 , n63752 , n63758 );
xor ( n63760 , n63749 , n63759 );
xor ( n63761 , n63760 , n62984 );
not ( n63762 , n52058 );
not ( n63763 , n63142 );
or ( n63764 , n63762 , n63763 );
not ( n63765 , n61951 );
not ( n63766 , n52222 );
or ( n63767 , n63765 , n63766 );
nand ( n63768 , n52893 , n61952 );
nand ( n63769 , n63767 , n63768 );
nand ( n63770 , n63769 , n50078 );
nand ( n63771 , n63764 , n63770 );
not ( n63772 , n46776 );
not ( n63773 , n63154 );
or ( n63774 , n63772 , n63773 );
not ( n63775 , n50263 );
not ( n63776 , n60357 );
or ( n63777 , n63775 , n63776 );
not ( n63778 , n61347 );
nand ( n63779 , n63778 , n48078 );
nand ( n63780 , n63777 , n63779 );
nand ( n63781 , n63780 , n50261 );
nand ( n63782 , n63774 , n63781 );
xor ( n63783 , n63771 , n63782 );
not ( n63784 , n50659 );
not ( n63785 , n63250 );
or ( n63786 , n63784 , n63785 );
not ( n63787 , n42652 );
and ( n63788 , n46072 , n63787 );
not ( n63789 , n46072 );
not ( n63790 , n831 );
not ( n63791 , n39432 );
or ( n63792 , n63790 , n63791 );
nand ( n63793 , n63792 , n42650 );
buf ( n63794 , n63793 );
and ( n63795 , n63789 , n63794 );
nor ( n63796 , n63788 , n63795 );
or ( n63797 , n63796 , n45861 );
nand ( n63798 , n63786 , n63797 );
xor ( n63799 , n63783 , n63798 );
xor ( n63800 , n63761 , n63799 );
xor ( n63801 , n63760 , n62984 );
and ( n63802 , n63801 , n63799 );
and ( n63803 , n63760 , n62984 );
or ( n63804 , n63802 , n63803 );
xor ( n63805 , n62871 , n62907 );
not ( n63806 , n46564 );
not ( n63807 , n62915 );
or ( n63808 , n63806 , n63807 );
not ( n63809 , n48952 );
not ( n63810 , n42398 );
or ( n63811 , n63809 , n63810 );
nand ( n63812 , n42397 , n52990 );
nand ( n63813 , n63811 , n63812 );
nand ( n63814 , n63813 , n49832 );
nand ( n63815 , n63808 , n63814 );
xor ( n63816 , n63805 , n63815 );
xor ( n63817 , n63816 , n63501 );
xor ( n63818 , n63817 , n63465 );
xor ( n63819 , n63816 , n63501 );
and ( n63820 , n63819 , n63465 );
and ( n63821 , n63816 , n63501 );
or ( n63822 , n63820 , n63821 );
xor ( n63823 , n63055 , n63595 );
xor ( n63824 , n63823 , n63519 );
xor ( n63825 , n63055 , n63595 );
and ( n63826 , n63825 , n63519 );
and ( n63827 , n63055 , n63595 );
or ( n63828 , n63826 , n63827 );
xor ( n63829 , n63609 , n63619 );
and ( n63830 , n63829 , n63630 );
and ( n63831 , n63609 , n63619 );
or ( n63832 , n63830 , n63831 );
xor ( n63833 , n63096 , n63633 );
xor ( n63834 , n63833 , n63238 );
xor ( n63835 , n63096 , n63633 );
and ( n63836 , n63835 , n63238 );
and ( n63837 , n63096 , n63633 );
or ( n63838 , n63836 , n63837 );
xor ( n63839 , n63165 , n63125 );
xor ( n63840 , n63839 , n63723 );
xor ( n63841 , n63165 , n63125 );
and ( n63842 , n63841 , n63723 );
and ( n63843 , n63165 , n63125 );
or ( n63844 , n63842 , n63843 );
xor ( n63845 , n63639 , n63260 );
xor ( n63846 , n63845 , n63266 );
xor ( n63847 , n63639 , n63260 );
and ( n63848 , n63847 , n63266 );
and ( n63849 , n63639 , n63260 );
or ( n63850 , n63848 , n63849 );
xor ( n63851 , n63818 , n63800 );
xor ( n63852 , n63851 , n63276 );
xor ( n63853 , n63818 , n63800 );
and ( n63854 , n63853 , n63276 );
and ( n63855 , n63818 , n63800 );
or ( n63856 , n63854 , n63855 );
xor ( n63857 , n63824 , n63282 );
xor ( n63858 , n63857 , n63840 );
xor ( n63859 , n63824 , n63282 );
and ( n63860 , n63859 , n63840 );
and ( n63861 , n63824 , n63282 );
or ( n63862 , n63860 , n63861 );
xor ( n63863 , n63288 , n63834 );
xor ( n63864 , n63863 , n63846 );
xor ( n63865 , n63288 , n63834 );
and ( n63866 , n63865 , n63846 );
and ( n63867 , n63288 , n63834 );
or ( n63868 , n63866 , n63867 );
xor ( n63869 , n63294 , n63852 );
xor ( n63870 , n63869 , n63300 );
xor ( n63871 , n63294 , n63852 );
and ( n63872 , n63871 , n63300 );
and ( n63873 , n63294 , n63852 );
or ( n63874 , n63872 , n63873 );
xor ( n63875 , n63858 , n63306 );
xor ( n63876 , n63875 , n63864 );
xor ( n63877 , n63858 , n63306 );
and ( n63878 , n63877 , n63864 );
and ( n63879 , n63858 , n63306 );
or ( n63880 , n63878 , n63879 );
xor ( n63881 , n63312 , n63870 );
xor ( n63882 , n63881 , n63318 );
xor ( n63883 , n63312 , n63870 );
and ( n63884 , n63883 , n63318 );
and ( n63885 , n63312 , n63870 );
or ( n63886 , n63884 , n63885 );
xor ( n63887 , n63876 , n63882 );
xor ( n63888 , n63887 , n63324 );
xor ( n63889 , n63876 , n63882 );
and ( n63890 , n63889 , n63324 );
and ( n63891 , n63876 , n63882 );
or ( n63892 , n63890 , n63891 );
xor ( n63893 , n63571 , n63581 );
and ( n63894 , n63893 , n63593 );
and ( n63895 , n63571 , n63581 );
or ( n63896 , n63894 , n63895 );
xor ( n63897 , n63534 , n63545 );
and ( n63898 , n63897 , n63559 );
and ( n63899 , n63534 , n63545 );
or ( n63900 , n63898 , n63899 );
xor ( n63901 , n63699 , n63710 );
and ( n63902 , n63901 , n63721 );
and ( n63903 , n63699 , n63710 );
or ( n63904 , n63902 , n63903 );
xor ( n63905 , n63738 , n63748 );
and ( n63906 , n63905 , n63759 );
and ( n63907 , n63738 , n63748 );
or ( n63908 , n63906 , n63907 );
xor ( n63909 , n63653 , n63664 );
and ( n63910 , n63909 , n63675 );
and ( n63911 , n63653 , n63664 );
or ( n63912 , n63910 , n63911 );
xor ( n63913 , n63771 , n63782 );
and ( n63914 , n63913 , n63798 );
and ( n63915 , n63771 , n63782 );
or ( n63916 , n63914 , n63915 );
xor ( n63917 , n62871 , n62907 );
and ( n63918 , n63917 , n63815 );
and ( n63919 , n62871 , n62907 );
or ( n63920 , n63918 , n63919 );
buf ( n63921 , n63389 );
buf ( n63922 , n63921 );
and ( n63923 , n63922 , n48689 );
not ( n63924 , n63366 );
not ( n63925 , n53170 );
or ( n63926 , n63924 , n63925 );
not ( n63927 , n41038 );
not ( n63928 , n51504 );
or ( n63929 , n63927 , n63928 );
not ( n63930 , n51891 );
nand ( n63931 , n63930 , n53549 );
nand ( n63932 , n63929 , n63931 );
nand ( n63933 , n51533 , n63932 );
nand ( n63934 , n63926 , n63933 );
xor ( n63935 , n63923 , n63934 );
not ( n63936 , n63376 );
not ( n63937 , n52482 );
or ( n63938 , n63936 , n63937 );
not ( n63939 , n56239 );
not ( n63940 , n52113 );
or ( n63941 , n63939 , n63940 );
nand ( n63942 , n52870 , n62861 );
nand ( n63943 , n63941 , n63942 );
not ( n63944 , n63943 );
or ( n63945 , n63944 , n62302 );
nand ( n63946 , n63938 , n63945 );
xor ( n63947 , n63935 , n63946 );
xor ( n63948 , n63923 , n63934 );
and ( n63949 , n63948 , n63946 );
and ( n63950 , n63923 , n63934 );
or ( n63951 , n63949 , n63950 );
not ( n63952 , n63396 );
not ( n63953 , n63409 );
not ( n63954 , n63953 );
or ( n63955 , n63952 , n63954 );
not ( n63956 , n63390 );
not ( n63957 , n46037 );
or ( n63958 , n63956 , n63957 );
not ( n63959 , n63393 );
nand ( n63960 , n63959 , n54721 );
nand ( n63961 , n63958 , n63960 );
nand ( n63962 , n63961 , n62843 );
nand ( n63963 , n63955 , n63962 );
not ( n63964 , n63434 );
not ( n63965 , n52853 );
or ( n63966 , n63964 , n63965 );
and ( n63967 , n49001 , n57253 );
not ( n63968 , n49001 );
and ( n63969 , n63968 , n55103 );
or ( n63970 , n63967 , n63969 );
nand ( n63971 , n63970 , n52469 );
nand ( n63972 , n63966 , n63971 );
xor ( n63973 , n63963 , n63972 );
not ( n63974 , n63445 );
or ( n63975 , n61329 , n63974 );
and ( n63976 , n53591 , n48486 );
and ( n63977 , n53590 , n48951 );
nor ( n63978 , n63976 , n63977 );
or ( n63979 , n63978 , n53618 );
nand ( n63980 , n63975 , n63979 );
xor ( n63981 , n63973 , n63980 );
xor ( n63982 , n63963 , n63972 );
and ( n63983 , n63982 , n63980 );
and ( n63984 , n63963 , n63972 );
or ( n63985 , n63983 , n63984 );
xor ( n63986 , n63463 , n63832 );
xor ( n63987 , n63986 , n63896 );
xor ( n63988 , n63463 , n63832 );
and ( n63989 , n63988 , n63896 );
and ( n63990 , n63463 , n63832 );
or ( n63991 , n63989 , n63990 );
not ( n63992 , n53675 );
not ( n63993 , n47803 );
not ( n63994 , n60874 );
or ( n63995 , n63993 , n63994 );
nand ( n63996 , n39056 , n50634 );
nand ( n63997 , n63995 , n63996 );
not ( n63998 , n63997 );
or ( n63999 , n63992 , n63998 );
nand ( n64000 , n63477 , n47407 );
nand ( n64001 , n63999 , n64000 );
xor ( n64002 , n63900 , n64001 );
not ( n64003 , n50659 );
not ( n64004 , n63796 );
not ( n64005 , n64004 );
or ( n64006 , n64003 , n64005 );
nand ( n64007 , n46072 , n44004 );
nand ( n64008 , n64006 , n64007 );
xor ( n64009 , n64002 , n64008 );
xor ( n64010 , n63900 , n64001 );
and ( n64011 , n64010 , n64008 );
and ( n64012 , n63900 , n64001 );
or ( n64013 , n64011 , n64012 );
not ( n64014 , n49252 );
not ( n64015 , n63487 );
or ( n64016 , n64014 , n64015 );
not ( n64017 , n49500 );
not ( n64018 , n60906 );
or ( n64019 , n64017 , n64018 );
nand ( n64020 , n39713 , n47979 );
nand ( n64021 , n64019 , n64020 );
nand ( n64022 , n64021 , n47384 );
nand ( n64023 , n64016 , n64022 );
not ( n64024 , n46267 );
not ( n64025 , n63498 );
or ( n64026 , n64024 , n64025 );
not ( n64027 , n46425 );
not ( n64028 , n61904 );
or ( n64029 , n64027 , n64028 );
nand ( n64030 , n62912 , n46422 );
nand ( n64031 , n64029 , n64030 );
nand ( n64032 , n64031 , n49026 );
nand ( n64033 , n64026 , n64032 );
xor ( n64034 , n64023 , n64033 );
not ( n64035 , n52267 );
not ( n64036 , n58047 );
or ( n64037 , n64035 , n64036 );
nand ( n64038 , n39779 , n48661 );
nand ( n64039 , n64037 , n64038 );
not ( n64040 , n64039 );
not ( n64041 , n51865 );
or ( n64042 , n64040 , n64041 );
or ( n64043 , n50057 , n63514 );
nand ( n64044 , n64042 , n64043 );
xor ( n64045 , n64034 , n64044 );
xor ( n64046 , n64023 , n64033 );
and ( n64047 , n64046 , n64044 );
and ( n64048 , n64023 , n64033 );
or ( n64049 , n64047 , n64048 );
xor ( n64050 , n63981 , n63947 );
not ( n64051 , n63456 );
not ( n64052 , n54315 );
or ( n64053 , n64051 , n64052 );
not ( n64054 , n54298 );
not ( n64055 , n58914 );
and ( n64056 , n64054 , n64055 );
not ( n64057 , n41668 );
and ( n64058 , n56274 , n64057 );
nor ( n64059 , n64056 , n64058 );
not ( n64060 , n64059 );
nand ( n64061 , n64060 , n56277 );
nand ( n64062 , n64053 , n64061 );
not ( n64063 , n55143 );
not ( n64064 , n63607 );
or ( n64065 , n64063 , n64064 );
not ( n64066 , n52379 );
not ( n64067 , n55148 );
or ( n64068 , n64066 , n64067 );
nand ( n64069 , n55582 , n58179 );
nand ( n64070 , n64068 , n64069 );
nand ( n64071 , n64070 , n54848 );
nand ( n64072 , n64065 , n64071 );
xor ( n64073 , n64062 , n64072 );
not ( n64074 , n55887 );
not ( n64075 , n63617 );
or ( n64076 , n64074 , n64075 );
not ( n64077 , n57186 );
not ( n64078 , n55892 );
or ( n64079 , n64077 , n64078 );
or ( n64080 , n55872 , n57186 );
nand ( n64081 , n64079 , n64080 );
nand ( n64082 , n64081 , n55459 );
nand ( n64083 , n64076 , n64082 );
xor ( n64084 , n64073 , n64083 );
xor ( n64085 , n64050 , n64084 );
xor ( n64086 , n63981 , n63947 );
and ( n64087 , n64086 , n64084 );
and ( n64088 , n63981 , n63947 );
or ( n64089 , n64087 , n64088 );
not ( n64090 , n63591 );
not ( n64091 , n60539 );
or ( n64092 , n64090 , n64091 );
not ( n64093 , n51204 );
not ( n64094 , n62510 );
or ( n64095 , n64093 , n64094 );
nand ( n64096 , n59935 , n48860 );
nand ( n64097 , n64095 , n64096 );
nand ( n64098 , n58908 , n64097 );
nand ( n64099 , n64092 , n64098 );
not ( n64100 , n63532 );
or ( n64101 , n60960 , n64100 );
not ( n64102 , n60285 );
and ( n64103 , n48898 , n64102 );
not ( n64104 , n48898 );
and ( n64105 , n64104 , n60285 );
nor ( n64106 , n64103 , n64105 );
or ( n64107 , n60963 , n64106 );
nand ( n64108 , n64101 , n64107 );
xor ( n64109 , n64099 , n64108 );
not ( n64110 , n63543 );
buf ( n64111 , n61548 );
not ( n64112 , n64111 );
or ( n64113 , n64110 , n64112 );
nand ( n64114 , n61537 , n47227 );
not ( n64115 , n64114 );
nand ( n64116 , n61416 , n47589 );
not ( n64117 , n64116 );
or ( n64118 , n64115 , n64117 );
nand ( n64119 , n64118 , n62428 );
nand ( n64120 , n64113 , n64119 );
xor ( n64121 , n64109 , n64120 );
not ( n64122 , n63628 );
not ( n64123 , n56776 );
or ( n64124 , n64122 , n64123 );
not ( n64125 , n48983 );
not ( n64126 , n58534 );
or ( n64127 , n64125 , n64126 );
nand ( n64128 , n57664 , n56348 );
nand ( n64129 , n64127 , n64128 );
nand ( n64130 , n56780 , n64129 );
nand ( n64131 , n64124 , n64130 );
not ( n64132 , n57628 );
not ( n64133 , n63569 );
or ( n64134 , n64132 , n64133 );
not ( n64135 , n55511 );
not ( n64136 , n62485 );
or ( n64137 , n64135 , n64136 );
nand ( n64138 , n57619 , n51670 );
nand ( n64139 , n64137 , n64138 );
nand ( n64140 , n59435 , n64139 );
nand ( n64141 , n64134 , n64140 );
xor ( n64142 , n64131 , n64141 );
not ( n64143 , n63080 );
not ( n64144 , n63579 );
or ( n64145 , n64143 , n64144 );
not ( n64146 , n61465 );
not ( n64147 , n51792 );
not ( n64148 , n62497 );
or ( n64149 , n64147 , n64148 );
nand ( n64150 , n58642 , n48829 );
nand ( n64151 , n64149 , n64150 );
not ( n64152 , n64151 );
or ( n64153 , n64146 , n64152 );
nand ( n64154 , n64145 , n64153 );
xor ( n64155 , n64142 , n64154 );
xor ( n64156 , n64121 , n64155 );
xor ( n64157 , n64156 , n63904 );
xor ( n64158 , n64121 , n64155 );
and ( n64159 , n64158 , n63904 );
and ( n64160 , n64121 , n64155 );
or ( n64161 , n64159 , n64160 );
xor ( n64162 , n63908 , n63912 );
not ( n64163 , n63552 );
not ( n64164 , n64163 );
or ( n64165 , n64164 , n63557 );
buf ( n64166 , n63551 );
not ( n64167 , n62451 );
and ( n64168 , n47646 , n64167 );
not ( n64169 , n47646 );
buf ( n64170 , n62451 );
and ( n64171 , n64169 , n64170 );
nor ( n64172 , n64168 , n64171 );
or ( n64173 , n64166 , n64172 );
nand ( n64174 , n64165 , n64173 );
not ( n64175 , n51223 );
not ( n64176 , n40691 );
not ( n64177 , n50946 );
or ( n64178 , n64176 , n64177 );
or ( n64179 , n50946 , n40691 );
nand ( n64180 , n64178 , n64179 );
not ( n64181 , n64180 );
or ( n64182 , n64175 , n64181 );
nand ( n64183 , n52526 , n63692 );
nand ( n64184 , n64182 , n64183 );
xor ( n64185 , n64174 , n64184 );
not ( n64186 , n52757 );
not ( n64187 , n50306 );
not ( n64188 , n59176 );
or ( n64189 , n64187 , n64188 );
buf ( n64190 , n50306 );
not ( n64191 , n64190 );
nand ( n64192 , n57332 , n64191 );
nand ( n64193 , n64189 , n64192 );
not ( n64194 , n64193 );
or ( n64195 , n64186 , n64194 );
nand ( n64196 , n63704 , n63708 );
nand ( n64197 , n64195 , n64196 );
xor ( n64198 , n64185 , n64197 );
xor ( n64199 , n64162 , n64198 );
xor ( n64200 , n63908 , n63912 );
and ( n64201 , n64200 , n64198 );
and ( n64202 , n63908 , n63912 );
or ( n64203 , n64201 , n64202 );
not ( n64204 , n60927 );
not ( n64205 , n49112 );
not ( n64206 , n54046 );
or ( n64207 , n64205 , n64206 );
nand ( n64208 , n40626 , n60289 );
nand ( n64209 , n64207 , n64208 );
not ( n64210 , n64209 );
or ( n64211 , n64204 , n64210 );
nand ( n64212 , n63673 , n62085 );
nand ( n64213 , n64211 , n64212 );
not ( n64214 , n52058 );
not ( n64215 , n63769 );
or ( n64216 , n64214 , n64215 );
not ( n64217 , n61951 );
not ( n64218 , n40527 );
or ( n64219 , n64217 , n64218 );
nand ( n64220 , n51916 , n61952 );
nand ( n64221 , n64219 , n64220 );
nand ( n64222 , n64221 , n62654 );
nand ( n64223 , n64216 , n64222 );
xor ( n64224 , n64213 , n64223 );
not ( n64225 , n52043 );
not ( n64226 , n48645 );
not ( n64227 , n39844 );
or ( n64228 , n64226 , n64227 );
nand ( n64229 , n58034 , n49679 );
nand ( n64230 , n64228 , n64229 );
not ( n64231 , n64230 );
or ( n64232 , n64225 , n64231 );
nand ( n64233 , n63718 , n50242 );
nand ( n64234 , n64232 , n64233 );
xor ( n64235 , n64224 , n64234 );
xor ( n64236 , n63916 , n64235 );
xor ( n64237 , n64236 , n63505 );
xor ( n64238 , n63916 , n64235 );
and ( n64239 , n64238 , n63505 );
and ( n64240 , n63916 , n64235 );
or ( n64241 , n64239 , n64240 );
xor ( n64242 , n63469 , n63920 );
not ( n64243 , n47873 );
not ( n64244 , n63757 );
or ( n64245 , n64243 , n64244 );
not ( n64246 , n51684 );
not ( n64247 , n56441 );
or ( n64248 , n64246 , n64247 );
nand ( n64249 , n54790 , n59174 );
nand ( n64250 , n64248 , n64249 );
nand ( n64251 , n64250 , n54623 );
nand ( n64252 , n64245 , n64251 );
not ( n64253 , n59633 );
not ( n64254 , n63649 );
or ( n64255 , n64253 , n64254 );
and ( n64256 , n53884 , n60602 );
not ( n64257 , n53884 );
and ( n64258 , n64257 , n62577 );
or ( n64259 , n64256 , n64258 );
nand ( n64260 , n64259 , n58977 );
nand ( n64261 , n64255 , n64260 );
xor ( n64262 , n64252 , n64261 );
not ( n64263 , n59950 );
not ( n64264 , n63660 );
or ( n64265 , n64263 , n64264 );
not ( n64266 , n59345 );
not ( n64267 , n56476 );
or ( n64268 , n64266 , n64267 );
nand ( n64269 , n40377 , n60617 );
nand ( n64270 , n64268 , n64269 );
nand ( n64271 , n64270 , n56639 );
nand ( n64272 , n64265 , n64271 );
xor ( n64273 , n64262 , n64272 );
xor ( n64274 , n64242 , n64273 );
xor ( n64275 , n63469 , n63920 );
and ( n64276 , n64275 , n64273 );
and ( n64277 , n63469 , n63920 );
or ( n64278 , n64276 , n64277 );
and ( n64279 , n63694 , n63683 );
not ( n64280 , n52421 );
not ( n64281 , n63734 );
or ( n64282 , n64280 , n64281 );
not ( n64283 , n51723 );
not ( n64284 , n56451 );
or ( n64285 , n64283 , n64284 );
nand ( n64286 , n40012 , n53228 );
nand ( n64287 , n64285 , n64286 );
nand ( n64288 , n64287 , n54875 );
nand ( n64289 , n64282 , n64288 );
xor ( n64290 , n64279 , n64289 );
not ( n64291 , n57314 );
not ( n64292 , n63744 );
or ( n64293 , n64291 , n64292 );
not ( n64294 , n52377 );
not ( n64295 , n56411 );
or ( n64296 , n64294 , n64295 );
nand ( n64297 , n40452 , n53973 );
nand ( n64298 , n64296 , n64297 );
nand ( n64299 , n64298 , n52004 );
nand ( n64300 , n64293 , n64299 );
xor ( n64301 , n64290 , n64300 );
xor ( n64302 , n64301 , n63523 );
xor ( n64303 , n64302 , n64045 );
xor ( n64304 , n64301 , n63523 );
and ( n64305 , n64304 , n64045 );
and ( n64306 , n64301 , n63523 );
or ( n64307 , n64305 , n64306 );
not ( n64308 , n46564 );
not ( n64309 , n63813 );
or ( n64310 , n64308 , n64309 );
and ( n64311 , n52990 , n42553 );
not ( n64312 , n52990 );
not ( n64313 , n63246 );
and ( n64314 , n64312 , n64313 );
nor ( n64315 , n64311 , n64314 );
nand ( n64316 , n64315 , n49832 );
nand ( n64317 , n64310 , n64316 );
xor ( n64318 , n64317 , n63425 );
not ( n64319 , n47827 );
and ( n64320 , n39331 , n46650 );
not ( n64321 , n39331 );
and ( n64322 , n64321 , n50087 );
or ( n64323 , n64320 , n64322 );
not ( n64324 , n64323 );
or ( n64325 , n64319 , n64324 );
nand ( n64326 , n63780 , n51157 );
nand ( n64327 , n64325 , n64326 );
xor ( n64328 , n64318 , n64327 );
xor ( n64329 , n63987 , n64328 );
xor ( n64330 , n64329 , n63599 );
xor ( n64331 , n63987 , n64328 );
and ( n64332 , n64331 , n63599 );
and ( n64333 , n63987 , n64328 );
or ( n64334 , n64332 , n64333 );
xor ( n64335 , n64062 , n64072 );
and ( n64336 , n64335 , n64083 );
and ( n64337 , n64062 , n64072 );
or ( n64338 , n64336 , n64337 );
xor ( n64339 , n64009 , n64157 );
xor ( n64340 , n64339 , n64085 );
xor ( n64341 , n64009 , n64157 );
and ( n64342 , n64341 , n64085 );
and ( n64343 , n64009 , n64157 );
or ( n64344 , n64342 , n64343 );
xor ( n64345 , n63637 , n64199 );
xor ( n64346 , n64345 , n63727 );
xor ( n64347 , n63637 , n64199 );
and ( n64348 , n64347 , n63727 );
and ( n64349 , n63637 , n64199 );
or ( n64350 , n64348 , n64349 );
xor ( n64351 , n63643 , n64237 );
xor ( n64352 , n64351 , n63804 );
xor ( n64353 , n63643 , n64237 );
and ( n64354 , n64353 , n63804 );
and ( n64355 , n63643 , n64237 );
or ( n64356 , n64354 , n64355 );
xor ( n64357 , n63822 , n64274 );
xor ( n64358 , n64357 , n63828 );
xor ( n64359 , n63822 , n64274 );
and ( n64360 , n64359 , n63828 );
and ( n64361 , n63822 , n64274 );
or ( n64362 , n64360 , n64361 );
xor ( n64363 , n64303 , n64330 );
xor ( n64364 , n64363 , n64340 );
xor ( n64365 , n64303 , n64330 );
and ( n64366 , n64365 , n64340 );
and ( n64367 , n64303 , n64330 );
or ( n64368 , n64366 , n64367 );
xor ( n64369 , n63838 , n63844 );
xor ( n64370 , n64369 , n63850 );
xor ( n64371 , n63838 , n63844 );
and ( n64372 , n64371 , n63850 );
and ( n64373 , n63838 , n63844 );
or ( n64374 , n64372 , n64373 );
xor ( n64375 , n64346 , n64358 );
xor ( n64376 , n64375 , n64352 );
xor ( n64377 , n64346 , n64358 );
and ( n64378 , n64377 , n64352 );
and ( n64379 , n64346 , n64358 );
or ( n64380 , n64378 , n64379 );
xor ( n64381 , n63856 , n64364 );
xor ( n64382 , n64381 , n63862 );
xor ( n64383 , n63856 , n64364 );
and ( n64384 , n64383 , n63862 );
and ( n64385 , n63856 , n64364 );
or ( n64386 , n64384 , n64385 );
xor ( n64387 , n64370 , n63868 );
xor ( n64388 , n64387 , n64376 );
xor ( n64389 , n64370 , n63868 );
and ( n64390 , n64389 , n64376 );
and ( n64391 , n64370 , n63868 );
or ( n64392 , n64390 , n64391 );
xor ( n64393 , n64382 , n63874 );
xor ( n64394 , n64393 , n63880 );
xor ( n64395 , n64382 , n63874 );
and ( n64396 , n64395 , n63880 );
and ( n64397 , n64382 , n63874 );
or ( n64398 , n64396 , n64397 );
xor ( n64399 , n64131 , n64141 );
and ( n64400 , n64399 , n64154 );
and ( n64401 , n64131 , n64141 );
or ( n64402 , n64400 , n64401 );
xor ( n64403 , n64388 , n64394 );
xor ( n64404 , n64403 , n63886 );
xor ( n64405 , n64388 , n64394 );
and ( n64406 , n64405 , n63886 );
and ( n64407 , n64388 , n64394 );
or ( n64408 , n64406 , n64407 );
xor ( n64409 , n64099 , n64108 );
and ( n64410 , n64409 , n64120 );
and ( n64411 , n64099 , n64108 );
or ( n64412 , n64410 , n64411 );
xor ( n64413 , n64174 , n64184 );
and ( n64414 , n64413 , n64197 );
and ( n64415 , n64174 , n64184 );
or ( n64416 , n64414 , n64415 );
xor ( n64417 , n64279 , n64289 );
and ( n64418 , n64417 , n64300 );
and ( n64419 , n64279 , n64289 );
or ( n64420 , n64418 , n64419 );
xor ( n64421 , n64252 , n64261 );
and ( n64422 , n64421 , n64272 );
and ( n64423 , n64252 , n64261 );
or ( n64424 , n64422 , n64423 );
xor ( n64425 , n64213 , n64223 );
and ( n64426 , n64425 , n64234 );
and ( n64427 , n64213 , n64223 );
or ( n64428 , n64426 , n64427 );
xor ( n64429 , n64317 , n63425 );
and ( n64430 , n64429 , n64327 );
and ( n64431 , n64317 , n63425 );
or ( n64432 , n64430 , n64431 );
not ( n64433 , n63932 );
not ( n64434 , n53543 );
or ( n64435 , n64433 , n64434 );
not ( n64436 , n53549 );
not ( n64437 , n53513 );
or ( n64438 , n64436 , n64437 );
nand ( n64439 , n41132 , n51566 );
nand ( n64440 , n64438 , n64439 );
nand ( n64441 , n64440 , n51145 );
nand ( n64442 , n64435 , n64441 );
buf ( n64443 , n63415 );
not ( n64444 , n64443 );
and ( n64445 , n64444 , n50914 );
xor ( n64446 , n64442 , n64445 );
not ( n64447 , n63943 );
not ( n64448 , n54266 );
or ( n64449 , n64447 , n64448 );
not ( n64450 , n52130 );
buf ( n64451 , n49809 );
not ( n64452 , n64451 );
not ( n64453 , n64452 );
or ( n64454 , n64450 , n64453 );
nand ( n64455 , n64451 , n52486 );
nand ( n64456 , n64454 , n64455 );
nand ( n64457 , n51766 , n64456 );
nand ( n64458 , n64449 , n64457 );
xor ( n64459 , n64446 , n64458 );
xor ( n64460 , n64442 , n64445 );
and ( n64461 , n64460 , n64458 );
and ( n64462 , n64442 , n64445 );
or ( n64463 , n64461 , n64462 );
not ( n64464 , n49832 );
not ( n64465 , n47508 );
not ( n64466 , n42651 );
not ( n64467 , n64466 );
or ( n64468 , n64465 , n64467 );
not ( n64469 , n42651 );
or ( n64470 , n64469 , n47508 );
nand ( n64471 , n64468 , n64470 );
not ( n64472 , n64471 );
or ( n64473 , n64464 , n64472 );
nand ( n64474 , n46564 , n64315 );
nand ( n64475 , n64473 , n64474 );
not ( n64476 , n51157 );
not ( n64477 , n64323 );
or ( n64478 , n64476 , n64477 );
not ( n64479 , n45951 );
not ( n64480 , n62715 );
or ( n64481 , n64479 , n64480 );
nand ( n64482 , n39253 , n50087 );
nand ( n64483 , n64481 , n64482 );
nand ( n64484 , n64483 , n45894 );
nand ( n64485 , n64478 , n64484 );
xor ( n64486 , n64475 , n64485 );
xor ( n64487 , n64486 , n63951 );
xor ( n64488 , n64475 , n64485 );
and ( n64489 , n64488 , n63951 );
and ( n64490 , n64475 , n64485 );
or ( n64491 , n64489 , n64490 );
xor ( n64492 , n63985 , n64338 );
xor ( n64493 , n64492 , n64402 );
xor ( n64494 , n63985 , n64338 );
and ( n64495 , n64494 , n64402 );
and ( n64496 , n63985 , n64338 );
or ( n64497 , n64495 , n64496 );
not ( n64498 , n61366 );
not ( n64499 , n64498 );
not ( n64500 , n63997 );
or ( n64501 , n64499 , n64500 );
not ( n64502 , n47803 );
not ( n64503 , n38497 );
or ( n64504 , n64502 , n64503 );
not ( n64505 , n47803 );
nand ( n64506 , n64505 , n38498 );
nand ( n64507 , n64504 , n64506 );
nand ( n64508 , n64507 , n53675 );
nand ( n64509 , n64501 , n64508 );
xor ( n64510 , n64509 , n64412 );
not ( n64511 , n53510 );
not ( n64512 , n49500 );
not ( n64513 , n59402 );
or ( n64514 , n64512 , n64513 );
nand ( n64515 , n39574 , n53997 );
nand ( n64516 , n64514 , n64515 );
not ( n64517 , n64516 );
or ( n64518 , n64511 , n64517 );
buf ( n64519 , n64021 );
nand ( n64520 , n64519 , n48989 );
nand ( n64521 , n64518 , n64520 );
xor ( n64522 , n64510 , n64521 );
xor ( n64523 , n64509 , n64412 );
and ( n64524 , n64523 , n64521 );
and ( n64525 , n64509 , n64412 );
or ( n64526 , n64524 , n64525 );
not ( n64527 , n49026 );
not ( n64528 , n46425 );
not ( n64529 , n62381 );
or ( n64530 , n64528 , n64529 );
nand ( n64531 , n62384 , n46422 );
nand ( n64532 , n64530 , n64531 );
not ( n64533 , n64532 );
or ( n64534 , n64527 , n64533 );
nand ( n64535 , n64031 , n46267 );
nand ( n64536 , n64534 , n64535 );
not ( n64537 , n51865 );
not ( n64538 , n52267 );
not ( n64539 , n58482 );
or ( n64540 , n64538 , n64539 );
nand ( n64541 , n58485 , n51351 );
nand ( n64542 , n64540 , n64541 );
not ( n64543 , n64542 );
or ( n64544 , n64537 , n64543 );
nand ( n64545 , n64039 , n49713 );
nand ( n64546 , n64544 , n64545 );
xor ( n64547 , n64536 , n64546 );
not ( n64548 , n63961 );
not ( n64549 , n63953 );
or ( n64550 , n64548 , n64549 );
and ( n64551 , n46273 , n63390 );
not ( n64552 , n46273 );
and ( n64553 , n64552 , n63921 );
or ( n64554 , n64551 , n64553 );
nand ( n64555 , n64554 , n62843 );
nand ( n64556 , n64550 , n64555 );
and ( n64557 , n57571 , n53946 );
not ( n64558 , n57571 );
and ( n64559 , n64558 , n52840 );
or ( n64560 , n64557 , n64559 );
not ( n64561 , n64560 );
not ( n64562 , n53571 );
or ( n64563 , n64561 , n64562 );
nand ( n64564 , n63970 , n52853 );
nand ( n64565 , n64563 , n64564 );
xor ( n64566 , n64556 , n64565 );
or ( n64567 , n61329 , n63978 );
and ( n64568 , n55918 , n52272 );
and ( n64569 , n53590 , n49190 );
nor ( n64570 , n64568 , n64569 );
or ( n64571 , n64570 , n53618 );
nand ( n64572 , n64567 , n64571 );
xor ( n64573 , n64566 , n64572 );
xor ( n64574 , n64547 , n64573 );
xor ( n64575 , n64536 , n64546 );
and ( n64576 , n64575 , n64573 );
and ( n64577 , n64536 , n64546 );
or ( n64578 , n64576 , n64577 );
or ( n64579 , n54314 , n64059 );
and ( n64580 , n63440 , n54322 );
not ( n64581 , n63440 );
and ( n64582 , n64581 , n54298 );
nor ( n64583 , n64580 , n64582 );
or ( n64584 , n64583 , n55866 );
nand ( n64585 , n64579 , n64584 );
not ( n64586 , n55143 );
not ( n64587 , n64070 );
or ( n64588 , n64586 , n64587 );
not ( n64589 , n58458 );
not ( n64590 , n55148 );
or ( n64591 , n64589 , n64590 );
nand ( n64592 , n55152 , n58459 );
nand ( n64593 , n64591 , n64592 );
nand ( n64594 , n64593 , n55155 );
nand ( n64595 , n64588 , n64594 );
xor ( n64596 , n64585 , n64595 );
not ( n64597 , n55887 );
not ( n64598 , n64081 );
or ( n64599 , n64597 , n64598 );
not ( n64600 , n47527 );
not ( n64601 , n55876 );
or ( n64602 , n64600 , n64601 );
not ( n64603 , n47527 );
nand ( n64604 , n55892 , n64603 );
nand ( n64605 , n64602 , n64604 );
nand ( n64606 , n64605 , n55458 );
nand ( n64607 , n64599 , n64606 );
xor ( n64608 , n64596 , n64607 );
xor ( n64609 , n64459 , n64608 );
not ( n64610 , n49624 );
not ( n64611 , n62510 );
or ( n64612 , n64610 , n64611 );
nand ( n64613 , n59935 , n49630 );
nand ( n64614 , n64612 , n64613 );
not ( n64615 , n64614 );
not ( n64616 , n58908 );
or ( n64617 , n64615 , n64616 );
nand ( n64618 , n64097 , n59570 );
nand ( n64619 , n64617 , n64618 );
or ( n64620 , n60960 , n64106 );
xnor ( n64621 , n47765 , n60285 );
or ( n64622 , n60963 , n64621 );
nand ( n64623 , n64620 , n64622 );
xor ( n64624 , n64619 , n64623 );
not ( n64625 , n61548 );
nand ( n64626 , n64114 , n64116 );
not ( n64627 , n64626 );
or ( n64628 , n64625 , n64627 );
not ( n64629 , n52165 );
not ( n64630 , n61416 );
not ( n64631 , n64630 );
or ( n64632 , n64629 , n64631 );
not ( n64633 , n61537 );
nand ( n64634 , n64633 , n47368 );
nand ( n64635 , n64632 , n64634 );
nand ( n64636 , n64635 , n61557 );
nand ( n64637 , n64628 , n64636 );
xor ( n64638 , n64624 , n64637 );
xor ( n64639 , n64609 , n64638 );
xor ( n64640 , n64459 , n64608 );
and ( n64641 , n64640 , n64638 );
and ( n64642 , n64459 , n64608 );
or ( n64643 , n64641 , n64642 );
not ( n64644 , n64129 );
not ( n64645 , n56775 );
or ( n64646 , n64644 , n64645 );
not ( n64647 , n56501 );
not ( n64648 , n47918 );
not ( n64649 , n58534 );
or ( n64650 , n64648 , n64649 );
nand ( n64651 , n56758 , n49245 );
nand ( n64652 , n64650 , n64651 );
nand ( n64653 , n64647 , n64652 );
nand ( n64654 , n64646 , n64653 );
not ( n64655 , n64139 );
not ( n64656 , n57628 );
or ( n64657 , n64655 , n64656 );
not ( n64658 , n57138 );
not ( n64659 , n54185 );
not ( n64660 , n57633 );
or ( n64661 , n64659 , n64660 );
nand ( n64662 , n57619 , n52712 );
nand ( n64663 , n64661 , n64662 );
nand ( n64664 , n64658 , n64663 );
nand ( n64665 , n64657 , n64664 );
xor ( n64666 , n64654 , n64665 );
not ( n64667 , n64151 );
not ( n64668 , n59445 );
or ( n64669 , n64667 , n64668 );
not ( n64670 , n52033 );
not ( n64671 , n58966 );
or ( n64672 , n64670 , n64671 );
nand ( n64673 , n58642 , n52038 );
nand ( n64674 , n64672 , n64673 );
nand ( n64675 , n61465 , n64674 );
nand ( n64676 , n64669 , n64675 );
xor ( n64677 , n64666 , n64676 );
xor ( n64678 , n64677 , n64424 );
xor ( n64679 , n64678 , n64416 );
xor ( n64680 , n64677 , n64424 );
and ( n64681 , n64680 , n64416 );
and ( n64682 , n64677 , n64424 );
or ( n64683 , n64681 , n64682 );
buf ( n64684 , n63552 );
or ( n64685 , n64684 , n64172 );
not ( n64686 , n49734 );
buf ( n64687 , n62456 );
not ( n64688 , n64687 );
or ( n64689 , n64686 , n64688 );
nand ( n64690 , n62449 , n47821 );
nand ( n64691 , n64689 , n64690 );
not ( n64692 , n64691 );
or ( n64693 , n64166 , n64692 );
nand ( n64694 , n64685 , n64693 );
not ( n64695 , n45861 );
not ( n64696 , n46474 );
not ( n64697 , n64696 );
or ( n64698 , n64695 , n64697 );
nand ( n64699 , n64698 , n46072 );
not ( n64700 , n64699 );
xor ( n64701 , n64694 , n64700 );
not ( n64702 , n50922 );
not ( n64703 , n50898 );
not ( n64704 , n50958 );
or ( n64705 , n64703 , n64704 );
nand ( n64706 , n40677 , n53904 );
nand ( n64707 , n64705 , n64706 );
not ( n64708 , n64707 );
or ( n64709 , n64702 , n64708 );
nand ( n64710 , n64180 , n50911 );
nand ( n64711 , n64709 , n64710 );
xor ( n64712 , n64701 , n64711 );
xor ( n64713 , n64420 , n64712 );
xor ( n64714 , n64713 , n64013 );
xor ( n64715 , n64420 , n64712 );
and ( n64716 , n64715 , n64013 );
and ( n64717 , n64420 , n64712 );
or ( n64718 , n64716 , n64717 );
not ( n64719 , n58168 );
not ( n64720 , n64209 );
or ( n64721 , n64719 , n64720 );
not ( n64722 , n49112 );
not ( n64723 , n53721 );
or ( n64724 , n64722 , n64723 );
nand ( n64725 , n40635 , n60289 );
nand ( n64726 , n64724 , n64725 );
nand ( n64727 , n64726 , n52191 );
nand ( n64728 , n64721 , n64727 );
not ( n64729 , n62654 );
not ( n64730 , n61951 );
not ( n64731 , n53730 );
or ( n64732 , n64730 , n64731 );
nand ( n64733 , n40591 , n61952 );
nand ( n64734 , n64732 , n64733 );
not ( n64735 , n64734 );
or ( n64736 , n64729 , n64735 );
not ( n64737 , n62663 );
nand ( n64738 , n64737 , n64221 );
nand ( n64739 , n64736 , n64738 );
xor ( n64740 , n64728 , n64739 );
not ( n64741 , n50242 );
not ( n64742 , n64230 );
or ( n64743 , n64741 , n64742 );
not ( n64744 , n50232 );
not ( n64745 , n63509 );
or ( n64746 , n64744 , n64745 );
not ( n64747 , n39893 );
nand ( n64748 , n64747 , n49679 );
nand ( n64749 , n64746 , n64748 );
nand ( n64750 , n64749 , n52962 );
nand ( n64751 , n64743 , n64750 );
xor ( n64752 , n64740 , n64751 );
xor ( n64753 , n64432 , n64752 );
xor ( n64754 , n64753 , n64428 );
xor ( n64755 , n64432 , n64752 );
and ( n64756 , n64755 , n64428 );
and ( n64757 , n64432 , n64752 );
or ( n64758 , n64756 , n64757 );
xor ( n64759 , n63991 , n64049 );
not ( n64760 , n52421 );
not ( n64761 , n64287 );
or ( n64762 , n64760 , n64761 );
not ( n64763 , n48856 );
not ( n64764 , n56962 );
or ( n64765 , n64763 , n64764 );
nand ( n64766 , n39962 , n53228 );
nand ( n64767 , n64765 , n64766 );
nand ( n64768 , n64767 , n54875 );
nand ( n64769 , n64762 , n64768 );
not ( n64770 , n63708 );
not ( n64771 , n64193 );
or ( n64772 , n64770 , n64771 );
not ( n64773 , n50304 );
not ( n64774 , n52222 );
or ( n64775 , n64773 , n64774 );
nand ( n64776 , n52223 , n50943 );
nand ( n64777 , n64775 , n64776 );
nand ( n64778 , n64777 , n52757 );
nand ( n64779 , n64772 , n64778 );
xor ( n64780 , n64769 , n64779 );
not ( n64781 , n57314 );
not ( n64782 , n64298 );
or ( n64783 , n64781 , n64782 );
not ( n64784 , n52377 );
not ( n64785 , n56975 );
or ( n64786 , n64784 , n64785 );
nand ( n64787 , n40512 , n53973 );
nand ( n64788 , n64786 , n64787 );
nand ( n64789 , n64788 , n52004 );
nand ( n64790 , n64783 , n64789 );
xor ( n64791 , n64780 , n64790 );
xor ( n64792 , n64759 , n64791 );
xor ( n64793 , n63991 , n64049 );
and ( n64794 , n64793 , n64791 );
and ( n64795 , n63991 , n64049 );
or ( n64796 , n64794 , n64795 );
not ( n64797 , n54623 );
not ( n64798 , n59174 );
not ( n64799 , n55199 );
or ( n64800 , n64798 , n64799 );
nand ( n64801 , n40381 , n55023 );
nand ( n64802 , n64800 , n64801 );
not ( n64803 , n64802 );
or ( n64804 , n64797 , n64803 );
nand ( n64805 , n64250 , n47873 );
nand ( n64806 , n64804 , n64805 );
not ( n64807 , n53104 );
not ( n64808 , n64259 );
or ( n64809 , n64807 , n64808 );
not ( n64810 , n60602 );
not ( n64811 , n40148 );
or ( n64812 , n64810 , n64811 );
nand ( n64813 , n54406 , n52728 );
nand ( n64814 , n64812 , n64813 );
nand ( n64815 , n64814 , n52723 );
nand ( n64816 , n64809 , n64815 );
xor ( n64817 , n64806 , n64816 );
not ( n64818 , n56639 );
not ( n64819 , n59345 );
not ( n64820 , n40225 );
or ( n64821 , n64819 , n64820 );
nand ( n64822 , n54432 , n60617 );
nand ( n64823 , n64821 , n64822 );
not ( n64824 , n64823 );
or ( n64825 , n64818 , n64824 );
nand ( n64826 , n64270 , n59950 );
nand ( n64827 , n64825 , n64826 );
xor ( n64828 , n64817 , n64827 );
xor ( n64829 , n64828 , n64487 );
xor ( n64830 , n64829 , n64493 );
xor ( n64831 , n64828 , n64487 );
and ( n64832 , n64831 , n64493 );
and ( n64833 , n64828 , n64487 );
or ( n64834 , n64832 , n64833 );
xor ( n64835 , n64556 , n64565 );
and ( n64836 , n64835 , n64572 );
and ( n64837 , n64556 , n64565 );
or ( n64838 , n64836 , n64837 );
xor ( n64839 , n64522 , n64574 );
xor ( n64840 , n64839 , n64089 );
xor ( n64841 , n64522 , n64574 );
and ( n64842 , n64841 , n64089 );
and ( n64843 , n64522 , n64574 );
or ( n64844 , n64842 , n64843 );
xor ( n64845 , n64161 , n64639 );
xor ( n64846 , n64845 , n64203 );
xor ( n64847 , n64161 , n64639 );
and ( n64848 , n64847 , n64203 );
and ( n64849 , n64161 , n64639 );
or ( n64850 , n64848 , n64849 );
xor ( n64851 , n64714 , n64679 );
xor ( n64852 , n64851 , n64278 );
xor ( n64853 , n64714 , n64679 );
and ( n64854 , n64853 , n64278 );
and ( n64855 , n64714 , n64679 );
or ( n64856 , n64854 , n64855 );
xor ( n64857 , n64241 , n64792 );
xor ( n64858 , n64857 , n64307 );
xor ( n64859 , n64241 , n64792 );
and ( n64860 , n64859 , n64307 );
and ( n64861 , n64241 , n64792 );
or ( n64862 , n64860 , n64861 );
xor ( n64863 , n64754 , n64334 );
xor ( n64864 , n64863 , n64344 );
xor ( n64865 , n64754 , n64334 );
and ( n64866 , n64865 , n64344 );
and ( n64867 , n64754 , n64334 );
or ( n64868 , n64866 , n64867 );
xor ( n64869 , n64840 , n64830 );
xor ( n64870 , n64869 , n64350 );
xor ( n64871 , n64840 , n64830 );
and ( n64872 , n64871 , n64350 );
and ( n64873 , n64840 , n64830 );
or ( n64874 , n64872 , n64873 );
xor ( n64875 , n64846 , n64356 );
xor ( n64876 , n64875 , n64852 );
xor ( n64877 , n64846 , n64356 );
and ( n64878 , n64877 , n64852 );
and ( n64879 , n64846 , n64356 );
or ( n64880 , n64878 , n64879 );
xor ( n64881 , n64362 , n64858 );
xor ( n64882 , n64881 , n64864 );
xor ( n64883 , n64362 , n64858 );
and ( n64884 , n64883 , n64864 );
and ( n64885 , n64362 , n64858 );
or ( n64886 , n64884 , n64885 );
xor ( n64887 , n64870 , n64368 );
xor ( n64888 , n64887 , n64374 );
xor ( n64889 , n64870 , n64368 );
and ( n64890 , n64889 , n64374 );
and ( n64891 , n64870 , n64368 );
or ( n64892 , n64890 , n64891 );
xor ( n64893 , n64380 , n64876 );
xor ( n64894 , n64893 , n64882 );
xor ( n64895 , n64380 , n64876 );
and ( n64896 , n64895 , n64882 );
and ( n64897 , n64380 , n64876 );
or ( n64898 , n64896 , n64897 );
xor ( n64899 , n64585 , n64595 );
and ( n64900 , n64899 , n64607 );
and ( n64901 , n64585 , n64595 );
or ( n64902 , n64900 , n64901 );
xor ( n64903 , n64888 , n64386 );
xor ( n64904 , n64903 , n64894 );
xor ( n64905 , n64888 , n64386 );
and ( n64906 , n64905 , n64894 );
and ( n64907 , n64888 , n64386 );
or ( n64908 , n64906 , n64907 );
xor ( n64909 , n64392 , n64398 );
xor ( n64910 , n64909 , n64904 );
xor ( n64911 , n64392 , n64398 );
and ( n64912 , n64911 , n64904 );
and ( n64913 , n64392 , n64398 );
or ( n64914 , n64912 , n64913 );
xor ( n64915 , n64654 , n64665 );
and ( n64916 , n64915 , n64676 );
and ( n64917 , n64654 , n64665 );
or ( n64918 , n64916 , n64917 );
xor ( n64919 , n64619 , n64623 );
and ( n64920 , n64919 , n64637 );
and ( n64921 , n64619 , n64623 );
or ( n64922 , n64920 , n64921 );
xor ( n64923 , n64694 , n64700 );
and ( n64924 , n64923 , n64711 );
and ( n64925 , n64694 , n64700 );
or ( n64926 , n64924 , n64925 );
xor ( n64927 , n64769 , n64779 );
and ( n64928 , n64927 , n64790 );
and ( n64929 , n64769 , n64779 );
or ( n64930 , n64928 , n64929 );
xor ( n64931 , n64806 , n64816 );
and ( n64932 , n64931 , n64827 );
and ( n64933 , n64806 , n64816 );
or ( n64934 , n64932 , n64933 );
xor ( n64935 , n64728 , n64739 );
and ( n64936 , n64935 , n64751 );
and ( n64937 , n64728 , n64739 );
or ( n64938 , n64936 , n64937 );
not ( n64939 , n64560 );
not ( n64940 , n52853 );
or ( n64941 , n64939 , n64940 );
not ( n64942 , n49545 );
not ( n64943 , n64942 );
not ( n64944 , n52837 );
or ( n64945 , n64943 , n64944 );
nand ( n64946 , n55481 , n50004 );
nand ( n64947 , n64945 , n64946 );
nand ( n64948 , n53571 , n64947 );
nand ( n64949 , n64941 , n64948 );
and ( n64950 , n63922 , n54722 );
xor ( n64951 , n64949 , n64950 );
not ( n64952 , n53609 );
not ( n64953 , n64570 );
not ( n64954 , n64953 );
or ( n64955 , n64952 , n64954 );
not ( n64956 , n49001 );
not ( n64957 , n53591 );
or ( n64958 , n64956 , n64957 );
not ( n64959 , n55917 );
nand ( n64960 , n64959 , n48997 );
nand ( n64961 , n64958 , n64960 );
nand ( n64962 , n64961 , n53326 );
nand ( n64963 , n64955 , n64962 );
xor ( n64964 , n64951 , n64963 );
xor ( n64965 , n64949 , n64950 );
and ( n64966 , n64965 , n64963 );
and ( n64967 , n64949 , n64950 );
or ( n64968 , n64966 , n64967 );
or ( n64969 , n62338 , n64583 );
not ( n64970 , n56274 );
and ( n64971 , n64970 , n48486 );
not ( n64972 , n48486 );
and ( n64973 , n54298 , n64972 );
nor ( n64974 , n64971 , n64973 );
or ( n64975 , n54326 , n64974 );
nand ( n64976 , n64969 , n64975 );
not ( n64977 , n64593 );
not ( n64978 , n55576 );
or ( n64979 , n64977 , n64978 );
not ( n64980 , n58915 );
not ( n64981 , n55148 );
or ( n64982 , n64980 , n64981 );
nand ( n64983 , n55118 , n58914 );
nand ( n64984 , n64982 , n64983 );
nand ( n64985 , n64984 , n55157 );
nand ( n64986 , n64979 , n64985 );
xor ( n64987 , n64976 , n64986 );
not ( n64988 , n56281 );
not ( n64989 , n64605 );
or ( n64990 , n64988 , n64989 );
not ( n64991 , n58180 );
not ( n64992 , n55893 );
or ( n64993 , n64991 , n64992 );
nand ( n64994 , n55892 , n41416 );
nand ( n64995 , n64993 , n64994 );
nand ( n64996 , n64995 , n59984 );
nand ( n64997 , n64990 , n64996 );
xor ( n64998 , n64987 , n64997 );
xor ( n64999 , n64976 , n64986 );
and ( n65000 , n64999 , n64997 );
and ( n65001 , n64976 , n64986 );
or ( n65002 , n65000 , n65001 );
xor ( n65003 , n64918 , n64922 );
not ( n65004 , n53510 );
not ( n65005 , n49500 );
not ( n65006 , n39056 );
not ( n65007 , n65006 );
or ( n65008 , n65005 , n65007 );
nand ( n65009 , n39056 , n47979 );
nand ( n65010 , n65008 , n65009 );
not ( n65011 , n65010 );
or ( n65012 , n65004 , n65011 );
nand ( n65013 , n64516 , n48989 );
nand ( n65014 , n65012 , n65013 );
xor ( n65015 , n65003 , n65014 );
xor ( n65016 , n64918 , n64922 );
and ( n65017 , n65016 , n65014 );
and ( n65018 , n64918 , n64922 );
or ( n65019 , n65017 , n65018 );
not ( n65020 , n54875 );
not ( n65021 , n48856 );
not ( n65022 , n39844 );
or ( n65023 , n65021 , n65022 );
nand ( n65024 , n61888 , n53228 );
nand ( n65025 , n65023 , n65024 );
not ( n65026 , n65025 );
or ( n65027 , n65020 , n65026 );
nand ( n65028 , n64767 , n52421 );
nand ( n65029 , n65027 , n65028 );
not ( n65030 , n45842 );
not ( n65031 , n64471 );
or ( n65032 , n65030 , n65031 );
nand ( n65033 , n47508 , n49832 );
nand ( n65034 , n65032 , n65033 );
xor ( n65035 , n65029 , n65034 );
not ( n65036 , n51865 );
not ( n65037 , n52267 );
not ( n65038 , n60906 );
or ( n65039 , n65037 , n65038 );
nand ( n65040 , n39714 , n51351 );
nand ( n65041 , n65039 , n65040 );
not ( n65042 , n65041 );
or ( n65043 , n65036 , n65042 );
nand ( n65044 , n64542 , n49713 );
nand ( n65045 , n65043 , n65044 );
xor ( n65046 , n65035 , n65045 );
xor ( n65047 , n65029 , n65034 );
and ( n65048 , n65047 , n65045 );
and ( n65049 , n65029 , n65034 );
or ( n65050 , n65048 , n65049 );
not ( n65051 , n48073 );
not ( n65052 , n50263 );
not ( n65053 , n62909 );
or ( n65054 , n65052 , n65053 );
nand ( n65055 , n62913 , n52080 );
nand ( n65056 , n65054 , n65055 );
not ( n65057 , n65056 );
or ( n65058 , n65051 , n65057 );
nand ( n65059 , n64483 , n48295 );
nand ( n65060 , n65058 , n65059 );
not ( n65061 , n50242 );
not ( n65062 , n64749 );
or ( n65063 , n65061 , n65062 );
not ( n65064 , n48645 );
not ( n65065 , n58047 );
or ( n65066 , n65064 , n65065 );
nand ( n65067 , n39779 , n49679 );
nand ( n65068 , n65066 , n65067 );
nand ( n65069 , n52962 , n65068 );
nand ( n65070 , n65063 , n65069 );
xor ( n65071 , n65060 , n65070 );
xor ( n65072 , n65071 , n64964 );
xor ( n65073 , n65060 , n65070 );
and ( n65074 , n65073 , n64964 );
and ( n65075 , n65060 , n65070 );
or ( n65076 , n65074 , n65075 );
not ( n65077 , n64691 );
not ( n65078 , n62463 );
or ( n65079 , n65077 , n65078 );
not ( n65080 , n47227 );
not ( n65081 , n64167 );
or ( n65082 , n65080 , n65081 );
not ( n65083 , n64687 );
nand ( n65084 , n65083 , n47589 );
nand ( n65085 , n65082 , n65084 );
nand ( n65086 , n65085 , n62467 );
nand ( n65087 , n65079 , n65086 );
not ( n65088 , n64554 );
not ( n65089 , n63411 );
not ( n65090 , n65089 );
or ( n65091 , n65088 , n65090 );
buf ( n65092 , n63398 );
not ( n65093 , n47646 );
not ( n65094 , n63922 );
not ( n65095 , n65094 );
or ( n65096 , n65093 , n65095 );
nand ( n65097 , n63922 , n47650 );
nand ( n65098 , n65096 , n65097 );
nand ( n65099 , n65092 , n65098 );
nand ( n65100 , n65091 , n65099 );
xor ( n65101 , n65087 , n65100 );
not ( n65102 , n51533 );
buf ( n65103 , n51505 );
not ( n65104 , n65103 );
not ( n65105 , n50654 );
or ( n65106 , n65104 , n65105 );
nand ( n65107 , n40692 , n53928 );
nand ( n65108 , n65106 , n65107 );
not ( n65109 , n65108 );
or ( n65110 , n65102 , n65109 );
not ( n65111 , n56355 );
not ( n65112 , n65111 );
nand ( n65113 , n65112 , n64440 );
nand ( n65114 , n65110 , n65113 );
xor ( n65115 , n65101 , n65114 );
xor ( n65116 , n64998 , n65115 );
not ( n65117 , n64614 );
not ( n65118 , n60539 );
or ( n65119 , n65117 , n65118 );
not ( n65120 , n51792 );
not ( n65121 , n62513 );
not ( n65122 , n65121 );
or ( n65123 , n65120 , n65122 );
nand ( n65124 , n59341 , n48829 );
nand ( n65125 , n65123 , n65124 );
nand ( n65126 , n59575 , n65125 );
nand ( n65127 , n65119 , n65126 );
not ( n65128 , n64621 );
not ( n65129 , n65128 );
not ( n65130 , n60960 );
not ( n65131 , n65130 );
or ( n65132 , n65129 , n65131 );
and ( n65133 , n51204 , n64102 );
not ( n65134 , n51204 );
and ( n65135 , n65134 , n60285 );
nor ( n65136 , n65133 , n65135 );
not ( n65137 , n65136 );
nand ( n65138 , n65137 , n60427 );
nand ( n65139 , n65132 , n65138 );
xor ( n65140 , n65127 , n65139 );
not ( n65141 , n64111 );
not ( n65142 , n64635 );
or ( n65143 , n65141 , n65142 );
not ( n65144 , n61557 );
not ( n65145 , n48898 );
not ( n65146 , n64630 );
or ( n65147 , n65145 , n65146 );
not ( n65148 , n61417 );
nand ( n65149 , n65148 , n48897 );
nand ( n65150 , n65147 , n65149 );
not ( n65151 , n65150 );
or ( n65152 , n65144 , n65151 );
nand ( n65153 , n65143 , n65152 );
xor ( n65154 , n65140 , n65153 );
xor ( n65155 , n65116 , n65154 );
xor ( n65156 , n64998 , n65115 );
and ( n65157 , n65156 , n65154 );
and ( n65158 , n64998 , n65115 );
or ( n65159 , n65157 , n65158 );
not ( n65160 , n56776 );
not ( n65161 , n64652 );
or ( n65162 , n65160 , n65161 );
and ( n65163 , n56785 , n57182 );
and ( n65164 , n56786 , n57186 );
nor ( n65165 , n65163 , n65164 );
not ( n65166 , n56780 );
or ( n65167 , n65165 , n65166 );
nand ( n65168 , n65162 , n65167 );
not ( n65169 , n57628 );
not ( n65170 , n64663 );
or ( n65171 , n65169 , n65170 );
not ( n65172 , n59435 );
and ( n65173 , n48983 , n57615 );
not ( n65174 , n48983 );
not ( n65175 , n59437 );
and ( n65176 , n65174 , n65175 );
nor ( n65177 , n65173 , n65176 );
or ( n65178 , n65172 , n65177 );
nand ( n65179 , n65171 , n65178 );
xor ( n65180 , n65168 , n65179 );
not ( n65181 , n64674 );
or ( n65182 , n64143 , n65181 );
buf ( n65183 , n58433 );
not ( n65184 , n65183 );
and ( n65185 , n51670 , n65184 );
not ( n65186 , n51670 );
not ( n65187 , n58642 );
and ( n65188 , n65186 , n65187 );
nor ( n65189 , n65185 , n65188 );
or ( n65190 , n64146 , n65189 );
nand ( n65191 , n65182 , n65190 );
xor ( n65192 , n65180 , n65191 );
xor ( n65193 , n65192 , n64926 );
xor ( n65194 , n65193 , n64930 );
xor ( n65195 , n65192 , n64926 );
and ( n65196 , n65195 , n64930 );
and ( n65197 , n65192 , n64926 );
or ( n65198 , n65196 , n65197 );
xor ( n65199 , n64934 , n64497 );
not ( n65200 , n51223 );
not ( n65201 , n50898 );
not ( n65202 , n59176 );
or ( n65203 , n65201 , n65202 );
nand ( n65204 , n40734 , n50894 );
nand ( n65205 , n65203 , n65204 );
not ( n65206 , n65205 );
or ( n65207 , n65200 , n65206 );
nand ( n65208 , n64707 , n52526 );
nand ( n65209 , n65207 , n65208 );
xor ( n65210 , n64699 , n65209 );
not ( n65211 , n64456 );
or ( n65212 , n52481 , n65211 );
not ( n65213 , n41037 );
not ( n65214 , n59999 );
or ( n65215 , n65213 , n65214 );
not ( n65216 , n50667 );
nand ( n65217 , n65216 , n52130 );
nand ( n65218 , n65215 , n65217 );
not ( n65219 , n65218 );
or ( n65220 , n62302 , n65219 );
nand ( n65221 , n65212 , n65220 );
not ( n65222 , n65221 );
xor ( n65223 , n65210 , n65222 );
xor ( n65224 , n65199 , n65223 );
xor ( n65225 , n64934 , n64497 );
and ( n65226 , n65225 , n65223 );
and ( n65227 , n64934 , n64497 );
or ( n65228 , n65226 , n65227 );
xor ( n65229 , n64938 , n64491 );
xor ( n65230 , n65229 , n64526 );
xor ( n65231 , n64938 , n64491 );
and ( n65232 , n65231 , n64526 );
and ( n65233 , n64938 , n64491 );
or ( n65234 , n65232 , n65233 );
not ( n65235 , n57314 );
not ( n65236 , n64788 );
or ( n65237 , n65235 , n65236 );
not ( n65238 , n52377 );
not ( n65239 , n56454 );
or ( n65240 , n65238 , n65239 );
nand ( n65241 , n40012 , n55013 );
nand ( n65242 , n65240 , n65241 );
nand ( n65243 , n65242 , n52004 );
nand ( n65244 , n65237 , n65243 );
not ( n65245 , n54623 );
not ( n65246 , n51680 );
not ( n65247 , n56411 );
or ( n65248 , n65246 , n65247 );
nand ( n65249 , n56412 , n51684 );
nand ( n65250 , n65248 , n65249 );
not ( n65251 , n65250 );
or ( n65252 , n65245 , n65251 );
nand ( n65253 , n64802 , n47873 );
nand ( n65254 , n65252 , n65253 );
xor ( n65255 , n65244 , n65254 );
not ( n65256 , n58977 );
not ( n65257 , n58982 );
not ( n65258 , n55641 );
or ( n65259 , n65257 , n65258 );
nand ( n65260 , n40389 , n52728 );
nand ( n65261 , n65259 , n65260 );
not ( n65262 , n65261 );
or ( n65263 , n65256 , n65262 );
nand ( n65264 , n64814 , n53104 );
nand ( n65265 , n65263 , n65264 );
xor ( n65266 , n65255 , n65265 );
not ( n65267 , n59950 );
not ( n65268 , n64823 );
or ( n65269 , n65267 , n65268 );
or ( n65270 , n59345 , n40363 );
nand ( n65271 , n59345 , n40363 );
nand ( n65272 , n65270 , n65271 , n56639 );
nand ( n65273 , n65269 , n65272 );
not ( n65274 , n64726 );
not ( n65275 , n58168 );
or ( n65276 , n65274 , n65275 );
not ( n65277 , n49112 );
not ( n65278 , n54020 );
or ( n65279 , n65277 , n65278 );
nand ( n65280 , n40377 , n60289 );
nand ( n65281 , n65279 , n65280 );
nand ( n65282 , n65281 , n52191 );
nand ( n65283 , n65276 , n65282 );
xor ( n65284 , n65273 , n65283 );
not ( n65285 , n62654 );
not ( n65286 , n61951 );
not ( n65287 , n54046 );
or ( n65288 , n65286 , n65287 );
nand ( n65289 , n40626 , n61947 );
nand ( n65290 , n65288 , n65289 );
not ( n65291 , n65290 );
or ( n65292 , n65285 , n65291 );
nand ( n65293 , n64734 , n62664 );
nand ( n65294 , n65292 , n65293 );
xor ( n65295 , n65284 , n65294 );
xor ( n65296 , n65266 , n65295 );
xor ( n65297 , n65296 , n64578 );
xor ( n65298 , n65266 , n65295 );
and ( n65299 , n65298 , n64578 );
and ( n65300 , n65266 , n65295 );
or ( n65301 , n65299 , n65300 );
not ( n65302 , n63708 );
not ( n65303 , n64777 );
or ( n65304 , n65302 , n65303 );
not ( n65305 , n64190 );
not ( n65306 , n61142 );
or ( n65307 , n65305 , n65306 );
nand ( n65308 , n51916 , n50943 );
nand ( n65309 , n65307 , n65308 );
nand ( n65310 , n65309 , n52757 );
nand ( n65311 , n65304 , n65310 );
not ( n65312 , n46267 );
not ( n65313 , n64532 );
or ( n65314 , n65312 , n65313 );
not ( n65315 , n46425 );
not ( n65316 , n63246 );
or ( n65317 , n65315 , n65316 );
not ( n65318 , n46425 );
nand ( n65319 , n65318 , n42554 );
nand ( n65320 , n65317 , n65319 );
nand ( n65321 , n65320 , n49026 );
nand ( n65322 , n65314 , n65321 );
xor ( n65323 , n65311 , n65322 );
xor ( n65324 , n65323 , n64463 );
xor ( n65325 , n65324 , n64643 );
xor ( n65326 , n65325 , n65046 );
xor ( n65327 , n65324 , n64643 );
and ( n65328 , n65327 , n65046 );
and ( n65329 , n65324 , n64643 );
or ( n65330 , n65328 , n65329 );
xor ( n65331 , n65015 , n65072 );
not ( n65332 , n47407 );
not ( n65333 , n64507 );
or ( n65334 , n65332 , n65333 );
and ( n65335 , n39330 , n48727 );
not ( n65336 , n39330 );
and ( n65337 , n65336 , n54028 );
or ( n65338 , n65335 , n65337 );
nand ( n65339 , n65338 , n53675 );
nand ( n65340 , n65334 , n65339 );
xor ( n65341 , n65340 , n64838 );
xor ( n65342 , n65341 , n64902 );
xor ( n65343 , n65331 , n65342 );
xor ( n65344 , n65015 , n65072 );
and ( n65345 , n65344 , n65342 );
and ( n65346 , n65015 , n65072 );
or ( n65347 , n65345 , n65346 );
xor ( n65348 , n65168 , n65179 );
and ( n65349 , n65348 , n65191 );
and ( n65350 , n65168 , n65179 );
or ( n65351 , n65349 , n65350 );
xor ( n65352 , n64683 , n65155 );
xor ( n65353 , n65352 , n64758 );
xor ( n65354 , n64683 , n65155 );
and ( n65355 , n65354 , n64758 );
and ( n65356 , n64683 , n65155 );
or ( n65357 , n65355 , n65356 );
xor ( n65358 , n64796 , n65194 );
xor ( n65359 , n65358 , n64718 );
xor ( n65360 , n64796 , n65194 );
and ( n65361 , n65360 , n64718 );
and ( n65362 , n64796 , n65194 );
or ( n65363 , n65361 , n65362 );
xor ( n65364 , n65224 , n65230 );
xor ( n65365 , n65364 , n64844 );
xor ( n65366 , n65224 , n65230 );
and ( n65367 , n65366 , n64844 );
and ( n65368 , n65224 , n65230 );
or ( n65369 , n65367 , n65368 );
xor ( n65370 , n65297 , n64834 );
xor ( n65371 , n65370 , n65343 );
xor ( n65372 , n65297 , n64834 );
and ( n65373 , n65372 , n65343 );
and ( n65374 , n65297 , n64834 );
or ( n65375 , n65373 , n65374 );
xor ( n65376 , n64850 , n65326 );
xor ( n65377 , n65376 , n65353 );
xor ( n65378 , n64850 , n65326 );
and ( n65379 , n65378 , n65353 );
and ( n65380 , n64850 , n65326 );
or ( n65381 , n65379 , n65380 );
xor ( n65382 , n64856 , n64862 );
xor ( n65383 , n65382 , n65359 );
xor ( n65384 , n64856 , n64862 );
and ( n65385 , n65384 , n65359 );
and ( n65386 , n64856 , n64862 );
or ( n65387 , n65385 , n65386 );
xor ( n65388 , n65371 , n64868 );
xor ( n65389 , n65388 , n65365 );
xor ( n65390 , n65371 , n64868 );
and ( n65391 , n65390 , n65365 );
and ( n65392 , n65371 , n64868 );
or ( n65393 , n65391 , n65392 );
xor ( n65394 , n65377 , n64874 );
xor ( n65395 , n65394 , n64880 );
xor ( n65396 , n65377 , n64874 );
and ( n65397 , n65396 , n64880 );
and ( n65398 , n65377 , n64874 );
or ( n65399 , n65397 , n65398 );
xor ( n65400 , n65383 , n64886 );
xor ( n65401 , n65400 , n65389 );
xor ( n65402 , n65383 , n64886 );
and ( n65403 , n65402 , n65389 );
and ( n65404 , n65383 , n64886 );
or ( n65405 , n65403 , n65404 );
xor ( n65406 , n64892 , n65395 );
xor ( n65407 , n65406 , n64898 );
xor ( n65408 , n64892 , n65395 );
and ( n65409 , n65408 , n64898 );
and ( n65410 , n64892 , n65395 );
or ( n65411 , n65409 , n65410 );
xor ( n65412 , n65127 , n65139 );
and ( n65413 , n65412 , n65153 );
and ( n65414 , n65127 , n65139 );
or ( n65415 , n65413 , n65414 );
xor ( n65416 , n65401 , n65407 );
xor ( n65417 , n65416 , n64908 );
xor ( n65418 , n65401 , n65407 );
and ( n65419 , n65418 , n64908 );
and ( n65420 , n65401 , n65407 );
or ( n65421 , n65419 , n65420 );
xor ( n65422 , n65087 , n65100 );
and ( n65423 , n65422 , n65114 );
and ( n65424 , n65087 , n65100 );
or ( n65425 , n65423 , n65424 );
xor ( n65426 , n64699 , n65209 );
and ( n65427 , n65426 , n65222 );
and ( n65428 , n64699 , n65209 );
or ( n65429 , n65427 , n65428 );
xor ( n65430 , n65244 , n65254 );
and ( n65431 , n65430 , n65265 );
and ( n65432 , n65244 , n65254 );
or ( n65433 , n65431 , n65432 );
xor ( n65434 , n65273 , n65283 );
and ( n65435 , n65434 , n65294 );
and ( n65436 , n65273 , n65283 );
or ( n65437 , n65435 , n65436 );
xor ( n65438 , n65311 , n65322 );
and ( n65439 , n65438 , n64463 );
and ( n65440 , n65311 , n65322 );
or ( n65441 , n65439 , n65440 );
xor ( n65442 , n65340 , n64838 );
and ( n65443 , n65442 , n64902 );
and ( n65444 , n65340 , n64838 );
or ( n65445 , n65443 , n65444 );
or ( n65446 , n46448 , n45748 );
nand ( n65447 , n65446 , n48952 );
not ( n65448 , n51765 );
not ( n65449 , n50403 );
not ( n65450 , n52870 );
or ( n65451 , n65449 , n65450 );
nand ( n65452 , n52113 , n41131 );
nand ( n65453 , n65451 , n65452 );
not ( n65454 , n65453 );
or ( n65455 , n65448 , n65454 );
nand ( n65456 , n65218 , n56310 );
nand ( n65457 , n65455 , n65456 );
xor ( n65458 , n65447 , n65457 );
not ( n65459 , n64947 );
not ( n65460 , n52852 );
or ( n65461 , n65459 , n65460 );
not ( n65462 , n50827 );
not ( n65463 , n57253 );
or ( n65464 , n65462 , n65463 );
nand ( n65465 , n55481 , n49806 );
nand ( n65466 , n65464 , n65465 );
nand ( n65467 , n53571 , n65466 );
nand ( n65468 , n65461 , n65467 );
xor ( n65469 , n65458 , n65468 );
xor ( n65470 , n65447 , n65457 );
and ( n65471 , n65470 , n65468 );
and ( n65472 , n65447 , n65457 );
or ( n65473 , n65471 , n65472 );
not ( n65474 , n65094 );
and ( n65475 , n65474 , n46273 );
not ( n65476 , n49838 );
not ( n65477 , n56802 );
or ( n65478 , n65476 , n65477 );
nand ( n65479 , n53590 , n49210 );
nand ( n65480 , n65478 , n65479 );
not ( n65481 , n65480 );
not ( n65482 , n53619 );
or ( n65483 , n65481 , n65482 );
not ( n65484 , n61329 );
nand ( n65485 , n65484 , n64961 );
nand ( n65486 , n65483 , n65485 );
xor ( n65487 , n65475 , n65486 );
not ( n65488 , n54315 );
or ( n65489 , n65488 , n64974 );
not ( n65490 , n55276 );
not ( n65491 , n49823 );
or ( n65492 , n65490 , n65491 );
not ( n65493 , n52272 );
nand ( n65494 , n65493 , n54298 );
nand ( n65495 , n65492 , n65494 );
not ( n65496 , n65495 );
or ( n65497 , n65496 , n55866 );
nand ( n65498 , n65489 , n65497 );
xor ( n65499 , n65487 , n65498 );
xor ( n65500 , n65475 , n65486 );
and ( n65501 , n65500 , n65498 );
and ( n65502 , n65475 , n65486 );
or ( n65503 , n65501 , n65502 );
not ( n65504 , n53675 );
not ( n65505 , n47803 );
not ( n65506 , n62715 );
or ( n65507 , n65505 , n65506 );
nand ( n65508 , n39253 , n48727 );
nand ( n65509 , n65507 , n65508 );
not ( n65510 , n65509 );
or ( n65511 , n65504 , n65510 );
nand ( n65512 , n65338 , n47407 );
nand ( n65513 , n65511 , n65512 );
xor ( n65514 , n65513 , n65351 );
xor ( n65515 , n65514 , n65415 );
xor ( n65516 , n65513 , n65351 );
and ( n65517 , n65516 , n65415 );
and ( n65518 , n65513 , n65351 );
or ( n65519 , n65517 , n65518 );
not ( n65520 , n53510 );
not ( n65521 , n49500 );
not ( n65522 , n62394 );
or ( n65523 , n65521 , n65522 );
nand ( n65524 , n38499 , n53997 );
nand ( n65525 , n65523 , n65524 );
not ( n65526 , n65525 );
or ( n65527 , n65520 , n65526 );
nand ( n65528 , n65010 , n49252 );
nand ( n65529 , n65527 , n65528 );
not ( n65530 , n51865 );
not ( n65531 , n49707 );
not ( n65532 , n39574 );
not ( n65533 , n65532 );
or ( n65534 , n65531 , n65533 );
nand ( n65535 , n39574 , n51351 );
nand ( n65536 , n65534 , n65535 );
not ( n65537 , n65536 );
or ( n65538 , n65530 , n65537 );
nand ( n65539 , n65041 , n49713 );
nand ( n65540 , n65538 , n65539 );
xor ( n65541 , n65529 , n65540 );
not ( n65542 , n65056 );
or ( n65543 , n65542 , n46775 );
and ( n65544 , n50263 , n42399 );
not ( n65545 , n50263 );
not ( n65546 , n42399 );
and ( n65547 , n65545 , n65546 );
or ( n65548 , n65544 , n65547 );
not ( n65549 , n65548 );
or ( n65550 , n65549 , n56080 );
nand ( n65551 , n65543 , n65550 );
xor ( n65552 , n65541 , n65551 );
xor ( n65553 , n65529 , n65540 );
and ( n65554 , n65553 , n65551 );
and ( n65555 , n65529 , n65540 );
or ( n65556 , n65554 , n65555 );
not ( n65557 , n52962 );
not ( n65558 , n48645 );
not ( n65559 , n58482 );
or ( n65560 , n65558 , n65559 );
nand ( n65561 , n39680 , n52048 );
nand ( n65562 , n65560 , n65561 );
not ( n65563 , n65562 );
or ( n65564 , n65557 , n65563 );
nand ( n65565 , n65068 , n52970 );
nand ( n65566 , n65564 , n65565 );
xor ( n65567 , n65566 , n65499 );
xor ( n65568 , n65567 , n65425 );
xor ( n65569 , n65566 , n65499 );
and ( n65570 , n65569 , n65425 );
and ( n65571 , n65566 , n65499 );
or ( n65572 , n65570 , n65571 );
not ( n65573 , n64984 );
not ( n65574 , n55143 );
or ( n65575 , n65573 , n65574 );
not ( n65576 , n41532 );
not ( n65577 , n55151 );
or ( n65578 , n65576 , n65577 );
nand ( n65579 , n55118 , n49233 );
nand ( n65580 , n65578 , n65579 );
nand ( n65581 , n65580 , n55933 );
nand ( n65582 , n65575 , n65581 );
not ( n65583 , n64995 );
not ( n65584 , n56281 );
or ( n65585 , n65583 , n65584 );
not ( n65586 , n58454 );
not ( n65587 , n55876 );
or ( n65588 , n65586 , n65587 );
nand ( n65589 , n59499 , n58459 );
nand ( n65590 , n65588 , n65589 );
nand ( n65591 , n65590 , n55458 );
nand ( n65592 , n65585 , n65591 );
xor ( n65593 , n65582 , n65592 );
not ( n65594 , n56776 );
or ( n65595 , n65594 , n65165 );
and ( n65596 , n57665 , n47527 );
and ( n65597 , n59045 , n59388 );
nor ( n65598 , n65596 , n65597 );
or ( n65599 , n65166 , n65598 );
nand ( n65600 , n65595 , n65599 );
xor ( n65601 , n65593 , n65600 );
xor ( n65602 , n65469 , n65601 );
or ( n65603 , n65136 , n60423 );
and ( n65604 , n64102 , n49624 );
and ( n65605 , n60969 , n49630 );
nor ( n65606 , n65604 , n65605 );
not ( n65607 , n59855 );
or ( n65608 , n65606 , n65607 );
nand ( n65609 , n65603 , n65608 );
not ( n65610 , n65150 );
not ( n65611 , n61548 );
or ( n65612 , n65610 , n65611 );
not ( n65613 , n47765 );
not ( n65614 , n61537 );
or ( n65615 , n65613 , n65614 );
nand ( n65616 , n61416 , n48589 );
nand ( n65617 , n65615 , n65616 );
nand ( n65618 , n65617 , n62428 );
nand ( n65619 , n65612 , n65618 );
xor ( n65620 , n65609 , n65619 );
not ( n65621 , n65085 );
not ( n65622 , n62463 );
or ( n65623 , n65621 , n65622 );
not ( n65624 , n49654 );
not ( n65625 , n62452 );
or ( n65626 , n65624 , n65625 );
nand ( n65627 , n62451 , n47368 );
nand ( n65628 , n65626 , n65627 );
nand ( n65629 , n65628 , n62467 );
nand ( n65630 , n65623 , n65629 );
xor ( n65631 , n65620 , n65630 );
xor ( n65632 , n65602 , n65631 );
xor ( n65633 , n65469 , n65601 );
and ( n65634 , n65633 , n65631 );
and ( n65635 , n65469 , n65601 );
or ( n65636 , n65634 , n65635 );
or ( n65637 , n65169 , n65177 );
not ( n65638 , n57631 );
and ( n65639 , n57615 , n56727 );
and ( n65640 , n57619 , n56731 );
nor ( n65641 , n65639 , n65640 );
or ( n65642 , n65638 , n65641 );
nand ( n65643 , n65637 , n65642 );
not ( n65644 , n65189 );
not ( n65645 , n65644 );
not ( n65646 , n63079 );
not ( n65647 , n65646 );
or ( n65648 , n65645 , n65647 );
not ( n65649 , n54185 );
not ( n65650 , n65183 );
or ( n65651 , n65649 , n65650 );
not ( n65652 , n58433 );
nand ( n65653 , n65652 , n52712 );
nand ( n65654 , n65651 , n65653 );
nand ( n65655 , n61465 , n65654 );
nand ( n65656 , n65648 , n65655 );
xor ( n65657 , n65643 , n65656 );
not ( n65658 , n65125 );
not ( n65659 , n62506 );
or ( n65660 , n65658 , n65659 );
not ( n65661 , n52033 );
not ( n65662 , n59340 );
or ( n65663 , n65661 , n65662 );
not ( n65664 , n63587 );
nand ( n65665 , n65664 , n52038 );
nand ( n65666 , n65663 , n65665 );
nand ( n65667 , n59575 , n65666 );
nand ( n65668 , n65660 , n65667 );
xor ( n65669 , n65657 , n65668 );
xor ( n65670 , n65669 , n65429 );
xor ( n65671 , n65670 , n65433 );
xor ( n65672 , n65669 , n65429 );
and ( n65673 , n65672 , n65433 );
and ( n65674 , n65669 , n65429 );
or ( n65675 , n65673 , n65674 );
xor ( n65676 , n65437 , n65050 );
xor ( n65677 , n65676 , n65441 );
xor ( n65678 , n65437 , n65050 );
and ( n65679 , n65678 , n65441 );
and ( n65680 , n65437 , n65050 );
or ( n65681 , n65679 , n65680 );
xor ( n65682 , n65445 , n65019 );
not ( n65683 , n62664 );
not ( n65684 , n65290 );
or ( n65685 , n65683 , n65684 );
not ( n65686 , n61951 );
not ( n65687 , n52906 );
or ( n65688 , n65686 , n65687 );
nand ( n65689 , n52907 , n61947 );
nand ( n65690 , n65688 , n65689 );
nand ( n65691 , n65690 , n62654 );
nand ( n65692 , n65685 , n65691 );
not ( n65693 , n52757 );
not ( n65694 , n53730 );
not ( n65695 , n64190 );
or ( n65696 , n65694 , n65695 );
nand ( n65697 , n52212 , n50943 );
nand ( n65698 , n65696 , n65697 );
not ( n65699 , n65698 );
or ( n65700 , n65693 , n65699 );
nand ( n65701 , n65309 , n63708 );
nand ( n65702 , n65700 , n65701 );
xor ( n65703 , n65692 , n65702 );
not ( n65704 , n54875 );
not ( n65705 , n51723 );
not ( n65706 , n39894 );
or ( n65707 , n65705 , n65706 );
not ( n65708 , n39893 );
nand ( n65709 , n65708 , n53228 );
nand ( n65710 , n65707 , n65709 );
not ( n65711 , n65710 );
or ( n65712 , n65704 , n65711 );
nand ( n65713 , n65025 , n52421 );
nand ( n65714 , n65712 , n65713 );
xor ( n65715 , n65703 , n65714 );
xor ( n65716 , n65682 , n65715 );
xor ( n65717 , n65445 , n65019 );
and ( n65718 , n65717 , n65715 );
and ( n65719 , n65445 , n65019 );
or ( n65720 , n65718 , n65719 );
not ( n65721 , n53104 );
not ( n65722 , n65261 );
or ( n65723 , n65721 , n65722 );
not ( n65724 , n60602 );
not ( n65725 , n40381 );
not ( n65726 , n65725 );
or ( n65727 , n65724 , n65726 );
not ( n65728 , n58982 );
nand ( n65729 , n65728 , n55203 );
nand ( n65730 , n65727 , n65729 );
nand ( n65731 , n65730 , n52723 );
nand ( n65732 , n65723 , n65731 );
not ( n65733 , n56639 );
not ( n65734 , n59345 );
not ( n65735 , n40148 );
or ( n65736 , n65734 , n65735 );
nand ( n65737 , n56010 , n60617 );
nand ( n65738 , n65736 , n65737 );
not ( n65739 , n65738 );
or ( n65740 , n65733 , n65739 );
and ( n65741 , n40363 , n59345 );
not ( n65742 , n40363 );
not ( n65743 , n59345 );
and ( n65744 , n65742 , n65743 );
nor ( n65745 , n65741 , n65744 );
nand ( n65746 , n65745 , n59950 );
nand ( n65747 , n65740 , n65746 );
xor ( n65748 , n65732 , n65747 );
not ( n65749 , n60927 );
not ( n65750 , n49112 );
not ( n65751 , n40225 );
or ( n65752 , n65750 , n65751 );
nand ( n65753 , n59601 , n60292 );
nand ( n65754 , n65752 , n65753 );
not ( n65755 , n65754 );
or ( n65756 , n65749 , n65755 );
nand ( n65757 , n65281 , n58168 );
nand ( n65758 , n65756 , n65757 );
xor ( n65759 , n65748 , n65758 );
not ( n65760 , n48894 );
not ( n65761 , n65242 );
or ( n65762 , n65760 , n65761 );
not ( n65763 , n52377 );
not ( n65764 , n57798 );
or ( n65765 , n65763 , n65764 );
nand ( n65766 , n57801 , n53973 );
nand ( n65767 , n65765 , n65766 );
nand ( n65768 , n52004 , n65767 );
nand ( n65769 , n65762 , n65768 );
not ( n65770 , n52151 );
not ( n65771 , n65205 );
or ( n65772 , n65770 , n65771 );
not ( n65773 , n50916 );
not ( n65774 , n65773 );
not ( n65775 , n52222 );
or ( n65776 , n65774 , n65775 );
nand ( n65777 , n52223 , n52781 );
nand ( n65778 , n65776 , n65777 );
nand ( n65779 , n65778 , n51223 );
nand ( n65780 , n65772 , n65779 );
xor ( n65781 , n65769 , n65780 );
not ( n65782 , n54623 );
not ( n65783 , n51680 );
not ( n65784 , n56020 );
or ( n65785 , n65783 , n65784 );
nand ( n65786 , n56976 , n51684 );
nand ( n65787 , n65785 , n65786 );
not ( n65788 , n65787 );
or ( n65789 , n65782 , n65788 );
nand ( n65790 , n65250 , n52022 );
nand ( n65791 , n65789 , n65790 );
xor ( n65792 , n65781 , n65791 );
xor ( n65793 , n65759 , n65792 );
not ( n65794 , n65098 );
not ( n65795 , n63411 );
not ( n65796 , n65795 );
or ( n65797 , n65794 , n65796 );
and ( n65798 , n47047 , n63412 );
not ( n65799 , n47047 );
and ( n65800 , n65799 , n63416 );
or ( n65801 , n65798 , n65800 );
nand ( n65802 , n65092 , n65801 );
nand ( n65803 , n65797 , n65802 );
not ( n65804 , n65108 );
not ( n65805 , n56355 );
or ( n65806 , n65804 , n65805 );
not ( n65807 , n53927 );
not ( n65808 , n65103 );
not ( n65809 , n52285 );
or ( n65810 , n65808 , n65809 );
nand ( n65811 , n40677 , n53928 );
nand ( n65812 , n65810 , n65811 );
nand ( n65813 , n65807 , n65812 );
nand ( n65814 , n65806 , n65813 );
xor ( n65815 , n65803 , n65814 );
xor ( n65816 , n65815 , n65221 );
xor ( n65817 , n65793 , n65816 );
xor ( n65818 , n65759 , n65792 );
and ( n65819 , n65818 , n65816 );
and ( n65820 , n65759 , n65792 );
or ( n65821 , n65819 , n65820 );
not ( n65822 , n49026 );
not ( n65823 , n46425 );
not ( n65824 , n63793 );
not ( n65825 , n65824 );
or ( n65826 , n65823 , n65825 );
nand ( n65827 , n46422 , n42651 );
nand ( n65828 , n65826 , n65827 );
not ( n65829 , n65828 );
or ( n65830 , n65822 , n65829 );
nand ( n65831 , n65320 , n46267 );
nand ( n65832 , n65830 , n65831 );
xor ( n65833 , n65832 , n64968 );
xor ( n65834 , n65833 , n65002 );
xor ( n65835 , n65834 , n65159 );
xor ( n65836 , n65835 , n65552 );
xor ( n65837 , n65834 , n65159 );
and ( n65838 , n65837 , n65552 );
and ( n65839 , n65834 , n65159 );
or ( n65840 , n65838 , n65839 );
xor ( n65841 , n65076 , n65515 );
xor ( n65842 , n65841 , n65568 );
xor ( n65843 , n65076 , n65515 );
and ( n65844 , n65843 , n65568 );
and ( n65845 , n65076 , n65515 );
or ( n65846 , n65844 , n65845 );
xor ( n65847 , n65582 , n65592 );
and ( n65848 , n65847 , n65600 );
and ( n65849 , n65582 , n65592 );
or ( n65850 , n65848 , n65849 );
xor ( n65851 , n65632 , n65198 );
xor ( n65852 , n65851 , n65671 );
xor ( n65853 , n65632 , n65198 );
and ( n65854 , n65853 , n65671 );
and ( n65855 , n65632 , n65198 );
or ( n65856 , n65854 , n65855 );
xor ( n65857 , n65234 , n65228 );
xor ( n65858 , n65857 , n65330 );
xor ( n65859 , n65234 , n65228 );
and ( n65860 , n65859 , n65330 );
and ( n65861 , n65234 , n65228 );
or ( n65862 , n65860 , n65861 );
xor ( n65863 , n65677 , n65716 );
xor ( n65864 , n65863 , n65347 );
xor ( n65865 , n65677 , n65716 );
and ( n65866 , n65865 , n65347 );
and ( n65867 , n65677 , n65716 );
or ( n65868 , n65866 , n65867 );
xor ( n65869 , n65817 , n65301 );
xor ( n65870 , n65869 , n65836 );
xor ( n65871 , n65817 , n65301 );
and ( n65872 , n65871 , n65836 );
and ( n65873 , n65817 , n65301 );
or ( n65874 , n65872 , n65873 );
xor ( n65875 , n65842 , n65363 );
xor ( n65876 , n65875 , n65357 );
xor ( n65877 , n65842 , n65363 );
and ( n65878 , n65877 , n65357 );
and ( n65879 , n65842 , n65363 );
or ( n65880 , n65878 , n65879 );
xor ( n65881 , n65852 , n65369 );
xor ( n65882 , n65881 , n65858 );
xor ( n65883 , n65852 , n65369 );
and ( n65884 , n65883 , n65858 );
and ( n65885 , n65852 , n65369 );
or ( n65886 , n65884 , n65885 );
xor ( n65887 , n65375 , n65864 );
xor ( n65888 , n65887 , n65870 );
xor ( n65889 , n65375 , n65864 );
and ( n65890 , n65889 , n65870 );
and ( n65891 , n65375 , n65864 );
or ( n65892 , n65890 , n65891 );
xor ( n65893 , n65381 , n65387 );
xor ( n65894 , n65893 , n65876 );
xor ( n65895 , n65381 , n65387 );
and ( n65896 , n65895 , n65876 );
and ( n65897 , n65381 , n65387 );
or ( n65898 , n65896 , n65897 );
xor ( n65899 , n65393 , n65882 );
xor ( n65900 , n65899 , n65888 );
xor ( n65901 , n65393 , n65882 );
and ( n65902 , n65901 , n65888 );
and ( n65903 , n65393 , n65882 );
or ( n65904 , n65902 , n65903 );
xor ( n65905 , n65399 , n65894 );
xor ( n65906 , n65905 , n65900 );
xor ( n65907 , n65399 , n65894 );
and ( n65908 , n65907 , n65900 );
and ( n65909 , n65399 , n65894 );
or ( n65910 , n65908 , n65909 );
xor ( n65911 , n65643 , n65656 );
and ( n65912 , n65911 , n65668 );
and ( n65913 , n65643 , n65656 );
or ( n65914 , n65912 , n65913 );
xor ( n65915 , n65405 , n65906 );
xor ( n65916 , n65915 , n65411 );
xor ( n65917 , n65405 , n65906 );
and ( n65918 , n65917 , n65411 );
and ( n65919 , n65405 , n65906 );
or ( n65920 , n65918 , n65919 );
xor ( n65921 , n65609 , n65619 );
and ( n65922 , n65921 , n65630 );
and ( n65923 , n65609 , n65619 );
or ( n65924 , n65922 , n65923 );
xor ( n65925 , n65803 , n65814 );
and ( n65926 , n65925 , n65221 );
and ( n65927 , n65803 , n65814 );
or ( n65928 , n65926 , n65927 );
xor ( n65929 , n65769 , n65780 );
and ( n65930 , n65929 , n65791 );
and ( n65931 , n65769 , n65780 );
or ( n65932 , n65930 , n65931 );
xor ( n65933 , n65732 , n65747 );
and ( n65934 , n65933 , n65758 );
and ( n65935 , n65732 , n65747 );
or ( n65936 , n65934 , n65935 );
xor ( n65937 , n65692 , n65702 );
and ( n65938 , n65937 , n65714 );
and ( n65939 , n65692 , n65702 );
or ( n65940 , n65938 , n65939 );
xor ( n65941 , n65832 , n64968 );
and ( n65942 , n65941 , n65002 );
and ( n65943 , n65832 , n64968 );
or ( n65944 , n65942 , n65943 );
not ( n65945 , n65480 );
not ( n65946 , n53609 );
or ( n65947 , n65945 , n65946 );
not ( n65948 , n64942 );
not ( n65949 , n55917 );
or ( n65950 , n65948 , n65949 );
nand ( n65951 , n53590 , n50004 );
nand ( n65952 , n65950 , n65951 );
nand ( n65953 , n65952 , n53326 );
nand ( n65954 , n65947 , n65953 );
not ( n65955 , n65495 );
not ( n65956 , n54315 );
or ( n65957 , n65955 , n65956 );
not ( n65958 , n49001 );
not ( n65959 , n64970 );
or ( n65960 , n65958 , n65959 );
nand ( n65961 , n56274 , n48997 );
nand ( n65962 , n65960 , n65961 );
nand ( n65963 , n55867 , n65962 );
nand ( n65964 , n65957 , n65963 );
xor ( n65965 , n65954 , n65964 );
not ( n65966 , n65580 );
not ( n65967 , n55576 );
or ( n65968 , n65966 , n65967 );
not ( n65969 , n50631 );
not ( n65970 , n65969 );
not ( n65971 , n55148 );
or ( n65972 , n65970 , n65971 );
nand ( n65973 , n55152 , n50084 );
nand ( n65974 , n65972 , n65973 );
nand ( n65975 , n65974 , n54848 );
nand ( n65976 , n65968 , n65975 );
xor ( n65977 , n65965 , n65976 );
xor ( n65978 , n65954 , n65964 );
and ( n65979 , n65978 , n65976 );
and ( n65980 , n65954 , n65964 );
or ( n65981 , n65979 , n65980 );
not ( n65982 , n58915 );
not ( n65983 , n55893 );
or ( n65984 , n65982 , n65983 );
nand ( n65985 , n55892 , n58914 );
nand ( n65986 , n65984 , n65985 );
not ( n65987 , n65986 );
not ( n65988 , n55459 );
or ( n65989 , n65987 , n65988 );
nand ( n65990 , n65590 , n56281 );
nand ( n65991 , n65989 , n65990 );
not ( n65992 , n65598 );
not ( n65993 , n65992 );
not ( n65994 , n56776 );
or ( n65995 , n65993 , n65994 );
not ( n65996 , n58994 );
not ( n65997 , n56759 );
or ( n65998 , n65996 , n65997 );
buf ( n65999 , n57664 );
nand ( n66000 , n65999 , n58179 );
nand ( n66001 , n65998 , n66000 );
nand ( n66002 , n56780 , n66001 );
nand ( n66003 , n65995 , n66002 );
xor ( n66004 , n65991 , n66003 );
buf ( n66005 , n59432 );
not ( n66006 , n66005 );
or ( n66007 , n66006 , n65641 );
and ( n66008 , n57615 , n57182 );
and ( n66009 , n57619 , n47332 );
nor ( n66010 , n66008 , n66009 );
or ( n66011 , n65638 , n66010 );
nand ( n66012 , n66007 , n66011 );
xor ( n66013 , n66004 , n66012 );
xor ( n66014 , n65991 , n66003 );
and ( n66015 , n66014 , n66012 );
and ( n66016 , n65991 , n66003 );
or ( n66017 , n66015 , n66016 );
not ( n66018 , n51865 );
not ( n66019 , n49707 );
not ( n66020 , n59891 );
or ( n66021 , n66019 , n66020 );
nand ( n66022 , n63152 , n52273 );
nand ( n66023 , n66021 , n66022 );
not ( n66024 , n66023 );
or ( n66025 , n66018 , n66024 );
nand ( n66026 , n65536 , n49713 );
nand ( n66027 , n66025 , n66026 );
xor ( n66028 , n65924 , n66027 );
not ( n66029 , n65828 );
not ( n66030 , n46267 );
or ( n66031 , n66029 , n66030 );
nand ( n66032 , n49026 , n46425 );
nand ( n66033 , n66031 , n66032 );
xor ( n66034 , n66028 , n66033 );
xor ( n66035 , n65924 , n66027 );
and ( n66036 , n66035 , n66033 );
and ( n66037 , n65924 , n66027 );
or ( n66038 , n66036 , n66037 );
not ( n66039 , n52970 );
not ( n66040 , n65562 );
or ( n66041 , n66039 , n66040 );
and ( n66042 , n60906 , n48645 );
not ( n66043 , n60906 );
and ( n66044 , n66043 , n52048 );
or ( n66045 , n66042 , n66044 );
nand ( n66046 , n66045 , n52962 );
nand ( n66047 , n66041 , n66046 );
not ( n66048 , n53675 );
not ( n66049 , n54028 );
not ( n66050 , n62909 );
or ( n66051 , n66049 , n66050 );
not ( n66052 , n62912 );
not ( n66053 , n66052 );
nand ( n66054 , n66053 , n50634 );
nand ( n66055 , n66051 , n66054 );
not ( n66056 , n66055 );
or ( n66057 , n66048 , n66056 );
nand ( n66058 , n65509 , n47407 );
nand ( n66059 , n66057 , n66058 );
xor ( n66060 , n66047 , n66059 );
not ( n66061 , n52421 );
not ( n66062 , n65710 );
or ( n66063 , n66061 , n66062 );
not ( n66064 , n51723 );
not ( n66065 , n59914 );
or ( n66066 , n66064 , n66065 );
nand ( n66067 , n59913 , n51724 );
nand ( n66068 , n66066 , n66067 );
nand ( n66069 , n66068 , n50767 );
nand ( n66070 , n66063 , n66069 );
xor ( n66071 , n66060 , n66070 );
xor ( n66072 , n66047 , n66059 );
and ( n66073 , n66072 , n66070 );
and ( n66074 , n66047 , n66059 );
or ( n66075 , n66073 , n66074 );
xor ( n66076 , n65977 , n66013 );
not ( n66077 , n65617 );
not ( n66078 , n61548 );
or ( n66079 , n66077 , n66078 );
not ( n66080 , n51204 );
not ( n66081 , n61537 );
or ( n66082 , n66080 , n66081 );
nand ( n66083 , n63541 , n48860 );
nand ( n66084 , n66082 , n66083 );
nand ( n66085 , n66084 , n61557 );
nand ( n66086 , n66079 , n66085 );
not ( n66087 , n65628 );
or ( n66088 , n64684 , n66087 );
not ( n66089 , n62449 );
and ( n66090 , n48898 , n66089 );
not ( n66091 , n48898 );
and ( n66092 , n66091 , n62451 );
nor ( n66093 , n66090 , n66092 );
or ( n66094 , n64166 , n66093 );
nand ( n66095 , n66088 , n66094 );
xor ( n66096 , n66086 , n66095 );
not ( n66097 , n65801 );
not ( n66098 , n65089 );
or ( n66099 , n66097 , n66098 );
not ( n66100 , n47227 );
not ( n66101 , n64443 );
or ( n66102 , n66100 , n66101 );
nand ( n66103 , n63416 , n47589 );
nand ( n66104 , n66102 , n66103 );
nand ( n66105 , n65092 , n66104 );
nand ( n66106 , n66099 , n66105 );
xor ( n66107 , n66096 , n66106 );
xor ( n66108 , n66076 , n66107 );
xor ( n66109 , n65977 , n66013 );
and ( n66110 , n66109 , n66107 );
and ( n66111 , n65977 , n66013 );
or ( n66112 , n66110 , n66111 );
not ( n66113 , n65654 );
not ( n66114 , n61961 );
or ( n66115 , n66113 , n66114 );
not ( n66116 , n48983 );
not ( n66117 , n65183 );
or ( n66118 , n66116 , n66117 );
nand ( n66119 , n65652 , n56348 );
nand ( n66120 , n66118 , n66119 );
nand ( n66121 , n61465 , n66120 );
nand ( n66122 , n66115 , n66121 );
not ( n66123 , n65666 );
not ( n66124 , n59571 );
or ( n66125 , n66123 , n66124 );
not ( n66126 , n55511 );
not ( n66127 , n59340 );
or ( n66128 , n66126 , n66127 );
nand ( n66129 , n59935 , n51670 );
nand ( n66130 , n66128 , n66129 );
nand ( n66131 , n59575 , n66130 );
nand ( n66132 , n66125 , n66131 );
xor ( n66133 , n66122 , n66132 );
not ( n66134 , n65606 );
not ( n66135 , n66134 );
not ( n66136 , n60960 );
not ( n66137 , n66136 );
or ( n66138 , n66135 , n66137 );
not ( n66139 , n51792 );
buf ( n66140 , n60285 );
not ( n66141 , n66140 );
not ( n66142 , n66141 );
or ( n66143 , n66139 , n66142 );
nand ( n66144 , n66140 , n48829 );
nand ( n66145 , n66143 , n66144 );
nand ( n66146 , n60427 , n66145 );
nand ( n66147 , n66138 , n66146 );
xor ( n66148 , n66133 , n66147 );
xor ( n66149 , n66148 , n65928 );
xor ( n66150 , n66149 , n65932 );
xor ( n66151 , n66148 , n65928 );
and ( n66152 , n66151 , n65932 );
and ( n66153 , n66148 , n65928 );
or ( n66154 , n66152 , n66153 );
not ( n66155 , n63415 );
and ( n66156 , n66155 , n47646 );
not ( n66157 , n51766 );
and ( n66158 , n40691 , n52110 );
not ( n66159 , n40691 );
and ( n66160 , n66159 , n53918 );
or ( n66161 , n66158 , n66160 );
not ( n66162 , n66161 );
or ( n66163 , n66157 , n66162 );
nand ( n66164 , n52482 , n65453 );
nand ( n66165 , n66163 , n66164 );
xor ( n66166 , n66156 , n66165 );
not ( n66167 , n51533 );
not ( n66168 , n65103 );
not ( n66169 , n51928 );
or ( n66170 , n66168 , n66169 );
nand ( n66171 , n51280 , n51508 );
nand ( n66172 , n66170 , n66171 );
not ( n66173 , n66172 );
or ( n66174 , n66167 , n66173 );
nand ( n66175 , n65812 , n56355 );
nand ( n66176 , n66174 , n66175 );
xor ( n66177 , n66166 , n66176 );
xor ( n66178 , n65936 , n66177 );
xor ( n66179 , n66178 , n65519 );
xor ( n66180 , n65936 , n66177 );
and ( n66181 , n66180 , n65519 );
and ( n66182 , n65936 , n66177 );
or ( n66183 , n66181 , n66182 );
xor ( n66184 , n65940 , n65944 );
xor ( n66185 , n66184 , n65556 );
xor ( n66186 , n65940 , n65944 );
and ( n66187 , n66186 , n65556 );
and ( n66188 , n65940 , n65944 );
or ( n66189 , n66187 , n66188 );
not ( n66190 , n52757 );
not ( n66191 , n50306 );
not ( n66192 , n40627 );
or ( n66193 , n66191 , n66192 );
nand ( n66194 , n50943 , n40626 );
nand ( n66195 , n66193 , n66194 );
not ( n66196 , n66195 );
or ( n66197 , n66190 , n66196 );
nand ( n66198 , n65698 , n63708 );
nand ( n66199 , n66197 , n66198 );
not ( n66200 , n52526 );
not ( n66201 , n65778 );
or ( n66202 , n66200 , n66201 );
not ( n66203 , n50895 );
not ( n66204 , n52570 );
or ( n66205 , n66203 , n66204 );
nand ( n66206 , n40526 , n51462 );
nand ( n66207 , n66205 , n66206 );
nand ( n66208 , n66207 , n51223 );
nand ( n66209 , n66202 , n66208 );
xor ( n66210 , n66199 , n66209 );
not ( n66211 , n52004 );
not ( n66212 , n52377 );
not ( n66213 , n39846 );
or ( n66214 , n66212 , n66213 );
not ( n66215 , n39844 );
nand ( n66216 , n66215 , n55013 );
nand ( n66217 , n66214 , n66216 );
not ( n66218 , n66217 );
or ( n66219 , n66211 , n66218 );
nand ( n66220 , n65767 , n48894 );
nand ( n66221 , n66219 , n66220 );
xor ( n66222 , n66210 , n66221 );
not ( n66223 , n56861 );
and ( n66224 , n54283 , n50020 );
not ( n66225 , n54283 );
not ( n66226 , n50020 );
and ( n66227 , n66225 , n66226 );
nor ( n66228 , n66224 , n66227 );
not ( n66229 , n66228 );
and ( n66230 , n66223 , n66229 );
not ( n66231 , n65466 );
nor ( n66232 , n66231 , n56853 );
nor ( n66233 , n66230 , n66232 );
buf ( n66234 , n49112 );
not ( n66235 , n66234 );
buf ( n66236 , n59194 );
not ( n66237 , n66236 );
or ( n66238 , n66235 , n66237 );
nand ( n66239 , n59195 , n60292 );
nand ( n66240 , n66238 , n66239 );
not ( n66241 , n66240 );
not ( n66242 , n52191 );
or ( n66243 , n66241 , n66242 );
nand ( n66244 , n65754 , n58168 );
nand ( n66245 , n66243 , n66244 );
xor ( n66246 , n66233 , n66245 );
not ( n66247 , n62664 );
not ( n66248 , n65690 );
or ( n66249 , n66247 , n66248 );
not ( n66250 , n61951 );
not ( n66251 , n56476 );
or ( n66252 , n66250 , n66251 );
nand ( n66253 , n53290 , n61952 );
nand ( n66254 , n66252 , n66253 );
nand ( n66255 , n66254 , n62654 );
nand ( n66256 , n66249 , n66255 );
xor ( n66257 , n66246 , n66256 );
xor ( n66258 , n66222 , n66257 );
not ( n66259 , n47873 );
not ( n66260 , n65787 );
or ( n66261 , n66259 , n66260 );
not ( n66262 , n51680 );
not ( n66263 , n56451 );
or ( n66264 , n66262 , n66263 );
nand ( n66265 , n51684 , n40012 );
nand ( n66266 , n66264 , n66265 );
nand ( n66267 , n66266 , n54623 );
nand ( n66268 , n66261 , n66267 );
not ( n66269 , n52723 );
not ( n66270 , n60602 );
not ( n66271 , n56411 );
or ( n66272 , n66270 , n66271 );
nand ( n66273 , n40452 , n62577 );
nand ( n66274 , n66272 , n66273 );
not ( n66275 , n66274 );
or ( n66276 , n66269 , n66275 );
nand ( n66277 , n65730 , n59633 );
nand ( n66278 , n66276 , n66277 );
xor ( n66279 , n66268 , n66278 );
not ( n66280 , n56639 );
not ( n66281 , n59345 );
not ( n66282 , n55641 );
or ( n66283 , n66281 , n66282 );
nand ( n66284 , n55645 , n60617 );
nand ( n66285 , n66283 , n66284 );
not ( n66286 , n66285 );
or ( n66287 , n66280 , n66286 );
nand ( n66288 , n65738 , n59950 );
nand ( n66289 , n66287 , n66288 );
xor ( n66290 , n66279 , n66289 );
xor ( n66291 , n66258 , n66290 );
xor ( n66292 , n66222 , n66257 );
and ( n66293 , n66292 , n66290 );
and ( n66294 , n66222 , n66257 );
or ( n66295 , n66293 , n66294 );
xor ( n66296 , n65636 , n65572 );
not ( n66297 , n51157 );
not ( n66298 , n65548 );
or ( n66299 , n66297 , n66298 );
not ( n66300 , n50263 );
not ( n66301 , n42554 );
not ( n66302 , n66301 );
or ( n66303 , n66300 , n66302 );
not ( n66304 , n63246 );
nand ( n66305 , n66304 , n52080 );
nand ( n66306 , n66303 , n66305 );
nand ( n66307 , n66306 , n48073 );
nand ( n66308 , n66299 , n66307 );
xor ( n66309 , n65473 , n66308 );
xor ( n66310 , n66309 , n65503 );
xor ( n66311 , n66296 , n66310 );
xor ( n66312 , n65636 , n65572 );
and ( n66313 , n66312 , n66310 );
and ( n66314 , n65636 , n65572 );
or ( n66315 , n66313 , n66314 );
not ( n66316 , n48989 );
not ( n66317 , n65525 );
or ( n66318 , n66316 , n66317 );
not ( n66319 , n49500 );
not ( n66320 , n60855 );
or ( n66321 , n66319 , n66320 );
nand ( n66322 , n62963 , n47979 );
nand ( n66323 , n66321 , n66322 );
nand ( n66324 , n66323 , n53510 );
nand ( n66325 , n66318 , n66324 );
xor ( n66326 , n65850 , n66325 );
xor ( n66327 , n66326 , n65914 );
xor ( n66328 , n66327 , n66071 );
xor ( n66329 , n66328 , n66034 );
xor ( n66330 , n66327 , n66071 );
and ( n66331 , n66330 , n66034 );
and ( n66332 , n66327 , n66071 );
or ( n66333 , n66331 , n66332 );
xor ( n66334 , n65675 , n66108 );
xor ( n66335 , n66334 , n66179 );
xor ( n66336 , n65675 , n66108 );
and ( n66337 , n66336 , n66179 );
and ( n66338 , n65675 , n66108 );
or ( n66339 , n66337 , n66338 );
xor ( n66340 , n66122 , n66132 );
and ( n66341 , n66340 , n66147 );
and ( n66342 , n66122 , n66132 );
or ( n66343 , n66341 , n66342 );
xor ( n66344 , n65821 , n66150 );
xor ( n66345 , n66344 , n65681 );
xor ( n66346 , n65821 , n66150 );
and ( n66347 , n66346 , n65681 );
and ( n66348 , n65821 , n66150 );
or ( n66349 , n66347 , n66348 );
xor ( n66350 , n65720 , n65840 );
xor ( n66351 , n66350 , n66185 );
xor ( n66352 , n65720 , n65840 );
and ( n66353 , n66352 , n66185 );
and ( n66354 , n65720 , n65840 );
or ( n66355 , n66353 , n66354 );
xor ( n66356 , n66291 , n65846 );
xor ( n66357 , n66356 , n66329 );
xor ( n66358 , n66291 , n65846 );
and ( n66359 , n66358 , n66329 );
and ( n66360 , n66291 , n65846 );
or ( n66361 , n66359 , n66360 );
xor ( n66362 , n66311 , n65856 );
xor ( n66363 , n66362 , n66335 );
xor ( n66364 , n66311 , n65856 );
and ( n66365 , n66364 , n66335 );
and ( n66366 , n66311 , n65856 );
or ( n66367 , n66365 , n66366 );
xor ( n66368 , n65868 , n65862 );
xor ( n66369 , n66368 , n66345 );
xor ( n66370 , n65868 , n65862 );
and ( n66371 , n66370 , n66345 );
and ( n66372 , n65868 , n65862 );
or ( n66373 , n66371 , n66372 );
xor ( n66374 , n66351 , n65874 );
xor ( n66375 , n66374 , n66357 );
xor ( n66376 , n66351 , n65874 );
and ( n66377 , n66376 , n66357 );
and ( n66378 , n66351 , n65874 );
or ( n66379 , n66377 , n66378 );
xor ( n66380 , n65880 , n66363 );
xor ( n66381 , n66380 , n65886 );
xor ( n66382 , n65880 , n66363 );
and ( n66383 , n66382 , n65886 );
and ( n66384 , n65880 , n66363 );
or ( n66385 , n66383 , n66384 );
xor ( n66386 , n66369 , n65892 );
xor ( n66387 , n66386 , n66375 );
xor ( n66388 , n66369 , n65892 );
and ( n66389 , n66388 , n66375 );
and ( n66390 , n66369 , n65892 );
or ( n66391 , n66389 , n66390 );
xor ( n66392 , n65898 , n66381 );
xor ( n66393 , n66392 , n65904 );
xor ( n66394 , n65898 , n66381 );
and ( n66395 , n66394 , n65904 );
and ( n66396 , n65898 , n66381 );
or ( n66397 , n66395 , n66396 );
xor ( n66398 , n66387 , n66393 );
xor ( n66399 , n66398 , n65910 );
xor ( n66400 , n66387 , n66393 );
and ( n66401 , n66400 , n65910 );
and ( n66402 , n66387 , n66393 );
or ( n66403 , n66401 , n66402 );
xor ( n66404 , n66086 , n66095 );
and ( n66405 , n66404 , n66106 );
and ( n66406 , n66086 , n66095 );
or ( n66407 , n66405 , n66406 );
xor ( n66408 , n66156 , n66165 );
and ( n66409 , n66408 , n66176 );
and ( n66410 , n66156 , n66165 );
or ( n66411 , n66409 , n66410 );
xor ( n66412 , n66268 , n66278 );
and ( n66413 , n66412 , n66289 );
and ( n66414 , n66268 , n66278 );
or ( n66415 , n66413 , n66414 );
xor ( n66416 , n66233 , n66245 );
and ( n66417 , n66416 , n66256 );
and ( n66418 , n66233 , n66245 );
or ( n66419 , n66417 , n66418 );
xor ( n66420 , n66199 , n66209 );
and ( n66421 , n66420 , n66221 );
and ( n66422 , n66199 , n66209 );
or ( n66423 , n66421 , n66422 );
xor ( n66424 , n65473 , n66308 );
and ( n66425 , n66424 , n65503 );
and ( n66426 , n65473 , n66308 );
or ( n66427 , n66425 , n66426 );
xor ( n66428 , n65850 , n66325 );
and ( n66429 , n66428 , n65914 );
and ( n66430 , n65850 , n66325 );
or ( n66431 , n66429 , n66430 );
or ( n66432 , n46267 , n46188 );
nand ( n66433 , n66432 , n46425 );
not ( n66434 , n66228 );
not ( n66435 , n66434 );
not ( n66436 , n52854 );
or ( n66437 , n66435 , n66436 );
not ( n66438 , n52841 );
not ( n66439 , n53513 );
or ( n66440 , n66438 , n66439 );
nand ( n66441 , n55104 , n52079 );
nand ( n66442 , n66440 , n66441 );
nand ( n66443 , n66442 , n52469 );
nand ( n66444 , n66437 , n66443 );
xor ( n66445 , n66433 , n66444 );
not ( n66446 , n65952 );
not ( n66447 , n53956 );
or ( n66448 , n66446 , n66447 );
not ( n66449 , n64451 );
not ( n66450 , n53615 );
or ( n66451 , n66449 , n66450 );
nand ( n66452 , n64452 , n53595 );
nand ( n66453 , n66451 , n66452 );
nand ( n66454 , n66453 , n54364 );
nand ( n66455 , n66448 , n66454 );
xor ( n66456 , n66445 , n66455 );
xor ( n66457 , n66433 , n66444 );
and ( n66458 , n66457 , n66455 );
and ( n66459 , n66433 , n66444 );
or ( n66460 , n66458 , n66459 );
not ( n66461 , n54077 );
not ( n66462 , n49209 );
not ( n66463 , n54467 );
or ( n66464 , n66462 , n66463 );
nand ( n66465 , n54298 , n49837 );
nand ( n66466 , n66464 , n66465 );
not ( n66467 , n66466 );
or ( n66468 , n66461 , n66467 );
nand ( n66469 , n65962 , n56810 );
nand ( n66470 , n66468 , n66469 );
not ( n66471 , n55934 );
not ( n66472 , n52272 );
not ( n66473 , n55125 );
or ( n66474 , n66472 , n66473 );
nand ( n66475 , n55152 , n49820 );
nand ( n66476 , n66474 , n66475 );
not ( n66477 , n66476 );
or ( n66478 , n66471 , n66477 );
nand ( n66479 , n55576 , n65974 );
nand ( n66480 , n66478 , n66479 );
xor ( n66481 , n66470 , n66480 );
not ( n66482 , n65986 );
not ( n66483 , n55887 );
or ( n66484 , n66482 , n66483 );
and ( n66485 , n41532 , n55846 );
not ( n66486 , n41532 );
and ( n66487 , n66486 , n55872 );
or ( n66488 , n66485 , n66487 );
nand ( n66489 , n66488 , n55458 );
nand ( n66490 , n66484 , n66489 );
xor ( n66491 , n66481 , n66490 );
xor ( n66492 , n66470 , n66480 );
and ( n66493 , n66492 , n66490 );
and ( n66494 , n66470 , n66480 );
or ( n66495 , n66493 , n66494 );
not ( n66496 , n48989 );
not ( n66497 , n66323 );
or ( n66498 , n66496 , n66497 );
not ( n66499 , n49500 );
not ( n66500 , n39253 );
not ( n66501 , n66500 );
or ( n66502 , n66499 , n66501 );
nand ( n66503 , n39253 , n47979 );
nand ( n66504 , n66502 , n66503 );
nand ( n66505 , n66504 , n47384 );
nand ( n66506 , n66498 , n66505 );
xor ( n66507 , n66506 , n66407 );
not ( n66508 , n49713 );
not ( n66509 , n66023 );
or ( n66510 , n66508 , n66509 );
not ( n66511 , n52267 );
not ( n66512 , n62394 );
or ( n66513 , n66511 , n66512 );
nand ( n66514 , n38499 , n51351 );
nand ( n66515 , n66513 , n66514 );
nand ( n66516 , n66515 , n51865 );
nand ( n66517 , n66510 , n66516 );
xor ( n66518 , n66507 , n66517 );
xor ( n66519 , n66506 , n66407 );
and ( n66520 , n66519 , n66517 );
and ( n66521 , n66506 , n66407 );
or ( n66522 , n66520 , n66521 );
not ( n66523 , n52962 );
and ( n66524 , n48645 , n59402 );
not ( n66525 , n48645 );
and ( n66526 , n66525 , n39574 );
or ( n66527 , n66524 , n66526 );
not ( n66528 , n66527 );
or ( n66529 , n66523 , n66528 );
nand ( n66530 , n66045 , n52970 );
nand ( n66531 , n66529 , n66530 );
not ( n66532 , n53675 );
not ( n66533 , n54028 );
not ( n66534 , n42399 );
or ( n66535 , n66533 , n66534 );
not ( n66536 , n42399 );
nand ( n66537 , n66536 , n50634 );
nand ( n66538 , n66535 , n66537 );
not ( n66539 , n66538 );
or ( n66540 , n66532 , n66539 );
nand ( n66541 , n66055 , n64498 );
nand ( n66542 , n66540 , n66541 );
xor ( n66543 , n66531 , n66542 );
not ( n66544 , n54875 );
not ( n66545 , n51723 );
buf ( n66546 , n39680 );
not ( n66547 , n66546 );
not ( n66548 , n66547 );
or ( n66549 , n66545 , n66548 );
nand ( n66550 , n58485 , n51724 );
nand ( n66551 , n66549 , n66550 );
not ( n66552 , n66551 );
or ( n66553 , n66544 , n66552 );
nand ( n66554 , n66068 , n52421 );
nand ( n66555 , n66553 , n66554 );
xor ( n66556 , n66543 , n66555 );
xor ( n66557 , n66531 , n66542 );
and ( n66558 , n66557 , n66555 );
and ( n66559 , n66531 , n66542 );
or ( n66560 , n66558 , n66559 );
or ( n66561 , n64164 , n66093 );
and ( n66562 , n47765 , n62452 );
not ( n66563 , n47765 );
and ( n66564 , n66563 , n64170 );
nor ( n66565 , n66562 , n66564 );
or ( n66566 , n64166 , n66565 );
nand ( n66567 , n66561 , n66566 );
not ( n66568 , n66104 );
buf ( n66569 , n63410 );
not ( n66570 , n66569 );
or ( n66571 , n66568 , n66570 );
not ( n66572 , n49654 );
not ( n66573 , n65094 );
or ( n66574 , n66572 , n66573 );
not ( n66575 , n63412 );
nand ( n66576 , n66575 , n47368 );
nand ( n66577 , n66574 , n66576 );
nand ( n66578 , n66577 , n65092 );
nand ( n66579 , n66571 , n66578 );
xor ( n66580 , n66567 , n66579 );
buf ( n66581 , n66575 );
and ( n66582 , n66581 , n47047 );
xor ( n66583 , n66580 , n66582 );
xor ( n66584 , n66456 , n66583 );
xor ( n66585 , n66584 , n66491 );
xor ( n66586 , n66456 , n66583 );
and ( n66587 , n66586 , n66491 );
and ( n66588 , n66456 , n66583 );
or ( n66589 , n66587 , n66588 );
not ( n66590 , n66130 );
not ( n66591 , n59571 );
or ( n66592 , n66590 , n66591 );
and ( n66593 , n52712 , n59578 );
not ( n66594 , n52712 );
and ( n66595 , n66594 , n59338 );
nor ( n66596 , n66593 , n66595 );
nand ( n66597 , n66596 , n59931 );
nand ( n66598 , n66592 , n66597 );
not ( n66599 , n66145 );
not ( n66600 , n65130 );
or ( n66601 , n66599 , n66600 );
not ( n66602 , n60963 );
not ( n66603 , n52033 );
not ( n66604 , n66141 );
or ( n66605 , n66603 , n66604 );
nand ( n66606 , n66140 , n52038 );
nand ( n66607 , n66605 , n66606 );
nand ( n66608 , n66602 , n66607 );
nand ( n66609 , n66601 , n66608 );
xor ( n66610 , n66598 , n66609 );
not ( n66611 , n66084 );
not ( n66612 , n61550 );
or ( n66613 , n66611 , n66612 );
not ( n66614 , n49624 );
buf ( n66615 , n64633 );
not ( n66616 , n66615 );
not ( n66617 , n66616 );
or ( n66618 , n66614 , n66617 );
not ( n66619 , n61537 );
nand ( n66620 , n66619 , n49630 );
nand ( n66621 , n66618 , n66620 );
nand ( n66622 , n61558 , n66621 );
nand ( n66623 , n66613 , n66622 );
xor ( n66624 , n66610 , n66623 );
not ( n66625 , n66001 );
not ( n66626 , n56776 );
or ( n66627 , n66625 , n66626 );
not ( n66628 , n58458 );
not ( n66629 , n56785 );
or ( n66630 , n66628 , n66629 );
nand ( n66631 , n56786 , n58459 );
nand ( n66632 , n66630 , n66631 );
nand ( n66633 , n56780 , n66632 );
nand ( n66634 , n66627 , n66633 );
not ( n66635 , n66010 );
not ( n66636 , n66635 );
not ( n66637 , n66005 );
or ( n66638 , n66636 , n66637 );
not ( n66639 , n47527 );
not ( n66640 , n59437 );
or ( n66641 , n66639 , n66640 );
buf ( n66642 , n57634 );
nand ( n66643 , n66642 , n64603 );
nand ( n66644 , n66641 , n66643 );
nand ( n66645 , n59435 , n66644 );
nand ( n66646 , n66638 , n66645 );
xor ( n66647 , n66634 , n66646 );
not ( n66648 , n66120 );
not ( n66649 , n63080 );
or ( n66650 , n66648 , n66649 );
not ( n66651 , n56727 );
buf ( n66652 , n58966 );
not ( n66653 , n66652 );
or ( n66654 , n66651 , n66653 );
not ( n66655 , n62497 );
nand ( n66656 , n66655 , n56731 );
nand ( n66657 , n66654 , n66656 );
nand ( n66658 , n61465 , n66657 );
nand ( n66659 , n66650 , n66658 );
xor ( n66660 , n66647 , n66659 );
xor ( n66661 , n66624 , n66660 );
xor ( n66662 , n66661 , n66411 );
xor ( n66663 , n66624 , n66660 );
and ( n66664 , n66663 , n66411 );
and ( n66665 , n66624 , n66660 );
or ( n66666 , n66664 , n66665 );
xor ( n66667 , n66415 , n66419 );
xor ( n66668 , n66667 , n66038 );
xor ( n66669 , n66415 , n66419 );
and ( n66670 , n66669 , n66038 );
and ( n66671 , n66415 , n66419 );
or ( n66672 , n66670 , n66671 );
xor ( n66673 , n66423 , n66427 );
xor ( n66674 , n66673 , n66431 );
xor ( n66675 , n66423 , n66427 );
and ( n66676 , n66675 , n66431 );
and ( n66677 , n66423 , n66427 );
or ( n66678 , n66676 , n66677 );
not ( n66679 , n58168 );
not ( n66680 , n66240 );
or ( n66681 , n66679 , n66680 );
not ( n66682 , n62077 );
not ( n66683 , n40148 );
or ( n66684 , n66682 , n66683 );
nand ( n66685 , n54406 , n60292 );
nand ( n66686 , n66684 , n66685 );
nand ( n66687 , n66686 , n60927 );
nand ( n66688 , n66681 , n66687 );
not ( n66689 , n62654 );
buf ( n66690 , n52740 );
or ( n66691 , n66690 , n59601 );
nand ( n66692 , n53660 , n66690 );
nand ( n66693 , n66691 , n66692 );
not ( n66694 , n66693 );
or ( n66695 , n66689 , n66694 );
buf ( n66696 , n52058 );
nand ( n66697 , n66254 , n66696 );
nand ( n66698 , n66695 , n66697 );
xor ( n66699 , n66688 , n66698 );
not ( n66700 , n52757 );
not ( n66701 , n50306 );
not ( n66702 , n59611 );
or ( n66703 , n66701 , n66702 );
not ( n66704 , n63656 );
not ( n66705 , n50306 );
nand ( n66706 , n66704 , n66705 );
nand ( n66707 , n66703 , n66706 );
not ( n66708 , n66707 );
or ( n66709 , n66700 , n66708 );
nand ( n66710 , n66195 , n63708 );
nand ( n66711 , n66709 , n66710 );
xor ( n66712 , n66699 , n66711 );
xor ( n66713 , n66075 , n66712 );
not ( n66714 , n51766 );
not ( n66715 , n53918 );
not ( n66716 , n50958 );
or ( n66717 , n66715 , n66716 );
nand ( n66718 , n40677 , n52113 );
nand ( n66719 , n66717 , n66718 );
not ( n66720 , n66719 );
or ( n66721 , n66714 , n66720 );
nand ( n66722 , n66161 , n52482 );
nand ( n66723 , n66721 , n66722 );
not ( n66724 , n66233 );
xor ( n66725 , n66723 , n66724 );
not ( n66726 , n54623 );
not ( n66727 , n59174 );
not ( n66728 , n39963 );
or ( n66729 , n66727 , n66728 );
nand ( n66730 , n57801 , n54628 );
nand ( n66731 , n66729 , n66730 );
not ( n66732 , n66731 );
or ( n66733 , n66726 , n66732 );
not ( n66734 , n66266 );
not ( n66735 , n47873 );
or ( n66736 , n66734 , n66735 );
nand ( n66737 , n66733 , n66736 );
xor ( n66738 , n66725 , n66737 );
xor ( n66739 , n66713 , n66738 );
xor ( n66740 , n66075 , n66712 );
and ( n66741 , n66740 , n66738 );
and ( n66742 , n66075 , n66712 );
or ( n66743 , n66741 , n66742 );
not ( n66744 , n51533 );
and ( n66745 , n52222 , n65103 );
not ( n66746 , n52222 );
and ( n66747 , n66746 , n51508 );
or ( n66748 , n66745 , n66747 );
not ( n66749 , n66748 );
or ( n66750 , n66744 , n66749 );
nand ( n66751 , n52139 , n66172 );
nand ( n66752 , n66750 , n66751 );
not ( n66753 , n53104 );
not ( n66754 , n66274 );
or ( n66755 , n66753 , n66754 );
not ( n66756 , n60602 );
not ( n66757 , n40513 );
or ( n66758 , n66756 , n66757 );
nand ( n66759 , n40514 , n62577 );
nand ( n66760 , n66758 , n66759 );
nand ( n66761 , n66760 , n58977 );
nand ( n66762 , n66755 , n66761 );
xor ( n66763 , n66752 , n66762 );
not ( n66764 , n56639 );
not ( n66765 , n59345 );
not ( n66766 , n59694 );
or ( n66767 , n66765 , n66766 );
not ( n66768 , n56058 );
nand ( n66769 , n66768 , n60617 );
nand ( n66770 , n66767 , n66769 );
not ( n66771 , n66770 );
or ( n66772 , n66764 , n66771 );
nand ( n66773 , n66285 , n59950 );
nand ( n66774 , n66772 , n66773 );
xor ( n66775 , n66763 , n66774 );
xor ( n66776 , n66775 , n66112 );
xor ( n66777 , n66776 , n66556 );
xor ( n66778 , n66775 , n66112 );
and ( n66779 , n66778 , n66556 );
and ( n66780 , n66775 , n66112 );
or ( n66781 , n66779 , n66780 );
not ( n66782 , n53631 );
not ( n66783 , n50263 );
not ( n66784 , n42652 );
not ( n66785 , n66784 );
or ( n66786 , n66783 , n66785 );
nand ( n66787 , n63794 , n52080 );
nand ( n66788 , n66786 , n66787 );
not ( n66789 , n66788 );
or ( n66790 , n66782 , n66789 );
nand ( n66791 , n66306 , n51157 );
nand ( n66792 , n66790 , n66791 );
xor ( n66793 , n66792 , n66017 );
xor ( n66794 , n66793 , n66343 );
xor ( n66795 , n66518 , n66794 );
not ( n66796 , n51223 );
not ( n66797 , n50895 );
buf ( n66798 , n54377 );
not ( n66799 , n66798 );
or ( n66800 , n66797 , n66799 );
nand ( n66801 , n40592 , n52781 );
nand ( n66802 , n66800 , n66801 );
not ( n66803 , n66802 );
or ( n66804 , n66796 , n66803 );
nand ( n66805 , n66207 , n52151 );
nand ( n66806 , n66804 , n66805 );
not ( n66807 , n57314 );
not ( n66808 , n66217 );
or ( n66809 , n66807 , n66808 );
not ( n66810 , n52377 );
not ( n66811 , n39894 );
or ( n66812 , n66810 , n66811 );
nand ( n66813 , n65708 , n55013 );
nand ( n66814 , n66812 , n66813 );
nand ( n66815 , n66814 , n52004 );
nand ( n66816 , n66809 , n66815 );
xor ( n66817 , n66806 , n66816 );
xor ( n66818 , n66817 , n65981 );
xor ( n66819 , n66795 , n66818 );
xor ( n66820 , n66518 , n66794 );
and ( n66821 , n66820 , n66818 );
and ( n66822 , n66518 , n66794 );
or ( n66823 , n66821 , n66822 );
xor ( n66824 , n66662 , n66154 );
xor ( n66825 , n66824 , n66585 );
xor ( n66826 , n66662 , n66154 );
and ( n66827 , n66826 , n66585 );
and ( n66828 , n66662 , n66154 );
or ( n66829 , n66827 , n66828 );
xor ( n66830 , n66634 , n66646 );
and ( n66831 , n66830 , n66659 );
and ( n66832 , n66634 , n66646 );
or ( n66833 , n66831 , n66832 );
xor ( n66834 , n66668 , n66295 );
xor ( n66835 , n66834 , n66183 );
xor ( n66836 , n66668 , n66295 );
and ( n66837 , n66836 , n66183 );
and ( n66838 , n66668 , n66295 );
or ( n66839 , n66837 , n66838 );
xor ( n66840 , n66189 , n66674 );
xor ( n66841 , n66840 , n66333 );
xor ( n66842 , n66189 , n66674 );
and ( n66843 , n66842 , n66333 );
and ( n66844 , n66189 , n66674 );
or ( n66845 , n66843 , n66844 );
xor ( n66846 , n66315 , n66739 );
xor ( n66847 , n66846 , n66819 );
xor ( n66848 , n66315 , n66739 );
and ( n66849 , n66848 , n66819 );
and ( n66850 , n66315 , n66739 );
or ( n66851 , n66849 , n66850 );
xor ( n66852 , n66777 , n66339 );
xor ( n66853 , n66852 , n66349 );
xor ( n66854 , n66777 , n66339 );
and ( n66855 , n66854 , n66349 );
and ( n66856 , n66777 , n66339 );
or ( n66857 , n66855 , n66856 );
xor ( n66858 , n66825 , n66355 );
xor ( n66859 , n66858 , n66835 );
xor ( n66860 , n66825 , n66355 );
and ( n66861 , n66860 , n66835 );
and ( n66862 , n66825 , n66355 );
or ( n66863 , n66861 , n66862 );
xor ( n66864 , n66847 , n66361 );
xor ( n66865 , n66864 , n66841 );
xor ( n66866 , n66847 , n66361 );
and ( n66867 , n66866 , n66841 );
and ( n66868 , n66847 , n66361 );
or ( n66869 , n66867 , n66868 );
xor ( n66870 , n66367 , n66373 );
xor ( n66871 , n66870 , n66853 );
xor ( n66872 , n66367 , n66373 );
and ( n66873 , n66872 , n66853 );
and ( n66874 , n66367 , n66373 );
or ( n66875 , n66873 , n66874 );
xor ( n66876 , n66859 , n66379 );
xor ( n66877 , n66876 , n66865 );
xor ( n66878 , n66859 , n66379 );
and ( n66879 , n66878 , n66865 );
and ( n66880 , n66859 , n66379 );
or ( n66881 , n66879 , n66880 );
xor ( n66882 , n66385 , n66871 );
xor ( n66883 , n66882 , n66391 );
xor ( n66884 , n66385 , n66871 );
and ( n66885 , n66884 , n66391 );
and ( n66886 , n66385 , n66871 );
or ( n66887 , n66885 , n66886 );
xor ( n66888 , n66877 , n66883 );
xor ( n66889 , n66888 , n66397 );
xor ( n66890 , n66877 , n66883 );
and ( n66891 , n66890 , n66397 );
and ( n66892 , n66877 , n66883 );
or ( n66893 , n66891 , n66892 );
xor ( n66894 , n66598 , n66609 );
and ( n66895 , n66894 , n66623 );
and ( n66896 , n66598 , n66609 );
or ( n66897 , n66895 , n66896 );
xor ( n66898 , n66567 , n66579 );
and ( n66899 , n66898 , n66582 );
and ( n66900 , n66567 , n66579 );
or ( n66901 , n66899 , n66900 );
xor ( n66902 , n66723 , n66724 );
and ( n66903 , n66902 , n66737 );
and ( n66904 , n66723 , n66724 );
or ( n66905 , n66903 , n66904 );
xor ( n66906 , n66752 , n66762 );
and ( n66907 , n66906 , n66774 );
and ( n66908 , n66752 , n66762 );
or ( n66909 , n66907 , n66908 );
xor ( n66910 , n66688 , n66698 );
and ( n66911 , n66910 , n66711 );
and ( n66912 , n66688 , n66698 );
or ( n66913 , n66911 , n66912 );
xor ( n66914 , n66806 , n66816 );
and ( n66915 , n66914 , n65981 );
and ( n66916 , n66806 , n66816 );
or ( n66917 , n66915 , n66916 );
xor ( n66918 , n66792 , n66017 );
and ( n66919 , n66918 , n66343 );
and ( n66920 , n66792 , n66017 );
or ( n66921 , n66919 , n66920 );
not ( n66922 , n66476 );
not ( n66923 , n55576 );
or ( n66924 , n66922 , n66923 );
and ( n66925 , n52592 , n55125 );
not ( n66926 , n52592 );
and ( n66927 , n66926 , n55152 );
or ( n66928 , n66925 , n66927 );
nand ( n66929 , n66928 , n54848 );
nand ( n66930 , n66924 , n66929 );
not ( n66931 , n66488 );
not ( n66932 , n56281 );
or ( n66933 , n66931 , n66932 );
not ( n66934 , n48486 );
not ( n66935 , n56285 );
or ( n66936 , n66934 , n66935 );
nand ( n66937 , n55891 , n50084 );
nand ( n66938 , n66936 , n66937 );
nand ( n66939 , n66938 , n59984 );
nand ( n66940 , n66933 , n66939 );
xor ( n66941 , n66930 , n66940 );
not ( n66942 , n66632 );
not ( n66943 , n56777 );
or ( n66944 , n66942 , n66943 );
not ( n66945 , n63059 );
buf ( n66946 , n48118 );
not ( n66947 , n66946 );
not ( n66948 , n66947 );
or ( n66949 , n66945 , n66948 );
nand ( n66950 , n56786 , n66946 );
nand ( n66951 , n66949 , n66950 );
nand ( n66952 , n56780 , n66951 );
nand ( n66953 , n66944 , n66952 );
xor ( n66954 , n66941 , n66953 );
xor ( n66955 , n66930 , n66940 );
and ( n66956 , n66955 , n66953 );
and ( n66957 , n66930 , n66940 );
or ( n66958 , n66956 , n66957 );
not ( n66959 , n66644 );
not ( n66960 , n66005 );
or ( n66961 , n66959 , n66960 );
not ( n66962 , n52379 );
not ( n66963 , n66642 );
not ( n66964 , n66963 );
or ( n66965 , n66962 , n66964 );
nand ( n66966 , n65175 , n41416 );
nand ( n66967 , n66965 , n66966 );
nand ( n66968 , n57631 , n66967 );
nand ( n66969 , n66961 , n66968 );
not ( n66970 , n66453 );
not ( n66971 , n53956 );
or ( n66972 , n66970 , n66971 );
and ( n66973 , n53615 , n50020 );
not ( n66974 , n53615 );
and ( n66975 , n66974 , n66226 );
or ( n66976 , n66973 , n66975 );
nand ( n66977 , n66976 , n53620 );
nand ( n66978 , n66972 , n66977 );
xor ( n66979 , n66969 , n66978 );
not ( n66980 , n59571 );
not ( n66981 , n66596 );
or ( n66982 , n66980 , n66981 );
buf ( n66983 , n65121 );
and ( n66984 , n66983 , n48983 );
not ( n66985 , n66983 );
and ( n66986 , n66985 , n56348 );
nor ( n66987 , n66984 , n66986 );
or ( n66988 , n59574 , n66987 );
nand ( n66989 , n66982 , n66988 );
xor ( n66990 , n66979 , n66989 );
xor ( n66991 , n66969 , n66978 );
and ( n66992 , n66991 , n66989 );
and ( n66993 , n66969 , n66978 );
or ( n66994 , n66992 , n66993 );
not ( n66995 , n52043 );
not ( n66996 , n48645 );
not ( n66997 , n65006 );
or ( n66998 , n66996 , n66997 );
nand ( n66999 , n39056 , n49679 );
nand ( n67000 , n66998 , n66999 );
not ( n67001 , n67000 );
or ( n67002 , n66995 , n67001 );
nand ( n67003 , n66527 , n52970 );
nand ( n67004 , n67002 , n67003 );
not ( n67005 , n46776 );
not ( n67006 , n66788 );
or ( n67007 , n67005 , n67006 );
nand ( n67008 , n47827 , n50263 );
nand ( n67009 , n67007 , n67008 );
xor ( n67010 , n67004 , n67009 );
not ( n67011 , n52421 );
not ( n67012 , n66551 );
or ( n67013 , n67011 , n67012 );
buf ( n67014 , n58933 );
and ( n67015 , n51723 , n67014 );
not ( n67016 , n51723 );
and ( n67017 , n67016 , n60905 );
or ( n67018 , n67015 , n67017 );
nand ( n67019 , n54875 , n67018 );
nand ( n67020 , n67013 , n67019 );
xor ( n67021 , n67010 , n67020 );
xor ( n67022 , n67004 , n67009 );
and ( n67023 , n67022 , n67020 );
and ( n67024 , n67004 , n67009 );
or ( n67025 , n67023 , n67024 );
not ( n67026 , n47384 );
and ( n67027 , n49500 , n66052 );
not ( n67028 , n49500 );
and ( n67029 , n67028 , n66053 );
or ( n67030 , n67027 , n67029 );
not ( n67031 , n67030 );
or ( n67032 , n67026 , n67031 );
nand ( n67033 , n66504 , n48989 );
nand ( n67034 , n67032 , n67033 );
not ( n67035 , n52004 );
not ( n67036 , n52377 );
not ( n67037 , n39779 );
not ( n67038 , n67037 );
or ( n67039 , n67036 , n67038 );
buf ( n67040 , n58047 );
not ( n67041 , n67040 );
nand ( n67042 , n67041 , n55013 );
nand ( n67043 , n67039 , n67042 );
not ( n67044 , n67043 );
or ( n67045 , n67035 , n67044 );
nand ( n67046 , n66814 , n57314 );
nand ( n67047 , n67045 , n67046 );
xor ( n67048 , n67034 , n67047 );
not ( n67049 , n66577 );
not ( n67050 , n65089 );
or ( n67051 , n67049 , n67050 );
not ( n67052 , n48898 );
not ( n67053 , n63412 );
or ( n67054 , n67052 , n67053 );
nand ( n67055 , n63922 , n48897 );
nand ( n67056 , n67054 , n67055 );
nand ( n67057 , n67056 , n65092 );
nand ( n67058 , n67051 , n67057 );
not ( n67059 , n66565 );
not ( n67060 , n67059 );
buf ( n67061 , n62463 );
not ( n67062 , n67061 );
or ( n67063 , n67060 , n67062 );
and ( n67064 , n66089 , n51204 );
and ( n67065 , n62451 , n48860 );
nor ( n67066 , n67064 , n67065 );
not ( n67067 , n67066 );
not ( n67068 , n62466 );
nand ( n67069 , n67067 , n67068 );
nand ( n67070 , n67063 , n67069 );
xor ( n67071 , n67058 , n67070 );
buf ( n67072 , n63922 );
and ( n67073 , n67072 , n47227 );
xor ( n67074 , n67071 , n67073 );
xor ( n67075 , n67048 , n67074 );
xor ( n67076 , n67034 , n67047 );
and ( n67077 , n67076 , n67074 );
and ( n67078 , n67034 , n67047 );
or ( n67079 , n67077 , n67078 );
not ( n67080 , n66607 );
not ( n67081 , n65130 );
or ( n67082 , n67080 , n67081 );
not ( n67083 , n54611 );
not ( n67084 , n66140 );
not ( n67085 , n67084 );
or ( n67086 , n67083 , n67085 );
nand ( n67087 , n66140 , n51670 );
nand ( n67088 , n67086 , n67087 );
nand ( n67089 , n60427 , n67088 );
nand ( n67090 , n67082 , n67089 );
not ( n67091 , n66621 );
not ( n67092 , n64111 );
or ( n67093 , n67091 , n67092 );
not ( n67094 , n65144 );
and ( n67095 , n51792 , n61537 );
not ( n67096 , n51792 );
and ( n67097 , n67096 , n66615 );
or ( n67098 , n67095 , n67097 );
nand ( n67099 , n67094 , n67098 );
nand ( n67100 , n67093 , n67099 );
xor ( n67101 , n67090 , n67100 );
not ( n67102 , n66657 );
not ( n67103 , n65646 );
or ( n67104 , n67102 , n67103 );
not ( n67105 , n57182 );
not ( n67106 , n66652 );
or ( n67107 , n67105 , n67106 );
nand ( n67108 , n65184 , n58195 );
nand ( n67109 , n67107 , n67108 );
nand ( n67110 , n61465 , n67109 );
nand ( n67111 , n67104 , n67110 );
xor ( n67112 , n67101 , n67111 );
xor ( n67113 , n66954 , n67112 );
xor ( n67114 , n67113 , n66990 );
xor ( n67115 , n66954 , n67112 );
and ( n67116 , n67115 , n66990 );
and ( n67117 , n66954 , n67112 );
or ( n67118 , n67116 , n67117 );
xor ( n67119 , n66905 , n66909 );
xor ( n67120 , n67119 , n66913 );
xor ( n67121 , n66905 , n66909 );
and ( n67122 , n67121 , n66913 );
and ( n67123 , n66905 , n66909 );
or ( n67124 , n67122 , n67123 );
xor ( n67125 , n66560 , n66917 );
xor ( n67126 , n67125 , n66921 );
xor ( n67127 , n66560 , n66917 );
and ( n67128 , n67127 , n66921 );
and ( n67129 , n66560 , n66917 );
or ( n67130 , n67128 , n67129 );
not ( n67131 , n62654 );
not ( n67132 , n61951 );
not ( n67133 , n66236 );
or ( n67134 , n67132 , n67133 );
nand ( n67135 , n40364 , n66690 );
nand ( n67136 , n67134 , n67135 );
not ( n67137 , n67136 );
or ( n67138 , n67131 , n67137 );
not ( n67139 , n66690 );
not ( n67140 , n67139 );
not ( n67141 , n40225 );
or ( n67142 , n67140 , n67141 );
nand ( n67143 , n67142 , n66692 );
nand ( n67144 , n67143 , n66696 );
nand ( n67145 , n67138 , n67144 );
not ( n67146 , n63708 );
not ( n67147 , n66707 );
or ( n67148 , n67146 , n67147 );
not ( n67149 , n50306 );
not ( n67150 , n53289 );
or ( n67151 , n67149 , n67150 );
nand ( n67152 , n54646 , n66705 );
nand ( n67153 , n67151 , n67152 );
nand ( n67154 , n67153 , n52757 );
nand ( n67155 , n67148 , n67154 );
xor ( n67156 , n67145 , n67155 );
not ( n67157 , n52151 );
not ( n67158 , n66802 );
or ( n67159 , n67157 , n67158 );
not ( n67160 , n51465 );
not ( n67161 , n53271 );
or ( n67162 , n67160 , n67161 );
nand ( n67163 , n40626 , n50899 );
nand ( n67164 , n67162 , n67163 );
nand ( n67165 , n67164 , n50922 );
nand ( n67166 , n67159 , n67165 );
xor ( n67167 , n67156 , n67166 );
xor ( n67168 , n66522 , n67167 );
not ( n67169 , n52469 );
not ( n67170 , n52980 );
not ( n67171 , n40692 );
or ( n67172 , n67170 , n67171 );
or ( n67173 , n40692 , n53189 );
nand ( n67174 , n67172 , n67173 );
not ( n67175 , n67174 );
or ( n67176 , n67169 , n67175 );
not ( n67177 , n56853 );
nand ( n67178 , n67177 , n66442 );
nand ( n67179 , n67176 , n67178 );
not ( n67180 , n51766 );
not ( n67181 , n53918 );
not ( n67182 , n59176 );
or ( n67183 , n67181 , n67182 );
nand ( n67184 , n59179 , n52110 );
nand ( n67185 , n67183 , n67184 );
not ( n67186 , n67185 );
or ( n67187 , n67180 , n67186 );
nand ( n67188 , n66719 , n53197 );
nand ( n67189 , n67187 , n67188 );
xor ( n67190 , n67179 , n67189 );
not ( n67191 , n58977 );
not ( n67192 , n60602 );
buf ( n67193 , n56454 );
not ( n67194 , n67193 );
or ( n67195 , n67192 , n67194 );
buf ( n67196 , n40012 );
nand ( n67197 , n67196 , n52728 );
nand ( n67198 , n67195 , n67197 );
not ( n67199 , n67198 );
or ( n67200 , n67191 , n67199 );
nand ( n67201 , n66760 , n53104 );
nand ( n67202 , n67200 , n67201 );
xor ( n67203 , n67190 , n67202 );
xor ( n67204 , n67168 , n67203 );
xor ( n67205 , n66522 , n67167 );
and ( n67206 , n67205 , n67203 );
and ( n67207 , n66522 , n67167 );
or ( n67208 , n67206 , n67207 );
not ( n67209 , n56639 );
not ( n67210 , n59345 );
not ( n67211 , n56407 );
or ( n67212 , n67210 , n67211 );
nand ( n67213 , n56412 , n60617 );
nand ( n67214 , n67212 , n67213 );
not ( n67215 , n67214 );
or ( n67216 , n67209 , n67215 );
nand ( n67217 , n66770 , n59950 );
nand ( n67218 , n67216 , n67217 );
not ( n67219 , n60927 );
not ( n67220 , n49112 );
not ( n67221 , n55641 );
or ( n67222 , n67220 , n67221 );
nand ( n67223 , n56441 , n60292 );
nand ( n67224 , n67222 , n67223 );
not ( n67225 , n67224 );
or ( n67226 , n67219 , n67225 );
nand ( n67227 , n66686 , n58168 );
nand ( n67228 , n67226 , n67227 );
xor ( n67229 , n67218 , n67228 );
not ( n67230 , n66466 );
or ( n67231 , n55161 , n67230 );
and ( n67232 , n62861 , n59078 );
not ( n67233 , n62861 );
and ( n67234 , n67233 , n54322 );
nor ( n67235 , n67232 , n67234 );
or ( n67236 , n54326 , n67235 );
nand ( n67237 , n67231 , n67236 );
not ( n67238 , n67237 );
xor ( n67239 , n67229 , n67238 );
not ( n67240 , n55066 );
not ( n67241 , n52816 );
not ( n67242 , n60138 );
or ( n67243 , n67241 , n67242 );
not ( n67244 , n52570 );
nand ( n67245 , n67244 , n53928 );
nand ( n67246 , n67243 , n67245 );
not ( n67247 , n67246 );
or ( n67248 , n67240 , n67247 );
nand ( n67249 , n66748 , n56355 );
nand ( n67250 , n67248 , n67249 );
not ( n67251 , n54623 );
not ( n67252 , n54625 );
not ( n67253 , n60167 );
or ( n67254 , n67252 , n67253 );
not ( n67255 , n62970 );
nand ( n67256 , n67255 , n55023 );
nand ( n67257 , n67254 , n67256 );
not ( n67258 , n67257 );
or ( n67259 , n67251 , n67258 );
nand ( n67260 , n66731 , n52022 );
nand ( n67261 , n67259 , n67260 );
xor ( n67262 , n67250 , n67261 );
xor ( n67263 , n67262 , n66460 );
xor ( n67264 , n67239 , n67263 );
not ( n67265 , n64498 );
not ( n67266 , n66538 );
or ( n67267 , n67265 , n67266 );
not ( n67268 , n54028 );
not ( n67269 , n66304 );
not ( n67270 , n67269 );
or ( n67271 , n67268 , n67270 );
nand ( n67272 , n42555 , n50634 );
nand ( n67273 , n67271 , n67272 );
nand ( n67274 , n67273 , n53675 );
nand ( n67275 , n67267 , n67274 );
xor ( n67276 , n66495 , n67275 );
xor ( n67277 , n67276 , n66833 );
xor ( n67278 , n67264 , n67277 );
xor ( n67279 , n67239 , n67263 );
and ( n67280 , n67279 , n67277 );
and ( n67281 , n67239 , n67263 );
or ( n67282 , n67280 , n67281 );
not ( n67283 , n51865 );
not ( n67284 , n52267 );
not ( n67285 , n39331 );
or ( n67286 , n67284 , n67285 );
nand ( n67287 , n39332 , n51351 );
nand ( n67288 , n67286 , n67287 );
not ( n67289 , n67288 );
or ( n67290 , n67283 , n67289 );
nand ( n67291 , n66515 , n49713 );
nand ( n67292 , n67290 , n67291 );
xor ( n67293 , n66897 , n67292 );
xor ( n67294 , n67293 , n66901 );
xor ( n67295 , n67294 , n66589 );
xor ( n67296 , n67295 , n67021 );
xor ( n67297 , n67294 , n66589 );
and ( n67298 , n67297 , n67021 );
and ( n67299 , n67294 , n66589 );
or ( n67300 , n67298 , n67299 );
xor ( n67301 , n67075 , n66666 );
xor ( n67302 , n67301 , n67114 );
xor ( n67303 , n67075 , n66666 );
and ( n67304 , n67303 , n67114 );
and ( n67305 , n67075 , n66666 );
or ( n67306 , n67304 , n67305 );
xor ( n67307 , n67120 , n66672 );
xor ( n67308 , n67307 , n66678 );
xor ( n67309 , n67120 , n66672 );
and ( n67310 , n67309 , n66678 );
and ( n67311 , n67120 , n66672 );
or ( n67312 , n67310 , n67311 );
xor ( n67313 , n67090 , n67100 );
and ( n67314 , n67313 , n67111 );
and ( n67315 , n67090 , n67100 );
or ( n67316 , n67314 , n67315 );
xor ( n67317 , n66743 , n67204 );
xor ( n67318 , n67317 , n67126 );
xor ( n67319 , n66743 , n67204 );
and ( n67320 , n67319 , n67126 );
and ( n67321 , n66743 , n67204 );
or ( n67322 , n67320 , n67321 );
xor ( n67323 , n66781 , n66823 );
xor ( n67324 , n67323 , n66829 );
xor ( n67325 , n66781 , n66823 );
and ( n67326 , n67325 , n66829 );
and ( n67327 , n66781 , n66823 );
or ( n67328 , n67326 , n67327 );
xor ( n67329 , n67278 , n67296 );
xor ( n67330 , n67329 , n67302 );
xor ( n67331 , n67278 , n67296 );
and ( n67332 , n67331 , n67302 );
and ( n67333 , n67278 , n67296 );
or ( n67334 , n67332 , n67333 );
xor ( n67335 , n66839 , n66845 );
xor ( n67336 , n67335 , n67308 );
xor ( n67337 , n66839 , n66845 );
and ( n67338 , n67337 , n67308 );
and ( n67339 , n66839 , n66845 );
or ( n67340 , n67338 , n67339 );
xor ( n67341 , n66851 , n67318 );
xor ( n67342 , n67341 , n67324 );
xor ( n67343 , n66851 , n67318 );
and ( n67344 , n67343 , n67324 );
and ( n67345 , n66851 , n67318 );
or ( n67346 , n67344 , n67345 );
xor ( n67347 , n66857 , n67330 );
xor ( n67348 , n67347 , n66863 );
xor ( n67349 , n66857 , n67330 );
and ( n67350 , n67349 , n66863 );
and ( n67351 , n66857 , n67330 );
or ( n67352 , n67350 , n67351 );
xor ( n67353 , n67336 , n66869 );
xor ( n67354 , n67353 , n67342 );
xor ( n67355 , n67336 , n66869 );
and ( n67356 , n67355 , n67342 );
and ( n67357 , n67336 , n66869 );
or ( n67358 , n67356 , n67357 );
xor ( n67359 , n66875 , n67348 );
xor ( n67360 , n67359 , n67354 );
xor ( n67361 , n66875 , n67348 );
and ( n67362 , n67361 , n67354 );
and ( n67363 , n66875 , n67348 );
or ( n67364 , n67362 , n67363 );
xor ( n67365 , n66881 , n67360 );
xor ( n67366 , n67365 , n66887 );
xor ( n67367 , n66881 , n67360 );
and ( n67368 , n67367 , n66887 );
and ( n67369 , n66881 , n67360 );
or ( n67370 , n67368 , n67369 );
xor ( n67371 , n67058 , n67070 );
and ( n67372 , n67371 , n67073 );
and ( n67373 , n67058 , n67070 );
or ( n67374 , n67372 , n67373 );
xor ( n67375 , n67179 , n67189 );
and ( n67376 , n67375 , n67202 );
and ( n67377 , n67179 , n67189 );
or ( n67378 , n67376 , n67377 );
xor ( n67379 , n67218 , n67228 );
and ( n67380 , n67379 , n67238 );
and ( n67381 , n67218 , n67228 );
or ( n67382 , n67380 , n67381 );
xor ( n67383 , n67145 , n67155 );
and ( n67384 , n67383 , n67166 );
and ( n67385 , n67145 , n67155 );
or ( n67386 , n67384 , n67385 );
xor ( n67387 , n67250 , n67261 );
and ( n67388 , n67387 , n66460 );
and ( n67389 , n67250 , n67261 );
or ( n67390 , n67388 , n67389 );
xor ( n67391 , n66495 , n67275 );
and ( n67392 , n67391 , n66833 );
and ( n67393 , n66495 , n67275 );
or ( n67394 , n67392 , n67393 );
xor ( n67395 , n66897 , n67292 );
and ( n67396 , n67395 , n66901 );
and ( n67397 , n66897 , n67292 );
or ( n67398 , n67396 , n67397 );
or ( n67399 , n48295 , n53631 );
nand ( n67400 , n67399 , n50263 );
not ( n67401 , n66976 );
not ( n67402 , n53956 );
or ( n67403 , n67401 , n67402 );
not ( n67404 , n53591 );
not ( n67405 , n52079 );
or ( n67406 , n67404 , n67405 );
not ( n67407 , n54249 );
nand ( n67408 , n67407 , n53615 );
nand ( n67409 , n67406 , n67408 );
nand ( n67410 , n67409 , n53619 );
nand ( n67411 , n67403 , n67410 );
xor ( n67412 , n67400 , n67411 );
or ( n67413 , n55161 , n67235 );
not ( n67414 , n64452 );
not ( n67415 , n55276 );
or ( n67416 , n67414 , n67415 );
not ( n67417 , n64970 );
nand ( n67418 , n67417 , n64451 );
nand ( n67419 , n67416 , n67418 );
not ( n67420 , n67419 );
or ( n67421 , n67420 , n54326 );
nand ( n67422 , n67413 , n67421 );
xor ( n67423 , n67412 , n67422 );
xor ( n67424 , n67400 , n67411 );
and ( n67425 , n67424 , n67422 );
and ( n67426 , n67400 , n67411 );
or ( n67427 , n67425 , n67426 );
not ( n67428 , n66928 );
not ( n67429 , n55144 );
or ( n67430 , n67428 , n67429 );
not ( n67431 , n49838 );
not ( n67432 , n55148 );
or ( n67433 , n67431 , n67432 );
nand ( n67434 , n55582 , n52796 );
nand ( n67435 , n67433 , n67434 );
nand ( n67436 , n55157 , n67435 );
nand ( n67437 , n67430 , n67436 );
not ( n67438 , n66938 );
not ( n67439 , n56281 );
or ( n67440 , n67438 , n67439 );
not ( n67441 , n49190 );
nand ( n67442 , n55846 , n67441 );
not ( n67443 , n67442 );
nand ( n67444 , n55892 , n49190 );
not ( n67445 , n67444 );
or ( n67446 , n67443 , n67445 );
nand ( n67447 , n67446 , n55458 );
nand ( n67448 , n67440 , n67447 );
xor ( n67449 , n67437 , n67448 );
not ( n67450 , n66951 );
not ( n67451 , n56777 );
or ( n67452 , n67450 , n67451 );
not ( n67453 , n41532 );
not ( n67454 , n65999 );
not ( n67455 , n67454 );
or ( n67456 , n67453 , n67455 );
nand ( n67457 , n56786 , n44112 );
nand ( n67458 , n67456 , n67457 );
nand ( n67459 , n60472 , n67458 );
nand ( n67460 , n67452 , n67459 );
xor ( n67461 , n67449 , n67460 );
xor ( n67462 , n67437 , n67448 );
and ( n67463 , n67462 , n67460 );
and ( n67464 , n67437 , n67448 );
or ( n67465 , n67463 , n67464 );
not ( n67466 , n49713 );
not ( n67467 , n67288 );
or ( n67468 , n67466 , n67467 );
not ( n67469 , n52267 );
not ( n67470 , n66500 );
or ( n67471 , n67469 , n67470 );
nand ( n67472 , n39253 , n48661 );
nand ( n67473 , n67471 , n67472 );
nand ( n67474 , n67473 , n51865 );
nand ( n67475 , n67468 , n67474 );
not ( n67476 , n52962 );
buf ( n67477 , n49679 );
not ( n67478 , n67477 );
not ( n67479 , n67478 );
not ( n67480 , n62394 );
or ( n67481 , n67479 , n67480 );
not ( n67482 , n62394 );
nand ( n67483 , n67482 , n52048 );
nand ( n67484 , n67481 , n67483 );
not ( n67485 , n67484 );
or ( n67486 , n67476 , n67485 );
nand ( n67487 , n67000 , n52970 );
nand ( n67488 , n67486 , n67487 );
xor ( n67489 , n67475 , n67488 );
not ( n67490 , n52421 );
not ( n67491 , n67018 );
or ( n67492 , n67490 , n67491 );
not ( n67493 , n51723 );
not ( n67494 , n59402 );
or ( n67495 , n67493 , n67494 );
not ( n67496 , n48856 );
nand ( n67497 , n67496 , n59403 );
nand ( n67498 , n67495 , n67497 );
nand ( n67499 , n67498 , n54875 );
nand ( n67500 , n67492 , n67499 );
xor ( n67501 , n67489 , n67500 );
xor ( n67502 , n67475 , n67488 );
and ( n67503 , n67502 , n67500 );
and ( n67504 , n67475 , n67488 );
or ( n67505 , n67503 , n67504 );
not ( n67506 , n47384 );
not ( n67507 , n49500 );
not ( n67508 , n42399 );
or ( n67509 , n67507 , n67508 );
nand ( n67510 , n65546 , n53997 );
nand ( n67511 , n67509 , n67510 );
not ( n67512 , n67511 );
or ( n67513 , n67506 , n67512 );
nand ( n67514 , n67030 , n48989 );
nand ( n67515 , n67513 , n67514 );
not ( n67516 , n52004 );
not ( n67517 , n52377 );
not ( n67518 , n60383 );
or ( n67519 , n67517 , n67518 );
nand ( n67520 , n66546 , n55013 );
nand ( n67521 , n67519 , n67520 );
not ( n67522 , n67521 );
or ( n67523 , n67516 , n67522 );
nand ( n67524 , n67043 , n57314 );
nand ( n67525 , n67523 , n67524 );
xor ( n67526 , n67515 , n67525 );
xor ( n67527 , n67526 , n67423 );
xor ( n67528 , n67515 , n67525 );
and ( n67529 , n67528 , n67423 );
and ( n67530 , n67515 , n67525 );
or ( n67531 , n67529 , n67530 );
not ( n67532 , n67088 );
not ( n67533 , n63029 );
or ( n67534 , n67532 , n67533 );
not ( n67535 , n54185 );
not ( n67536 , n67084 );
or ( n67537 , n67535 , n67536 );
nand ( n67538 , n66140 , n54184 );
nand ( n67539 , n67537 , n67538 );
nand ( n67540 , n66602 , n67539 );
nand ( n67541 , n67534 , n67540 );
not ( n67542 , n67098 );
not ( n67543 , n64111 );
or ( n67544 , n67542 , n67543 );
not ( n67545 , n52033 );
not ( n67546 , n61537 );
or ( n67547 , n67545 , n67546 );
nand ( n67548 , n66619 , n55959 );
nand ( n67549 , n67547 , n67548 );
nand ( n67550 , n61557 , n67549 );
nand ( n67551 , n67544 , n67550 );
xor ( n67552 , n67541 , n67551 );
or ( n67553 , n64164 , n67066 );
and ( n67554 , n66089 , n49624 );
not ( n67555 , n64167 );
and ( n67556 , n67555 , n49630 );
nor ( n67557 , n67554 , n67556 );
or ( n67558 , n64166 , n67557 );
nand ( n67559 , n67553 , n67558 );
xor ( n67560 , n67552 , n67559 );
xor ( n67561 , n67560 , n67461 );
not ( n67562 , n66967 );
not ( n67563 , n60482 );
or ( n67564 , n67562 , n67563 );
not ( n67565 , n58458 );
not ( n67566 , n66963 );
or ( n67567 , n67565 , n67566 );
buf ( n67568 , n66642 );
nand ( n67569 , n67568 , n58459 );
nand ( n67570 , n67567 , n67569 );
nand ( n67571 , n57631 , n67570 );
nand ( n67572 , n67564 , n67571 );
not ( n67573 , n67109 );
not ( n67574 , n63080 );
or ( n67575 , n67573 , n67574 );
not ( n67576 , n47527 );
not ( n67577 , n65187 );
or ( n67578 , n67576 , n67577 );
nand ( n67579 , n58642 , n59388 );
nand ( n67580 , n67578 , n67579 );
nand ( n67581 , n61465 , n67580 );
nand ( n67582 , n67575 , n67581 );
xor ( n67583 , n67572 , n67582 );
not ( n67584 , n62506 );
or ( n67585 , n67584 , n66987 );
not ( n67586 , n60542 );
and ( n67587 , n56731 , n65664 );
not ( n67588 , n56731 );
and ( n67589 , n67588 , n63587 );
nor ( n67590 , n67587 , n67589 );
or ( n67591 , n67586 , n67590 );
nand ( n67592 , n67585 , n67591 );
xor ( n67593 , n67583 , n67592 );
xor ( n67594 , n67561 , n67593 );
xor ( n67595 , n67560 , n67461 );
and ( n67596 , n67595 , n67593 );
and ( n67597 , n67560 , n67461 );
or ( n67598 , n67596 , n67597 );
xor ( n67599 , n67378 , n67382 );
xor ( n67600 , n67599 , n67386 );
xor ( n67601 , n67378 , n67382 );
and ( n67602 , n67601 , n67386 );
and ( n67603 , n67378 , n67382 );
or ( n67604 , n67602 , n67603 );
not ( n67605 , n67056 );
not ( n67606 , n65795 );
or ( n67607 , n67605 , n67606 );
not ( n67608 , n47765 );
not ( n67609 , n63412 );
or ( n67610 , n67608 , n67609 );
nand ( n67611 , n66575 , n48589 );
nand ( n67612 , n67610 , n67611 );
nand ( n67613 , n65092 , n67612 );
nand ( n67614 , n67607 , n67613 );
not ( n67615 , n66581 );
nor ( n67616 , n67615 , n47368 );
xor ( n67617 , n67614 , n67616 );
not ( n67618 , n53571 );
not ( n67619 , n54283 );
not ( n67620 , n51574 );
or ( n67621 , n67619 , n67620 );
nand ( n67622 , n52284 , n52980 );
nand ( n67623 , n67621 , n67622 );
not ( n67624 , n67623 );
or ( n67625 , n67618 , n67624 );
nand ( n67626 , n67174 , n52854 );
nand ( n67627 , n67625 , n67626 );
xor ( n67628 , n67617 , n67627 );
xor ( n67629 , n67628 , n67394 );
xor ( n67630 , n67629 , n67398 );
xor ( n67631 , n67628 , n67394 );
and ( n67632 , n67631 , n67398 );
and ( n67633 , n67628 , n67394 );
or ( n67634 , n67632 , n67633 );
not ( n67635 , n51223 );
not ( n67636 , n51465 );
not ( n67637 , n63656 );
or ( n67638 , n67636 , n67637 );
not ( n67639 , n65773 );
nand ( n67640 , n59612 , n67639 );
nand ( n67641 , n67638 , n67640 );
not ( n67642 , n67641 );
or ( n67643 , n67635 , n67642 );
nand ( n67644 , n67164 , n52151 );
nand ( n67645 , n67643 , n67644 );
not ( n67646 , n55066 );
not ( n67647 , n65103 );
not ( n67648 , n53730 );
or ( n67649 , n67647 , n67648 );
nand ( n67650 , n40592 , n51566 );
nand ( n67651 , n67649 , n67650 );
not ( n67652 , n67651 );
or ( n67653 , n67646 , n67652 );
nand ( n67654 , n67246 , n56355 );
nand ( n67655 , n67653 , n67654 );
xor ( n67656 , n67645 , n67655 );
xor ( n67657 , n67656 , n67237 );
xor ( n67658 , n67025 , n67657 );
not ( n67659 , n60927 );
not ( n67660 , n62077 );
not ( n67661 , n65725 );
or ( n67662 , n67660 , n67661 );
nand ( n67663 , n59697 , n60292 );
nand ( n67664 , n67662 , n67663 );
not ( n67665 , n67664 );
or ( n67666 , n67659 , n67665 );
nand ( n67667 , n62085 , n67224 );
nand ( n67668 , n67666 , n67667 );
not ( n67669 , n52058 );
not ( n67670 , n67136 );
or ( n67671 , n67669 , n67670 );
not ( n67672 , n61951 );
not ( n67673 , n62626 );
or ( n67674 , n67672 , n67673 );
buf ( n67675 , n54406 );
nand ( n67676 , n67675 , n61952 );
nand ( n67677 , n67674 , n67676 );
nand ( n67678 , n67677 , n62654 );
nand ( n67679 , n67671 , n67678 );
xor ( n67680 , n67668 , n67679 );
not ( n67681 , n67153 );
not ( n67682 , n63708 );
or ( n67683 , n67681 , n67682 );
and ( n67684 , n64191 , n54433 );
not ( n67685 , n64191 );
and ( n67686 , n67685 , n56074 );
nor ( n67687 , n67684 , n67686 );
or ( n67688 , n67687 , n59828 );
nand ( n67689 , n67683 , n67688 );
xor ( n67690 , n67680 , n67689 );
xor ( n67691 , n67658 , n67690 );
xor ( n67692 , n67025 , n67657 );
and ( n67693 , n67692 , n67690 );
and ( n67694 , n67025 , n67657 );
or ( n67695 , n67693 , n67694 );
not ( n67696 , n53104 );
not ( n67697 , n67198 );
or ( n67698 , n67696 , n67697 );
not ( n67699 , n58982 );
not ( n67700 , n59651 );
or ( n67701 , n67699 , n67700 );
not ( n67702 , n59651 );
nand ( n67703 , n67702 , n52728 );
nand ( n67704 , n67701 , n67703 );
nand ( n67705 , n67704 , n58977 );
nand ( n67706 , n67698 , n67705 );
not ( n67707 , n52490 );
not ( n67708 , n51602 );
or ( n67709 , n67707 , n67708 );
nand ( n67710 , n51601 , n52110 );
nand ( n67711 , n67709 , n67710 );
not ( n67712 , n67711 );
not ( n67713 , n51766 );
or ( n67714 , n67712 , n67713 );
nand ( n67715 , n67185 , n52482 );
nand ( n67716 , n67714 , n67715 );
xor ( n67717 , n67706 , n67716 );
not ( n67718 , n59345 );
not ( n67719 , n56020 );
or ( n67720 , n67718 , n67719 );
not ( n67721 , n40513 );
nand ( n67722 , n67721 , n65743 );
nand ( n67723 , n67720 , n67722 );
nand ( n67724 , n67723 , n56639 );
nand ( n67725 , n67214 , n59950 );
nand ( n67726 , n67724 , n67725 );
xor ( n67727 , n67717 , n67726 );
xor ( n67728 , n67727 , n67390 );
xor ( n67729 , n67728 , n67079 );
xor ( n67730 , n67727 , n67390 );
and ( n67731 , n67730 , n67079 );
and ( n67732 , n67727 , n67390 );
or ( n67733 , n67731 , n67732 );
not ( n67734 , n52022 );
not ( n67735 , n67257 );
or ( n67736 , n67734 , n67735 );
not ( n67737 , n54625 );
not ( n67738 , n39893 );
or ( n67739 , n67737 , n67738 );
nand ( n67740 , n57787 , n54628 );
nand ( n67741 , n67739 , n67740 );
nand ( n67742 , n67741 , n54623 );
nand ( n67743 , n67736 , n67742 );
xor ( n67744 , n67743 , n66958 );
xor ( n67745 , n67744 , n66994 );
xor ( n67746 , n67118 , n67745 );
not ( n67747 , n64498 );
not ( n67748 , n67273 );
or ( n67749 , n67747 , n67748 );
not ( n67750 , n47803 );
not ( n67751 , n42653 );
or ( n67752 , n67750 , n67751 );
nand ( n67753 , n63794 , n48727 );
nand ( n67754 , n67752 , n67753 );
nand ( n67755 , n67754 , n53675 );
nand ( n67756 , n67749 , n67755 );
xor ( n67757 , n67756 , n67316 );
xor ( n67758 , n67757 , n67374 );
xor ( n67759 , n67746 , n67758 );
xor ( n67760 , n67118 , n67745 );
and ( n67761 , n67760 , n67758 );
and ( n67762 , n67118 , n67745 );
or ( n67763 , n67761 , n67762 );
xor ( n67764 , n67501 , n67527 );
xor ( n67765 , n67764 , n67594 );
xor ( n67766 , n67501 , n67527 );
and ( n67767 , n67766 , n67594 );
and ( n67768 , n67501 , n67527 );
or ( n67769 , n67767 , n67768 );
xor ( n67770 , n67124 , n67600 );
xor ( n67771 , n67770 , n67130 );
xor ( n67772 , n67124 , n67600 );
and ( n67773 , n67772 , n67130 );
and ( n67774 , n67124 , n67600 );
or ( n67775 , n67773 , n67774 );
xor ( n67776 , n67572 , n67582 );
and ( n67777 , n67776 , n67592 );
and ( n67778 , n67572 , n67582 );
or ( n67779 , n67777 , n67778 );
xor ( n67780 , n67208 , n67300 );
xor ( n67781 , n67780 , n67729 );
xor ( n67782 , n67208 , n67300 );
and ( n67783 , n67782 , n67729 );
and ( n67784 , n67208 , n67300 );
or ( n67785 , n67783 , n67784 );
xor ( n67786 , n67630 , n67282 );
xor ( n67787 , n67786 , n67691 );
xor ( n67788 , n67630 , n67282 );
and ( n67789 , n67788 , n67691 );
and ( n67790 , n67630 , n67282 );
or ( n67791 , n67789 , n67790 );
xor ( n67792 , n67306 , n67765 );
xor ( n67793 , n67792 , n67759 );
xor ( n67794 , n67306 , n67765 );
and ( n67795 , n67794 , n67759 );
and ( n67796 , n67306 , n67765 );
or ( n67797 , n67795 , n67796 );
xor ( n67798 , n67312 , n67771 );
xor ( n67799 , n67798 , n67322 );
xor ( n67800 , n67312 , n67771 );
and ( n67801 , n67800 , n67322 );
and ( n67802 , n67312 , n67771 );
or ( n67803 , n67801 , n67802 );
xor ( n67804 , n67328 , n67787 );
xor ( n67805 , n67804 , n67781 );
xor ( n67806 , n67328 , n67787 );
and ( n67807 , n67806 , n67781 );
and ( n67808 , n67328 , n67787 );
or ( n67809 , n67807 , n67808 );
xor ( n67810 , n67793 , n67334 );
xor ( n67811 , n67810 , n67340 );
xor ( n67812 , n67793 , n67334 );
and ( n67813 , n67812 , n67340 );
and ( n67814 , n67793 , n67334 );
or ( n67815 , n67813 , n67814 );
xor ( n67816 , n67799 , n67346 );
xor ( n67817 , n67816 , n67805 );
xor ( n67818 , n67799 , n67346 );
and ( n67819 , n67818 , n67805 );
and ( n67820 , n67799 , n67346 );
or ( n67821 , n67819 , n67820 );
xor ( n67822 , n67811 , n67352 );
xor ( n67823 , n67822 , n67358 );
xor ( n67824 , n67811 , n67352 );
and ( n67825 , n67824 , n67358 );
and ( n67826 , n67811 , n67352 );
or ( n67827 , n67825 , n67826 );
xor ( n67828 , n67817 , n67823 );
xor ( n67829 , n67828 , n67364 );
xor ( n67830 , n67817 , n67823 );
and ( n67831 , n67830 , n67364 );
and ( n67832 , n67817 , n67823 );
or ( n67833 , n67831 , n67832 );
xor ( n67834 , n67541 , n67551 );
and ( n67835 , n67834 , n67559 );
and ( n67836 , n67541 , n67551 );
or ( n67837 , n67835 , n67836 );
xor ( n67838 , n67614 , n67616 );
and ( n67839 , n67838 , n67627 );
and ( n67840 , n67614 , n67616 );
or ( n67841 , n67839 , n67840 );
xor ( n67842 , n67706 , n67716 );
and ( n67843 , n67842 , n67726 );
and ( n67844 , n67706 , n67716 );
or ( n67845 , n67843 , n67844 );
xor ( n67846 , n67668 , n67679 );
and ( n67847 , n67846 , n67689 );
and ( n67848 , n67668 , n67679 );
or ( n67849 , n67847 , n67848 );
xor ( n67850 , n67645 , n67655 );
and ( n67851 , n67850 , n67237 );
and ( n67852 , n67645 , n67655 );
or ( n67853 , n67851 , n67852 );
xor ( n67854 , n67743 , n66958 );
and ( n67855 , n67854 , n66994 );
and ( n67856 , n67743 , n66958 );
or ( n67857 , n67855 , n67856 );
xor ( n67858 , n67756 , n67316 );
and ( n67859 , n67858 , n67374 );
and ( n67860 , n67756 , n67316 );
or ( n67861 , n67859 , n67860 );
buf ( n67862 , n55887 );
not ( n67863 , n67862 );
nand ( n67864 , n67444 , n67442 );
not ( n67865 , n67864 );
or ( n67866 , n67863 , n67865 );
not ( n67867 , n52592 );
not ( n67868 , n58604 );
or ( n67869 , n67867 , n67868 );
nand ( n67870 , n56749 , n41287 );
nand ( n67871 , n67869 , n67870 );
nand ( n67872 , n55458 , n67871 );
nand ( n67873 , n67866 , n67872 );
not ( n67874 , n67458 );
not ( n67875 , n56777 );
or ( n67876 , n67874 , n67875 );
not ( n67877 , n41407 );
not ( n67878 , n67454 );
or ( n67879 , n67877 , n67878 );
nand ( n67880 , n56679 , n64972 );
nand ( n67881 , n67879 , n67880 );
nand ( n67882 , n56780 , n67881 );
nand ( n67883 , n67876 , n67882 );
xor ( n67884 , n67873 , n67883 );
not ( n67885 , n60482 );
not ( n67886 , n67570 );
or ( n67887 , n67885 , n67886 );
and ( n67888 , n66946 , n66642 );
not ( n67889 , n66946 );
buf ( n67890 , n59437 );
and ( n67891 , n67889 , n67890 );
nor ( n67892 , n67888 , n67891 );
or ( n67893 , n65638 , n67892 );
nand ( n67894 , n67887 , n67893 );
xor ( n67895 , n67884 , n67894 );
xor ( n67896 , n67873 , n67883 );
and ( n67897 , n67896 , n67894 );
and ( n67898 , n67873 , n67883 );
or ( n67899 , n67897 , n67898 );
not ( n67900 , n67580 );
not ( n67901 , n59445 );
or ( n67902 , n67900 , n67901 );
not ( n67903 , n58994 );
not ( n67904 , n58966 );
or ( n67905 , n67903 , n67904 );
not ( n67906 , n58994 );
nand ( n67907 , n58642 , n67906 );
nand ( n67908 , n67905 , n67907 );
nand ( n67909 , n61465 , n67908 );
nand ( n67910 , n67902 , n67909 );
not ( n67911 , n67419 );
not ( n67912 , n54316 );
or ( n67913 , n67911 , n67912 );
not ( n67914 , n50020 );
not ( n67915 , n59078 );
or ( n67916 , n67914 , n67915 );
not ( n67917 , n67417 );
nand ( n67918 , n67917 , n51891 );
nand ( n67919 , n67916 , n67918 );
nand ( n67920 , n54077 , n67919 );
nand ( n67921 , n67913 , n67920 );
xor ( n67922 , n67910 , n67921 );
not ( n67923 , n67539 );
not ( n67924 , n66136 );
or ( n67925 , n67923 , n67924 );
not ( n67926 , n48983 );
not ( n67927 , n66141 );
or ( n67928 , n67926 , n67927 );
nand ( n67929 , n66140 , n56348 );
nand ( n67930 , n67928 , n67929 );
nand ( n67931 , n66602 , n67930 );
nand ( n67932 , n67925 , n67931 );
xor ( n67933 , n67922 , n67932 );
xor ( n67934 , n67910 , n67921 );
and ( n67935 , n67934 , n67932 );
and ( n67936 , n67910 , n67921 );
or ( n67937 , n67935 , n67936 );
not ( n67938 , n49713 );
not ( n67939 , n67473 );
or ( n67940 , n67938 , n67939 );
not ( n67941 , n52267 );
not ( n67942 , n66052 );
or ( n67943 , n67941 , n67942 );
nand ( n67944 , n61907 , n51351 );
nand ( n67945 , n67943 , n67944 );
nand ( n67946 , n67945 , n51865 );
nand ( n67947 , n67940 , n67946 );
not ( n67948 , n52022 );
not ( n67949 , n67741 );
or ( n67950 , n67948 , n67949 );
nor ( n67951 , n54628 , n54622 );
nand ( n67952 , n67951 , n67037 );
not ( n67953 , n54622 );
nand ( n67954 , n67953 , n59913 , n54628 );
and ( n67955 , n67952 , n67954 );
nand ( n67956 , n67950 , n67955 );
xor ( n67957 , n67947 , n67956 );
xor ( n67958 , n67957 , n67427 );
xor ( n67959 , n67947 , n67956 );
and ( n67960 , n67959 , n67427 );
and ( n67961 , n67947 , n67956 );
or ( n67962 , n67960 , n67961 );
and ( n67963 , n67072 , n48898 );
not ( n67964 , n67612 );
not ( n67965 , n65089 );
or ( n67966 , n67964 , n67965 );
and ( n67967 , n51204 , n63415 );
not ( n67968 , n51204 );
not ( n67969 , n63412 );
and ( n67970 , n67968 , n67969 );
or ( n67971 , n67967 , n67970 );
nand ( n67972 , n65092 , n67971 );
nand ( n67973 , n67966 , n67972 );
xor ( n67974 , n67963 , n67973 );
not ( n67975 , n54364 );
and ( n67976 , n40691 , n53591 );
not ( n67977 , n40691 );
and ( n67978 , n67977 , n53596 );
or ( n67979 , n67976 , n67978 );
not ( n67980 , n67979 );
or ( n67981 , n67975 , n67980 );
not ( n67982 , n61329 );
nand ( n67983 , n67982 , n67409 );
nand ( n67984 , n67981 , n67983 );
xor ( n67985 , n67974 , n67984 );
not ( n67986 , n67549 );
not ( n67987 , n61548 );
or ( n67988 , n67986 , n67987 );
not ( n67989 , n55511 );
not ( n67990 , n61537 );
or ( n67991 , n67989 , n67990 );
nand ( n67992 , n63541 , n51670 );
nand ( n67993 , n67991 , n67992 );
nand ( n67994 , n62428 , n67993 );
nand ( n67995 , n67988 , n67994 );
or ( n67996 , n64164 , n67557 );
not ( n67997 , n51792 );
not ( n67998 , n62452 );
or ( n67999 , n67997 , n67998 );
nand ( n68000 , n62451 , n48829 );
nand ( n68001 , n67999 , n68000 );
not ( n68002 , n68001 );
or ( n68003 , n64166 , n68002 );
nand ( n68004 , n67996 , n68003 );
xor ( n68005 , n67995 , n68004 );
not ( n68006 , n59575 );
not ( n68007 , n57182 );
not ( n68008 , n63587 );
or ( n68009 , n68007 , n68008 );
nand ( n68010 , n62513 , n47332 );
nand ( n68011 , n68009 , n68010 );
not ( n68012 , n68011 );
or ( n68013 , n68006 , n68012 );
or ( n68014 , n66980 , n67590 );
nand ( n68015 , n68013 , n68014 );
xor ( n68016 , n68005 , n68015 );
xor ( n68017 , n67985 , n68016 );
xor ( n68018 , n68017 , n67895 );
xor ( n68019 , n67985 , n68016 );
and ( n68020 , n68019 , n67895 );
and ( n68021 , n67985 , n68016 );
or ( n68022 , n68020 , n68021 );
xor ( n68023 , n67933 , n67841 );
xor ( n68024 , n68023 , n67845 );
xor ( n68025 , n67933 , n67841 );
and ( n68026 , n68025 , n67845 );
and ( n68027 , n67933 , n67841 );
or ( n68028 , n68026 , n68027 );
xor ( n68029 , n67849 , n67853 );
xor ( n68030 , n68029 , n67861 );
xor ( n68031 , n67849 , n67853 );
and ( n68032 , n68031 , n67861 );
and ( n68033 , n67849 , n67853 );
or ( n68034 , n68032 , n68033 );
not ( n68035 , n52151 );
not ( n68036 , n67641 );
or ( n68037 , n68035 , n68036 );
not ( n68038 , n50898 );
not ( n68039 , n53289 );
or ( n68040 , n68038 , n68039 );
nand ( n68041 , n54646 , n67639 );
nand ( n68042 , n68040 , n68041 );
nand ( n68043 , n68042 , n51223 );
nand ( n68044 , n68037 , n68043 );
not ( n68045 , n51533 );
not ( n68046 , n65103 );
not ( n68047 , n40627 );
or ( n68048 , n68046 , n68047 );
buf ( n68049 , n40626 );
nand ( n68050 , n68049 , n53928 );
nand ( n68051 , n68048 , n68050 );
not ( n68052 , n68051 );
or ( n68053 , n68045 , n68052 );
nand ( n68054 , n67651 , n56355 );
nand ( n68055 , n68053 , n68054 );
xor ( n68056 , n68044 , n68055 );
not ( n68057 , n53197 );
not ( n68058 , n67711 );
or ( n68059 , n68057 , n68058 );
not ( n68060 , n52114 );
not ( n68061 , n60138 );
or ( n68062 , n68060 , n68061 );
nand ( n68063 , n51916 , n52110 );
nand ( n68064 , n68062 , n68063 );
nand ( n68065 , n68064 , n51766 );
nand ( n68066 , n68059 , n68065 );
xor ( n68067 , n68056 , n68066 );
xor ( n68068 , n67505 , n68067 );
not ( n68069 , n66696 );
not ( n68070 , n67677 );
or ( n68071 , n68069 , n68070 );
not ( n68072 , n61951 );
not ( n68073 , n40389 );
not ( n68074 , n68073 );
or ( n68075 , n68072 , n68074 );
nand ( n68076 , n40389 , n61952 );
nand ( n68077 , n68075 , n68076 );
nand ( n68078 , n68077 , n62654 );
nand ( n68079 , n68071 , n68078 );
not ( n68080 , n67435 );
not ( n68081 , n55144 );
or ( n68082 , n68080 , n68081 );
and ( n68083 , n40854 , n55125 );
not ( n68084 , n40854 );
and ( n68085 , n68084 , n55120 );
nor ( n68086 , n68083 , n68085 );
not ( n68087 , n68086 );
nand ( n68088 , n68087 , n54848 );
nand ( n68089 , n68082 , n68088 );
not ( n68090 , n68089 );
xor ( n68091 , n68079 , n68090 );
or ( n68092 , n67687 , n59820 );
not ( n68093 , n50306 );
not ( n68094 , n54811 );
or ( n68095 , n68093 , n68094 );
nand ( n68096 , n40364 , n50943 );
nand ( n68097 , n68095 , n68096 );
not ( n68098 , n68097 );
or ( n68099 , n68098 , n59828 );
nand ( n68100 , n68092 , n68099 );
xor ( n68101 , n68091 , n68100 );
xor ( n68102 , n68068 , n68101 );
xor ( n68103 , n67505 , n68067 );
and ( n68104 , n68103 , n68101 );
and ( n68105 , n67505 , n68067 );
or ( n68106 , n68104 , n68105 );
not ( n68107 , n52854 );
not ( n68108 , n67623 );
or ( n68109 , n68107 , n68108 );
not ( n68110 , n40733 );
not ( n68111 , n53190 );
or ( n68112 , n68110 , n68111 );
nand ( n68113 , n59179 , n53947 );
nand ( n68114 , n68112 , n68113 );
nand ( n68115 , n53571 , n68114 );
nand ( n68116 , n68109 , n68115 );
not ( n68117 , n59950 );
not ( n68118 , n67723 );
or ( n68119 , n68117 , n68118 );
not ( n68120 , n59345 );
not ( n68121 , n67193 );
or ( n68122 , n68120 , n68121 );
nand ( n68123 , n67196 , n65743 );
nand ( n68124 , n68122 , n68123 );
nand ( n68125 , n68124 , n56639 );
nand ( n68126 , n68119 , n68125 );
xor ( n68127 , n68116 , n68126 );
not ( n68128 , n62085 );
not ( n68129 , n67664 );
or ( n68130 , n68128 , n68129 );
not ( n68131 , n62077 );
not ( n68132 , n56411 );
or ( n68133 , n68131 , n68132 );
nand ( n68134 , n40452 , n60289 );
nand ( n68135 , n68133 , n68134 );
nand ( n68136 , n68135 , n60927 );
nand ( n68137 , n68130 , n68136 );
xor ( n68138 , n68127 , n68137 );
xor ( n68139 , n67857 , n68138 );
not ( n68140 , n58977 );
not ( n68141 , n60602 );
not ( n68142 , n58034 );
not ( n68143 , n68142 );
or ( n68144 , n68141 , n68143 );
not ( n68145 , n39844 );
nand ( n68146 , n68145 , n62577 );
nand ( n68147 , n68144 , n68146 );
not ( n68148 , n68147 );
or ( n68149 , n68140 , n68148 );
nand ( n68150 , n67704 , n59633 );
nand ( n68151 , n68149 , n68150 );
xor ( n68152 , n68151 , n67465 );
xor ( n68153 , n68152 , n67779 );
xor ( n68154 , n68139 , n68153 );
xor ( n68155 , n67857 , n68138 );
and ( n68156 , n68155 , n68153 );
and ( n68157 , n67857 , n68138 );
or ( n68158 , n68156 , n68157 );
xor ( n68159 , n67598 , n67958 );
not ( n68160 , n49252 );
not ( n68161 , n67511 );
or ( n68162 , n68160 , n68161 );
and ( n68163 , n49500 , n66301 );
not ( n68164 , n49500 );
and ( n68165 , n68164 , n42555 );
or ( n68166 , n68163 , n68165 );
nand ( n68167 , n68166 , n47384 );
nand ( n68168 , n68162 , n68167 );
xor ( n68169 , n68168 , n67837 );
not ( n68170 , n52962 );
not ( n68171 , n67478 );
not ( n68172 , n60855 );
or ( n68173 , n68171 , n68172 );
or ( n68174 , n60855 , n48645 );
nand ( n68175 , n68173 , n68174 );
not ( n68176 , n68175 );
or ( n68177 , n68170 , n68176 );
nand ( n68178 , n67484 , n52970 );
nand ( n68179 , n68177 , n68178 );
xor ( n68180 , n68169 , n68179 );
xor ( n68181 , n68159 , n68180 );
xor ( n68182 , n67598 , n67958 );
and ( n68183 , n68182 , n68180 );
and ( n68184 , n67598 , n67958 );
or ( n68185 , n68183 , n68184 );
not ( n68186 , n54875 );
not ( n68187 , n51723 );
not ( n68188 , n60874 );
or ( n68189 , n68187 , n68188 );
nand ( n68190 , n39056 , n53228 );
nand ( n68191 , n68189 , n68190 );
not ( n68192 , n68191 );
or ( n68193 , n68186 , n68192 );
nand ( n68194 , n67498 , n52421 );
nand ( n68195 , n68193 , n68194 );
not ( n68196 , n47407 );
not ( n68197 , n67754 );
or ( n68198 , n68196 , n68197 );
nand ( n68199 , n53675 , n54028 );
nand ( n68200 , n68198 , n68199 );
xor ( n68201 , n68195 , n68200 );
not ( n68202 , n48894 );
not ( n68203 , n67521 );
or ( n68204 , n68202 , n68203 );
not ( n68205 , n52377 );
buf ( n68206 , n60906 );
not ( n68207 , n68206 );
or ( n68208 , n68205 , n68207 );
nand ( n68209 , n39714 , n55013 );
nand ( n68210 , n68208 , n68209 );
nand ( n68211 , n68210 , n52004 );
nand ( n68212 , n68204 , n68211 );
xor ( n68213 , n68201 , n68212 );
xor ( n68214 , n67531 , n68213 );
xor ( n68215 , n68214 , n68018 );
xor ( n68216 , n67531 , n68213 );
and ( n68217 , n68216 , n68018 );
and ( n68218 , n67531 , n68213 );
or ( n68219 , n68217 , n68218 );
xor ( n68220 , n67604 , n67695 );
xor ( n68221 , n68220 , n68024 );
xor ( n68222 , n67604 , n67695 );
and ( n68223 , n68222 , n68024 );
and ( n68224 , n67604 , n67695 );
or ( n68225 , n68223 , n68224 );
xor ( n68226 , n67634 , n68030 );
xor ( n68227 , n68226 , n67763 );
xor ( n68228 , n67634 , n68030 );
and ( n68229 , n68228 , n67763 );
and ( n68230 , n67634 , n68030 );
or ( n68231 , n68229 , n68230 );
xor ( n68232 , n67995 , n68004 );
and ( n68233 , n68232 , n68015 );
and ( n68234 , n67995 , n68004 );
or ( n68235 , n68233 , n68234 );
xor ( n68236 , n67733 , n68154 );
xor ( n68237 , n68236 , n68102 );
xor ( n68238 , n67733 , n68154 );
and ( n68239 , n68238 , n68102 );
and ( n68240 , n67733 , n68154 );
or ( n68241 , n68239 , n68240 );
xor ( n68242 , n67769 , n68215 );
xor ( n68243 , n68242 , n68181 );
xor ( n68244 , n67769 , n68215 );
and ( n68245 , n68244 , n68181 );
and ( n68246 , n67769 , n68215 );
or ( n68247 , n68245 , n68246 );
xor ( n68248 , n67775 , n67791 );
xor ( n68249 , n68248 , n67785 );
xor ( n68250 , n67775 , n67791 );
and ( n68251 , n68250 , n67785 );
and ( n68252 , n67775 , n67791 );
or ( n68253 , n68251 , n68252 );
xor ( n68254 , n68221 , n68227 );
xor ( n68255 , n68254 , n68237 );
xor ( n68256 , n68221 , n68227 );
and ( n68257 , n68256 , n68237 );
and ( n68258 , n68221 , n68227 );
or ( n68259 , n68257 , n68258 );
xor ( n68260 , n67797 , n68243 );
xor ( n68261 , n68260 , n67803 );
xor ( n68262 , n67797 , n68243 );
and ( n68263 , n68262 , n67803 );
and ( n68264 , n67797 , n68243 );
or ( n68265 , n68263 , n68264 );
xor ( n68266 , n67809 , n68255 );
xor ( n68267 , n68266 , n68249 );
xor ( n68268 , n67809 , n68255 );
and ( n68269 , n68268 , n68249 );
and ( n68270 , n67809 , n68255 );
or ( n68271 , n68269 , n68270 );
xor ( n68272 , n68261 , n67815 );
xor ( n68273 , n68272 , n67821 );
xor ( n68274 , n68261 , n67815 );
and ( n68275 , n68274 , n67821 );
and ( n68276 , n68261 , n67815 );
or ( n68277 , n68275 , n68276 );
xor ( n68278 , n68267 , n68273 );
xor ( n68279 , n68278 , n67827 );
xor ( n68280 , n68267 , n68273 );
and ( n68281 , n68280 , n67827 );
and ( n68282 , n68267 , n68273 );
or ( n68283 , n68281 , n68282 );
xor ( n68284 , n67963 , n67973 );
and ( n68285 , n68284 , n67984 );
and ( n68286 , n67963 , n67973 );
or ( n68287 , n68285 , n68286 );
xor ( n68288 , n68116 , n68126 );
and ( n68289 , n68288 , n68137 );
and ( n68290 , n68116 , n68126 );
or ( n68291 , n68289 , n68290 );
xor ( n68292 , n68079 , n68090 );
and ( n68293 , n68292 , n68100 );
and ( n68294 , n68079 , n68090 );
or ( n68295 , n68293 , n68294 );
xor ( n68296 , n68044 , n68055 );
and ( n68297 , n68296 , n68066 );
and ( n68298 , n68044 , n68055 );
or ( n68299 , n68297 , n68298 );
xor ( n68300 , n68151 , n67465 );
and ( n68301 , n68300 , n67779 );
and ( n68302 , n68151 , n67465 );
or ( n68303 , n68301 , n68302 );
xor ( n68304 , n68168 , n67837 );
and ( n68305 , n68304 , n68179 );
and ( n68306 , n68168 , n67837 );
or ( n68307 , n68305 , n68306 );
xor ( n68308 , n68195 , n68200 );
and ( n68309 , n68308 , n68212 );
and ( n68310 , n68195 , n68200 );
or ( n68311 , n68309 , n68310 );
or ( n68312 , n47407 , n48929 );
nand ( n68313 , n68312 , n54028 );
not ( n68314 , n67919 );
not ( n68315 , n54316 );
or ( n68316 , n68314 , n68315 );
not ( n68317 , n56274 );
not ( n68318 , n53513 );
or ( n68319 , n68317 , n68318 );
nand ( n68320 , n55276 , n54249 );
nand ( n68321 , n68319 , n68320 );
nand ( n68322 , n68321 , n54077 );
nand ( n68323 , n68316 , n68322 );
xor ( n68324 , n68313 , n68323 );
not ( n68325 , n64452 );
not ( n68326 , n55148 );
or ( n68327 , n68325 , n68326 );
not ( n68328 , n52916 );
nand ( n68329 , n68328 , n55582 );
nand ( n68330 , n68327 , n68329 );
not ( n68331 , n68330 );
not ( n68332 , n54848 );
or ( n68333 , n68331 , n68332 );
not ( n68334 , n55576 );
or ( n68335 , n68334 , n68086 );
nand ( n68336 , n68333 , n68335 );
xor ( n68337 , n68324 , n68336 );
xor ( n68338 , n68313 , n68323 );
and ( n68339 , n68338 , n68336 );
and ( n68340 , n68313 , n68323 );
or ( n68341 , n68339 , n68340 );
not ( n68342 , n67871 );
not ( n68343 , n56281 );
or ( n68344 , n68342 , n68343 );
not ( n68345 , n49838 );
not ( n68346 , n55873 );
or ( n68347 , n68345 , n68346 );
nand ( n68348 , n56749 , n52796 );
nand ( n68349 , n68347 , n68348 );
nand ( n68350 , n68349 , n55458 );
nand ( n68351 , n68344 , n68350 );
not ( n68352 , n67881 );
not ( n68353 , n56777 );
or ( n68354 , n68352 , n68353 );
not ( n68355 , n56785 );
not ( n68356 , n52272 );
or ( n68357 , n68355 , n68356 );
nand ( n68358 , n52271 , n56758 );
nand ( n68359 , n68357 , n68358 );
nand ( n68360 , n56780 , n68359 );
nand ( n68361 , n68354 , n68360 );
xor ( n68362 , n68351 , n68361 );
or ( n68363 , n66006 , n67892 );
not ( n68364 , n41532 );
not ( n68365 , n62485 );
or ( n68366 , n68364 , n68365 );
nand ( n68367 , n57619 , n49233 );
nand ( n68368 , n68366 , n68367 );
not ( n68369 , n68368 );
or ( n68370 , n65638 , n68369 );
nand ( n68371 , n68363 , n68370 );
xor ( n68372 , n68362 , n68371 );
xor ( n68373 , n68351 , n68361 );
and ( n68374 , n68373 , n68371 );
and ( n68375 , n68351 , n68361 );
or ( n68376 , n68374 , n68375 );
not ( n68377 , n51865 );
not ( n68378 , n49707 );
not ( n68379 , n42399 );
or ( n68380 , n68378 , n68379 );
not ( n68381 , n62381 );
nand ( n68382 , n68381 , n48661 );
nand ( n68383 , n68380 , n68382 );
not ( n68384 , n68383 );
or ( n68385 , n68377 , n68384 );
nand ( n68386 , n67945 , n49713 );
nand ( n68387 , n68385 , n68386 );
not ( n68388 , n54625 );
not ( n68389 , n58482 );
or ( n68390 , n68388 , n68389 );
nand ( n68391 , n39680 , n55023 );
nand ( n68392 , n68390 , n68391 );
not ( n68393 , n68392 );
not ( n68394 , n54623 );
or ( n68395 , n68393 , n68394 );
or ( n68396 , n67037 , n54628 );
not ( n68397 , n59913 );
nand ( n68398 , n68397 , n54628 );
nand ( n68399 , n68396 , n68398 , n52022 );
nand ( n68400 , n68395 , n68399 );
xor ( n68401 , n68387 , n68400 );
xor ( n68402 , n68401 , n67899 );
xor ( n68403 , n68387 , n68400 );
and ( n68404 , n68403 , n67899 );
and ( n68405 , n68387 , n68400 );
or ( n68406 , n68404 , n68405 );
xor ( n68407 , n68287 , n68337 );
not ( n68408 , n67993 );
not ( n68409 , n61548 );
or ( n68410 , n68408 , n68409 );
not ( n68411 , n52712 );
not ( n68412 , n64633 );
or ( n68413 , n68411 , n68412 );
not ( n68414 , n63541 );
nand ( n68415 , n68414 , n54185 );
nand ( n68416 , n68413 , n68415 );
nand ( n68417 , n68416 , n61557 );
nand ( n68418 , n68410 , n68417 );
not ( n68419 , n68001 );
not ( n68420 , n62463 );
or ( n68421 , n68419 , n68420 );
not ( n68422 , n52038 );
not ( n68423 , n62449 );
or ( n68424 , n68422 , n68423 );
not ( n68425 , n62451 );
nand ( n68426 , n68425 , n52033 );
nand ( n68427 , n68424 , n68426 );
nand ( n68428 , n62467 , n68427 );
nand ( n68429 , n68421 , n68428 );
xor ( n68430 , n68418 , n68429 );
not ( n68431 , n67971 );
not ( n68432 , n65089 );
or ( n68433 , n68431 , n68432 );
not ( n68434 , n66575 );
nand ( n68435 , n68434 , n49624 );
not ( n68436 , n68435 );
nand ( n68437 , n63922 , n49630 );
not ( n68438 , n68437 );
or ( n68439 , n68436 , n68438 );
nand ( n68440 , n68439 , n65092 );
nand ( n68441 , n68433 , n68440 );
xor ( n68442 , n68430 , n68441 );
xor ( n68443 , n68407 , n68442 );
xor ( n68444 , n68287 , n68337 );
and ( n68445 , n68444 , n68442 );
and ( n68446 , n68287 , n68337 );
or ( n68447 , n68445 , n68446 );
not ( n68448 , n67908 );
not ( n68449 , n61961 );
or ( n68450 , n68448 , n68449 );
not ( n68451 , n58454 );
not ( n68452 , n58966 );
or ( n68453 , n68451 , n68452 );
nand ( n68454 , n58642 , n58459 );
nand ( n68455 , n68453 , n68454 );
nand ( n68456 , n60400 , n68455 );
nand ( n68457 , n68450 , n68456 );
not ( n68458 , n68011 );
not ( n68459 , n60539 );
or ( n68460 , n68458 , n68459 );
not ( n68461 , n47527 );
not ( n68462 , n59578 );
or ( n68463 , n68461 , n68462 );
nand ( n68464 , n62513 , n51360 );
nand ( n68465 , n68463 , n68464 );
nand ( n68466 , n68465 , n59931 );
nand ( n68467 , n68460 , n68466 );
xor ( n68468 , n68457 , n68467 );
not ( n68469 , n67930 );
not ( n68470 , n63029 );
or ( n68471 , n68469 , n68470 );
not ( n68472 , n56727 );
not ( n68473 , n66141 );
or ( n68474 , n68472 , n68473 );
nand ( n68475 , n66140 , n56731 );
nand ( n68476 , n68474 , n68475 );
nand ( n68477 , n66602 , n68476 );
nand ( n68478 , n68471 , n68477 );
xor ( n68479 , n68468 , n68478 );
xor ( n68480 , n68479 , n68372 );
xor ( n68481 , n68480 , n68291 );
xor ( n68482 , n68479 , n68372 );
and ( n68483 , n68482 , n68291 );
and ( n68484 , n68479 , n68372 );
or ( n68485 , n68483 , n68484 );
xor ( n68486 , n68295 , n68299 );
xor ( n68487 , n68486 , n68303 );
xor ( n68488 , n68295 , n68299 );
and ( n68489 , n68488 , n68303 );
and ( n68490 , n68295 , n68299 );
or ( n68491 , n68489 , n68490 );
xor ( n68492 , n68311 , n67962 );
not ( n68493 , n52125 );
not ( n68494 , n68064 );
or ( n68495 , n68493 , n68494 );
not ( n68496 , n52490 );
not ( n68497 , n53730 );
or ( n68498 , n68496 , n68497 );
not ( n68499 , n53918 );
nand ( n68500 , n68499 , n54380 );
nand ( n68501 , n68498 , n68500 );
nand ( n68502 , n68501 , n51766 );
nand ( n68503 , n68495 , n68502 );
xor ( n68504 , n68503 , n68089 );
not ( n68505 , n58977 );
not ( n68506 , n60602 );
not ( n68507 , n59417 );
not ( n68508 , n68507 );
or ( n68509 , n68506 , n68508 );
not ( n68510 , n39894 );
nand ( n68511 , n68510 , n52728 );
nand ( n68512 , n68509 , n68511 );
not ( n68513 , n68512 );
or ( n68514 , n68505 , n68513 );
nand ( n68515 , n68147 , n53104 );
nand ( n68516 , n68514 , n68515 );
xor ( n68517 , n68504 , n68516 );
xor ( n68518 , n68492 , n68517 );
xor ( n68519 , n68311 , n67962 );
and ( n68520 , n68519 , n68517 );
and ( n68521 , n68311 , n67962 );
or ( n68522 , n68520 , n68521 );
not ( n68523 , n52757 );
not ( n68524 , n50304 );
not ( n68525 , n54405 );
or ( n68526 , n68524 , n68525 );
nand ( n68527 , n56010 , n50943 );
nand ( n68528 , n68526 , n68527 );
not ( n68529 , n68528 );
or ( n68530 , n68523 , n68529 );
nand ( n68531 , n68097 , n63708 );
nand ( n68532 , n68530 , n68531 );
not ( n68533 , n51223 );
not ( n68534 , n51465 );
not ( n68535 , n40225 );
or ( n68536 , n68534 , n68535 );
nand ( n68537 , n53660 , n50916 );
nand ( n68538 , n68536 , n68537 );
not ( n68539 , n68538 );
or ( n68540 , n68533 , n68539 );
nand ( n68541 , n68042 , n52151 );
nand ( n68542 , n68540 , n68541 );
xor ( n68543 , n68532 , n68542 );
not ( n68544 , n55066 );
not ( n68545 , n65103 );
not ( n68546 , n59611 );
or ( n68547 , n68545 , n68546 );
nand ( n68548 , n59612 , n53928 );
nand ( n68549 , n68547 , n68548 );
not ( n68550 , n68549 );
or ( n68551 , n68544 , n68550 );
nand ( n68552 , n68051 , n56355 );
nand ( n68553 , n68551 , n68552 );
xor ( n68554 , n68543 , n68553 );
not ( n68555 , n53182 );
not ( n68556 , n68114 );
or ( n68557 , n68555 , n68556 );
not ( n68558 , n53190 );
not ( n68559 , n52894 );
or ( n68560 , n68558 , n68559 );
nand ( n68561 , n51601 , n53947 );
nand ( n68562 , n68560 , n68561 );
nand ( n68563 , n68562 , n52469 );
nand ( n68564 , n68557 , n68563 );
not ( n68565 , n60927 );
not ( n68566 , n66234 );
not ( n68567 , n40513 );
or ( n68568 , n68566 , n68567 );
nand ( n68569 , n56023 , n60289 );
nand ( n68570 , n68568 , n68569 );
not ( n68571 , n68570 );
or ( n68572 , n68565 , n68571 );
nand ( n68573 , n68135 , n58168 );
nand ( n68574 , n68572 , n68573 );
xor ( n68575 , n68564 , n68574 );
not ( n68576 , n62654 );
not ( n68577 , n67139 );
not ( n68578 , n59694 );
or ( n68579 , n68577 , n68578 );
nand ( n68580 , n40382 , n61952 );
nand ( n68581 , n68579 , n68580 );
not ( n68582 , n68581 );
or ( n68583 , n68576 , n68582 );
nand ( n68584 , n68077 , n62664 );
nand ( n68585 , n68583 , n68584 );
xor ( n68586 , n68575 , n68585 );
xor ( n68587 , n68554 , n68586 );
xor ( n68588 , n68587 , n68307 );
xor ( n68589 , n68554 , n68586 );
and ( n68590 , n68589 , n68307 );
and ( n68591 , n68554 , n68586 );
or ( n68592 , n68590 , n68591 );
and ( n68593 , n66155 , n47765 );
not ( n68594 , n54364 );
not ( n68595 , n53596 );
not ( n68596 , n51574 );
or ( n68597 , n68595 , n68596 );
not ( n68598 , n51574 );
nand ( n68599 , n68598 , n53591 );
nand ( n68600 , n68597 , n68599 );
not ( n68601 , n68600 );
or ( n68602 , n68594 , n68601 );
buf ( n68603 , n53956 );
nand ( n68604 , n67979 , n68603 );
nand ( n68605 , n68602 , n68604 );
xor ( n68606 , n68593 , n68605 );
not ( n68607 , n59950 );
not ( n68608 , n68124 );
or ( n68609 , n68607 , n68608 );
not ( n68610 , n59345 );
not ( n68611 , n59654 );
not ( n68612 , n68611 );
or ( n68613 , n68610 , n68612 );
nand ( n68614 , n57801 , n60617 );
nand ( n68615 , n68613 , n68614 );
nand ( n68616 , n68615 , n56639 );
nand ( n68617 , n68609 , n68616 );
xor ( n68618 , n68606 , n68617 );
xor ( n68619 , n67937 , n68235 );
not ( n68620 , n68166 );
or ( n68621 , n68620 , n48988 );
not ( n68622 , n63794 );
not ( n68623 , n47979 );
or ( n68624 , n68622 , n68623 );
nand ( n68625 , n65824 , n49500 );
nand ( n68626 , n68624 , n68625 );
not ( n68627 , n68626 );
or ( n68628 , n68627 , n53509 );
nand ( n68629 , n68621 , n68628 );
xor ( n68630 , n68619 , n68629 );
xor ( n68631 , n68618 , n68630 );
xor ( n68632 , n68631 , n68402 );
xor ( n68633 , n68618 , n68630 );
and ( n68634 , n68633 , n68402 );
and ( n68635 , n68618 , n68630 );
or ( n68636 , n68634 , n68635 );
not ( n68637 , n52970 );
not ( n68638 , n68175 );
or ( n68639 , n68637 , n68638 );
not ( n68640 , n67478 );
not ( n68641 , n39254 );
or ( n68642 , n68640 , n68641 );
buf ( n68643 , n39253 );
nand ( n68644 , n68643 , n52048 );
nand ( n68645 , n68642 , n68644 );
nand ( n68646 , n68645 , n52962 );
nand ( n68647 , n68639 , n68646 );
not ( n68648 , n52421 );
not ( n68649 , n68191 );
or ( n68650 , n68648 , n68649 );
not ( n68651 , n51723 );
not ( n68652 , n38499 );
not ( n68653 , n68652 );
or ( n68654 , n68651 , n68653 );
not ( n68655 , n62394 );
nand ( n68656 , n68655 , n51724 );
nand ( n68657 , n68654 , n68656 );
nand ( n68658 , n68657 , n54875 );
nand ( n68659 , n68650 , n68658 );
xor ( n68660 , n68647 , n68659 );
not ( n68661 , n57314 );
not ( n68662 , n68210 );
or ( n68663 , n68661 , n68662 );
not ( n68664 , n52377 );
not ( n68665 , n59399 );
or ( n68666 , n68664 , n68665 );
not ( n68667 , n65532 );
nand ( n68668 , n68667 , n55013 );
nand ( n68669 , n68666 , n68668 );
nand ( n68670 , n68669 , n52004 );
nand ( n68671 , n68663 , n68670 );
xor ( n68672 , n68660 , n68671 );
xor ( n68673 , n68022 , n68672 );
xor ( n68674 , n68673 , n68481 );
xor ( n68675 , n68022 , n68672 );
and ( n68676 , n68675 , n68481 );
and ( n68677 , n68022 , n68672 );
or ( n68678 , n68676 , n68677 );
xor ( n68679 , n68028 , n68443 );
xor ( n68680 , n68679 , n68487 );
xor ( n68681 , n68028 , n68443 );
and ( n68682 , n68681 , n68487 );
and ( n68683 , n68028 , n68443 );
or ( n68684 , n68682 , n68683 );
xor ( n68685 , n68034 , n68106 );
xor ( n68686 , n68685 , n68185 );
xor ( n68687 , n68034 , n68106 );
and ( n68688 , n68687 , n68185 );
and ( n68689 , n68034 , n68106 );
or ( n68690 , n68688 , n68689 );
xor ( n68691 , n68457 , n68467 );
and ( n68692 , n68691 , n68478 );
and ( n68693 , n68457 , n68467 );
or ( n68694 , n68692 , n68693 );
xor ( n68695 , n68588 , n68158 );
xor ( n68696 , n68695 , n68518 );
xor ( n68697 , n68588 , n68158 );
and ( n68698 , n68697 , n68518 );
and ( n68699 , n68588 , n68158 );
or ( n68700 , n68698 , n68699 );
xor ( n68701 , n68674 , n68219 );
xor ( n68702 , n68701 , n68632 );
xor ( n68703 , n68674 , n68219 );
and ( n68704 , n68703 , n68632 );
and ( n68705 , n68674 , n68219 );
or ( n68706 , n68704 , n68705 );
xor ( n68707 , n68225 , n68680 );
xor ( n68708 , n68707 , n68241 );
xor ( n68709 , n68225 , n68680 );
and ( n68710 , n68709 , n68241 );
and ( n68711 , n68225 , n68680 );
or ( n68712 , n68710 , n68711 );
xor ( n68713 , n68686 , n68231 );
xor ( n68714 , n68713 , n68696 );
xor ( n68715 , n68686 , n68231 );
and ( n68716 , n68715 , n68696 );
and ( n68717 , n68686 , n68231 );
or ( n68718 , n68716 , n68717 );
xor ( n68719 , n68247 , n68702 );
xor ( n68720 , n68719 , n68253 );
xor ( n68721 , n68247 , n68702 );
and ( n68722 , n68721 , n68253 );
and ( n68723 , n68247 , n68702 );
or ( n68724 , n68722 , n68723 );
xor ( n68725 , n68708 , n68259 );
xor ( n68726 , n68725 , n68714 );
xor ( n68727 , n68708 , n68259 );
and ( n68728 , n68727 , n68714 );
and ( n68729 , n68708 , n68259 );
or ( n68730 , n68728 , n68729 );
xor ( n68731 , n68720 , n68265 );
xor ( n68732 , n68731 , n68271 );
xor ( n68733 , n68720 , n68265 );
and ( n68734 , n68733 , n68271 );
and ( n68735 , n68720 , n68265 );
or ( n68736 , n68734 , n68735 );
xor ( n68737 , n68726 , n68732 );
xor ( n68738 , n68737 , n68277 );
xor ( n68739 , n68726 , n68732 );
and ( n68740 , n68739 , n68277 );
and ( n68741 , n68726 , n68732 );
or ( n68742 , n68740 , n68741 );
xor ( n68743 , n68418 , n68429 );
and ( n68744 , n68743 , n68441 );
and ( n68745 , n68418 , n68429 );
or ( n68746 , n68744 , n68745 );
xor ( n68747 , n68593 , n68605 );
and ( n68748 , n68747 , n68617 );
and ( n68749 , n68593 , n68605 );
or ( n68750 , n68748 , n68749 );
xor ( n68751 , n68564 , n68574 );
and ( n68752 , n68751 , n68585 );
and ( n68753 , n68564 , n68574 );
or ( n68754 , n68752 , n68753 );
xor ( n68755 , n68532 , n68542 );
and ( n68756 , n68755 , n68553 );
and ( n68757 , n68532 , n68542 );
or ( n68758 , n68756 , n68757 );
xor ( n68759 , n68503 , n68089 );
and ( n68760 , n68759 , n68516 );
and ( n68761 , n68503 , n68089 );
or ( n68762 , n68760 , n68761 );
xor ( n68763 , n67937 , n68235 );
and ( n68764 , n68763 , n68629 );
and ( n68765 , n67937 , n68235 );
or ( n68766 , n68764 , n68765 );
xor ( n68767 , n68647 , n68659 );
and ( n68768 , n68767 , n68671 );
and ( n68769 , n68647 , n68659 );
or ( n68770 , n68768 , n68769 );
not ( n68771 , n68359 );
not ( n68772 , n56776 );
or ( n68773 , n68771 , n68772 );
not ( n68774 , n49001 );
not ( n68775 , n56785 );
or ( n68776 , n68774 , n68775 );
nand ( n68777 , n52589 , n59045 );
nand ( n68778 , n68776 , n68777 );
nand ( n68779 , n56780 , n68778 );
nand ( n68780 , n68773 , n68779 );
not ( n68781 , n68368 );
not ( n68782 , n66005 );
or ( n68783 , n68781 , n68782 );
not ( n68784 , n65969 );
not ( n68785 , n62485 );
or ( n68786 , n68784 , n68785 );
nand ( n68787 , n57619 , n50084 );
nand ( n68788 , n68786 , n68787 );
nand ( n68789 , n57631 , n68788 );
nand ( n68790 , n68783 , n68789 );
xor ( n68791 , n68780 , n68790 );
not ( n68792 , n68455 );
not ( n68793 , n63080 );
or ( n68794 , n68792 , n68793 );
not ( n68795 , n58915 );
not ( n68796 , n62497 );
or ( n68797 , n68795 , n68796 );
nand ( n68798 , n65652 , n66946 );
nand ( n68799 , n68797 , n68798 );
nand ( n68800 , n61465 , n68799 );
nand ( n68801 , n68794 , n68800 );
xor ( n68802 , n68791 , n68801 );
xor ( n68803 , n68780 , n68790 );
and ( n68804 , n68803 , n68801 );
and ( n68805 , n68780 , n68790 );
or ( n68806 , n68804 , n68805 );
not ( n68807 , n68465 );
not ( n68808 , n60539 );
or ( n68809 , n68807 , n68808 );
not ( n68810 , n59574 );
not ( n68811 , n58994 );
not ( n68812 , n63587 );
or ( n68813 , n68811 , n68812 );
nand ( n68814 , n59338 , n58179 );
nand ( n68815 , n68813 , n68814 );
nand ( n68816 , n68810 , n68815 );
nand ( n68817 , n68809 , n68816 );
not ( n68818 , n68330 );
not ( n68819 , n55144 );
or ( n68820 , n68818 , n68819 );
not ( n68821 , n66226 );
not ( n68822 , n55119 );
or ( n68823 , n68821 , n68822 );
not ( n68824 , n65216 );
nand ( n68825 , n68824 , n55152 );
nand ( n68826 , n68823 , n68825 );
nand ( n68827 , n68826 , n55934 );
nand ( n68828 , n68820 , n68827 );
xor ( n68829 , n68817 , n68828 );
not ( n68830 , n68416 );
not ( n68831 , n64111 );
or ( n68832 , n68830 , n68831 );
not ( n68833 , n48983 );
not ( n68834 , n66616 );
or ( n68835 , n68833 , n68834 );
nand ( n68836 , n66615 , n56348 );
nand ( n68837 , n68835 , n68836 );
nand ( n68838 , n68837 , n61558 );
nand ( n68839 , n68832 , n68838 );
xor ( n68840 , n68829 , n68839 );
xor ( n68841 , n68817 , n68828 );
and ( n68842 , n68841 , n68839 );
and ( n68843 , n68817 , n68828 );
or ( n68844 , n68842 , n68843 );
xor ( n68845 , n68341 , n68376 );
not ( n68846 , n68427 );
not ( n68847 , n62463 );
or ( n68848 , n68846 , n68847 );
not ( n68849 , n62449 );
not ( n68850 , n51670 );
and ( n68851 , n68849 , n68850 );
and ( n68852 , n62451 , n51670 );
nor ( n68853 , n68851 , n68852 );
not ( n68854 , n68853 );
nand ( n68855 , n68854 , n67068 );
nand ( n68856 , n68848 , n68855 );
not ( n68857 , n49624 );
not ( n68858 , n64443 );
or ( n68859 , n68857 , n68858 );
nand ( n68860 , n68859 , n68437 );
not ( n68861 , n68860 );
not ( n68862 , n65089 );
or ( n68863 , n68861 , n68862 );
not ( n68864 , n51792 );
not ( n68865 , n63415 );
or ( n68866 , n68864 , n68865 );
nand ( n68867 , n63922 , n48829 );
nand ( n68868 , n68866 , n68867 );
nand ( n68869 , n68868 , n65092 );
nand ( n68870 , n68863 , n68869 );
xor ( n68871 , n68856 , n68870 );
not ( n68872 , n68476 );
not ( n68873 , n66136 );
or ( n68874 , n68872 , n68873 );
not ( n68875 , n57182 );
not ( n68876 , n67084 );
or ( n68877 , n68875 , n68876 );
not ( n68878 , n60286 );
nand ( n68879 , n68878 , n58195 );
nand ( n68880 , n68877 , n68879 );
nand ( n68881 , n60427 , n68880 );
nand ( n68882 , n68874 , n68881 );
xor ( n68883 , n68871 , n68882 );
xor ( n68884 , n68845 , n68883 );
xor ( n68885 , n68341 , n68376 );
and ( n68886 , n68885 , n68883 );
and ( n68887 , n68341 , n68376 );
or ( n68888 , n68886 , n68887 );
xor ( n68889 , n68840 , n68802 );
xor ( n68890 , n68889 , n68750 );
xor ( n68891 , n68840 , n68802 );
and ( n68892 , n68891 , n68750 );
and ( n68893 , n68840 , n68802 );
or ( n68894 , n68892 , n68893 );
xor ( n68895 , n68754 , n68758 );
and ( n68896 , n66581 , n51204 );
not ( n68897 , n54327 );
and ( n68898 , n40691 , n54322 );
not ( n68899 , n40691 );
and ( n68900 , n68899 , n59078 );
or ( n68901 , n68898 , n68900 );
not ( n68902 , n68901 );
or ( n68903 , n68897 , n68902 );
not ( n68904 , n55161 );
nand ( n68905 , n68904 , n68321 );
nand ( n68906 , n68903 , n68905 );
xor ( n68907 , n68896 , n68906 );
not ( n68908 , n53956 );
not ( n68909 , n68600 );
or ( n68910 , n68908 , n68909 );
not ( n68911 , n53615 );
not ( n68912 , n53259 );
or ( n68913 , n68911 , n68912 );
nand ( n68914 , n54032 , n53591 );
nand ( n68915 , n68913 , n68914 );
nand ( n68916 , n68915 , n53620 );
nand ( n68917 , n68910 , n68916 );
xor ( n68918 , n68907 , n68917 );
xor ( n68919 , n68895 , n68918 );
xor ( n68920 , n68754 , n68758 );
and ( n68921 , n68920 , n68918 );
and ( n68922 , n68754 , n68758 );
or ( n68923 , n68921 , n68922 );
xor ( n68924 , n68762 , n68766 );
xor ( n68925 , n68924 , n68770 );
xor ( n68926 , n68762 , n68766 );
and ( n68927 , n68926 , n68770 );
and ( n68928 , n68762 , n68766 );
or ( n68929 , n68927 , n68928 );
not ( n68930 , n51766 );
not ( n68931 , n52130 );
not ( n68932 , n68931 );
not ( n68933 , n53271 );
or ( n68934 , n68932 , n68933 );
nand ( n68935 , n40626 , n52110 );
nand ( n68936 , n68934 , n68935 );
not ( n68937 , n68936 );
or ( n68938 , n68930 , n68937 );
nand ( n68939 , n68501 , n52482 );
nand ( n68940 , n68938 , n68939 );
not ( n68941 , n52854 );
not ( n68942 , n68562 );
or ( n68943 , n68941 , n68942 );
not ( n68944 , n52841 );
not ( n68945 , n40527 );
or ( n68946 , n68944 , n68945 );
nand ( n68947 , n51912 , n52980 );
nand ( n68948 , n68946 , n68947 );
nand ( n68949 , n68948 , n53571 );
nand ( n68950 , n68943 , n68949 );
xor ( n68951 , n68940 , n68950 );
not ( n68952 , n59950 );
not ( n68953 , n68615 );
or ( n68954 , n68952 , n68953 );
not ( n68955 , n59345 );
not ( n68956 , n39844 );
or ( n68957 , n68955 , n68956 );
nand ( n68958 , n68145 , n60617 );
nand ( n68959 , n68957 , n68958 );
not ( n68960 , n68959 );
not ( n68961 , n56639 );
or ( n68962 , n68960 , n68961 );
nand ( n68963 , n68954 , n68962 );
xor ( n68964 , n68951 , n68963 );
xor ( n68965 , n68406 , n68964 );
not ( n68966 , n58168 );
not ( n68967 , n68570 );
or ( n68968 , n68966 , n68967 );
not ( n68969 , n62077 );
not ( n68970 , n63180 );
or ( n68971 , n68969 , n68970 );
nand ( n68972 , n67196 , n60292 );
nand ( n68973 , n68971 , n68972 );
nand ( n68974 , n68973 , n60927 );
nand ( n68975 , n68968 , n68974 );
not ( n68976 , n62654 );
not ( n68977 , n61951 );
not ( n68978 , n55630 );
or ( n68979 , n68977 , n68978 );
not ( n68980 , n56407 );
nand ( n68981 , n68980 , n61952 );
nand ( n68982 , n68979 , n68981 );
not ( n68983 , n68982 );
or ( n68984 , n68976 , n68983 );
nand ( n68985 , n68581 , n66696 );
nand ( n68986 , n68984 , n68985 );
xor ( n68987 , n68975 , n68986 );
not ( n68988 , n52757 );
not ( n68989 , n64190 );
buf ( n68990 , n55645 );
not ( n68991 , n68990 );
not ( n68992 , n68991 );
or ( n68993 , n68989 , n68992 );
not ( n68994 , n68073 );
nand ( n68995 , n68994 , n66705 );
nand ( n68996 , n68993 , n68995 );
not ( n68997 , n68996 );
or ( n68998 , n68988 , n68997 );
nand ( n68999 , n68528 , n63708 );
nand ( n69000 , n68998 , n68999 );
xor ( n69001 , n68987 , n69000 );
xor ( n69002 , n68965 , n69001 );
xor ( n69003 , n68406 , n68964 );
and ( n69004 , n69003 , n69001 );
and ( n69005 , n68406 , n68964 );
or ( n69006 , n69004 , n69005 );
not ( n69007 , n50922 );
not ( n69008 , n65773 );
not ( n69009 , n66236 );
or ( n69010 , n69008 , n69009 );
nand ( n69011 , n63204 , n52781 );
nand ( n69012 , n69010 , n69011 );
not ( n69013 , n69012 );
or ( n69014 , n69007 , n69013 );
nand ( n69015 , n68538 , n52151 );
nand ( n69016 , n69014 , n69015 );
not ( n69017 , n56355 );
not ( n69018 , n68549 );
or ( n69019 , n69017 , n69018 );
not ( n69020 , n53931 );
not ( n69021 , n56476 );
or ( n69022 , n69020 , n69021 );
nand ( n69023 , n63217 , n53928 );
nand ( n69024 , n69022 , n69023 );
nand ( n69025 , n69024 , n51533 );
nand ( n69026 , n69019 , n69025 );
xor ( n69027 , n69016 , n69026 );
not ( n69028 , n55887 );
not ( n69029 , n68349 );
or ( n69030 , n69028 , n69029 );
not ( n69031 , n40855 );
not ( n69032 , n55872 );
or ( n69033 , n69031 , n69032 );
not ( n69034 , n55892 );
nand ( n69035 , n69034 , n56239 );
nand ( n69036 , n69033 , n69035 );
not ( n69037 , n69036 );
or ( n69038 , n69037 , n58066 );
nand ( n69039 , n69030 , n69038 );
not ( n69040 , n69039 );
xor ( n69041 , n69027 , n69040 );
xor ( n69042 , n69041 , n68884 );
xor ( n69043 , n69042 , n68447 );
xor ( n69044 , n69041 , n68884 );
and ( n69045 , n69044 , n68447 );
and ( n69046 , n69041 , n68884 );
or ( n69047 , n69045 , n69046 );
xor ( n69048 , n68694 , n68746 );
not ( n69049 , n49713 );
not ( n69050 , n68383 );
or ( n69051 , n69049 , n69050 );
not ( n69052 , n52267 );
not ( n69053 , n67269 );
or ( n69054 , n69052 , n69053 );
nand ( n69055 , n42555 , n51351 );
nand ( n69056 , n69054 , n69055 );
nand ( n69057 , n69056 , n51865 );
nand ( n69058 , n69051 , n69057 );
xor ( n69059 , n69048 , n69058 );
not ( n69060 , n54875 );
not ( n69061 , n51723 );
not ( n69062 , n60855 );
or ( n69063 , n69061 , n69062 );
nand ( n69064 , n62963 , n51724 );
nand ( n69065 , n69063 , n69064 );
not ( n69066 , n69065 );
or ( n69067 , n69060 , n69066 );
nand ( n69068 , n68657 , n52421 );
nand ( n69069 , n69067 , n69068 );
not ( n69070 , n52004 );
not ( n69071 , n52377 );
not ( n69072 , n39056 );
not ( n69073 , n69072 );
or ( n69074 , n69071 , n69073 );
nand ( n69075 , n39056 , n55013 );
nand ( n69076 , n69074 , n69075 );
not ( n69077 , n69076 );
or ( n69078 , n69070 , n69077 );
nand ( n69079 , n68669 , n57314 );
nand ( n69080 , n69078 , n69079 );
xor ( n69081 , n69069 , n69080 );
not ( n69082 , n59633 );
not ( n69083 , n68512 );
or ( n69084 , n69082 , n69083 );
not ( n69085 , n58982 );
not ( n69086 , n67040 );
or ( n69087 , n69085 , n69086 );
nand ( n69088 , n59913 , n62577 );
nand ( n69089 , n69087 , n69088 );
nand ( n69090 , n69089 , n58977 );
nand ( n69091 , n69084 , n69090 );
xor ( n69092 , n69081 , n69091 );
xor ( n69093 , n69059 , n69092 );
not ( n69094 , n48989 );
not ( n69095 , n68626 );
or ( n69096 , n69094 , n69095 );
nand ( n69097 , n47384 , n49500 );
nand ( n69098 , n69096 , n69097 );
not ( n69099 , n54623 );
not ( n69100 , n59174 );
not ( n69101 , n60906 );
or ( n69102 , n69100 , n69101 );
nand ( n69103 , n39714 , n54628 );
nand ( n69104 , n69102 , n69103 );
not ( n69105 , n69104 );
or ( n69106 , n69099 , n69105 );
nand ( n69107 , n52022 , n68392 );
nand ( n69108 , n69106 , n69107 );
xor ( n69109 , n69098 , n69108 );
not ( n69110 , n52970 );
not ( n69111 , n68645 );
or ( n69112 , n69110 , n69111 );
not ( n69113 , n67478 );
not ( n69114 , n66052 );
or ( n69115 , n69113 , n69114 );
nand ( n69116 , n61907 , n67477 );
nand ( n69117 , n69115 , n69116 );
nand ( n69118 , n69117 , n52962 );
nand ( n69119 , n69112 , n69118 );
xor ( n69120 , n69109 , n69119 );
xor ( n69121 , n69093 , n69120 );
xor ( n69122 , n69059 , n69092 );
and ( n69123 , n69122 , n69120 );
and ( n69124 , n69059 , n69092 );
or ( n69125 , n69123 , n69124 );
xor ( n69126 , n68890 , n68485 );
xor ( n69127 , n69126 , n68491 );
xor ( n69128 , n68890 , n68485 );
and ( n69129 , n69128 , n68491 );
and ( n69130 , n68890 , n68485 );
or ( n69131 , n69129 , n69130 );
xor ( n69132 , n68919 , n68522 );
xor ( n69133 , n69132 , n68592 );
xor ( n69134 , n68919 , n68522 );
and ( n69135 , n69134 , n68592 );
and ( n69136 , n68919 , n68522 );
or ( n69137 , n69135 , n69136 );
xor ( n69138 , n68925 , n69002 );
xor ( n69139 , n69138 , n68636 );
xor ( n69140 , n68925 , n69002 );
and ( n69141 , n69140 , n68636 );
and ( n69142 , n68925 , n69002 );
or ( n69143 , n69141 , n69142 );
xor ( n69144 , n68856 , n68870 );
and ( n69145 , n69144 , n68882 );
and ( n69146 , n68856 , n68870 );
or ( n69147 , n69145 , n69146 );
xor ( n69148 , n68678 , n69121 );
xor ( n69149 , n69148 , n69043 );
xor ( n69150 , n68678 , n69121 );
and ( n69151 , n69150 , n69043 );
and ( n69152 , n68678 , n69121 );
or ( n69153 , n69151 , n69152 );
xor ( n69154 , n68684 , n69127 );
xor ( n69155 , n69154 , n68690 );
xor ( n69156 , n68684 , n69127 );
and ( n69157 , n69156 , n68690 );
and ( n69158 , n68684 , n69127 );
or ( n69159 , n69157 , n69158 );
xor ( n69160 , n69133 , n68700 );
xor ( n69161 , n69160 , n69139 );
xor ( n69162 , n69133 , n68700 );
and ( n69163 , n69162 , n69139 );
and ( n69164 , n69133 , n68700 );
or ( n69165 , n69163 , n69164 );
xor ( n69166 , n68706 , n69149 );
xor ( n69167 , n69166 , n68712 );
xor ( n69168 , n68706 , n69149 );
and ( n69169 , n69168 , n68712 );
and ( n69170 , n68706 , n69149 );
or ( n69171 , n69169 , n69170 );
xor ( n69172 , n69155 , n69161 );
xor ( n69173 , n69172 , n68718 );
xor ( n69174 , n69155 , n69161 );
and ( n69175 , n69174 , n68718 );
and ( n69176 , n69155 , n69161 );
or ( n69177 , n69175 , n69176 );
xor ( n69178 , n68724 , n69167 );
xor ( n69179 , n69178 , n68730 );
xor ( n69180 , n68724 , n69167 );
and ( n69181 , n69180 , n68730 );
and ( n69182 , n68724 , n69167 );
or ( n69183 , n69181 , n69182 );
xor ( n69184 , n69173 , n69179 );
xor ( n69185 , n69184 , n68736 );
xor ( n69186 , n69173 , n69179 );
and ( n69187 , n69186 , n68736 );
and ( n69188 , n69173 , n69179 );
or ( n69189 , n69187 , n69188 );
xor ( n69190 , n68896 , n68906 );
and ( n69191 , n69190 , n68917 );
and ( n69192 , n68896 , n68906 );
or ( n69193 , n69191 , n69192 );
xor ( n69194 , n68975 , n68986 );
and ( n69195 , n69194 , n69000 );
and ( n69196 , n68975 , n68986 );
or ( n69197 , n69195 , n69196 );
xor ( n69198 , n69016 , n69026 );
and ( n69199 , n69198 , n69040 );
and ( n69200 , n69016 , n69026 );
or ( n69201 , n69199 , n69200 );
xor ( n69202 , n68940 , n68950 );
and ( n69203 , n69202 , n68963 );
and ( n69204 , n68940 , n68950 );
or ( n69205 , n69203 , n69204 );
xor ( n69206 , n68694 , n68746 );
and ( n69207 , n69206 , n69058 );
and ( n69208 , n68694 , n68746 );
or ( n69209 , n69207 , n69208 );
xor ( n69210 , n69069 , n69080 );
and ( n69211 , n69210 , n69091 );
and ( n69212 , n69069 , n69080 );
or ( n69213 , n69211 , n69212 );
xor ( n69214 , n69098 , n69108 );
and ( n69215 , n69214 , n69119 );
and ( n69216 , n69098 , n69108 );
or ( n69217 , n69215 , n69216 );
not ( n69218 , n53509 );
not ( n69219 , n48988 );
or ( n69220 , n69218 , n69219 );
nand ( n69221 , n69220 , n49500 );
not ( n69222 , n68826 );
not ( n69223 , n55576 );
or ( n69224 , n69222 , n69223 );
not ( n69225 , n55582 );
not ( n69226 , n52076 );
or ( n69227 , n69225 , n69226 );
nand ( n69228 , n55125 , n50404 );
nand ( n69229 , n69227 , n69228 );
nand ( n69230 , n69229 , n55934 );
nand ( n69231 , n69224 , n69230 );
xor ( n69232 , n69221 , n69231 );
not ( n69233 , n69036 );
not ( n69234 , n56281 );
or ( n69235 , n69233 , n69234 );
not ( n69236 , n52916 );
not ( n69237 , n55891 );
not ( n69238 , n69237 );
or ( n69239 , n69236 , n69238 );
nand ( n69240 , n55872 , n64451 );
nand ( n69241 , n69239 , n69240 );
nand ( n69242 , n69241 , n59984 );
nand ( n69243 , n69235 , n69242 );
xor ( n69244 , n69232 , n69243 );
xor ( n69245 , n69221 , n69231 );
and ( n69246 , n69245 , n69243 );
and ( n69247 , n69221 , n69231 );
or ( n69248 , n69246 , n69247 );
not ( n69249 , n68778 );
or ( n69250 , n65594 , n69249 );
and ( n69251 , n57665 , n57571 );
and ( n69252 , n49837 , n61518 );
nor ( n69253 , n69251 , n69252 );
or ( n69254 , n65166 , n69253 );
nand ( n69255 , n69250 , n69254 );
not ( n69256 , n68788 );
not ( n69257 , n66005 );
or ( n69258 , n69256 , n69257 );
not ( n69259 , n57619 );
not ( n69260 , n48679 );
and ( n69261 , n69259 , n69260 );
and ( n69262 , n65175 , n48679 );
nor ( n69263 , n69261 , n69262 );
not ( n69264 , n69263 );
nand ( n69265 , n69264 , n57631 );
nand ( n69266 , n69258 , n69265 );
xor ( n69267 , n69255 , n69266 );
not ( n69268 , n68799 );
or ( n69269 , n64143 , n69268 );
not ( n69270 , n41532 );
and ( n69271 , n69270 , n65184 );
not ( n69272 , n69270 );
and ( n69273 , n69272 , n62497 );
nor ( n69274 , n69271 , n69273 );
or ( n69275 , n69274 , n64146 );
nand ( n69276 , n69269 , n69275 );
xor ( n69277 , n69267 , n69276 );
xor ( n69278 , n69255 , n69266 );
and ( n69279 , n69278 , n69276 );
and ( n69280 , n69255 , n69266 );
or ( n69281 , n69279 , n69280 );
xor ( n69282 , n68806 , n68844 );
xor ( n69283 , n69282 , n69244 );
xor ( n69284 , n68806 , n68844 );
and ( n69285 , n69284 , n69244 );
and ( n69286 , n68806 , n68844 );
or ( n69287 , n69285 , n69286 );
or ( n69288 , n64684 , n68853 );
and ( n69289 , n64167 , n54185 );
and ( n69290 , n62451 , n52712 );
nor ( n69291 , n69289 , n69290 );
or ( n69292 , n64166 , n69291 );
nand ( n69293 , n69288 , n69292 );
not ( n69294 , n68868 );
not ( n69295 , n66569 );
or ( n69296 , n69294 , n69295 );
not ( n69297 , n52033 );
not ( n69298 , n63415 );
or ( n69299 , n69297 , n69298 );
nand ( n69300 , n63922 , n55959 );
nand ( n69301 , n69299 , n69300 );
nand ( n69302 , n65092 , n69301 );
nand ( n69303 , n69296 , n69302 );
xor ( n69304 , n69293 , n69303 );
not ( n69305 , n63412 );
and ( n69306 , n69305 , n49624 );
xor ( n69307 , n69304 , n69306 );
not ( n69308 , n68815 );
not ( n69309 , n62506 );
or ( n69310 , n69308 , n69309 );
not ( n69311 , n58458 );
not ( n69312 , n65121 );
or ( n69313 , n69311 , n69312 );
not ( n69314 , n63587 );
nand ( n69315 , n69314 , n58459 );
nand ( n69316 , n69313 , n69315 );
nand ( n69317 , n59575 , n69316 );
nand ( n69318 , n69310 , n69317 );
not ( n69319 , n68880 );
not ( n69320 , n65130 );
or ( n69321 , n69319 , n69320 );
not ( n69322 , n47527 );
not ( n69323 , n66141 );
or ( n69324 , n69322 , n69323 );
nand ( n69325 , n66140 , n64603 );
nand ( n69326 , n69324 , n69325 );
nand ( n69327 , n60427 , n69326 );
nand ( n69328 , n69321 , n69327 );
xor ( n69329 , n69318 , n69328 );
not ( n69330 , n68837 );
not ( n69331 , n64111 );
or ( n69332 , n69330 , n69331 );
not ( n69333 , n66615 );
and ( n69334 , n56727 , n69333 );
not ( n69335 , n56727 );
and ( n69336 , n69335 , n66615 );
or ( n69337 , n69334 , n69336 );
nand ( n69338 , n62428 , n69337 );
nand ( n69339 , n69332 , n69338 );
xor ( n69340 , n69329 , n69339 );
xor ( n69341 , n69307 , n69340 );
xor ( n69342 , n69341 , n69277 );
xor ( n69343 , n69307 , n69340 );
and ( n69344 , n69343 , n69277 );
and ( n69345 , n69307 , n69340 );
or ( n69346 , n69344 , n69345 );
xor ( n69347 , n69193 , n69197 );
xor ( n69348 , n69347 , n69201 );
xor ( n69349 , n69193 , n69197 );
and ( n69350 , n69349 , n69201 );
and ( n69351 , n69193 , n69197 );
or ( n69352 , n69350 , n69351 );
xor ( n69353 , n69205 , n69209 );
xor ( n69354 , n69353 , n69213 );
xor ( n69355 , n69205 , n69209 );
and ( n69356 , n69355 , n69213 );
and ( n69357 , n69205 , n69209 );
or ( n69358 , n69356 , n69357 );
not ( n69359 , n52139 );
not ( n69360 , n69024 );
or ( n69361 , n69359 , n69360 );
not ( n69362 , n51146 );
not ( n69363 , n65103 );
not ( n69364 , n40225 );
or ( n69365 , n69363 , n69364 );
or ( n69366 , n40225 , n65103 );
nand ( n69367 , n69365 , n69366 );
nand ( n69368 , n69362 , n69367 );
nand ( n69369 , n69361 , n69368 );
not ( n69370 , n51766 );
and ( n69371 , n54415 , n52114 );
not ( n69372 , n54415 );
and ( n69373 , n69372 , n52110 );
or ( n69374 , n69371 , n69373 );
not ( n69375 , n69374 );
or ( n69376 , n69370 , n69375 );
nand ( n69377 , n53197 , n68936 );
nand ( n69378 , n69376 , n69377 );
xor ( n69379 , n69369 , n69378 );
xor ( n69380 , n69379 , n69039 );
xor ( n69381 , n69217 , n69380 );
not ( n69382 , n66696 );
not ( n69383 , n68982 );
or ( n69384 , n69382 , n69383 );
not ( n69385 , n61951 );
not ( n69386 , n56020 );
or ( n69387 , n69385 , n69386 );
nand ( n69388 , n56023 , n61952 );
nand ( n69389 , n69387 , n69388 );
nand ( n69390 , n69389 , n62654 );
nand ( n69391 , n69384 , n69390 );
not ( n69392 , n63708 );
not ( n69393 , n68996 );
or ( n69394 , n69392 , n69393 );
not ( n69395 , n50304 );
not ( n69396 , n65725 );
or ( n69397 , n69395 , n69396 );
nand ( n69398 , n55203 , n66705 );
nand ( n69399 , n69397 , n69398 );
nand ( n69400 , n69399 , n52757 );
nand ( n69401 , n69394 , n69400 );
xor ( n69402 , n69391 , n69401 );
not ( n69403 , n52151 );
not ( n69404 , n69012 );
or ( n69405 , n69403 , n69404 );
not ( n69406 , n65773 );
not ( n69407 , n54402 );
or ( n69408 , n69406 , n69407 );
not ( n69409 , n62626 );
nand ( n69410 , n69409 , n67639 );
nand ( n69411 , n69408 , n69410 );
nand ( n69412 , n50922 , n69411 );
nand ( n69413 , n69405 , n69412 );
xor ( n69414 , n69402 , n69413 );
xor ( n69415 , n69381 , n69414 );
xor ( n69416 , n69217 , n69380 );
and ( n69417 , n69416 , n69414 );
and ( n69418 , n69217 , n69380 );
or ( n69419 , n69417 , n69418 );
not ( n69420 , n54327 );
not ( n69421 , n54298 );
not ( n69422 , n52285 );
or ( n69423 , n69421 , n69422 );
nand ( n69424 , n40677 , n54322 );
nand ( n69425 , n69423 , n69424 );
not ( n69426 , n69425 );
or ( n69427 , n69420 , n69426 );
nand ( n69428 , n68901 , n54316 );
nand ( n69429 , n69427 , n69428 );
not ( n69430 , n62085 );
not ( n69431 , n68973 );
or ( n69432 , n69430 , n69431 );
not ( n69433 , n62077 );
not ( n69434 , n57798 );
or ( n69435 , n69433 , n69434 );
nand ( n69436 , n59654 , n60292 );
nand ( n69437 , n69435 , n69436 );
nand ( n69438 , n69437 , n60927 );
nand ( n69439 , n69432 , n69438 );
xor ( n69440 , n69429 , n69439 );
not ( n69441 , n53620 );
buf ( n69442 , n52893 );
not ( n69443 , n69442 );
not ( n69444 , n53596 );
not ( n69445 , n69444 );
or ( n69446 , n69443 , n69445 );
nand ( n69447 , n53615 , n52222 );
nand ( n69448 , n69446 , n69447 );
not ( n69449 , n69448 );
or ( n69450 , n69441 , n69449 );
nand ( n69451 , n68915 , n68603 );
nand ( n69452 , n69450 , n69451 );
xor ( n69453 , n69440 , n69452 );
xor ( n69454 , n69453 , n69283 );
not ( n69455 , n52854 );
not ( n69456 , n68948 );
or ( n69457 , n69455 , n69456 );
not ( n69458 , n55104 );
not ( n69459 , n69458 );
not ( n69460 , n54377 );
or ( n69461 , n69459 , n69460 );
nand ( n69462 , n54380 , n52837 );
nand ( n69463 , n69461 , n69462 );
nand ( n69464 , n69463 , n53571 );
nand ( n69465 , n69457 , n69464 );
not ( n69466 , n59950 );
not ( n69467 , n68959 );
or ( n69468 , n69466 , n69467 );
not ( n69469 , n59345 );
not ( n69470 , n39894 );
or ( n69471 , n69469 , n69470 );
nand ( n69472 , n59413 , n60617 );
nand ( n69473 , n69471 , n69472 );
nand ( n69474 , n69473 , n56639 );
nand ( n69475 , n69468 , n69474 );
xor ( n69476 , n69465 , n69475 );
xor ( n69477 , n69476 , n69147 );
xor ( n69478 , n69454 , n69477 );
xor ( n69479 , n69453 , n69283 );
and ( n69480 , n69479 , n69477 );
and ( n69481 , n69453 , n69283 );
or ( n69482 , n69480 , n69481 );
not ( n69483 , n52022 );
not ( n69484 , n69104 );
or ( n69485 , n69483 , n69484 );
not ( n69486 , n54625 );
not ( n69487 , n59402 );
or ( n69488 , n69486 , n69487 );
nand ( n69489 , n39574 , n55023 );
nand ( n69490 , n69488 , n69489 );
nand ( n69491 , n69490 , n54623 );
nand ( n69492 , n69485 , n69491 );
not ( n69493 , n52970 );
not ( n69494 , n69117 );
or ( n69495 , n69493 , n69494 );
not ( n69496 , n57810 );
not ( n69497 , n42399 );
or ( n69498 , n69496 , n69497 );
nand ( n69499 , n65546 , n67477 );
nand ( n69500 , n69498 , n69499 );
nand ( n69501 , n69500 , n52043 );
nand ( n69502 , n69495 , n69501 );
xor ( n69503 , n69492 , n69502 );
not ( n69504 , n58977 );
not ( n69505 , n60602 );
not ( n69506 , n62357 );
or ( n69507 , n69505 , n69506 );
nand ( n69508 , n66546 , n52728 );
nand ( n69509 , n69507 , n69508 );
not ( n69510 , n69509 );
or ( n69511 , n69504 , n69510 );
nand ( n69512 , n69089 , n53104 );
nand ( n69513 , n69511 , n69512 );
xor ( n69514 , n69503 , n69513 );
xor ( n69515 , n68888 , n69514 );
not ( n69516 , n51865 );
not ( n69517 , n52267 );
not ( n69518 , n65824 );
or ( n69519 , n69517 , n69518 );
not ( n69520 , n63787 );
nand ( n69521 , n69520 , n51351 );
nand ( n69522 , n69519 , n69521 );
not ( n69523 , n69522 );
or ( n69524 , n69516 , n69523 );
nand ( n69525 , n69056 , n49713 );
nand ( n69526 , n69524 , n69525 );
not ( n69527 , n52421 );
not ( n69528 , n69065 );
or ( n69529 , n69527 , n69528 );
buf ( n69530 , n39253 );
not ( n69531 , n69530 );
not ( n69532 , n51724 );
or ( n69533 , n69531 , n69532 );
not ( n69534 , n69530 );
nand ( n69535 , n69534 , n51723 );
nand ( n69536 , n69533 , n69535 );
nand ( n69537 , n69536 , n54875 );
nand ( n69538 , n69529 , n69537 );
xor ( n69539 , n69526 , n69538 );
not ( n69540 , n69076 );
or ( n69541 , n69540 , n56515 );
and ( n69542 , n68652 , n52377 );
not ( n69543 , n68652 );
and ( n69544 , n69543 , n55013 );
or ( n69545 , n69542 , n69544 );
not ( n69546 , n69545 );
or ( n69547 , n69546 , n56523 );
nand ( n69548 , n69541 , n69547 );
xor ( n69549 , n69539 , n69548 );
xor ( n69550 , n69515 , n69549 );
xor ( n69551 , n68888 , n69514 );
and ( n69552 , n69551 , n69549 );
and ( n69553 , n68888 , n69514 );
or ( n69554 , n69552 , n69553 );
xor ( n69555 , n68923 , n69342 );
xor ( n69556 , n69555 , n68894 );
xor ( n69557 , n68923 , n69342 );
and ( n69558 , n69557 , n68894 );
and ( n69559 , n68923 , n69342 );
or ( n69560 , n69558 , n69559 );
xor ( n69561 , n69348 , n68929 );
xor ( n69562 , n69561 , n69006 );
xor ( n69563 , n69348 , n68929 );
and ( n69564 , n69563 , n69006 );
and ( n69565 , n69348 , n68929 );
or ( n69566 , n69564 , n69565 );
xor ( n69567 , n69354 , n69125 );
xor ( n69568 , n69567 , n69047 );
xor ( n69569 , n69354 , n69125 );
and ( n69570 , n69569 , n69047 );
and ( n69571 , n69354 , n69125 );
or ( n69572 , n69570 , n69571 );
xor ( n69573 , n69318 , n69328 );
and ( n69574 , n69573 , n69339 );
and ( n69575 , n69318 , n69328 );
or ( n69576 , n69574 , n69575 );
xor ( n69577 , n69415 , n69550 );
xor ( n69578 , n69577 , n69478 );
xor ( n69579 , n69415 , n69550 );
and ( n69580 , n69579 , n69478 );
and ( n69581 , n69415 , n69550 );
or ( n69582 , n69580 , n69581 );
xor ( n69583 , n69137 , n69556 );
xor ( n69584 , n69583 , n69131 );
xor ( n69585 , n69137 , n69556 );
and ( n69586 , n69585 , n69131 );
and ( n69587 , n69137 , n69556 );
or ( n69588 , n69586 , n69587 );
xor ( n69589 , n69143 , n69562 );
xor ( n69590 , n69589 , n69568 );
xor ( n69591 , n69143 , n69562 );
and ( n69592 , n69591 , n69568 );
and ( n69593 , n69143 , n69562 );
or ( n69594 , n69592 , n69593 );
xor ( n69595 , n69153 , n69578 );
xor ( n69596 , n69595 , n69159 );
xor ( n69597 , n69153 , n69578 );
and ( n69598 , n69597 , n69159 );
and ( n69599 , n69153 , n69578 );
or ( n69600 , n69598 , n69599 );
xor ( n69601 , n69584 , n69165 );
xor ( n69602 , n69601 , n69590 );
xor ( n69603 , n69584 , n69165 );
and ( n69604 , n69603 , n69590 );
and ( n69605 , n69584 , n69165 );
or ( n69606 , n69604 , n69605 );
xor ( n69607 , n69171 , n69596 );
xor ( n69608 , n69607 , n69177 );
xor ( n69609 , n69171 , n69596 );
and ( n69610 , n69609 , n69177 );
and ( n69611 , n69171 , n69596 );
or ( n69612 , n69610 , n69611 );
xor ( n69613 , n69602 , n69608 );
xor ( n69614 , n69613 , n69183 );
xor ( n69615 , n69602 , n69608 );
and ( n69616 , n69615 , n69183 );
and ( n69617 , n69602 , n69608 );
or ( n69618 , n69616 , n69617 );
xor ( n69619 , n69293 , n69303 );
and ( n69620 , n69619 , n69306 );
and ( n69621 , n69293 , n69303 );
or ( n69622 , n69620 , n69621 );
xor ( n69623 , n69429 , n69439 );
and ( n69624 , n69623 , n69452 );
and ( n69625 , n69429 , n69439 );
or ( n69626 , n69624 , n69625 );
xor ( n69627 , n69391 , n69401 );
and ( n69628 , n69627 , n69413 );
and ( n69629 , n69391 , n69401 );
or ( n69630 , n69628 , n69629 );
xor ( n69631 , n69369 , n69378 );
and ( n69632 , n69631 , n69039 );
and ( n69633 , n69369 , n69378 );
or ( n69634 , n69632 , n69633 );
xor ( n69635 , n69465 , n69475 );
and ( n69636 , n69635 , n69147 );
and ( n69637 , n69465 , n69475 );
or ( n69638 , n69636 , n69637 );
xor ( n69639 , n69526 , n69538 );
and ( n69640 , n69639 , n69548 );
and ( n69641 , n69526 , n69538 );
or ( n69642 , n69640 , n69641 );
xor ( n69643 , n69492 , n69502 );
and ( n69644 , n69643 , n69513 );
and ( n69645 , n69492 , n69502 );
or ( n69646 , n69644 , n69645 );
or ( n69647 , n67885 , n69263 );
not ( n69648 , n57631 );
and ( n69649 , n52592 , n62485 );
not ( n69650 , n52592 );
and ( n69651 , n69650 , n65175 );
nor ( n69652 , n69649 , n69651 );
or ( n69653 , n69648 , n69652 );
nand ( n69654 , n69647 , n69653 );
not ( n69655 , n69274 );
not ( n69656 , n69655 );
not ( n69657 , n65646 );
or ( n69658 , n69656 , n69657 );
not ( n69659 , n48486 );
not ( n69660 , n66652 );
or ( n69661 , n69659 , n69660 );
nand ( n69662 , n65184 , n48951 );
nand ( n69663 , n69661 , n69662 );
nand ( n69664 , n61465 , n69663 );
nand ( n69665 , n69658 , n69664 );
xor ( n69666 , n69654 , n69665 );
not ( n69667 , n69316 );
or ( n69668 , n66980 , n69667 );
and ( n69669 , n66947 , n66983 );
not ( n69670 , n66947 );
and ( n69671 , n69670 , n65664 );
nor ( n69672 , n69669 , n69671 );
or ( n69673 , n67586 , n69672 );
nand ( n69674 , n69668 , n69673 );
xor ( n69675 , n69666 , n69674 );
xor ( n69676 , n69654 , n69665 );
and ( n69677 , n69676 , n69674 );
and ( n69678 , n69654 , n69665 );
or ( n69679 , n69677 , n69678 );
not ( n69680 , n69326 );
not ( n69681 , n65130 );
or ( n69682 , n69680 , n69681 );
and ( n69683 , n58180 , n66141 );
not ( n69684 , n58180 );
and ( n69685 , n69684 , n66140 );
nor ( n69686 , n69683 , n69685 );
or ( n69687 , n60963 , n69686 );
nand ( n69688 , n69682 , n69687 );
not ( n69689 , n69241 );
not ( n69690 , n56281 );
or ( n69691 , n69689 , n69690 );
not ( n69692 , n50021 );
not ( n69693 , n55873 );
or ( n69694 , n69692 , n69693 );
not ( n69695 , n55846 );
nand ( n69696 , n50020 , n69695 );
nand ( n69697 , n69694 , n69696 );
nand ( n69698 , n59984 , n69697 );
nand ( n69699 , n69691 , n69698 );
xor ( n69700 , n69688 , n69699 );
or ( n69701 , n64164 , n69291 );
not ( n69702 , n64166 );
not ( n69703 , n69702 );
not ( n69704 , n64170 );
and ( n69705 , n48983 , n69704 );
not ( n69706 , n48983 );
not ( n69707 , n62452 );
and ( n69708 , n69706 , n69707 );
nor ( n69709 , n69705 , n69708 );
or ( n69710 , n69703 , n69709 );
nand ( n69711 , n69701 , n69710 );
xor ( n69712 , n69700 , n69711 );
xor ( n69713 , n69688 , n69699 );
and ( n69714 , n69713 , n69711 );
and ( n69715 , n69688 , n69699 );
or ( n69716 , n69714 , n69715 );
not ( n69717 , n69301 );
not ( n69718 , n65089 );
or ( n69719 , n69717 , n69718 );
and ( n69720 , n54611 , n65094 );
not ( n69721 , n54611 );
and ( n69722 , n69721 , n65474 );
or ( n69723 , n69720 , n69722 );
nand ( n69724 , n69723 , n65092 );
nand ( n69725 , n69719 , n69724 );
and ( n69726 , n67072 , n51792 );
xor ( n69727 , n69725 , n69726 );
buf ( n69728 , n61549 );
not ( n69729 , n69337 );
or ( n69730 , n69728 , n69729 );
not ( n69731 , n61558 );
and ( n69732 , n57182 , n61537 );
not ( n69733 , n57182 );
and ( n69734 , n69733 , n61540 );
or ( n69735 , n69732 , n69734 );
not ( n69736 , n69735 );
or ( n69737 , n69731 , n69736 );
nand ( n69738 , n69730 , n69737 );
xor ( n69739 , n69727 , n69738 );
xor ( n69740 , n69576 , n69739 );
xor ( n69741 , n69740 , n69712 );
xor ( n69742 , n69576 , n69739 );
and ( n69743 , n69742 , n69712 );
and ( n69744 , n69576 , n69739 );
or ( n69745 , n69743 , n69744 );
xor ( n69746 , n69675 , n69626 );
xor ( n69747 , n69746 , n69630 );
xor ( n69748 , n69675 , n69626 );
and ( n69749 , n69748 , n69630 );
and ( n69750 , n69675 , n69626 );
or ( n69751 , n69749 , n69750 );
xor ( n69752 , n69634 , n69638 );
xor ( n69753 , n69752 , n69642 );
xor ( n69754 , n69634 , n69638 );
and ( n69755 , n69754 , n69642 );
and ( n69756 , n69634 , n69638 );
or ( n69757 , n69755 , n69756 );
not ( n69758 , n52139 );
not ( n69759 , n69367 );
or ( n69760 , n69758 , n69759 );
nand ( n69761 , n59195 , n51566 );
not ( n69762 , n69761 );
nand ( n69763 , n66236 , n65103 );
not ( n69764 , n69763 );
or ( n69765 , n69762 , n69764 );
nand ( n69766 , n69765 , n51533 );
nand ( n69767 , n69760 , n69766 );
not ( n69768 , n52125 );
not ( n69769 , n69374 );
or ( n69770 , n69768 , n69769 );
not ( n69771 , n52114 );
not ( n69772 , n53286 );
or ( n69773 , n69771 , n69772 );
not ( n69774 , n54020 );
nand ( n69775 , n69774 , n52110 );
nand ( n69776 , n69773 , n69775 );
nand ( n69777 , n69776 , n51766 );
nand ( n69778 , n69770 , n69777 );
xor ( n69779 , n69767 , n69778 );
not ( n69780 , n53571 );
and ( n69781 , n53271 , n52840 );
not ( n69782 , n53271 );
and ( n69783 , n69782 , n55104 );
or ( n69784 , n69781 , n69783 );
not ( n69785 , n69784 );
or ( n69786 , n69780 , n69785 );
nand ( n69787 , n69463 , n52854 );
nand ( n69788 , n69786 , n69787 );
xor ( n69789 , n69779 , n69788 );
xor ( n69790 , n69646 , n69789 );
not ( n69791 , n52757 );
not ( n69792 , n55630 );
not ( n69793 , n64190 );
or ( n69794 , n69792 , n69793 );
nand ( n69795 , n56412 , n64191 );
nand ( n69796 , n69794 , n69795 );
not ( n69797 , n69796 );
or ( n69798 , n69791 , n69797 );
nand ( n69799 , n69399 , n63708 );
nand ( n69800 , n69798 , n69799 );
not ( n69801 , n52151 );
not ( n69802 , n69411 );
or ( n69803 , n69801 , n69802 );
not ( n69804 , n51461 );
not ( n69805 , n56438 );
or ( n69806 , n69804 , n69805 );
nand ( n69807 , n54791 , n52781 );
nand ( n69808 , n69806 , n69807 );
nand ( n69809 , n69808 , n50922 );
nand ( n69810 , n69803 , n69809 );
xor ( n69811 , n69800 , n69810 );
not ( n69812 , n69253 );
not ( n69813 , n69812 );
not ( n69814 , n56777 );
or ( n69815 , n69813 , n69814 );
not ( n69816 , n51740 );
not ( n69817 , n56785 );
or ( n69818 , n69816 , n69817 );
buf ( n69819 , n56759 );
not ( n69820 , n69819 );
nand ( n69821 , n69820 , n40855 );
nand ( n69822 , n69818 , n69821 );
nand ( n69823 , n56780 , n69822 );
nand ( n69824 , n69815 , n69823 );
not ( n69825 , n69824 );
xor ( n69826 , n69811 , n69825 );
xor ( n69827 , n69790 , n69826 );
xor ( n69828 , n69646 , n69789 );
and ( n69829 , n69828 , n69826 );
and ( n69830 , n69646 , n69789 );
or ( n69831 , n69829 , n69830 );
not ( n69832 , n54848 );
not ( n69833 , n55124 );
not ( n69834 , n50654 );
or ( n69835 , n69833 , n69834 );
nand ( n69836 , n40692 , n55119 );
nand ( n69837 , n69835 , n69836 );
not ( n69838 , n69837 );
or ( n69839 , n69832 , n69838 );
nand ( n69840 , n55576 , n69229 );
nand ( n69841 , n69839 , n69840 );
not ( n69842 , n54327 );
not ( n69843 , n54323 );
not ( n69844 , n40735 );
or ( n69845 , n69843 , n69844 );
not ( n69846 , n59078 );
nand ( n69847 , n69846 , n57332 );
nand ( n69848 , n69845 , n69847 );
not ( n69849 , n69848 );
or ( n69850 , n69842 , n69849 );
nand ( n69851 , n69425 , n54316 );
nand ( n69852 , n69850 , n69851 );
xor ( n69853 , n69841 , n69852 );
not ( n69854 , n66696 );
not ( n69855 , n69389 );
or ( n69856 , n69854 , n69855 );
xor ( n69857 , n61951 , n67196 );
nand ( n69858 , n62654 , n69857 );
nand ( n69859 , n69856 , n69858 );
xor ( n69860 , n69853 , n69859 );
not ( n69861 , n56639 );
not ( n69862 , n59345 );
not ( n69863 , n67037 );
or ( n69864 , n69862 , n69863 );
nand ( n69865 , n59913 , n60617 );
nand ( n69866 , n69864 , n69865 );
not ( n69867 , n69866 );
or ( n69868 , n69861 , n69867 );
nand ( n69869 , n69473 , n59950 );
nand ( n69870 , n69868 , n69869 );
xor ( n69871 , n69870 , n69248 );
xor ( n69872 , n69871 , n69281 );
xor ( n69873 , n69860 , n69872 );
xor ( n69874 , n69873 , n69287 );
xor ( n69875 , n69860 , n69872 );
and ( n69876 , n69875 , n69287 );
and ( n69877 , n69860 , n69872 );
or ( n69878 , n69876 , n69877 );
not ( n69879 , n53956 );
not ( n69880 , n69448 );
or ( n69881 , n69879 , n69880 );
not ( n69882 , n55089 );
not ( n69883 , n40527 );
or ( n69884 , n69882 , n69883 );
nand ( n69885 , n51916 , n69444 );
nand ( n69886 , n69884 , n69885 );
nand ( n69887 , n69886 , n53620 );
nand ( n69888 , n69881 , n69887 );
not ( n69889 , n60927 );
not ( n69890 , n66234 );
not ( n69891 , n62970 );
or ( n69892 , n69890 , n69891 );
not ( n69893 , n66234 );
nand ( n69894 , n39845 , n69893 );
nand ( n69895 , n69892 , n69894 );
not ( n69896 , n69895 );
or ( n69897 , n69889 , n69896 );
nand ( n69898 , n69437 , n58168 );
nand ( n69899 , n69897 , n69898 );
xor ( n69900 , n69888 , n69899 );
xor ( n69901 , n69900 , n69622 );
xor ( n69902 , n69901 , n69346 );
not ( n69903 , n52962 );
not ( n69904 , n67477 );
not ( n69905 , n42555 );
or ( n69906 , n69904 , n69905 );
nand ( n69907 , n57810 , n67269 );
nand ( n69908 , n69906 , n69907 );
not ( n69909 , n69908 );
or ( n69910 , n69903 , n69909 );
nand ( n69911 , n69500 , n52970 );
nand ( n69912 , n69910 , n69911 );
not ( n69913 , n57314 );
not ( n69914 , n69545 );
or ( n69915 , n69913 , n69914 );
not ( n69916 , n52377 );
not ( n69917 , n39333 );
or ( n69918 , n69916 , n69917 );
not ( n69919 , n60855 );
nand ( n69920 , n69919 , n55013 );
nand ( n69921 , n69918 , n69920 );
nand ( n69922 , n69921 , n52004 );
nand ( n69923 , n69915 , n69922 );
xor ( n69924 , n69912 , n69923 );
not ( n69925 , n54623 );
not ( n69926 , n59174 );
not ( n69927 , n60874 );
or ( n69928 , n69926 , n69927 );
nand ( n69929 , n63152 , n54628 );
nand ( n69930 , n69928 , n69929 );
not ( n69931 , n69930 );
or ( n69932 , n69925 , n69931 );
nand ( n69933 , n69490 , n52022 );
nand ( n69934 , n69932 , n69933 );
xor ( n69935 , n69924 , n69934 );
xor ( n69936 , n69902 , n69935 );
xor ( n69937 , n69901 , n69346 );
and ( n69938 , n69937 , n69935 );
and ( n69939 , n69901 , n69346 );
or ( n69940 , n69938 , n69939 );
not ( n69941 , n49713 );
not ( n69942 , n69522 );
or ( n69943 , n69941 , n69942 );
nand ( n69944 , n51865 , n49707 );
nand ( n69945 , n69943 , n69944 );
not ( n69946 , n53104 );
not ( n69947 , n69509 );
or ( n69948 , n69946 , n69947 );
not ( n69949 , n60602 );
not ( n69950 , n62931 );
or ( n69951 , n69949 , n69950 );
nand ( n69952 , n39714 , n62577 );
nand ( n69953 , n69951 , n69952 );
nand ( n69954 , n69953 , n58977 );
nand ( n69955 , n69948 , n69954 );
xor ( n69956 , n69945 , n69955 );
not ( n69957 , n54875 );
not ( n69958 , n51723 );
not ( n69959 , n62909 );
or ( n69960 , n69958 , n69959 );
buf ( n69961 , n62909 );
not ( n69962 , n69961 );
nand ( n69963 , n69962 , n51724 );
nand ( n69964 , n69960 , n69963 );
not ( n69965 , n69964 );
or ( n69966 , n69957 , n69965 );
nand ( n69967 , n52421 , n69536 );
nand ( n69968 , n69966 , n69967 );
xor ( n69969 , n69956 , n69968 );
xor ( n69970 , n69969 , n69741 );
xor ( n69971 , n69970 , n69352 );
xor ( n69972 , n69969 , n69741 );
and ( n69973 , n69972 , n69352 );
and ( n69974 , n69969 , n69741 );
or ( n69975 , n69973 , n69974 );
xor ( n69976 , n69358 , n69419 );
xor ( n69977 , n69976 , n69747 );
xor ( n69978 , n69358 , n69419 );
and ( n69979 , n69978 , n69747 );
and ( n69980 , n69358 , n69419 );
or ( n69981 , n69979 , n69980 );
xor ( n69982 , n69482 , n69753 );
xor ( n69983 , n69982 , n69554 );
xor ( n69984 , n69482 , n69753 );
and ( n69985 , n69984 , n69554 );
and ( n69986 , n69482 , n69753 );
or ( n69987 , n69985 , n69986 );
xor ( n69988 , n69827 , n69560 );
xor ( n69989 , n69988 , n69936 );
xor ( n69990 , n69827 , n69560 );
and ( n69991 , n69990 , n69936 );
and ( n69992 , n69827 , n69560 );
or ( n69993 , n69991 , n69992 );
xor ( n69994 , n69725 , n69726 );
and ( n69995 , n69994 , n69738 );
and ( n69996 , n69725 , n69726 );
or ( n69997 , n69995 , n69996 );
xor ( n69998 , n69874 , n69566 );
xor ( n69999 , n69998 , n69971 );
xor ( n70000 , n69874 , n69566 );
and ( n70001 , n70000 , n69971 );
and ( n70002 , n69874 , n69566 );
or ( n70003 , n70001 , n70002 );
xor ( n70004 , n69977 , n69572 );
xor ( n70005 , n70004 , n69983 );
xor ( n70006 , n69977 , n69572 );
and ( n70007 , n70006 , n69983 );
and ( n70008 , n69977 , n69572 );
or ( n70009 , n70007 , n70008 );
xor ( n70010 , n69582 , n69989 );
xor ( n70011 , n70010 , n69588 );
xor ( n70012 , n69582 , n69989 );
and ( n70013 , n70012 , n69588 );
and ( n70014 , n69582 , n69989 );
or ( n70015 , n70013 , n70014 );
xor ( n70016 , n69999 , n70005 );
xor ( n70017 , n70016 , n69594 );
xor ( n70018 , n69999 , n70005 );
and ( n70019 , n70018 , n69594 );
and ( n70020 , n69999 , n70005 );
or ( n70021 , n70019 , n70020 );
xor ( n70022 , n70011 , n69600 );
xor ( n70023 , n70022 , n69606 );
xor ( n70024 , n70011 , n69600 );
and ( n70025 , n70024 , n69606 );
and ( n70026 , n70011 , n69600 );
or ( n70027 , n70025 , n70026 );
xor ( n70028 , n70017 , n70023 );
xor ( n70029 , n70028 , n69612 );
xor ( n70030 , n70017 , n70023 );
and ( n70031 , n70030 , n69612 );
and ( n70032 , n70017 , n70023 );
or ( n70033 , n70031 , n70032 );
xor ( n70034 , n69841 , n69852 );
and ( n70035 , n70034 , n69859 );
and ( n70036 , n69841 , n69852 );
or ( n70037 , n70035 , n70036 );
xor ( n70038 , n69800 , n69810 );
and ( n70039 , n70038 , n69825 );
and ( n70040 , n69800 , n69810 );
or ( n70041 , n70039 , n70040 );
xor ( n70042 , n69767 , n69778 );
and ( n70043 , n70042 , n69788 );
and ( n70044 , n69767 , n69778 );
or ( n70045 , n70043 , n70044 );
xor ( n70046 , n69888 , n69899 );
and ( n70047 , n70046 , n69622 );
and ( n70048 , n69888 , n69899 );
or ( n70049 , n70047 , n70048 );
xor ( n70050 , n69912 , n69923 );
and ( n70051 , n70050 , n69934 );
and ( n70052 , n69912 , n69923 );
or ( n70053 , n70051 , n70052 );
xor ( n70054 , n69945 , n69955 );
and ( n70055 , n70054 , n69968 );
and ( n70056 , n69945 , n69955 );
or ( n70057 , n70055 , n70056 );
xor ( n70058 , n69870 , n69248 );
and ( n70059 , n70058 , n69281 );
and ( n70060 , n69870 , n69248 );
or ( n70061 , n70059 , n70060 );
not ( n70062 , n60633 );
not ( n70063 , n50057 );
or ( n70064 , n70062 , n70063 );
nand ( n70065 , n70064 , n52267 );
not ( n70066 , n69697 );
not ( n70067 , n56281 );
or ( n70068 , n70066 , n70067 );
not ( n70069 , n55872 );
not ( n70070 , n53513 );
or ( n70071 , n70069 , n70070 );
nand ( n70072 , n52079 , n69237 );
nand ( n70073 , n70071 , n70072 );
nand ( n70074 , n70073 , n55458 );
nand ( n70075 , n70068 , n70074 );
xor ( n70076 , n70065 , n70075 );
not ( n70077 , n69822 );
not ( n70078 , n56777 );
or ( n70079 , n70077 , n70078 );
not ( n70080 , n65999 );
not ( n70081 , n64451 );
or ( n70082 , n70080 , n70081 );
buf ( n70083 , n52916 );
nand ( n70084 , n69819 , n70083 );
nand ( n70085 , n70082 , n70084 );
nand ( n70086 , n56780 , n70085 );
nand ( n70087 , n70079 , n70086 );
xor ( n70088 , n70076 , n70087 );
xor ( n70089 , n70065 , n70075 );
and ( n70090 , n70089 , n70087 );
and ( n70091 , n70065 , n70075 );
or ( n70092 , n70090 , n70091 );
or ( n70093 , n65169 , n69652 );
and ( n70094 , n57615 , n53706 );
not ( n70095 , n57571 );
and ( n70096 , n57619 , n70095 );
nor ( n70097 , n70094 , n70096 );
or ( n70098 , n65638 , n70097 );
nand ( n70099 , n70093 , n70098 );
not ( n70100 , n69663 );
not ( n70101 , n65646 );
or ( n70102 , n70100 , n70101 );
not ( n70103 , n62496 );
not ( n70104 , n49820 );
and ( n70105 , n70103 , n70104 );
and ( n70106 , n52271 , n65652 );
nor ( n70107 , n70105 , n70106 );
not ( n70108 , n70107 );
nand ( n70109 , n70108 , n61465 );
nand ( n70110 , n70102 , n70109 );
xor ( n70111 , n70099 , n70110 );
not ( n70112 , n69672 );
not ( n70113 , n70112 );
not ( n70114 , n62506 );
or ( n70115 , n70113 , n70114 );
not ( n70116 , n41532 );
not ( n70117 , n65121 );
or ( n70118 , n70116 , n70117 );
nand ( n70119 , n65664 , n44112 );
nand ( n70120 , n70118 , n70119 );
nand ( n70121 , n70120 , n59575 );
nand ( n70122 , n70115 , n70121 );
xor ( n70123 , n70111 , n70122 );
xor ( n70124 , n70099 , n70110 );
and ( n70125 , n70124 , n70122 );
and ( n70126 , n70099 , n70110 );
or ( n70127 , n70125 , n70126 );
xor ( n70128 , n69997 , n70088 );
or ( n70129 , n60960 , n69686 );
and ( n70130 , n60286 , n58458 );
and ( n70131 , n66140 , n58459 );
nor ( n70132 , n70130 , n70131 );
or ( n70133 , n60963 , n70132 );
nand ( n70134 , n70129 , n70133 );
not ( n70135 , n69735 );
not ( n70136 , n64111 );
or ( n70137 , n70135 , n70136 );
not ( n70138 , n47527 );
not ( n70139 , n64630 );
or ( n70140 , n70138 , n70139 );
nand ( n70141 , n61540 , n64603 );
nand ( n70142 , n70140 , n70141 );
nand ( n70143 , n61558 , n70142 );
nand ( n70144 , n70137 , n70143 );
xor ( n70145 , n70134 , n70144 );
not ( n70146 , n69709 );
not ( n70147 , n70146 );
not ( n70148 , n67061 );
or ( n70149 , n70147 , n70148 );
not ( n70150 , n62449 );
not ( n70151 , n56731 );
and ( n70152 , n70150 , n70151 );
and ( n70153 , n69707 , n56731 );
nor ( n70154 , n70152 , n70153 );
not ( n70155 , n70154 );
nand ( n70156 , n70155 , n67068 );
nand ( n70157 , n70149 , n70156 );
xor ( n70158 , n70145 , n70157 );
xor ( n70159 , n70128 , n70158 );
xor ( n70160 , n69997 , n70088 );
and ( n70161 , n70160 , n70158 );
and ( n70162 , n69997 , n70088 );
or ( n70163 , n70161 , n70162 );
xor ( n70164 , n70123 , n70037 );
xor ( n70165 , n70164 , n70041 );
xor ( n70166 , n70123 , n70037 );
and ( n70167 , n70166 , n70041 );
and ( n70168 , n70123 , n70037 );
or ( n70169 , n70167 , n70168 );
not ( n70170 , n69723 );
not ( n70171 , n65795 );
or ( n70172 , n70170 , n70171 );
not ( n70173 , n52712 );
not ( n70174 , n70173 );
not ( n70175 , n63412 );
or ( n70176 , n70174 , n70175 );
nand ( n70177 , n69305 , n52712 );
nand ( n70178 , n70176 , n70177 );
nand ( n70179 , n70178 , n65092 );
nand ( n70180 , n70172 , n70179 );
and ( n70181 , n64444 , n52033 );
xor ( n70182 , n70180 , n70181 );
buf ( n70183 , n54848 );
not ( n70184 , n70183 );
not ( n70185 , n55582 );
not ( n70186 , n52289 );
not ( n70187 , n70186 );
or ( n70188 , n70185 , n70187 );
nand ( n70189 , n52289 , n55148 );
nand ( n70190 , n70188 , n70189 );
not ( n70191 , n70190 );
or ( n70192 , n70184 , n70191 );
not ( n70193 , n68334 );
nand ( n70194 , n69837 , n70193 );
nand ( n70195 , n70192 , n70194 );
xor ( n70196 , n70182 , n70195 );
xor ( n70197 , n70045 , n70196 );
xor ( n70198 , n70197 , n70053 );
xor ( n70199 , n70045 , n70196 );
and ( n70200 , n70199 , n70053 );
and ( n70201 , n70045 , n70196 );
or ( n70202 , n70200 , n70201 );
xor ( n70203 , n70057 , n70061 );
not ( n70204 , n51223 );
not ( n70205 , n51461 );
not ( n70206 , n59694 );
or ( n70207 , n70205 , n70206 );
nand ( n70208 , n59697 , n53904 );
nand ( n70209 , n70207 , n70208 );
not ( n70210 , n70209 );
or ( n70211 , n70204 , n70210 );
nand ( n70212 , n69808 , n52526 );
nand ( n70213 , n70211 , n70212 );
not ( n70214 , n51533 );
not ( n70215 , n52816 );
not ( n70216 , n54402 );
or ( n70217 , n70215 , n70216 );
nand ( n70218 , n40149 , n53928 );
nand ( n70219 , n70217 , n70218 );
not ( n70220 , n70219 );
or ( n70221 , n70214 , n70220 );
not ( n70222 , n69763 );
not ( n70223 , n69761 );
or ( n70224 , n70222 , n70223 );
nand ( n70225 , n70224 , n56355 );
nand ( n70226 , n70221 , n70225 );
xor ( n70227 , n70213 , n70226 );
not ( n70228 , n51766 );
not ( n70229 , n52114 );
not ( n70230 , n55242 );
or ( n70231 , n70229 , n70230 );
nand ( n70232 , n53660 , n52110 );
nand ( n70233 , n70231 , n70232 );
not ( n70234 , n70233 );
or ( n70235 , n70228 , n70234 );
nand ( n70236 , n52482 , n69776 );
nand ( n70237 , n70235 , n70236 );
xor ( n70238 , n70227 , n70237 );
xor ( n70239 , n70203 , n70238 );
xor ( n70240 , n70057 , n70061 );
and ( n70241 , n70240 , n70238 );
and ( n70242 , n70057 , n70061 );
or ( n70243 , n70241 , n70242 );
not ( n70244 , n52469 );
not ( n70245 , n52840 );
not ( n70246 , n59611 );
or ( n70247 , n70245 , n70246 );
nand ( n70248 , n59612 , n53947 );
nand ( n70249 , n70247 , n70248 );
not ( n70250 , n70249 );
or ( n70251 , n70244 , n70250 );
nand ( n70252 , n69784 , n52854 );
nand ( n70253 , n70251 , n70252 );
xor ( n70254 , n70253 , n69824 );
not ( n70255 , n69886 );
not ( n70256 , n68603 );
or ( n70257 , n70255 , n70256 );
not ( n70258 , n55089 );
not ( n70259 , n53730 );
or ( n70260 , n70258 , n70259 );
nand ( n70261 , n40592 , n69444 );
nand ( n70262 , n70260 , n70261 );
nand ( n70263 , n54364 , n70262 );
nand ( n70264 , n70257 , n70263 );
xor ( n70265 , n70254 , n70264 );
not ( n70266 , n66696 );
not ( n70267 , n69857 );
or ( n70268 , n70266 , n70267 );
not ( n70269 , n61951 );
not ( n70270 , n59651 );
or ( n70271 , n70269 , n70270 );
nand ( n70272 , n59654 , n61952 );
nand ( n70273 , n70271 , n70272 );
nand ( n70274 , n70273 , n62654 );
nand ( n70275 , n70268 , n70274 );
not ( n70276 , n54327 );
not ( n70277 , n54323 );
not ( n70278 , n69442 );
not ( n70279 , n70278 );
or ( n70280 , n70277 , n70279 );
nand ( n70281 , n69442 , n54468 );
nand ( n70282 , n70280 , n70281 );
not ( n70283 , n70282 );
or ( n70284 , n70276 , n70283 );
nand ( n70285 , n69848 , n54316 );
nand ( n70286 , n70284 , n70285 );
xor ( n70287 , n70275 , n70286 );
not ( n70288 , n52757 );
not ( n70289 , n64190 );
not ( n70290 , n67721 );
not ( n70291 , n70290 );
or ( n70292 , n70289 , n70291 );
nand ( n70293 , n67721 , n66705 );
nand ( n70294 , n70292 , n70293 );
not ( n70295 , n70294 );
or ( n70296 , n70288 , n70295 );
nand ( n70297 , n69796 , n52749 );
nand ( n70298 , n70296 , n70297 );
xor ( n70299 , n70287 , n70298 );
xor ( n70300 , n70265 , n70299 );
xor ( n70301 , n70300 , n70049 );
xor ( n70302 , n70265 , n70299 );
and ( n70303 , n70302 , n70049 );
and ( n70304 , n70265 , n70299 );
or ( n70305 , n70303 , n70304 );
not ( n70306 , n56639 );
not ( n70307 , n59345 );
not ( n70308 , n66547 );
or ( n70309 , n70307 , n70308 );
nand ( n70310 , n66546 , n65743 );
nand ( n70311 , n70309 , n70310 );
not ( n70312 , n70311 );
or ( n70313 , n70306 , n70312 );
nand ( n70314 , n69866 , n59950 );
nand ( n70315 , n70313 , n70314 );
xor ( n70316 , n70315 , n69679 );
xor ( n70317 , n70316 , n69716 );
xor ( n70318 , n70317 , n69745 );
not ( n70319 , n58168 );
not ( n70320 , n69895 );
or ( n70321 , n70319 , n70320 );
not ( n70322 , n62077 );
not ( n70323 , n39895 );
or ( n70324 , n70322 , n70323 );
nand ( n70325 , n68510 , n60289 );
nand ( n70326 , n70324 , n70325 );
nand ( n70327 , n70326 , n52191 );
nand ( n70328 , n70321 , n70327 );
not ( n70329 , n52962 );
not ( n70330 , n67478 );
not ( n70331 , n66784 );
or ( n70332 , n70330 , n70331 );
not ( n70333 , n42653 );
nand ( n70334 , n70333 , n67477 );
nand ( n70335 , n70332 , n70334 );
not ( n70336 , n70335 );
or ( n70337 , n70329 , n70336 );
nand ( n70338 , n69908 , n52970 );
nand ( n70339 , n70337 , n70338 );
xor ( n70340 , n70328 , n70339 );
not ( n70341 , n52004 );
nand ( n70342 , n69530 , n55013 );
nand ( n70343 , n69534 , n52377 );
nand ( n70344 , n70342 , n70343 );
not ( n70345 , n70344 );
or ( n70346 , n70341 , n70345 );
nand ( n70347 , n69921 , n57314 );
nand ( n70348 , n70346 , n70347 );
xor ( n70349 , n70340 , n70348 );
xor ( n70350 , n70318 , n70349 );
xor ( n70351 , n70317 , n69745 );
and ( n70352 , n70351 , n70349 );
and ( n70353 , n70317 , n69745 );
or ( n70354 , n70352 , n70353 );
buf ( n70355 , n47873 );
not ( n70356 , n70355 );
not ( n70357 , n69930 );
or ( n70358 , n70356 , n70357 );
not ( n70359 , n59174 );
not ( n70360 , n62394 );
or ( n70361 , n70359 , n70360 );
nand ( n70362 , n38499 , n55023 );
nand ( n70363 , n70361 , n70362 );
nand ( n70364 , n54623 , n70363 );
nand ( n70365 , n70358 , n70364 );
not ( n70366 , n58977 );
and ( n70367 , n58982 , n39574 );
not ( n70368 , n58982 );
and ( n70369 , n70368 , n59402 );
nor ( n70370 , n70367 , n70369 );
not ( n70371 , n70370 );
or ( n70372 , n70366 , n70371 );
nand ( n70373 , n69953 , n53104 );
nand ( n70374 , n70372 , n70373 );
xor ( n70375 , n70365 , n70374 );
not ( n70376 , n52421 );
not ( n70377 , n69964 );
or ( n70378 , n70376 , n70377 );
not ( n70379 , n51723 );
not ( n70380 , n62381 );
or ( n70381 , n70379 , n70380 );
nand ( n70382 , n66536 , n51724 );
nand ( n70383 , n70381 , n70382 );
nand ( n70384 , n70383 , n54875 );
nand ( n70385 , n70378 , n70384 );
xor ( n70386 , n70375 , n70385 );
xor ( n70387 , n70386 , n70159 );
xor ( n70388 , n70387 , n69751 );
xor ( n70389 , n70386 , n70159 );
and ( n70390 , n70389 , n69751 );
and ( n70391 , n70386 , n70159 );
or ( n70392 , n70390 , n70391 );
xor ( n70393 , n69757 , n70198 );
xor ( n70394 , n70393 , n69831 );
xor ( n70395 , n69757 , n70198 );
and ( n70396 , n70395 , n69831 );
and ( n70397 , n69757 , n70198 );
or ( n70398 , n70396 , n70397 );
xor ( n70399 , n70165 , n69878 );
xor ( n70400 , n70399 , n69940 );
xor ( n70401 , n70165 , n69878 );
and ( n70402 , n70401 , n69940 );
and ( n70403 , n70165 , n69878 );
or ( n70404 , n70402 , n70403 );
xor ( n70405 , n70301 , n70239 );
xor ( n70406 , n70405 , n69975 );
xor ( n70407 , n70301 , n70239 );
and ( n70408 , n70407 , n69975 );
and ( n70409 , n70301 , n70239 );
or ( n70410 , n70408 , n70409 );
xor ( n70411 , n70134 , n70144 );
and ( n70412 , n70411 , n70157 );
and ( n70413 , n70134 , n70144 );
or ( n70414 , n70412 , n70413 );
xor ( n70415 , n70350 , n69981 );
xor ( n70416 , n70415 , n70388 );
xor ( n70417 , n70350 , n69981 );
and ( n70418 , n70417 , n70388 );
and ( n70419 , n70350 , n69981 );
or ( n70420 , n70418 , n70419 );
xor ( n70421 , n70394 , n69987 );
xor ( n70422 , n70421 , n70400 );
xor ( n70423 , n70394 , n69987 );
and ( n70424 , n70423 , n70400 );
and ( n70425 , n70394 , n69987 );
or ( n70426 , n70424 , n70425 );
xor ( n70427 , n69993 , n70406 );
xor ( n70428 , n70427 , n70003 );
xor ( n70429 , n69993 , n70406 );
and ( n70430 , n70429 , n70003 );
and ( n70431 , n69993 , n70406 );
or ( n70432 , n70430 , n70431 );
xor ( n70433 , n70416 , n70009 );
xor ( n70434 , n70433 , n70422 );
xor ( n70435 , n70416 , n70009 );
and ( n70436 , n70435 , n70422 );
and ( n70437 , n70416 , n70009 );
or ( n70438 , n70436 , n70437 );
xor ( n70439 , n70428 , n70015 );
xor ( n70440 , n70439 , n70021 );
xor ( n70441 , n70428 , n70015 );
and ( n70442 , n70441 , n70021 );
and ( n70443 , n70428 , n70015 );
or ( n70444 , n70442 , n70443 );
xor ( n70445 , n70434 , n70440 );
xor ( n70446 , n70445 , n70027 );
xor ( n70447 , n70434 , n70440 );
and ( n70448 , n70447 , n70027 );
and ( n70449 , n70434 , n70440 );
or ( n70450 , n70448 , n70449 );
xor ( n70451 , n70180 , n70181 );
and ( n70452 , n70451 , n70195 );
and ( n70453 , n70180 , n70181 );
or ( n70454 , n70452 , n70453 );
xor ( n70455 , n70275 , n70286 );
and ( n70456 , n70455 , n70298 );
and ( n70457 , n70275 , n70286 );
or ( n70458 , n70456 , n70457 );
xor ( n70459 , n70213 , n70226 );
and ( n70460 , n70459 , n70237 );
and ( n70461 , n70213 , n70226 );
or ( n70462 , n70460 , n70461 );
xor ( n70463 , n70253 , n69824 );
and ( n70464 , n70463 , n70264 );
and ( n70465 , n70253 , n69824 );
or ( n70466 , n70464 , n70465 );
xor ( n70467 , n70328 , n70339 );
and ( n70468 , n70467 , n70348 );
and ( n70469 , n70328 , n70339 );
or ( n70470 , n70468 , n70469 );
xor ( n70471 , n70365 , n70374 );
and ( n70472 , n70471 , n70385 );
and ( n70473 , n70365 , n70374 );
or ( n70474 , n70472 , n70473 );
xor ( n70475 , n70315 , n69679 );
and ( n70476 , n70475 , n69716 );
and ( n70477 , n70315 , n69679 );
or ( n70478 , n70476 , n70477 );
not ( n70479 , n61961 );
or ( n70480 , n70479 , n70107 );
and ( n70481 , n65183 , n41288 );
and ( n70482 , n65652 , n41287 );
nor ( n70483 , n70481 , n70482 );
or ( n70484 , n64146 , n70483 );
nand ( n70485 , n70480 , n70484 );
not ( n70486 , n70120 );
buf ( n70487 , n59571 );
not ( n70488 , n70487 );
or ( n70489 , n70486 , n70488 );
not ( n70490 , n48486 );
not ( n70491 , n66983 );
or ( n70492 , n70490 , n70491 );
nand ( n70493 , n65664 , n48951 );
nand ( n70494 , n70492 , n70493 );
nand ( n70495 , n59575 , n70494 );
nand ( n70496 , n70489 , n70495 );
xor ( n70497 , n70485 , n70496 );
not ( n70498 , n70132 );
not ( n70499 , n70498 );
buf ( n70500 , n65130 );
not ( n70501 , n70500 );
or ( n70502 , n70499 , n70501 );
not ( n70503 , n58915 );
not ( n70504 , n60286 );
or ( n70505 , n70503 , n70504 );
buf ( n70506 , n66140 );
nand ( n70507 , n70506 , n66946 );
nand ( n70508 , n70505 , n70507 );
nand ( n70509 , n60427 , n70508 );
nand ( n70510 , n70502 , n70509 );
xor ( n70511 , n70497 , n70510 );
xor ( n70512 , n70485 , n70496 );
and ( n70513 , n70512 , n70510 );
and ( n70514 , n70485 , n70496 );
or ( n70515 , n70513 , n70514 );
not ( n70516 , n61550 );
not ( n70517 , n70142 );
or ( n70518 , n70516 , n70517 );
not ( n70519 , n52379 );
not ( n70520 , n61537 );
or ( n70521 , n70519 , n70520 );
nand ( n70522 , n66615 , n67906 );
nand ( n70523 , n70521 , n70522 );
nand ( n70524 , n67094 , n70523 );
nand ( n70525 , n70518 , n70524 );
not ( n70526 , n70085 );
not ( n70527 , n56777 );
or ( n70528 , n70526 , n70527 );
not ( n70529 , n50020 );
not ( n70530 , n65999 );
or ( n70531 , n70529 , n70530 );
nand ( n70532 , n69819 , n50021 );
nand ( n70533 , n70531 , n70532 );
nand ( n70534 , n60472 , n70533 );
nand ( n70535 , n70528 , n70534 );
xor ( n70536 , n70525 , n70535 );
or ( n70537 , n64684 , n70154 );
and ( n70538 , n58195 , n69707 );
not ( n70539 , n58195 );
and ( n70540 , n70539 , n66089 );
nor ( n70541 , n70538 , n70540 );
or ( n70542 , n64166 , n70541 );
nand ( n70543 , n70537 , n70542 );
xor ( n70544 , n70536 , n70543 );
xor ( n70545 , n70525 , n70535 );
and ( n70546 , n70545 , n70543 );
and ( n70547 , n70525 , n70535 );
or ( n70548 , n70546 , n70547 );
xor ( n70549 , n70544 , n70511 );
xor ( n70550 , n70549 , n70458 );
xor ( n70551 , n70544 , n70511 );
and ( n70552 , n70551 , n70458 );
and ( n70553 , n70544 , n70511 );
or ( n70554 , n70552 , n70553 );
xor ( n70555 , n70462 , n70466 );
xor ( n70556 , n70555 , n70454 );
xor ( n70557 , n70462 , n70466 );
and ( n70558 , n70557 , n70454 );
and ( n70559 , n70462 , n70466 );
or ( n70560 , n70558 , n70559 );
xor ( n70561 , n70474 , n70478 );
not ( n70562 , n55066 );
not ( n70563 , n65103 );
not ( n70564 , n57390 );
or ( n70565 , n70563 , n70564 );
nand ( n70566 , n68990 , n53928 );
nand ( n70567 , n70565 , n70566 );
not ( n70568 , n70567 );
or ( n70569 , n70562 , n70568 );
nand ( n70570 , n70219 , n56355 );
nand ( n70571 , n70569 , n70570 );
not ( n70572 , n52125 );
not ( n70573 , n70233 );
or ( n70574 , n70572 , n70573 );
not ( n70575 , n52490 );
not ( n70576 , n54811 );
or ( n70577 , n70575 , n70576 );
not ( n70578 , n63201 );
nand ( n70579 , n70578 , n52110 );
nand ( n70580 , n70577 , n70579 );
nand ( n70581 , n70580 , n51766 );
nand ( n70582 , n70574 , n70581 );
xor ( n70583 , n70571 , n70582 );
not ( n70584 , n70249 );
not ( n70585 , n52854 );
or ( n70586 , n70584 , n70585 );
not ( n70587 , n52841 );
not ( n70588 , n54020 );
or ( n70589 , n70587 , n70588 );
nand ( n70590 , n53290 , n52837 );
nand ( n70591 , n70589 , n70590 );
not ( n70592 , n70591 );
or ( n70593 , n70592 , n56861 );
nand ( n70594 , n70586 , n70593 );
xor ( n70595 , n70583 , n70594 );
xor ( n70596 , n70561 , n70595 );
xor ( n70597 , n70474 , n70478 );
and ( n70598 , n70597 , n70595 );
and ( n70599 , n70474 , n70478 );
or ( n70600 , n70598 , n70599 );
not ( n70601 , n67885 );
not ( n70602 , n70097 );
and ( n70603 , n70601 , n70602 );
buf ( n70604 , n57631 );
not ( n70605 , n70604 );
and ( n70606 , n40855 , n67568 );
not ( n70607 , n40855 );
not ( n70608 , n67568 );
and ( n70609 , n70607 , n70608 );
nor ( n70610 , n70606 , n70609 );
nor ( n70611 , n70605 , n70610 );
nor ( n70612 , n70603 , n70611 );
not ( n70613 , n68603 );
not ( n70614 , n70262 );
or ( n70615 , n70613 , n70614 );
not ( n70616 , n55089 );
not ( n70617 , n40627 );
or ( n70618 , n70616 , n70617 );
nand ( n70619 , n40628 , n53591 );
nand ( n70620 , n70618 , n70619 );
nand ( n70621 , n70620 , n53620 );
nand ( n70622 , n70615 , n70621 );
xor ( n70623 , n70612 , n70622 );
not ( n70624 , n54316 );
not ( n70625 , n70282 );
or ( n70626 , n70624 , n70625 );
not ( n70627 , n54468 );
not ( n70628 , n70627 );
not ( n70629 , n60138 );
or ( n70630 , n70628 , n70629 );
nand ( n70631 , n53347 , n55276 );
nand ( n70632 , n70630 , n70631 );
nand ( n70633 , n70632 , n54327 );
nand ( n70634 , n70626 , n70633 );
xor ( n70635 , n70623 , n70634 );
not ( n70636 , n70183 );
not ( n70637 , n55120 );
buf ( n70638 , n40733 );
not ( n70639 , n70638 );
or ( n70640 , n70637 , n70639 );
nand ( n70641 , n57332 , n55148 );
nand ( n70642 , n70640 , n70641 );
not ( n70643 , n70642 );
or ( n70644 , n70636 , n70643 );
nand ( n70645 , n70190 , n55144 );
nand ( n70646 , n70644 , n70645 );
not ( n70647 , n63708 );
not ( n70648 , n70294 );
or ( n70649 , n70647 , n70648 );
not ( n70650 , n64190 );
not ( n70651 , n63180 );
or ( n70652 , n70650 , n70651 );
buf ( n70653 , n67196 );
nand ( n70654 , n70653 , n66705 );
nand ( n70655 , n70652 , n70654 );
nand ( n70656 , n70655 , n52757 );
nand ( n70657 , n70649 , n70656 );
xor ( n70658 , n70646 , n70657 );
not ( n70659 , n50922 );
not ( n70660 , n50895 );
not ( n70661 , n40451 );
not ( n70662 , n70661 );
or ( n70663 , n70660 , n70662 );
nand ( n70664 , n68980 , n67639 );
nand ( n70665 , n70663 , n70664 );
not ( n70666 , n70665 );
or ( n70667 , n70659 , n70666 );
nand ( n70668 , n70209 , n52151 );
nand ( n70669 , n70667 , n70668 );
xor ( n70670 , n70658 , n70669 );
xor ( n70671 , n70635 , n70670 );
xor ( n70672 , n70671 , n70470 );
xor ( n70673 , n70635 , n70670 );
and ( n70674 , n70673 , n70470 );
and ( n70675 , n70635 , n70670 );
or ( n70676 , n70674 , n70675 );
xor ( n70677 , n70127 , n70414 );
not ( n70678 , n70178 );
not ( n70679 , n65795 );
or ( n70680 , n70678 , n70679 );
not ( n70681 , n48983 );
not ( n70682 , n64443 );
or ( n70683 , n70681 , n70682 );
nand ( n70684 , n63416 , n56348 );
nand ( n70685 , n70683 , n70684 );
nand ( n70686 , n70685 , n65092 );
nand ( n70687 , n70680 , n70686 );
and ( n70688 , n67072 , n54611 );
xor ( n70689 , n70687 , n70688 );
not ( n70690 , n59984 );
and ( n70691 , n40691 , n55873 );
not ( n70692 , n40691 );
and ( n70693 , n70692 , n69695 );
or ( n70694 , n70691 , n70693 );
not ( n70695 , n70694 );
or ( n70696 , n70690 , n70695 );
nand ( n70697 , n55887 , n70073 );
nand ( n70698 , n70696 , n70697 );
xor ( n70699 , n70689 , n70698 );
xor ( n70700 , n70677 , n70699 );
xor ( n70701 , n70700 , n70163 );
not ( n70702 , n62654 );
not ( n70703 , n61951 );
not ( n70704 , n39844 );
or ( n70705 , n70703 , n70704 );
nand ( n70706 , n58034 , n61952 );
nand ( n70707 , n70705 , n70706 );
not ( n70708 , n70707 );
or ( n70709 , n70702 , n70708 );
nand ( n70710 , n70273 , n62664 );
nand ( n70711 , n70709 , n70710 );
not ( n70712 , n52421 );
not ( n70713 , n70383 );
or ( n70714 , n70712 , n70713 );
not ( n70715 , n51723 );
not ( n70716 , n66301 );
or ( n70717 , n70715 , n70716 );
nand ( n70718 , n42555 , n51724 );
nand ( n70719 , n70717 , n70718 );
nand ( n70720 , n70719 , n54875 );
nand ( n70721 , n70714 , n70720 );
xor ( n70722 , n70711 , n70721 );
not ( n70723 , n54623 );
not ( n70724 , n59174 );
not ( n70725 , n39333 );
or ( n70726 , n70724 , n70725 );
nand ( n70727 , n39332 , n54628 );
nand ( n70728 , n70726 , n70727 );
not ( n70729 , n70728 );
or ( n70730 , n70723 , n70729 );
nand ( n70731 , n70363 , n52022 );
nand ( n70732 , n70730 , n70731 );
xor ( n70733 , n70722 , n70732 );
xor ( n70734 , n70701 , n70733 );
xor ( n70735 , n70700 , n70163 );
and ( n70736 , n70735 , n70733 );
and ( n70737 , n70700 , n70163 );
or ( n70738 , n70736 , n70737 );
not ( n70739 , n59950 );
not ( n70740 , n70311 );
or ( n70741 , n70739 , n70740 );
not ( n70742 , n59345 );
not ( n70743 , n68206 );
or ( n70744 , n70742 , n70743 );
nand ( n70745 , n39714 , n65743 );
nand ( n70746 , n70744 , n70745 );
nand ( n70747 , n70746 , n56639 );
nand ( n70748 , n70741 , n70747 );
not ( n70749 , n60927 );
not ( n70750 , n66234 );
not ( n70751 , n67040 );
or ( n70752 , n70750 , n70751 );
nand ( n70753 , n59913 , n69893 );
nand ( n70754 , n70752 , n70753 );
not ( n70755 , n70754 );
or ( n70756 , n70749 , n70755 );
nand ( n70757 , n70326 , n62085 );
nand ( n70758 , n70756 , n70757 );
xor ( n70759 , n70748 , n70758 );
xor ( n70760 , n70759 , n70092 );
not ( n70761 , n58977 );
not ( n70762 , n60602 );
not ( n70763 , n60874 );
or ( n70764 , n70762 , n70763 );
nand ( n70765 , n39056 , n62577 );
nand ( n70766 , n70764 , n70765 );
not ( n70767 , n70766 );
or ( n70768 , n70761 , n70767 );
nand ( n70769 , n70370 , n59633 );
nand ( n70770 , n70768 , n70769 );
not ( n70771 , n57314 );
not ( n70772 , n70344 );
or ( n70773 , n70771 , n70772 );
not ( n70774 , n52377 );
not ( n70775 , n66052 );
or ( n70776 , n70774 , n70775 );
nand ( n70777 , n66053 , n55013 );
nand ( n70778 , n70776 , n70777 );
nand ( n70779 , n70778 , n52004 );
nand ( n70780 , n70773 , n70779 );
xor ( n70781 , n70770 , n70780 );
not ( n70782 , n70335 );
or ( n70783 , n70782 , n50241 );
or ( n70784 , n50239 , n67477 );
nand ( n70785 , n70783 , n70784 );
xor ( n70786 , n70781 , n70785 );
xor ( n70787 , n70760 , n70786 );
xor ( n70788 , n70787 , n70169 );
xor ( n70789 , n70760 , n70786 );
and ( n70790 , n70789 , n70169 );
and ( n70791 , n70760 , n70786 );
or ( n70792 , n70790 , n70791 );
xor ( n70793 , n70550 , n70305 );
xor ( n70794 , n70793 , n70243 );
xor ( n70795 , n70550 , n70305 );
and ( n70796 , n70795 , n70243 );
and ( n70797 , n70550 , n70305 );
or ( n70798 , n70796 , n70797 );
xor ( n70799 , n70556 , n70202 );
xor ( n70800 , n70799 , n70354 );
xor ( n70801 , n70556 , n70202 );
and ( n70802 , n70801 , n70354 );
and ( n70803 , n70556 , n70202 );
or ( n70804 , n70802 , n70803 );
xor ( n70805 , n70672 , n70596 );
xor ( n70806 , n70805 , n70788 );
xor ( n70807 , n70672 , n70596 );
and ( n70808 , n70807 , n70788 );
and ( n70809 , n70672 , n70596 );
or ( n70810 , n70808 , n70809 );
xor ( n70811 , n70392 , n70734 );
xor ( n70812 , n70811 , n70398 );
xor ( n70813 , n70392 , n70734 );
and ( n70814 , n70813 , n70398 );
and ( n70815 , n70392 , n70734 );
or ( n70816 , n70814 , n70815 );
xor ( n70817 , n70687 , n70688 );
and ( n70818 , n70817 , n70698 );
and ( n70819 , n70687 , n70688 );
or ( n70820 , n70818 , n70819 );
xor ( n70821 , n70404 , n70794 );
xor ( n70822 , n70821 , n70800 );
xor ( n70823 , n70404 , n70794 );
and ( n70824 , n70823 , n70800 );
and ( n70825 , n70404 , n70794 );
or ( n70826 , n70824 , n70825 );
xor ( n70827 , n70806 , n70410 );
xor ( n70828 , n70827 , n70812 );
xor ( n70829 , n70806 , n70410 );
and ( n70830 , n70829 , n70812 );
and ( n70831 , n70806 , n70410 );
or ( n70832 , n70830 , n70831 );
xor ( n70833 , n70420 , n70426 );
xor ( n70834 , n70833 , n70822 );
xor ( n70835 , n70420 , n70426 );
and ( n70836 , n70835 , n70822 );
and ( n70837 , n70420 , n70426 );
or ( n70838 , n70836 , n70837 );
xor ( n70839 , n70828 , n70432 );
xor ( n70840 , n70839 , n70438 );
xor ( n70841 , n70828 , n70432 );
and ( n70842 , n70841 , n70438 );
and ( n70843 , n70828 , n70432 );
or ( n70844 , n70842 , n70843 );
xor ( n70845 , n70834 , n70840 );
xor ( n70846 , n70845 , n70444 );
xor ( n70847 , n70834 , n70840 );
and ( n70848 , n70847 , n70444 );
and ( n70849 , n70834 , n70840 );
or ( n70850 , n70848 , n70849 );
xor ( n70851 , n70646 , n70657 );
and ( n70852 , n70851 , n70669 );
and ( n70853 , n70646 , n70657 );
or ( n70854 , n70852 , n70853 );
xor ( n70855 , n70571 , n70582 );
and ( n70856 , n70855 , n70594 );
and ( n70857 , n70571 , n70582 );
or ( n70858 , n70856 , n70857 );
xor ( n70859 , n70612 , n70622 );
and ( n70860 , n70859 , n70634 );
and ( n70861 , n70612 , n70622 );
or ( n70862 , n70860 , n70861 );
xor ( n70863 , n70711 , n70721 );
and ( n70864 , n70863 , n70732 );
and ( n70865 , n70711 , n70721 );
or ( n70866 , n70864 , n70865 );
xor ( n70867 , n70770 , n70780 );
and ( n70868 , n70867 , n70785 );
and ( n70869 , n70770 , n70780 );
or ( n70870 , n70868 , n70869 );
xor ( n70871 , n70748 , n70758 );
and ( n70872 , n70871 , n70092 );
and ( n70873 , n70748 , n70758 );
or ( n70874 , n70872 , n70873 );
xor ( n70875 , n70127 , n70414 );
and ( n70876 , n70875 , n70699 );
and ( n70877 , n70127 , n70414 );
or ( n70878 , n70876 , n70877 );
not ( n70879 , n50239 );
not ( n70880 , n50241 );
or ( n70881 , n70879 , n70880 );
nand ( n70882 , n70881 , n48645 );
not ( n70883 , n70533 );
not ( n70884 , n56777 );
or ( n70885 , n70883 , n70884 );
not ( n70886 , n69820 );
not ( n70887 , n52076 );
or ( n70888 , n70886 , n70887 );
not ( n70889 , n52076 );
nand ( n70890 , n70889 , n67454 );
nand ( n70891 , n70888 , n70890 );
nand ( n70892 , n56780 , n70891 );
nand ( n70893 , n70885 , n70892 );
xor ( n70894 , n70882 , n70893 );
or ( n70895 , n70610 , n66006 );
and ( n70896 , n64452 , n66963 );
not ( n70897 , n64452 );
and ( n70898 , n70897 , n67568 );
nor ( n70899 , n70896 , n70898 );
or ( n70900 , n69648 , n70899 );
nand ( n70901 , n70895 , n70900 );
xor ( n70902 , n70894 , n70901 );
xor ( n70903 , n70882 , n70893 );
and ( n70904 , n70903 , n70901 );
and ( n70905 , n70882 , n70893 );
or ( n70906 , n70904 , n70905 );
or ( n70907 , n64143 , n70483 );
not ( n70908 , n41216 );
and ( n70909 , n66652 , n70908 );
and ( n70910 , n58642 , n70095 );
nor ( n70911 , n70909 , n70910 );
or ( n70912 , n64146 , n70911 );
nand ( n70913 , n70907 , n70912 );
not ( n70914 , n70494 );
not ( n70915 , n66980 );
not ( n70916 , n70915 );
or ( n70917 , n70914 , n70916 );
and ( n70918 , n49190 , n66985 );
not ( n70919 , n49190 );
buf ( n70920 , n63587 );
and ( n70921 , n70919 , n70920 );
nor ( n70922 , n70918 , n70921 );
not ( n70923 , n70922 );
nand ( n70924 , n70923 , n60542 );
nand ( n70925 , n70917 , n70924 );
xor ( n70926 , n70913 , n70925 );
not ( n70927 , n70508 );
not ( n70928 , n70500 );
or ( n70929 , n70927 , n70928 );
buf ( n70930 , n66602 );
not ( n70931 , n41532 );
not ( n70932 , n66141 );
or ( n70933 , n70931 , n70932 );
nand ( n70934 , n68878 , n69270 );
nand ( n70935 , n70933 , n70934 );
nand ( n70936 , n70930 , n70935 );
nand ( n70937 , n70929 , n70936 );
xor ( n70938 , n70926 , n70937 );
xor ( n70939 , n70913 , n70925 );
and ( n70940 , n70939 , n70937 );
and ( n70941 , n70913 , n70925 );
or ( n70942 , n70940 , n70941 );
not ( n70943 , n70523 );
not ( n70944 , n61550 );
or ( n70945 , n70943 , n70944 );
not ( n70946 , n58458 );
not ( n70947 , n61537 );
or ( n70948 , n70946 , n70947 );
nand ( n70949 , n66615 , n58459 );
nand ( n70950 , n70948 , n70949 );
nand ( n70951 , n67094 , n70950 );
nand ( n70952 , n70945 , n70951 );
or ( n70953 , n64684 , n70541 );
and ( n70954 , n47527 , n62452 );
not ( n70955 , n47527 );
and ( n70956 , n70955 , n64170 );
nor ( n70957 , n70954 , n70956 );
or ( n70958 , n69703 , n70957 );
nand ( n70959 , n70953 , n70958 );
xor ( n70960 , n70952 , n70959 );
not ( n70961 , n65795 );
not ( n70962 , n70685 );
or ( n70963 , n70961 , n70962 );
buf ( n70964 , n63398 );
not ( n70965 , n70964 );
not ( n70966 , n63922 );
not ( n70967 , n56731 );
and ( n70968 , n70966 , n70967 );
and ( n70969 , n63922 , n56731 );
nor ( n70970 , n70968 , n70969 );
or ( n70971 , n70965 , n70970 );
nand ( n70972 , n70963 , n70971 );
xor ( n70973 , n70960 , n70972 );
xor ( n70974 , n70973 , n70938 );
xor ( n70975 , n70974 , n70820 );
xor ( n70976 , n70973 , n70938 );
and ( n70977 , n70976 , n70820 );
and ( n70978 , n70973 , n70938 );
or ( n70979 , n70977 , n70978 );
xor ( n70980 , n70858 , n70862 );
xor ( n70981 , n70980 , n70854 );
xor ( n70982 , n70858 , n70862 );
and ( n70983 , n70982 , n70854 );
and ( n70984 , n70858 , n70862 );
or ( n70985 , n70983 , n70984 );
xor ( n70986 , n70866 , n70874 );
not ( n70987 , n54364 );
not ( n70988 , n53596 );
not ( n70989 , n63656 );
or ( n70990 , n70988 , n70989 );
not ( n70991 , n53615 );
nand ( n70992 , n59612 , n70991 );
nand ( n70993 , n70990 , n70992 );
not ( n70994 , n70993 );
or ( n70995 , n70987 , n70994 );
nand ( n70996 , n70620 , n68603 );
nand ( n70997 , n70995 , n70996 );
not ( n70998 , n54327 );
not ( n70999 , n54323 );
not ( n71000 , n66798 );
or ( n71001 , n70999 , n71000 );
nand ( n71002 , n40592 , n54468 );
nand ( n71003 , n71001 , n71002 );
not ( n71004 , n71003 );
or ( n71005 , n70998 , n71004 );
nand ( n71006 , n70632 , n54316 );
nand ( n71007 , n71005 , n71006 );
xor ( n71008 , n70997 , n71007 );
not ( n71009 , n62654 );
not ( n71010 , n61951 );
not ( n71011 , n59414 );
or ( n71012 , n71010 , n71011 );
not ( n71013 , n39895 );
nand ( n71014 , n71013 , n66690 );
nand ( n71015 , n71012 , n71014 );
not ( n71016 , n71015 );
or ( n71017 , n71009 , n71016 );
nand ( n71018 , n70707 , n66696 );
nand ( n71019 , n71017 , n71018 );
xor ( n71020 , n71008 , n71019 );
xor ( n71021 , n70986 , n71020 );
xor ( n71022 , n70866 , n70874 );
and ( n71023 , n71022 , n71020 );
and ( n71024 , n70866 , n70874 );
or ( n71025 , n71023 , n71024 );
not ( n71026 , n70183 );
not ( n71027 , n55582 );
not ( n71028 , n70278 );
or ( n71029 , n71027 , n71028 );
nand ( n71030 , n69442 , n55148 );
nand ( n71031 , n71029 , n71030 );
not ( n71032 , n71031 );
or ( n71033 , n71026 , n71032 );
nand ( n71034 , n70642 , n70193 );
nand ( n71035 , n71033 , n71034 );
not ( n71036 , n52151 );
not ( n71037 , n70665 );
or ( n71038 , n71036 , n71037 );
not ( n71039 , n51465 );
not ( n71040 , n70290 );
or ( n71041 , n71039 , n71040 );
not ( n71042 , n50895 );
nand ( n71043 , n67721 , n71042 );
nand ( n71044 , n71041 , n71043 );
nand ( n71045 , n71044 , n51223 );
nand ( n71046 , n71038 , n71045 );
xor ( n71047 , n71035 , n71046 );
not ( n71048 , n51533 );
not ( n71049 , n53931 );
not ( n71050 , n59694 );
or ( n71051 , n71049 , n71050 );
not ( n71052 , n65725 );
not ( n71053 , n53931 );
nand ( n71054 , n71052 , n71053 );
nand ( n71055 , n71051 , n71054 );
not ( n71056 , n71055 );
or ( n71057 , n71048 , n71056 );
nand ( n71058 , n70567 , n56355 );
nand ( n71059 , n71057 , n71058 );
xor ( n71060 , n71047 , n71059 );
not ( n71061 , n53197 );
not ( n71062 , n70580 );
or ( n71063 , n71061 , n71062 );
not ( n71064 , n68931 );
not ( n71065 , n40148 );
or ( n71066 , n71064 , n71065 );
not ( n71067 , n54402 );
nand ( n71068 , n71067 , n52113 );
nand ( n71069 , n71066 , n71068 );
nand ( n71070 , n71069 , n51766 );
nand ( n71071 , n71063 , n71070 );
not ( n71072 , n55104 );
not ( n71073 , n56074 );
not ( n71074 , n71073 );
or ( n71075 , n71072 , n71074 );
not ( n71076 , n59601 );
nand ( n71077 , n71076 , n52840 );
nand ( n71078 , n71075 , n71077 );
not ( n71079 , n71078 );
not ( n71080 , n52469 );
or ( n71081 , n71079 , n71080 );
nand ( n71082 , n53182 , n70591 );
nand ( n71083 , n71081 , n71082 );
xor ( n71084 , n71071 , n71083 );
not ( n71085 , n70612 );
xor ( n71086 , n71084 , n71085 );
xor ( n71087 , n71060 , n71086 );
and ( n71088 , n67072 , n70173 );
not ( n71089 , n59984 );
not ( n71090 , n55872 );
not ( n71091 , n52286 );
or ( n71092 , n71090 , n71091 );
not ( n71093 , n52286 );
not ( n71094 , n55872 );
nand ( n71095 , n71093 , n71094 );
nand ( n71096 , n71092 , n71095 );
not ( n71097 , n71096 );
or ( n71098 , n71089 , n71097 );
not ( n71099 , n69028 );
nand ( n71100 , n70694 , n71099 );
nand ( n71101 , n71098 , n71100 );
xor ( n71102 , n71088 , n71101 );
not ( n71103 , n52749 );
not ( n71104 , n70655 );
or ( n71105 , n71103 , n71104 );
not ( n71106 , n59651 );
not ( n71107 , n50306 );
or ( n71108 , n71106 , n71107 );
nand ( n71109 , n39964 , n66705 );
nand ( n71110 , n71108 , n71109 );
nand ( n71111 , n71110 , n52757 );
nand ( n71112 , n71105 , n71111 );
xor ( n71113 , n71102 , n71112 );
xor ( n71114 , n71087 , n71113 );
xor ( n71115 , n71060 , n71086 );
and ( n71116 , n71115 , n71113 );
and ( n71117 , n71060 , n71086 );
or ( n71118 , n71116 , n71117 );
xor ( n71119 , n70515 , n70548 );
xor ( n71120 , n71119 , n70902 );
xor ( n71121 , n70870 , n71120 );
xor ( n71122 , n71121 , n70878 );
xor ( n71123 , n70870 , n71120 );
and ( n71124 , n71123 , n70878 );
and ( n71125 , n70870 , n71120 );
or ( n71126 , n71124 , n71125 );
not ( n71127 , n56639 );
not ( n71128 , n59345 );
not ( n71129 , n65532 );
or ( n71130 , n71128 , n71129 );
nand ( n71131 , n39574 , n60617 );
nand ( n71132 , n71130 , n71131 );
not ( n71133 , n71132 );
or ( n71134 , n71127 , n71133 );
nand ( n71135 , n70746 , n59950 );
nand ( n71136 , n71134 , n71135 );
not ( n71137 , n52004 );
not ( n71138 , n52377 );
not ( n71139 , n68381 );
not ( n71140 , n71139 );
or ( n71141 , n71138 , n71140 );
nand ( n71142 , n68381 , n55013 );
nand ( n71143 , n71141 , n71142 );
not ( n71144 , n71143 );
or ( n71145 , n71137 , n71144 );
nand ( n71146 , n70778 , n48894 );
nand ( n71147 , n71145 , n71146 );
xor ( n71148 , n71136 , n71147 );
not ( n71149 , n52191 );
not ( n71150 , n62077 );
not ( n71151 , n58482 );
or ( n71152 , n71150 , n71151 );
nand ( n71153 , n60386 , n60289 );
nand ( n71154 , n71152 , n71153 );
not ( n71155 , n71154 );
or ( n71156 , n71149 , n71155 );
nand ( n71157 , n70754 , n58168 );
nand ( n71158 , n71156 , n71157 );
xor ( n71159 , n71148 , n71158 );
not ( n71160 , n54875 );
not ( n71161 , n51723 );
buf ( n71162 , n42651 );
not ( n71163 , n71162 );
not ( n71164 , n71163 );
or ( n71165 , n71161 , n71164 );
nand ( n71166 , n71162 , n51724 );
nand ( n71167 , n71165 , n71166 );
not ( n71168 , n71167 );
or ( n71169 , n71160 , n71168 );
nand ( n71170 , n70719 , n52421 );
nand ( n71171 , n71169 , n71170 );
not ( n71172 , n52022 );
not ( n71173 , n70728 );
or ( n71174 , n71172 , n71173 );
not ( n71175 , n59174 );
not ( n71176 , n69530 );
not ( n71177 , n71176 );
or ( n71178 , n71175 , n71177 );
nand ( n71179 , n69530 , n54628 );
nand ( n71180 , n71178 , n71179 );
nand ( n71181 , n71180 , n54623 );
nand ( n71182 , n71174 , n71181 );
xor ( n71183 , n71171 , n71182 );
not ( n71184 , n58977 );
and ( n71185 , n60602 , n38499 );
not ( n71186 , n60602 );
and ( n71187 , n71186 , n68652 );
nor ( n71188 , n71185 , n71187 );
not ( n71189 , n71188 );
or ( n71190 , n71184 , n71189 );
nand ( n71191 , n70766 , n53104 );
nand ( n71192 , n71190 , n71191 );
xor ( n71193 , n71183 , n71192 );
xor ( n71194 , n71159 , n71193 );
xor ( n71195 , n71194 , n70560 );
xor ( n71196 , n71159 , n71193 );
and ( n71197 , n71196 , n70560 );
and ( n71198 , n71159 , n71193 );
or ( n71199 , n71197 , n71198 );
xor ( n71200 , n70554 , n70975 );
xor ( n71201 , n71200 , n70600 );
xor ( n71202 , n70554 , n70975 );
and ( n71203 , n71202 , n70600 );
and ( n71204 , n70554 , n70975 );
or ( n71205 , n71203 , n71204 );
xor ( n71206 , n70676 , n70981 );
xor ( n71207 , n71206 , n71114 );
xor ( n71208 , n70676 , n70981 );
and ( n71209 , n71208 , n71114 );
and ( n71210 , n70676 , n70981 );
or ( n71211 , n71209 , n71210 );
xor ( n71212 , n71021 , n70738 );
xor ( n71213 , n71212 , n70792 );
xor ( n71214 , n71021 , n70738 );
and ( n71215 , n71214 , n70792 );
and ( n71216 , n71021 , n70738 );
or ( n71217 , n71215 , n71216 );
xor ( n71218 , n71195 , n71122 );
xor ( n71219 , n71218 , n70798 );
xor ( n71220 , n71195 , n71122 );
and ( n71221 , n71220 , n70798 );
and ( n71222 , n71195 , n71122 );
or ( n71223 , n71221 , n71222 );
xor ( n71224 , n70952 , n70959 );
and ( n71225 , n71224 , n70972 );
and ( n71226 , n70952 , n70959 );
or ( n71227 , n71225 , n71226 );
xor ( n71228 , n71201 , n70804 );
xor ( n71229 , n71228 , n71207 );
xor ( n71230 , n71201 , n70804 );
and ( n71231 , n71230 , n71207 );
and ( n71232 , n71201 , n70804 );
or ( n71233 , n71231 , n71232 );
xor ( n71234 , n70810 , n71213 );
xor ( n71235 , n71234 , n71219 );
xor ( n71236 , n70810 , n71213 );
and ( n71237 , n71236 , n71219 );
and ( n71238 , n70810 , n71213 );
or ( n71239 , n71237 , n71238 );
xor ( n71240 , n70816 , n70826 );
xor ( n71241 , n71240 , n71229 );
xor ( n71242 , n70816 , n70826 );
and ( n71243 , n71242 , n71229 );
and ( n71244 , n70816 , n70826 );
or ( n71245 , n71243 , n71244 );
xor ( n71246 , n71235 , n70832 );
xor ( n71247 , n71246 , n70838 );
xor ( n71248 , n71235 , n70832 );
and ( n71249 , n71248 , n70838 );
and ( n71250 , n71235 , n70832 );
or ( n71251 , n71249 , n71250 );
xor ( n71252 , n71241 , n71247 );
xor ( n71253 , n71252 , n70844 );
xor ( n71254 , n71241 , n71247 );
and ( n71255 , n71254 , n70844 );
and ( n71256 , n71241 , n71247 );
or ( n71257 , n71255 , n71256 );
xor ( n71258 , n71088 , n71101 );
and ( n71259 , n71258 , n71112 );
and ( n71260 , n71088 , n71101 );
or ( n71261 , n71259 , n71260 );
xor ( n71262 , n71035 , n71046 );
and ( n71263 , n71262 , n71059 );
and ( n71264 , n71035 , n71046 );
or ( n71265 , n71263 , n71264 );
xor ( n71266 , n71071 , n71083 );
and ( n71267 , n71266 , n71085 );
and ( n71268 , n71071 , n71083 );
or ( n71269 , n71267 , n71268 );
xor ( n71270 , n70997 , n71007 );
and ( n71271 , n71270 , n71019 );
and ( n71272 , n70997 , n71007 );
or ( n71273 , n71271 , n71272 );
xor ( n71274 , n71171 , n71182 );
and ( n71275 , n71274 , n71192 );
and ( n71276 , n71171 , n71182 );
or ( n71277 , n71275 , n71276 );
xor ( n71278 , n71136 , n71147 );
and ( n71279 , n71278 , n71158 );
and ( n71280 , n71136 , n71147 );
or ( n71281 , n71279 , n71280 );
xor ( n71282 , n70515 , n70548 );
and ( n71283 , n71282 , n70902 );
and ( n71284 , n70515 , n70548 );
or ( n71285 , n71283 , n71284 );
or ( n71286 , n67584 , n70922 );
and ( n71287 , n41286 , n63587 );
not ( n71288 , n41286 );
and ( n71289 , n71288 , n62513 );
nor ( n71290 , n71287 , n71289 );
or ( n71291 , n67586 , n71290 );
nand ( n71292 , n71286 , n71291 );
not ( n71293 , n70935 );
not ( n71294 , n70500 );
or ( n71295 , n71293 , n71294 );
not ( n71296 , n48486 );
not ( n71297 , n60286 );
or ( n71298 , n71296 , n71297 );
nand ( n71299 , n70506 , n64972 );
nand ( n71300 , n71298 , n71299 );
nand ( n71301 , n70930 , n71300 );
nand ( n71302 , n71295 , n71301 );
xor ( n71303 , n71292 , n71302 );
not ( n71304 , n64111 );
not ( n71305 , n70950 );
or ( n71306 , n71304 , n71305 );
not ( n71307 , n61540 );
and ( n71308 , n71307 , n58915 );
not ( n71309 , n64630 );
and ( n71310 , n71309 , n58914 );
nor ( n71311 , n71308 , n71310 );
or ( n71312 , n65144 , n71311 );
nand ( n71313 , n71306 , n71312 );
xor ( n71314 , n71303 , n71313 );
xor ( n71315 , n71292 , n71302 );
and ( n71316 , n71315 , n71313 );
and ( n71317 , n71292 , n71302 );
or ( n71318 , n71316 , n71317 );
or ( n71319 , n64164 , n70957 );
and ( n71320 , n58994 , n69704 );
not ( n71321 , n58994 );
and ( n71322 , n71321 , n62449 );
nor ( n71323 , n71320 , n71322 );
or ( n71324 , n64166 , n71323 );
nand ( n71325 , n71319 , n71324 );
not ( n71326 , n70899 );
not ( n71327 , n71326 );
not ( n71328 , n60482 );
or ( n71329 , n71327 , n71328 );
not ( n71330 , n51891 );
not ( n71331 , n71330 );
not ( n71332 , n71331 );
not ( n71333 , n70608 );
or ( n71334 , n71332 , n71333 );
nand ( n71335 , n66642 , n50020 );
nand ( n71336 , n71334 , n71335 );
nand ( n71337 , n70604 , n71336 );
nand ( n71338 , n71329 , n71337 );
xor ( n71339 , n71325 , n71338 );
not ( n71340 , n70970 );
not ( n71341 , n71340 );
not ( n71342 , n65089 );
or ( n71343 , n71341 , n71342 );
not ( n71344 , n57182 );
not ( n71345 , n63412 );
or ( n71346 , n71344 , n71345 );
nand ( n71347 , n67072 , n57186 );
nand ( n71348 , n71346 , n71347 );
nand ( n71349 , n70964 , n71348 );
nand ( n71350 , n71343 , n71349 );
xor ( n71351 , n71339 , n71350 );
xor ( n71352 , n71325 , n71338 );
and ( n71353 , n71352 , n71350 );
and ( n71354 , n71325 , n71338 );
or ( n71355 , n71353 , n71354 );
and ( n71356 , n64444 , n48983 );
not ( n71357 , n60472 );
not ( n71358 , n56786 );
not ( n71359 , n50654 );
or ( n71360 , n71358 , n71359 );
not ( n71361 , n51841 );
buf ( n71362 , n67454 );
nand ( n71363 , n71361 , n71362 );
nand ( n71364 , n71360 , n71363 );
not ( n71365 , n71364 );
or ( n71366 , n71357 , n71365 );
nand ( n71367 , n56777 , n70891 );
nand ( n71368 , n71366 , n71367 );
xor ( n71369 , n71356 , n71368 );
not ( n71370 , n59984 );
not ( n71371 , n55873 );
not ( n71372 , n71371 );
not ( n71373 , n40735 );
or ( n71374 , n71372 , n71373 );
nand ( n71375 , n54032 , n69237 );
nand ( n71376 , n71374 , n71375 );
not ( n71377 , n71376 );
or ( n71378 , n71370 , n71377 );
nand ( n71379 , n71096 , n67862 );
nand ( n71380 , n71378 , n71379 );
xor ( n71381 , n71369 , n71380 );
xor ( n71382 , n71269 , n71381 );
xor ( n71383 , n71382 , n71261 );
xor ( n71384 , n71269 , n71381 );
and ( n71385 , n71384 , n71261 );
and ( n71386 , n71269 , n71381 );
or ( n71387 , n71385 , n71386 );
xor ( n71388 , n71265 , n71273 );
xor ( n71389 , n71388 , n71277 );
xor ( n71390 , n71265 , n71273 );
and ( n71391 , n71390 , n71277 );
and ( n71392 , n71265 , n71273 );
or ( n71393 , n71391 , n71392 );
not ( n71394 , n54327 );
not ( n71395 , n54302 );
not ( n71396 , n71395 );
not ( n71397 , n52432 );
or ( n71398 , n71396 , n71397 );
nand ( n71399 , n68049 , n55276 );
nand ( n71400 , n71398 , n71399 );
not ( n71401 , n71400 );
or ( n71402 , n71394 , n71401 );
nand ( n71403 , n71003 , n54316 );
nand ( n71404 , n71402 , n71403 );
not ( n71405 , n70183 );
not ( n71406 , n55582 );
not ( n71407 , n52570 );
or ( n71408 , n71406 , n71407 );
not ( n71409 , n55120 );
nand ( n71410 , n51916 , n71409 );
nand ( n71411 , n71408 , n71410 );
not ( n71412 , n71411 );
or ( n71413 , n71405 , n71412 );
nand ( n71414 , n71031 , n70193 );
nand ( n71415 , n71413 , n71414 );
xor ( n71416 , n71404 , n71415 );
not ( n71417 , n52757 );
buf ( n71418 , n39844 );
and ( n71419 , n71418 , n64190 );
not ( n71420 , n71418 );
and ( n71421 , n71420 , n66705 );
or ( n71422 , n71419 , n71421 );
not ( n71423 , n71422 );
or ( n71424 , n71417 , n71423 );
nand ( n71425 , n71110 , n52749 );
nand ( n71426 , n71424 , n71425 );
xor ( n71427 , n71416 , n71426 );
not ( n71428 , n52151 );
not ( n71429 , n71044 );
or ( n71430 , n71428 , n71429 );
not ( n71431 , n65773 );
not ( n71432 , n63180 );
or ( n71433 , n71431 , n71432 );
nand ( n71434 , n70653 , n50916 );
nand ( n71435 , n71433 , n71434 );
nand ( n71436 , n71435 , n50922 );
nand ( n71437 , n71430 , n71436 );
not ( n71438 , n56355 );
not ( n71439 , n71055 );
or ( n71440 , n71438 , n71439 );
not ( n71441 , n53931 );
not ( n71442 , n68980 );
not ( n71443 , n71442 );
or ( n71444 , n71441 , n71443 );
not ( n71445 , n65103 );
nand ( n71446 , n68980 , n71445 );
nand ( n71447 , n71444 , n71446 );
nand ( n71448 , n71447 , n51533 );
nand ( n71449 , n71440 , n71448 );
xor ( n71450 , n71437 , n71449 );
not ( n71451 , n51766 );
not ( n71452 , n68931 );
not ( n71453 , n68991 );
or ( n71454 , n71452 , n71453 );
nand ( n71455 , n68994 , n52130 );
nand ( n71456 , n71454 , n71455 );
not ( n71457 , n71456 );
or ( n71458 , n71451 , n71457 );
nand ( n71459 , n71069 , n53197 );
nand ( n71460 , n71458 , n71459 );
xor ( n71461 , n71450 , n71460 );
xor ( n71462 , n71427 , n71461 );
not ( n71463 , n63079 );
not ( n71464 , n70911 );
and ( n71465 , n71463 , n71464 );
buf ( n71466 , n61465 );
not ( n71467 , n71466 );
and ( n71468 , n40854 , n65183 );
not ( n71469 , n40854 );
and ( n71470 , n71469 , n58642 );
nor ( n71471 , n71468 , n71470 );
nor ( n71472 , n71467 , n71471 );
nor ( n71473 , n71465 , n71472 );
not ( n71474 , n52469 );
not ( n71475 , n54283 );
buf ( n71476 , n63201 );
not ( n71477 , n71476 );
or ( n71478 , n71475 , n71477 );
buf ( n71479 , n59195 );
nand ( n71480 , n71479 , n55104 );
nand ( n71481 , n71478 , n71480 );
not ( n71482 , n71481 );
or ( n71483 , n71474 , n71482 );
nand ( n71484 , n71078 , n52854 );
nand ( n71485 , n71483 , n71484 );
xor ( n71486 , n71473 , n71485 );
not ( n71487 , n68603 );
not ( n71488 , n70993 );
or ( n71489 , n71487 , n71488 );
not ( n71490 , n53596 );
not ( n71491 , n54020 );
or ( n71492 , n71490 , n71491 );
nand ( n71493 , n54646 , n70991 );
nand ( n71494 , n71492 , n71493 );
nand ( n71495 , n71494 , n53620 );
nand ( n71496 , n71489 , n71495 );
xor ( n71497 , n71486 , n71496 );
xor ( n71498 , n71462 , n71497 );
xor ( n71499 , n71427 , n71461 );
and ( n71500 , n71499 , n71497 );
and ( n71501 , n71427 , n71461 );
or ( n71502 , n71500 , n71501 );
not ( n71503 , n66696 );
not ( n71504 , n71015 );
or ( n71505 , n71503 , n71504 );
not ( n71506 , n61951 );
not ( n71507 , n67040 );
or ( n71508 , n71506 , n71507 );
not ( n71509 , n67037 );
nand ( n71510 , n71509 , n61952 );
nand ( n71511 , n71508 , n71510 );
nand ( n71512 , n71511 , n62654 );
nand ( n71513 , n71505 , n71512 );
xor ( n71514 , n70906 , n71513 );
xor ( n71515 , n71514 , n70942 );
xor ( n71516 , n71281 , n71515 );
xor ( n71517 , n71516 , n70979 );
xor ( n71518 , n71281 , n71515 );
and ( n71519 , n71518 , n70979 );
and ( n71520 , n71281 , n71515 );
or ( n71521 , n71519 , n71520 );
not ( n71522 , n52004 );
and ( n71523 , n55013 , n67269 );
not ( n71524 , n55013 );
not ( n71525 , n67269 );
and ( n71526 , n71524 , n71525 );
nor ( n71527 , n71523 , n71526 );
not ( n71528 , n71527 );
or ( n71529 , n71522 , n71528 );
nand ( n71530 , n71143 , n48894 );
nand ( n71531 , n71529 , n71530 );
not ( n71532 , n59633 );
not ( n71533 , n71188 );
or ( n71534 , n71532 , n71533 );
not ( n71535 , n60602 );
not ( n71536 , n60855 );
or ( n71537 , n71535 , n71536 );
nand ( n71538 , n39332 , n52728 );
nand ( n71539 , n71537 , n71538 );
nand ( n71540 , n71539 , n58977 );
nand ( n71541 , n71534 , n71540 );
xor ( n71542 , n71531 , n71541 );
not ( n71543 , n56639 );
not ( n71544 , n59345 );
not ( n71545 , n59891 );
or ( n71546 , n71544 , n71545 );
not ( n71547 , n59891 );
nand ( n71548 , n71547 , n65743 );
nand ( n71549 , n71546 , n71548 );
not ( n71550 , n71549 );
or ( n71551 , n71543 , n71550 );
nand ( n71552 , n71132 , n59950 );
nand ( n71553 , n71551 , n71552 );
xor ( n71554 , n71542 , n71553 );
xor ( n71555 , n71285 , n71554 );
not ( n71556 , n52421 );
not ( n71557 , n71167 );
or ( n71558 , n71556 , n71557 );
nand ( n71559 , n54875 , n51723 );
nand ( n71560 , n71558 , n71559 );
not ( n71561 , n62085 );
not ( n71562 , n71154 );
or ( n71563 , n71561 , n71562 );
not ( n71564 , n66234 );
not ( n71565 , n68206 );
or ( n71566 , n71564 , n71565 );
not ( n71567 , n68206 );
nand ( n71568 , n71567 , n69893 );
nand ( n71569 , n71566 , n71568 );
nand ( n71570 , n71569 , n52191 );
nand ( n71571 , n71563 , n71570 );
xor ( n71572 , n71560 , n71571 );
not ( n71573 , n54623 );
not ( n71574 , n59174 );
not ( n71575 , n69961 );
or ( n71576 , n71574 , n71575 );
not ( n71577 , n62909 );
nand ( n71578 , n71577 , n54628 );
nand ( n71579 , n71576 , n71578 );
not ( n71580 , n71579 );
or ( n71581 , n71573 , n71580 );
nand ( n71582 , n71180 , n52022 );
nand ( n71583 , n71581 , n71582 );
xor ( n71584 , n71572 , n71583 );
xor ( n71585 , n71555 , n71584 );
xor ( n71586 , n71285 , n71554 );
and ( n71587 , n71586 , n71584 );
and ( n71588 , n71285 , n71554 );
or ( n71589 , n71587 , n71588 );
xor ( n71590 , n71227 , n71351 );
xor ( n71591 , n71590 , n71314 );
xor ( n71592 , n70985 , n71591 );
xor ( n71593 , n71592 , n71118 );
xor ( n71594 , n70985 , n71591 );
and ( n71595 , n71594 , n71118 );
and ( n71596 , n70985 , n71591 );
or ( n71597 , n71595 , n71596 );
xor ( n71598 , n71025 , n71383 );
xor ( n71599 , n71598 , n71389 );
xor ( n71600 , n71025 , n71383 );
and ( n71601 , n71600 , n71389 );
and ( n71602 , n71025 , n71383 );
or ( n71603 , n71601 , n71602 );
xor ( n71604 , n71126 , n71498 );
xor ( n71605 , n71604 , n71199 );
xor ( n71606 , n71126 , n71498 );
and ( n71607 , n71606 , n71199 );
and ( n71608 , n71126 , n71498 );
or ( n71609 , n71607 , n71608 );
xor ( n71610 , n71585 , n71517 );
xor ( n71611 , n71610 , n71205 );
xor ( n71612 , n71585 , n71517 );
and ( n71613 , n71612 , n71205 );
and ( n71614 , n71585 , n71517 );
or ( n71615 , n71613 , n71614 );
xor ( n71616 , n71593 , n71599 );
xor ( n71617 , n71616 , n71211 );
xor ( n71618 , n71593 , n71599 );
and ( n71619 , n71618 , n71211 );
and ( n71620 , n71593 , n71599 );
or ( n71621 , n71619 , n71620 );
xor ( n71622 , n71356 , n71368 );
and ( n71623 , n71622 , n71380 );
and ( n71624 , n71356 , n71368 );
or ( n71625 , n71623 , n71624 );
xor ( n71626 , n71217 , n71605 );
xor ( n71627 , n71626 , n71223 );
xor ( n71628 , n71217 , n71605 );
and ( n71629 , n71628 , n71223 );
and ( n71630 , n71217 , n71605 );
or ( n71631 , n71629 , n71630 );
xor ( n71632 , n71611 , n71233 );
xor ( n71633 , n71632 , n71617 );
xor ( n71634 , n71611 , n71233 );
and ( n71635 , n71634 , n71617 );
and ( n71636 , n71611 , n71233 );
or ( n71637 , n71635 , n71636 );
xor ( n71638 , n71627 , n71239 );
xor ( n71639 , n71638 , n71245 );
xor ( n71640 , n71627 , n71239 );
and ( n71641 , n71640 , n71245 );
and ( n71642 , n71627 , n71239 );
or ( n71643 , n71641 , n71642 );
xor ( n71644 , n71633 , n71639 );
xor ( n71645 , n71644 , n71251 );
xor ( n71646 , n71633 , n71639 );
and ( n71647 , n71646 , n71251 );
and ( n71648 , n71633 , n71639 );
or ( n71649 , n71647 , n71648 );
xor ( n71650 , n71437 , n71449 );
and ( n71651 , n71650 , n71460 );
and ( n71652 , n71437 , n71449 );
or ( n71653 , n71651 , n71652 );
xor ( n71654 , n71473 , n71485 );
and ( n71655 , n71654 , n71496 );
and ( n71656 , n71473 , n71485 );
or ( n71657 , n71655 , n71656 );
xor ( n71658 , n71404 , n71415 );
and ( n71659 , n71658 , n71426 );
and ( n71660 , n71404 , n71415 );
or ( n71661 , n71659 , n71660 );
xor ( n71662 , n71531 , n71541 );
and ( n71663 , n71662 , n71553 );
and ( n71664 , n71531 , n71541 );
or ( n71665 , n71663 , n71664 );
xor ( n71666 , n71560 , n71571 );
and ( n71667 , n71666 , n71583 );
and ( n71668 , n71560 , n71571 );
or ( n71669 , n71667 , n71668 );
xor ( n71670 , n70906 , n71513 );
and ( n71671 , n71670 , n70942 );
and ( n71672 , n70906 , n71513 );
or ( n71673 , n71671 , n71672 );
xor ( n71674 , n71227 , n71351 );
and ( n71675 , n71674 , n71314 );
and ( n71676 , n71227 , n71351 );
or ( n71677 , n71675 , n71676 );
or ( n71678 , n52421 , n54875 );
nand ( n71679 , n71678 , n51723 );
not ( n71680 , n71336 );
or ( n71681 , n67885 , n71680 );
and ( n71682 , n67890 , n52079 );
not ( n71683 , n67890 );
and ( n71684 , n71683 , n53513 );
nor ( n71685 , n71682 , n71684 );
or ( n71686 , n71685 , n65638 );
nand ( n71687 , n71681 , n71686 );
xor ( n71688 , n71679 , n71687 );
not ( n71689 , n65646 );
or ( n71690 , n71689 , n71471 );
buf ( n71691 , n52916 );
and ( n71692 , n71691 , n65183 );
not ( n71693 , n71691 );
and ( n71694 , n71693 , n62496 );
or ( n71695 , n71692 , n71694 );
not ( n71696 , n71695 );
or ( n71697 , n64146 , n71696 );
nand ( n71698 , n71690 , n71697 );
xor ( n71699 , n71688 , n71698 );
xor ( n71700 , n71679 , n71687 );
and ( n71701 , n71700 , n71698 );
and ( n71702 , n71679 , n71687 );
or ( n71703 , n71701 , n71702 );
not ( n71704 , n71290 );
not ( n71705 , n71704 );
not ( n71706 , n62506 );
or ( n71707 , n71705 , n71706 );
not ( n71708 , n70908 );
not ( n71709 , n66983 );
or ( n71710 , n71708 , n71709 );
not ( n71711 , n59340 );
nand ( n71712 , n71711 , n50387 );
nand ( n71713 , n71710 , n71712 );
nand ( n71714 , n59575 , n71713 );
nand ( n71715 , n71707 , n71714 );
not ( n71716 , n71300 );
not ( n71717 , n70500 );
or ( n71718 , n71716 , n71717 );
not ( n71719 , n67441 );
not ( n71720 , n67084 );
or ( n71721 , n71719 , n71720 );
nand ( n71722 , n70506 , n49820 );
nand ( n71723 , n71721 , n71722 );
nand ( n71724 , n60427 , n71723 );
nand ( n71725 , n71718 , n71724 );
xor ( n71726 , n71715 , n71725 );
or ( n71727 , n69728 , n71311 );
and ( n71728 , n41532 , n61939 );
not ( n71729 , n41532 );
and ( n71730 , n71729 , n71309 );
or ( n71731 , n71728 , n71730 );
not ( n71732 , n71731 );
or ( n71733 , n65144 , n71732 );
nand ( n71734 , n71727 , n71733 );
xor ( n71735 , n71726 , n71734 );
xor ( n71736 , n71715 , n71725 );
and ( n71737 , n71736 , n71734 );
and ( n71738 , n71715 , n71725 );
or ( n71739 , n71737 , n71738 );
xor ( n71740 , n71735 , n71625 );
xor ( n71741 , n71740 , n71653 );
xor ( n71742 , n71735 , n71625 );
and ( n71743 , n71742 , n71653 );
and ( n71744 , n71735 , n71625 );
or ( n71745 , n71743 , n71744 );
xor ( n71746 , n71657 , n71661 );
xor ( n71747 , n71746 , n71665 );
xor ( n71748 , n71657 , n71661 );
and ( n71749 , n71748 , n71665 );
and ( n71750 , n71657 , n71661 );
or ( n71751 , n71749 , n71750 );
not ( n71752 , n53620 );
not ( n71753 , n55089 );
not ( n71754 , n40225 );
or ( n71755 , n71753 , n71754 );
not ( n71756 , n53596 );
nand ( n71757 , n53660 , n71756 );
nand ( n71758 , n71755 , n71757 );
not ( n71759 , n71758 );
or ( n71760 , n71752 , n71759 );
nand ( n71761 , n68603 , n71494 );
nand ( n71762 , n71760 , n71761 );
not ( n71763 , n71473 );
xor ( n71764 , n71762 , n71763 );
not ( n71765 , n54327 );
not ( n71766 , n70627 );
not ( n71767 , n66704 );
not ( n71768 , n71767 );
or ( n71769 , n71766 , n71768 );
not ( n71770 , n59611 );
nand ( n71771 , n71770 , n54302 );
nand ( n71772 , n71769 , n71771 );
not ( n71773 , n71772 );
or ( n71774 , n71765 , n71773 );
nand ( n71775 , n71400 , n54316 );
nand ( n71776 , n71774 , n71775 );
xor ( n71777 , n71764 , n71776 );
xor ( n71778 , n71669 , n71777 );
not ( n71779 , n60472 );
not ( n71780 , n69820 );
not ( n71781 , n70186 );
or ( n71782 , n71780 , n71781 );
nand ( n71783 , n52289 , n56785 );
nand ( n71784 , n71782 , n71783 );
not ( n71785 , n71784 );
or ( n71786 , n71779 , n71785 );
nand ( n71787 , n71364 , n56777 );
nand ( n71788 , n71786 , n71787 );
not ( n71789 , n52151 );
not ( n71790 , n71435 );
or ( n71791 , n71789 , n71790 );
not ( n71792 , n50895 );
not ( n71793 , n68611 );
or ( n71794 , n71792 , n71793 );
nand ( n71795 , n62618 , n50946 );
nand ( n71796 , n71794 , n71795 );
nand ( n71797 , n71796 , n51223 );
nand ( n71798 , n71791 , n71797 );
xor ( n71799 , n71788 , n71798 );
not ( n71800 , n59984 );
and ( n71801 , n71094 , n51602 );
not ( n71802 , n71094 );
and ( n71803 , n71802 , n69442 );
nor ( n71804 , n71801 , n71803 );
not ( n71805 , n71804 );
or ( n71806 , n71800 , n71805 );
nand ( n71807 , n71376 , n67862 );
nand ( n71808 , n71806 , n71807 );
xor ( n71809 , n71799 , n71808 );
xor ( n71810 , n71778 , n71809 );
xor ( n71811 , n71669 , n71777 );
and ( n71812 , n71811 , n71809 );
and ( n71813 , n71669 , n71777 );
or ( n71814 , n71812 , n71813 );
not ( n71815 , n56355 );
not ( n71816 , n71447 );
or ( n71817 , n71815 , n71816 );
not ( n71818 , n53931 );
not ( n71819 , n70290 );
or ( n71820 , n71818 , n71819 );
nand ( n71821 , n67721 , n71445 );
nand ( n71822 , n71820 , n71821 );
nand ( n71823 , n71822 , n51533 );
nand ( n71824 , n71817 , n71823 );
not ( n71825 , n51766 );
not ( n71826 , n68931 );
not ( n71827 , n59694 );
or ( n71828 , n71826 , n71827 );
not ( n71829 , n59694 );
nand ( n71830 , n71829 , n52487 );
nand ( n71831 , n71828 , n71830 );
not ( n71832 , n71831 );
or ( n71833 , n71825 , n71832 );
nand ( n71834 , n71456 , n53197 );
nand ( n71835 , n71833 , n71834 );
xor ( n71836 , n71824 , n71835 );
not ( n71837 , n52854 );
not ( n71838 , n71481 );
or ( n71839 , n71837 , n71838 );
not ( n71840 , n54283 );
not ( n71841 , n62626 );
or ( n71842 , n71840 , n71841 );
nand ( n71843 , n71067 , n55104 );
nand ( n71844 , n71842 , n71843 );
nand ( n71845 , n71844 , n53571 );
nand ( n71846 , n71839 , n71845 );
xor ( n71847 , n71836 , n71846 );
xor ( n71848 , n71847 , n71673 );
not ( n71849 , n70193 );
not ( n71850 , n71411 );
or ( n71851 , n71849 , n71850 );
not ( n71852 , n55120 );
not ( n71853 , n52208 );
or ( n71854 , n71852 , n71853 );
nand ( n71855 , n40592 , n71409 );
nand ( n71856 , n71854 , n71855 );
nand ( n71857 , n71856 , n70183 );
nand ( n71858 , n71851 , n71857 );
not ( n71859 , n52757 );
not ( n71860 , n64190 );
not ( n71861 , n59414 );
or ( n71862 , n71860 , n71861 );
not ( n71863 , n59414 );
nand ( n71864 , n71863 , n64191 );
nand ( n71865 , n71862 , n71864 );
not ( n71866 , n71865 );
or ( n71867 , n71859 , n71866 );
nand ( n71868 , n71422 , n52749 );
nand ( n71869 , n71867 , n71868 );
xor ( n71870 , n71858 , n71869 );
not ( n71871 , n57314 );
not ( n71872 , n71527 );
or ( n71873 , n71871 , n71872 );
not ( n71874 , n55013 );
buf ( n71875 , n63794 );
not ( n71876 , n71875 );
not ( n71877 , n71876 );
or ( n71878 , n71874 , n71877 );
not ( n71879 , n71162 );
or ( n71880 , n71879 , n55013 );
nand ( n71881 , n71878 , n71880 );
not ( n71882 , n71881 );
nand ( n71883 , n71882 , n52004 );
nand ( n71884 , n71873 , n71883 );
xor ( n71885 , n71870 , n71884 );
xor ( n71886 , n71848 , n71885 );
xor ( n71887 , n71847 , n71673 );
and ( n71888 , n71887 , n71885 );
and ( n71889 , n71847 , n71673 );
or ( n71890 , n71888 , n71889 );
not ( n71891 , n52022 );
not ( n71892 , n71579 );
or ( n71893 , n71891 , n71892 );
not ( n71894 , n59174 );
not ( n71895 , n71139 );
or ( n71896 , n71894 , n71895 );
nand ( n71897 , n68381 , n54628 );
nand ( n71898 , n71896 , n71897 );
nand ( n71899 , n71898 , n54623 );
nand ( n71900 , n71893 , n71899 );
xor ( n71901 , n71900 , n71318 );
not ( n71902 , n62654 );
not ( n71903 , n61951 );
not ( n71904 , n60386 );
not ( n71905 , n71904 );
or ( n71906 , n71903 , n71905 );
nand ( n71907 , n39681 , n66690 );
nand ( n71908 , n71906 , n71907 );
not ( n71909 , n71908 );
or ( n71910 , n71902 , n71909 );
nand ( n71911 , n71511 , n66696 );
nand ( n71912 , n71910 , n71911 );
xor ( n71913 , n71901 , n71912 );
xor ( n71914 , n71677 , n71913 );
not ( n71915 , n59633 );
not ( n71916 , n71539 );
or ( n71917 , n71915 , n71916 );
not ( n71918 , n60602 );
not ( n71919 , n39254 );
or ( n71920 , n71918 , n71919 );
nand ( n71921 , n69530 , n52728 );
nand ( n71922 , n71920 , n71921 );
nand ( n71923 , n71922 , n58977 );
nand ( n71924 , n71917 , n71923 );
not ( n71925 , n59950 );
not ( n71926 , n71549 );
or ( n71927 , n71925 , n71926 );
and ( n71928 , n62394 , n59345 );
not ( n71929 , n62394 );
and ( n71930 , n71929 , n65743 );
or ( n71931 , n71928 , n71930 );
nand ( n71932 , n71931 , n56639 );
nand ( n71933 , n71927 , n71932 );
xor ( n71934 , n71924 , n71933 );
not ( n71935 , n52191 );
not ( n71936 , n66234 );
not ( n71937 , n65532 );
or ( n71938 , n71936 , n71937 );
nand ( n71939 , n39575 , n60289 );
nand ( n71940 , n71938 , n71939 );
not ( n71941 , n71940 );
or ( n71942 , n71935 , n71941 );
nand ( n71943 , n71569 , n62085 );
nand ( n71944 , n71942 , n71943 );
xor ( n71945 , n71934 , n71944 );
xor ( n71946 , n71914 , n71945 );
xor ( n71947 , n71677 , n71913 );
and ( n71948 , n71947 , n71945 );
and ( n71949 , n71677 , n71913 );
or ( n71950 , n71948 , n71949 );
or ( n71951 , n64164 , n71323 );
and ( n71952 , n58459 , n64170 );
not ( n71953 , n58459 );
and ( n71954 , n71953 , n66089 );
nor ( n71955 , n71952 , n71954 );
or ( n71956 , n64166 , n71955 );
nand ( n71957 , n71951 , n71956 );
not ( n71958 , n71348 );
not ( n71959 , n66569 );
not ( n71960 , n71959 );
not ( n71961 , n71960 );
or ( n71962 , n71958 , n71961 );
not ( n71963 , n47527 );
not ( n71964 , n63412 );
or ( n71965 , n71963 , n71964 );
nand ( n71966 , n67072 , n59388 );
nand ( n71967 , n71965 , n71966 );
nand ( n71968 , n70964 , n71967 );
nand ( n71969 , n71962 , n71968 );
xor ( n71970 , n71957 , n71969 );
not ( n71971 , n63415 );
and ( n71972 , n71971 , n56727 );
xor ( n71973 , n71970 , n71972 );
xor ( n71974 , n71355 , n71973 );
xor ( n71975 , n71974 , n71699 );
xor ( n71976 , n71387 , n71975 );
xor ( n71977 , n71976 , n71741 );
xor ( n71978 , n71387 , n71975 );
and ( n71979 , n71978 , n71741 );
and ( n71980 , n71387 , n71975 );
or ( n71981 , n71979 , n71980 );
xor ( n71982 , n71393 , n71502 );
xor ( n71983 , n71982 , n71589 );
xor ( n71984 , n71393 , n71502 );
and ( n71985 , n71984 , n71589 );
and ( n71986 , n71393 , n71502 );
or ( n71987 , n71985 , n71986 );
xor ( n71988 , n71521 , n71886 );
xor ( n71989 , n71988 , n71810 );
xor ( n71990 , n71521 , n71886 );
and ( n71991 , n71990 , n71810 );
and ( n71992 , n71521 , n71886 );
or ( n71993 , n71991 , n71992 );
xor ( n71994 , n71747 , n71946 );
xor ( n71995 , n71994 , n71977 );
xor ( n71996 , n71747 , n71946 );
and ( n71997 , n71996 , n71977 );
and ( n71998 , n71747 , n71946 );
or ( n71999 , n71997 , n71998 );
xor ( n72000 , n71597 , n71983 );
xor ( n72001 , n72000 , n71603 );
xor ( n72002 , n71597 , n71983 );
and ( n72003 , n72002 , n71603 );
and ( n72004 , n71597 , n71983 );
or ( n72005 , n72003 , n72004 );
xor ( n72006 , n71957 , n71969 );
and ( n72007 , n72006 , n71972 );
and ( n72008 , n71957 , n71969 );
or ( n72009 , n72007 , n72008 );
xor ( n72010 , n71609 , n71989 );
xor ( n72011 , n72010 , n71615 );
xor ( n72012 , n71609 , n71989 );
and ( n72013 , n72012 , n71615 );
and ( n72014 , n71609 , n71989 );
or ( n72015 , n72013 , n72014 );
xor ( n72016 , n71995 , n71621 );
xor ( n72017 , n72016 , n72001 );
xor ( n72018 , n71995 , n71621 );
and ( n72019 , n72018 , n72001 );
and ( n72020 , n71995 , n71621 );
or ( n72021 , n72019 , n72020 );
xor ( n72022 , n72011 , n71631 );
xor ( n72023 , n72022 , n71637 );
xor ( n72024 , n72011 , n71631 );
and ( n72025 , n72024 , n71637 );
and ( n72026 , n72011 , n71631 );
or ( n72027 , n72025 , n72026 );
xor ( n72028 , n72017 , n72023 );
xor ( n72029 , n72028 , n71643 );
xor ( n72030 , n72017 , n72023 );
and ( n72031 , n72030 , n71643 );
and ( n72032 , n72017 , n72023 );
or ( n72033 , n72031 , n72032 );
xor ( n72034 , n71788 , n71798 );
and ( n72035 , n72034 , n71808 );
and ( n72036 , n71788 , n71798 );
or ( n72037 , n72035 , n72036 );
xor ( n72038 , n71824 , n71835 );
and ( n72039 , n72038 , n71846 );
and ( n72040 , n71824 , n71835 );
or ( n72041 , n72039 , n72040 );
xor ( n72042 , n71762 , n71763 );
and ( n72043 , n72042 , n71776 );
and ( n72044 , n71762 , n71763 );
or ( n72045 , n72043 , n72044 );
xor ( n72046 , n71858 , n71869 );
and ( n72047 , n72046 , n71884 );
and ( n72048 , n71858 , n71869 );
or ( n72049 , n72047 , n72048 );
xor ( n72050 , n71924 , n71933 );
and ( n72051 , n72050 , n71944 );
and ( n72052 , n71924 , n71933 );
or ( n72053 , n72051 , n72052 );
xor ( n72054 , n71900 , n71318 );
and ( n72055 , n72054 , n71912 );
and ( n72056 , n71900 , n71318 );
or ( n72057 , n72055 , n72056 );
xor ( n72058 , n71355 , n71973 );
and ( n72059 , n72058 , n71699 );
and ( n72060 , n71355 , n71973 );
or ( n72061 , n72059 , n72060 );
not ( n72062 , n71723 );
not ( n72063 , n65130 );
or ( n72064 , n72062 , n72063 );
not ( n72065 , n41288 );
not ( n72066 , n66141 );
or ( n72067 , n72065 , n72066 );
nand ( n72068 , n66140 , n48997 );
nand ( n72069 , n72067 , n72068 );
nand ( n72070 , n60427 , n72069 );
nand ( n72071 , n72064 , n72070 );
not ( n72072 , n71731 );
not ( n72073 , n64111 );
or ( n72074 , n72072 , n72073 );
and ( n72075 , n48486 , n69333 );
not ( n72076 , n48486 );
and ( n72077 , n72076 , n71309 );
or ( n72078 , n72075 , n72077 );
nand ( n72079 , n67094 , n72078 );
nand ( n72080 , n72074 , n72079 );
xor ( n72081 , n72071 , n72080 );
or ( n72082 , n64164 , n71955 );
not ( n72083 , n66089 );
and ( n72084 , n66946 , n72083 );
not ( n72085 , n66946 );
and ( n72086 , n72085 , n69704 );
nor ( n72087 , n72084 , n72086 );
or ( n72088 , n69703 , n72087 );
nand ( n72089 , n72082 , n72088 );
xor ( n72090 , n72081 , n72089 );
xor ( n72091 , n72071 , n72080 );
and ( n72092 , n72091 , n72089 );
and ( n72093 , n72071 , n72080 );
or ( n72094 , n72092 , n72093 );
not ( n72095 , n71967 );
not ( n72096 , n65795 );
or ( n72097 , n72095 , n72096 );
not ( n72098 , n42127 );
not ( n72099 , n63415 );
or ( n72100 , n72098 , n72099 );
nand ( n72101 , n65474 , n41416 );
nand ( n72102 , n72100 , n72101 );
nand ( n72103 , n65092 , n72102 );
nand ( n72104 , n72097 , n72103 );
not ( n72105 , n71695 );
buf ( n72106 , n63080 );
not ( n72107 , n72106 );
or ( n72108 , n72105 , n72107 );
not ( n72109 , n50021 );
not ( n72110 , n65187 );
or ( n72111 , n72109 , n72110 );
nand ( n72112 , n58642 , n55674 );
nand ( n72113 , n72111 , n72112 );
nand ( n72114 , n61465 , n72113 );
nand ( n72115 , n72108 , n72114 );
xor ( n72116 , n72104 , n72115 );
and ( n72117 , n66581 , n57182 );
xor ( n72118 , n72116 , n72117 );
xor ( n72119 , n72104 , n72115 );
and ( n72120 , n72119 , n72117 );
and ( n72121 , n72104 , n72115 );
or ( n72122 , n72120 , n72121 );
xor ( n72123 , n72037 , n72041 );
xor ( n72124 , n72123 , n72049 );
xor ( n72125 , n72037 , n72041 );
and ( n72126 , n72125 , n72049 );
and ( n72127 , n72037 , n72041 );
or ( n72128 , n72126 , n72127 );
xor ( n72129 , n72053 , n72057 );
not ( n72130 , n71713 );
buf ( n72131 , n62506 );
not ( n72132 , n72131 );
or ( n72133 , n72130 , n72132 );
not ( n72134 , n70920 );
not ( n72135 , n40856 );
or ( n72136 , n72134 , n72135 );
nand ( n72137 , n59341 , n40855 );
nand ( n72138 , n72136 , n72137 );
nand ( n72139 , n60542 , n72138 );
nand ( n72140 , n72133 , n72139 );
not ( n72141 , n72140 );
not ( n72142 , n55161 );
not ( n72143 , n72142 );
not ( n72144 , n71772 );
or ( n72145 , n72143 , n72144 );
and ( n72146 , n70627 , n56476 );
not ( n72147 , n70627 );
not ( n72148 , n53286 );
and ( n72149 , n72147 , n72148 );
or ( n72150 , n72146 , n72149 );
nand ( n72151 , n72150 , n54327 );
nand ( n72152 , n72145 , n72151 );
xor ( n72153 , n72141 , n72152 );
not ( n72154 , n70193 );
not ( n72155 , n71856 );
or ( n72156 , n72154 , n72155 );
not ( n72157 , n40628 );
not ( n72158 , n71409 );
and ( n72159 , n72157 , n72158 );
not ( n72160 , n53271 );
and ( n72161 , n72160 , n71409 );
nor ( n72162 , n72159 , n72161 );
not ( n72163 , n72162 );
nand ( n72164 , n72163 , n70183 );
nand ( n72165 , n72156 , n72164 );
xor ( n72166 , n72153 , n72165 );
xor ( n72167 , n72129 , n72166 );
xor ( n72168 , n72053 , n72057 );
and ( n72169 , n72168 , n72166 );
and ( n72170 , n72053 , n72057 );
or ( n72171 , n72169 , n72170 );
not ( n72172 , n70604 );
not ( n72173 , n66963 );
not ( n72174 , n40691 );
or ( n72175 , n72173 , n72174 );
not ( n72176 , n71361 );
nand ( n72177 , n72176 , n67568 );
nand ( n72178 , n72175 , n72177 );
not ( n72179 , n72178 );
or ( n72180 , n72172 , n72179 );
not ( n72181 , n71685 );
not ( n72182 , n67885 );
nand ( n72183 , n72181 , n72182 );
nand ( n72184 , n72180 , n72183 );
buf ( n72185 , n60472 );
not ( n72186 , n72185 );
not ( n72187 , n69820 );
not ( n72188 , n70638 );
or ( n72189 , n72187 , n72188 );
nand ( n72190 , n40736 , n56785 );
nand ( n72191 , n72189 , n72190 );
not ( n72192 , n72191 );
or ( n72193 , n72186 , n72192 );
nand ( n72194 , n71784 , n56777 );
nand ( n72195 , n72193 , n72194 );
xor ( n72196 , n72184 , n72195 );
not ( n72197 , n56355 );
not ( n72198 , n72197 );
not ( n72199 , n72198 );
not ( n72200 , n71822 );
or ( n72201 , n72199 , n72200 );
not ( n72202 , n53931 );
not ( n72203 , n67193 );
or ( n72204 , n72202 , n72203 );
not ( n72205 , n63180 );
nand ( n72206 , n72205 , n71053 );
nand ( n72207 , n72204 , n72206 );
nand ( n72208 , n72207 , n51533 );
nand ( n72209 , n72201 , n72208 );
xor ( n72210 , n72196 , n72209 );
not ( n72211 , n52125 );
not ( n72212 , n71831 );
or ( n72213 , n72211 , n72212 );
not ( n72214 , n52114 );
not ( n72215 , n70661 );
or ( n72216 , n72214 , n72215 );
not ( n72217 , n70661 );
nand ( n72218 , n72217 , n52130 );
nand ( n72219 , n72216 , n72218 );
buf ( n72220 , n51766 );
nand ( n72221 , n72219 , n72220 );
nand ( n72222 , n72213 , n72221 );
not ( n72223 , n52854 );
not ( n72224 , n71844 );
or ( n72225 , n72223 , n72224 );
not ( n72226 , n69458 );
not ( n72227 , n57390 );
or ( n72228 , n72226 , n72227 );
nand ( n72229 , n68990 , n55104 );
nand ( n72230 , n72228 , n72229 );
nand ( n72231 , n72230 , n52469 );
nand ( n72232 , n72225 , n72231 );
xor ( n72233 , n72222 , n72232 );
not ( n72234 , n54364 );
not ( n72235 , n55089 );
not ( n72236 , n66236 );
or ( n72237 , n72235 , n72236 );
not ( n72238 , n55089 );
nand ( n72239 , n71479 , n72238 );
nand ( n72240 , n72237 , n72239 );
not ( n72241 , n72240 );
or ( n72242 , n72234 , n72241 );
nand ( n72243 , n71758 , n68603 );
nand ( n72244 , n72242 , n72243 );
xor ( n72245 , n72233 , n72244 );
xor ( n72246 , n72210 , n72245 );
or ( n72247 , n71881 , n56515 );
or ( n72248 , n55013 , n56523 );
nand ( n72249 , n72247 , n72248 );
not ( n72250 , n58977 );
not ( n72251 , n58982 );
buf ( n72252 , n66052 );
not ( n72253 , n72252 );
or ( n72254 , n72251 , n72253 );
not ( n72255 , n60602 );
nand ( n72256 , n72255 , n71577 );
nand ( n72257 , n72254 , n72256 );
not ( n72258 , n72257 );
or ( n72259 , n72250 , n72258 );
nand ( n72260 , n53104 , n71922 );
nand ( n72261 , n72259 , n72260 );
xor ( n72262 , n72249 , n72261 );
xor ( n72263 , n72262 , n71703 );
xor ( n72264 , n72246 , n72263 );
xor ( n72265 , n72210 , n72245 );
and ( n72266 , n72265 , n72263 );
and ( n72267 , n72210 , n72245 );
or ( n72268 , n72266 , n72267 );
not ( n72269 , n63708 );
not ( n72270 , n71865 );
or ( n72271 , n72269 , n72270 );
not ( n72272 , n64190 );
not ( n72273 , n67037 );
or ( n72274 , n72272 , n72273 );
buf ( n72275 , n59913 );
nand ( n72276 , n72275 , n64191 );
nand ( n72277 , n72274 , n72276 );
nand ( n72278 , n72277 , n52757 );
nand ( n72279 , n72271 , n72278 );
xor ( n72280 , n71739 , n72279 );
xor ( n72281 , n72280 , n72009 );
not ( n72282 , n71099 );
not ( n72283 , n71804 );
or ( n72284 , n72282 , n72283 );
not ( n72285 , n69695 );
not ( n72286 , n51913 );
or ( n72287 , n72285 , n72286 );
not ( n72288 , n55846 );
not ( n72289 , n72288 );
nand ( n72290 , n51916 , n72289 );
nand ( n72291 , n72287 , n72290 );
nand ( n72292 , n72291 , n59984 );
nand ( n72293 , n72284 , n72292 );
not ( n72294 , n50922 );
not ( n72295 , n50895 );
not ( n72296 , n71418 );
or ( n72297 , n72295 , n72296 );
not ( n72298 , n60167 );
nand ( n72299 , n72298 , n67639 );
nand ( n72300 , n72297 , n72299 );
not ( n72301 , n72300 );
or ( n72302 , n72294 , n72301 );
nand ( n72303 , n71796 , n52151 );
nand ( n72304 , n72302 , n72303 );
xor ( n72305 , n72293 , n72304 );
not ( n72306 , n54623 );
not ( n72307 , n71525 );
and ( n72308 , n72307 , n59174 );
not ( n72309 , n72307 );
buf ( n72310 , n54628 );
and ( n72311 , n72309 , n72310 );
or ( n72312 , n72308 , n72311 );
not ( n72313 , n72312 );
or ( n72314 , n72306 , n72313 );
nand ( n72315 , n71898 , n52022 );
nand ( n72316 , n72314 , n72315 );
xor ( n72317 , n72305 , n72316 );
xor ( n72318 , n72281 , n72317 );
xor ( n72319 , n72318 , n72061 );
xor ( n72320 , n72281 , n72317 );
and ( n72321 , n72320 , n72061 );
and ( n72322 , n72281 , n72317 );
or ( n72323 , n72321 , n72322 );
not ( n72324 , n59950 );
not ( n72325 , n71931 );
or ( n72326 , n72324 , n72325 );
not ( n72327 , n59345 );
not ( n72328 , n39331 );
or ( n72329 , n72327 , n72328 );
nand ( n72330 , n69919 , n65743 );
nand ( n72331 , n72329 , n72330 );
nand ( n72332 , n72331 , n56639 );
nand ( n72333 , n72326 , n72332 );
not ( n72334 , n52191 );
not ( n72335 , n39056 );
not ( n72336 , n69893 );
and ( n72337 , n72335 , n72336 );
and ( n72338 , n71547 , n60289 );
nor ( n72339 , n72337 , n72338 );
not ( n72340 , n72339 );
not ( n72341 , n72340 );
or ( n72342 , n72334 , n72341 );
nand ( n72343 , n71940 , n58168 );
nand ( n72344 , n72342 , n72343 );
xor ( n72345 , n72333 , n72344 );
not ( n72346 , n66696 );
not ( n72347 , n71908 );
or ( n72348 , n72346 , n72347 );
not ( n72349 , n61951 );
not ( n72350 , n68206 );
or ( n72351 , n72349 , n72350 );
nand ( n72352 , n39714 , n66690 );
nand ( n72353 , n72351 , n72352 );
nand ( n72354 , n72353 , n62654 );
nand ( n72355 , n72348 , n72354 );
xor ( n72356 , n72345 , n72355 );
xor ( n72357 , n72356 , n71745 );
xor ( n72358 , n72118 , n72090 );
xor ( n72359 , n72358 , n72045 );
xor ( n72360 , n72357 , n72359 );
xor ( n72361 , n72356 , n71745 );
and ( n72362 , n72361 , n72359 );
and ( n72363 , n72356 , n71745 );
or ( n72364 , n72362 , n72363 );
xor ( n72365 , n71814 , n71751 );
xor ( n72366 , n72365 , n72124 );
xor ( n72367 , n71814 , n71751 );
and ( n72368 , n72367 , n72124 );
and ( n72369 , n71814 , n71751 );
or ( n72370 , n72368 , n72369 );
xor ( n72371 , n71950 , n72264 );
xor ( n72372 , n72371 , n72167 );
xor ( n72373 , n71950 , n72264 );
and ( n72374 , n72373 , n72167 );
and ( n72375 , n71950 , n72264 );
or ( n72376 , n72374 , n72375 );
xor ( n72377 , n71890 , n72319 );
xor ( n72378 , n72377 , n71981 );
xor ( n72379 , n71890 , n72319 );
and ( n72380 , n72379 , n71981 );
and ( n72381 , n71890 , n72319 );
or ( n72382 , n72380 , n72381 );
xor ( n72383 , n72360 , n71987 );
xor ( n72384 , n72383 , n72366 );
xor ( n72385 , n72360 , n71987 );
and ( n72386 , n72385 , n72366 );
and ( n72387 , n72360 , n71987 );
or ( n72388 , n72386 , n72387 );
xor ( n72389 , n71993 , n72372 );
xor ( n72390 , n72389 , n71999 );
xor ( n72391 , n71993 , n72372 );
and ( n72392 , n72391 , n71999 );
and ( n72393 , n71993 , n72372 );
or ( n72394 , n72392 , n72393 );
xor ( n72395 , n72184 , n72195 );
and ( n72396 , n72395 , n72209 );
and ( n72397 , n72184 , n72195 );
or ( n72398 , n72396 , n72397 );
xor ( n72399 , n72378 , n72005 );
xor ( n72400 , n72399 , n72384 );
xor ( n72401 , n72378 , n72005 );
and ( n72402 , n72401 , n72384 );
and ( n72403 , n72378 , n72005 );
or ( n72404 , n72402 , n72403 );
xor ( n72405 , n72390 , n72015 );
xor ( n72406 , n72405 , n72400 );
xor ( n72407 , n72390 , n72015 );
and ( n72408 , n72407 , n72400 );
and ( n72409 , n72390 , n72015 );
or ( n72410 , n72408 , n72409 );
xor ( n72411 , n72021 , n72406 );
xor ( n72412 , n72411 , n72027 );
xor ( n72413 , n72021 , n72406 );
and ( n72414 , n72413 , n72027 );
and ( n72415 , n72021 , n72406 );
or ( n72416 , n72414 , n72415 );
xor ( n72417 , n72222 , n72232 );
and ( n72418 , n72417 , n72244 );
and ( n72419 , n72222 , n72232 );
or ( n72420 , n72418 , n72419 );
xor ( n72421 , n72141 , n72152 );
and ( n72422 , n72421 , n72165 );
and ( n72423 , n72141 , n72152 );
or ( n72424 , n72422 , n72423 );
xor ( n72425 , n72293 , n72304 );
and ( n72426 , n72425 , n72316 );
and ( n72427 , n72293 , n72304 );
or ( n72428 , n72426 , n72427 );
xor ( n72429 , n72333 , n72344 );
and ( n72430 , n72429 , n72355 );
and ( n72431 , n72333 , n72344 );
or ( n72432 , n72430 , n72431 );
xor ( n72433 , n72249 , n72261 );
and ( n72434 , n72433 , n71703 );
and ( n72435 , n72249 , n72261 );
or ( n72436 , n72434 , n72435 );
xor ( n72437 , n71739 , n72279 );
and ( n72438 , n72437 , n72009 );
and ( n72439 , n71739 , n72279 );
or ( n72440 , n72438 , n72439 );
xor ( n72441 , n72118 , n72090 );
and ( n72442 , n72441 , n72045 );
and ( n72443 , n72118 , n72090 );
or ( n72444 , n72442 , n72443 );
or ( n72445 , n48894 , n52004 );
nand ( n72446 , n72445 , n52377 );
not ( n72447 , n72113 );
not ( n72448 , n65646 );
or ( n72449 , n72447 , n72448 );
not ( n72450 , n65183 );
not ( n72451 , n41132 );
or ( n72452 , n72450 , n72451 );
not ( n72453 , n52079 );
nand ( n72454 , n72453 , n62496 );
nand ( n72455 , n72452 , n72454 );
nand ( n72456 , n71466 , n72455 );
nand ( n72457 , n72449 , n72456 );
xor ( n72458 , n72446 , n72457 );
not ( n72459 , n70487 );
not ( n72460 , n72138 );
or ( n72461 , n72459 , n72460 );
and ( n72462 , n71691 , n66983 );
not ( n72463 , n71691 );
not ( n72464 , n70920 );
and ( n72465 , n72463 , n72464 );
nor ( n72466 , n72462 , n72465 );
or ( n72467 , n67586 , n72466 );
nand ( n72468 , n72461 , n72467 );
xor ( n72469 , n72458 , n72468 );
xor ( n72470 , n72446 , n72457 );
and ( n72471 , n72470 , n72468 );
and ( n72472 , n72446 , n72457 );
or ( n72473 , n72471 , n72472 );
not ( n72474 , n70500 );
not ( n72475 , n72069 );
or ( n72476 , n72474 , n72475 );
not ( n72477 , n66140 );
and ( n72478 , n72477 , n41217 );
and ( n72479 , n66140 , n50387 );
nor ( n72480 , n72478 , n72479 );
or ( n72481 , n60963 , n72480 );
nand ( n72482 , n72476 , n72481 );
not ( n72483 , n72078 );
not ( n72484 , n69728 );
not ( n72485 , n72484 );
or ( n72486 , n72483 , n72485 );
not ( n72487 , n67441 );
not ( n72488 , n61537 );
or ( n72489 , n72487 , n72488 );
nand ( n72490 , n61416 , n49190 );
nand ( n72491 , n72489 , n72490 );
nand ( n72492 , n61558 , n72491 );
nand ( n72493 , n72486 , n72492 );
xor ( n72494 , n72482 , n72493 );
buf ( n72495 , n64164 );
or ( n72496 , n72495 , n72087 );
not ( n72497 , n48306 );
not ( n72498 , n69704 );
or ( n72499 , n72497 , n72498 );
nand ( n72500 , n64170 , n69270 );
nand ( n72501 , n72499 , n72500 );
not ( n72502 , n72501 );
or ( n72503 , n64166 , n72502 );
nand ( n72504 , n72496 , n72503 );
xor ( n72505 , n72494 , n72504 );
xor ( n72506 , n72482 , n72493 );
and ( n72507 , n72506 , n72504 );
and ( n72508 , n72482 , n72493 );
or ( n72509 , n72507 , n72508 );
xor ( n72510 , n72398 , n72420 );
xor ( n72511 , n72510 , n72424 );
xor ( n72512 , n72398 , n72420 );
and ( n72513 , n72512 , n72424 );
and ( n72514 , n72398 , n72420 );
or ( n72515 , n72513 , n72514 );
xor ( n72516 , n72432 , n72436 );
xor ( n72517 , n72516 , n72440 );
xor ( n72518 , n72432 , n72436 );
and ( n72519 , n72518 , n72440 );
and ( n72520 , n72432 , n72436 );
or ( n72521 , n72519 , n72520 );
not ( n72522 , n52854 );
not ( n72523 , n72230 );
or ( n72524 , n72522 , n72523 );
not ( n72525 , n69458 );
not ( n72526 , n59694 );
or ( n72527 , n72525 , n72526 );
nand ( n72528 , n71052 , n55104 );
nand ( n72529 , n72527 , n72528 );
nand ( n72530 , n72529 , n52469 );
nand ( n72531 , n72524 , n72530 );
not ( n72532 , n54364 );
and ( n72533 , n53596 , n54402 );
not ( n72534 , n53596 );
and ( n72535 , n72534 , n69409 );
or ( n72536 , n72533 , n72535 );
not ( n72537 , n72536 );
or ( n72538 , n72532 , n72537 );
nand ( n72539 , n72240 , n68603 );
nand ( n72540 , n72538 , n72539 );
xor ( n72541 , n72531 , n72540 );
not ( n72542 , n54327 );
not ( n72543 , n54725 );
not ( n72544 , n59601 );
not ( n72545 , n72544 );
or ( n72546 , n72543 , n72545 );
nand ( n72547 , n40226 , n54302 );
nand ( n72548 , n72546 , n72547 );
not ( n72549 , n72548 );
or ( n72550 , n72542 , n72549 );
not ( n72551 , n55161 );
nand ( n72552 , n72551 , n72150 );
nand ( n72553 , n72550 , n72552 );
xor ( n72554 , n72541 , n72553 );
or ( n72555 , n72162 , n68334 );
not ( n72556 , n55120 );
not ( n72557 , n59611 );
or ( n72558 , n72556 , n72557 );
nand ( n72559 , n71770 , n71409 );
nand ( n72560 , n72558 , n72559 );
not ( n72561 , n72560 );
not ( n72562 , n70183 );
or ( n72563 , n72561 , n72562 );
nand ( n72564 , n72555 , n72563 );
xor ( n72565 , n72140 , n72564 );
not ( n72566 , n59984 );
not ( n72567 , n71371 );
not ( n72568 , n66798 );
or ( n72569 , n72567 , n72568 );
nand ( n72570 , n40592 , n71094 );
nand ( n72571 , n72569 , n72570 );
not ( n72572 , n72571 );
or ( n72573 , n72566 , n72572 );
nand ( n72574 , n72291 , n71099 );
nand ( n72575 , n72573 , n72574 );
xor ( n72576 , n72565 , n72575 );
xor ( n72577 , n72554 , n72576 );
not ( n72578 , n56355 );
not ( n72579 , n72207 );
or ( n72580 , n72578 , n72579 );
not ( n72581 , n53931 );
not ( n72582 , n59651 );
or ( n72583 , n72581 , n72582 );
nand ( n72584 , n39964 , n71053 );
nand ( n72585 , n72583 , n72584 );
nand ( n72586 , n72585 , n51533 );
nand ( n72587 , n72580 , n72586 );
not ( n72588 , n72185 );
not ( n72589 , n71362 );
not ( n72590 , n72589 );
not ( n72591 , n51602 );
or ( n72592 , n72590 , n72591 );
buf ( n72593 , n69819 );
nand ( n72594 , n69442 , n72593 );
nand ( n72595 , n72592 , n72594 );
not ( n72596 , n72595 );
or ( n72597 , n72588 , n72596 );
nand ( n72598 , n72191 , n56777 );
nand ( n72599 , n72597 , n72598 );
xor ( n72600 , n72587 , n72599 );
not ( n72601 , n53197 );
not ( n72602 , n72219 );
or ( n72603 , n72601 , n72602 );
and ( n72604 , n52487 , n70290 );
not ( n72605 , n52487 );
not ( n72606 , n40514 );
not ( n72607 , n72606 );
and ( n72608 , n72605 , n72607 );
or ( n72609 , n72604 , n72608 );
not ( n72610 , n72609 );
nand ( n72611 , n72610 , n72220 );
nand ( n72612 , n72603 , n72611 );
xor ( n72613 , n72600 , n72612 );
xor ( n72614 , n72577 , n72613 );
xor ( n72615 , n72554 , n72576 );
and ( n72616 , n72615 , n72613 );
and ( n72617 , n72554 , n72576 );
or ( n72618 , n72616 , n72617 );
or ( n72619 , n72339 , n58167 );
and ( n72620 , n66234 , n68652 );
not ( n72621 , n66234 );
not ( n72622 , n62394 );
and ( n72623 , n72621 , n72622 );
nor ( n72624 , n72620 , n72623 );
or ( n72625 , n72624 , n59811 );
nand ( n72626 , n72619 , n72625 );
not ( n72627 , n72353 );
not ( n72628 , n66696 );
or ( n72629 , n72627 , n72628 );
not ( n72630 , n61951 );
not ( n72631 , n59399 );
or ( n72632 , n72630 , n72631 );
nand ( n72633 , n68667 , n61952 );
nand ( n72634 , n72632 , n72633 );
not ( n72635 , n72634 );
not ( n72636 , n62654 );
or ( n72637 , n72635 , n72636 );
nand ( n72638 , n72629 , n72637 );
xor ( n72639 , n72626 , n72638 );
not ( n72640 , n72257 );
or ( n72641 , n72640 , n59632 );
buf ( n72642 , n42399 );
and ( n72643 , n60602 , n72642 );
not ( n72644 , n60602 );
and ( n72645 , n72644 , n68381 );
nor ( n72646 , n72643 , n72645 );
or ( n72647 , n72646 , n59630 );
nand ( n72648 , n72641 , n72647 );
xor ( n72649 , n72639 , n72648 );
xor ( n72650 , n72428 , n72649 );
xor ( n72651 , n72094 , n72122 );
not ( n72652 , n72277 );
or ( n72653 , n72652 , n59820 );
not ( n72654 , n66546 );
not ( n72655 , n64191 );
and ( n72656 , n72654 , n72655 );
and ( n72657 , n39681 , n66705 );
nor ( n72658 , n72656 , n72657 );
or ( n72659 , n72658 , n59828 );
nand ( n72660 , n72653 , n72659 );
xor ( n72661 , n72651 , n72660 );
xor ( n72662 , n72650 , n72661 );
xor ( n72663 , n72428 , n72649 );
and ( n72664 , n72663 , n72661 );
and ( n72665 , n72428 , n72649 );
or ( n72666 , n72664 , n72665 );
not ( n72667 , n52151 );
not ( n72668 , n72300 );
or ( n72669 , n72667 , n72668 );
not ( n72670 , n51465 );
not ( n72671 , n59414 );
or ( n72672 , n72670 , n72671 );
nand ( n72673 , n71013 , n67639 );
nand ( n72674 , n72672 , n72673 );
nand ( n72675 , n72674 , n50922 );
nand ( n72676 , n72669 , n72675 );
not ( n72677 , n52022 );
not ( n72678 , n72312 );
or ( n72679 , n72677 , n72678 );
not ( n72680 , n59174 );
not ( n72681 , n71876 );
or ( n72682 , n72680 , n72681 );
nand ( n72683 , n71875 , n54628 );
nand ( n72684 , n72682 , n72683 );
nand ( n72685 , n72684 , n54623 );
nand ( n72686 , n72679 , n72685 );
xor ( n72687 , n72676 , n72686 );
not ( n72688 , n56639 );
not ( n72689 , n59345 );
not ( n72690 , n71176 );
or ( n72691 , n72689 , n72690 );
nand ( n72692 , n69530 , n60617 );
nand ( n72693 , n72691 , n72692 );
not ( n72694 , n72693 );
or ( n72695 , n72688 , n72694 );
nand ( n72696 , n72331 , n59950 );
nand ( n72697 , n72695 , n72696 );
xor ( n72698 , n72687 , n72697 );
xor ( n72699 , n72698 , n72444 );
xor ( n72700 , n72505 , n72469 );
not ( n72701 , n72102 );
or ( n72702 , n63411 , n72701 );
xor ( n72703 , n58459 , n66575 );
not ( n72704 , n65092 );
or ( n72705 , n72703 , n72704 );
nand ( n72706 , n72702 , n72705 );
not ( n72707 , n64444 );
nor ( n72708 , n72707 , n59388 );
xor ( n72709 , n72706 , n72708 );
not ( n72710 , n69648 );
not ( n72711 , n72710 );
not ( n72712 , n52289 );
not ( n72713 , n70608 );
and ( n72714 , n72712 , n72713 );
and ( n72715 , n52289 , n70608 );
nor ( n72716 , n72714 , n72715 );
not ( n72717 , n72716 );
not ( n72718 , n72717 );
or ( n72719 , n72711 , n72718 );
nand ( n72720 , n72178 , n72182 );
nand ( n72721 , n72719 , n72720 );
xor ( n72722 , n72709 , n72721 );
xor ( n72723 , n72700 , n72722 );
xor ( n72724 , n72699 , n72723 );
xor ( n72725 , n72698 , n72444 );
and ( n72726 , n72725 , n72723 );
and ( n72727 , n72698 , n72444 );
or ( n72728 , n72726 , n72727 );
xor ( n72729 , n72128 , n72511 );
xor ( n72730 , n72729 , n72171 );
xor ( n72731 , n72128 , n72511 );
and ( n72732 , n72731 , n72171 );
and ( n72733 , n72128 , n72511 );
or ( n72734 , n72732 , n72733 );
xor ( n72735 , n72517 , n72614 );
xor ( n72736 , n72735 , n72323 );
xor ( n72737 , n72517 , n72614 );
and ( n72738 , n72737 , n72323 );
and ( n72739 , n72517 , n72614 );
or ( n72740 , n72738 , n72739 );
xor ( n72741 , n72268 , n72364 );
xor ( n72742 , n72741 , n72662 );
xor ( n72743 , n72268 , n72364 );
and ( n72744 , n72743 , n72662 );
and ( n72745 , n72268 , n72364 );
or ( n72746 , n72744 , n72745 );
xor ( n72747 , n72370 , n72724 );
xor ( n72748 , n72747 , n72730 );
xor ( n72749 , n72370 , n72724 );
and ( n72750 , n72749 , n72730 );
and ( n72751 , n72370 , n72724 );
or ( n72752 , n72750 , n72751 );
xor ( n72753 , n72376 , n72736 );
xor ( n72754 , n72753 , n72742 );
xor ( n72755 , n72376 , n72736 );
and ( n72756 , n72755 , n72742 );
and ( n72757 , n72376 , n72736 );
or ( n72758 , n72756 , n72757 );
xor ( n72759 , n72706 , n72708 );
and ( n72760 , n72759 , n72721 );
and ( n72761 , n72706 , n72708 );
or ( n72762 , n72760 , n72761 );
xor ( n72763 , n72382 , n72388 );
xor ( n72764 , n72763 , n72748 );
xor ( n72765 , n72382 , n72388 );
and ( n72766 , n72765 , n72748 );
and ( n72767 , n72382 , n72388 );
or ( n72768 , n72766 , n72767 );
xor ( n72769 , n72754 , n72394 );
xor ( n72770 , n72769 , n72404 );
xor ( n72771 , n72754 , n72394 );
and ( n72772 , n72771 , n72404 );
and ( n72773 , n72754 , n72394 );
or ( n72774 , n72772 , n72773 );
xor ( n72775 , n72764 , n72770 );
xor ( n72776 , n72775 , n72410 );
xor ( n72777 , n72764 , n72770 );
and ( n72778 , n72777 , n72410 );
and ( n72779 , n72764 , n72770 );
or ( n72780 , n72778 , n72779 );
xor ( n72781 , n72587 , n72599 );
and ( n72782 , n72781 , n72612 );
and ( n72783 , n72587 , n72599 );
or ( n72784 , n72782 , n72783 );
xor ( n72785 , n72531 , n72540 );
and ( n72786 , n72785 , n72553 );
and ( n72787 , n72531 , n72540 );
or ( n72788 , n72786 , n72787 );
xor ( n72789 , n72140 , n72564 );
and ( n72790 , n72789 , n72575 );
and ( n72791 , n72140 , n72564 );
or ( n72792 , n72790 , n72791 );
xor ( n72793 , n72676 , n72686 );
and ( n72794 , n72793 , n72697 );
and ( n72795 , n72676 , n72686 );
or ( n72796 , n72794 , n72795 );
xor ( n72797 , n72626 , n72638 );
and ( n72798 , n72797 , n72648 );
and ( n72799 , n72626 , n72638 );
or ( n72800 , n72798 , n72799 );
xor ( n72801 , n72094 , n72122 );
and ( n72802 , n72801 , n72660 );
and ( n72803 , n72094 , n72122 );
or ( n72804 , n72802 , n72803 );
xor ( n72805 , n72505 , n72469 );
and ( n72806 , n72805 , n72722 );
and ( n72807 , n72505 , n72469 );
or ( n72808 , n72806 , n72807 );
not ( n72809 , n72491 );
not ( n72810 , n69728 );
not ( n72811 , n72810 );
or ( n72812 , n72809 , n72811 );
not ( n72813 , n61540 );
not ( n72814 , n48997 );
or ( n72815 , n72813 , n72814 );
not ( n72816 , n66615 );
nand ( n72817 , n72816 , n41286 );
nand ( n72818 , n72815 , n72817 );
nand ( n72819 , n61558 , n72818 );
nand ( n72820 , n72812 , n72819 );
not ( n72821 , n72501 );
not ( n72822 , n67061 );
or ( n72823 , n72821 , n72822 );
not ( n72824 , n48486 );
not ( n72825 , n69704 );
or ( n72826 , n72824 , n72825 );
nand ( n72827 , n69707 , n48951 );
nand ( n72828 , n72826 , n72827 );
nand ( n72829 , n67068 , n72828 );
nand ( n72830 , n72823 , n72829 );
xor ( n72831 , n72820 , n72830 );
or ( n72832 , n71959 , n72703 );
not ( n72833 , n64444 );
not ( n72834 , n66946 );
and ( n72835 , n72833 , n72834 );
and ( n72836 , n63922 , n66946 );
nor ( n72837 , n72835 , n72836 );
not ( n72838 , n70964 );
or ( n72839 , n72837 , n72838 );
nand ( n72840 , n72832 , n72839 );
xor ( n72841 , n72831 , n72840 );
xor ( n72842 , n72820 , n72830 );
and ( n72843 , n72842 , n72840 );
and ( n72844 , n72820 , n72830 );
or ( n72845 , n72843 , n72844 );
buf ( n72846 , n65474 );
and ( n72847 , n72846 , n42127 );
not ( n72848 , n60542 );
not ( n72849 , n55674 );
not ( n72850 , n72464 );
or ( n72851 , n72849 , n72850 );
or ( n72852 , n62513 , n50020 );
nand ( n72853 , n72851 , n72852 );
not ( n72854 , n72853 );
or ( n72855 , n72848 , n72854 );
not ( n72856 , n72466 );
nand ( n72857 , n72856 , n70487 );
nand ( n72858 , n72855 , n72857 );
xor ( n72859 , n72847 , n72858 );
not ( n72860 , n71466 );
not ( n72861 , n65183 );
not ( n72862 , n71361 );
or ( n72863 , n72861 , n72862 );
or ( n72864 , n71361 , n65187 );
nand ( n72865 , n72863 , n72864 );
not ( n72866 , n72865 );
or ( n72867 , n72860 , n72866 );
nand ( n72868 , n65646 , n72455 );
nand ( n72869 , n72867 , n72868 );
xor ( n72870 , n72859 , n72869 );
xor ( n72871 , n72847 , n72858 );
and ( n72872 , n72871 , n72869 );
and ( n72873 , n72847 , n72858 );
or ( n72874 , n72872 , n72873 );
xor ( n72875 , n72792 , n72800 );
xor ( n72876 , n72875 , n72804 );
xor ( n72877 , n72792 , n72800 );
and ( n72878 , n72877 , n72804 );
and ( n72879 , n72792 , n72800 );
or ( n72880 , n72878 , n72879 );
not ( n72881 , n68603 );
not ( n72882 , n72536 );
or ( n72883 , n72881 , n72882 );
not ( n72884 , n53596 );
not ( n72885 , n68991 );
or ( n72886 , n72884 , n72885 );
nand ( n72887 , n68994 , n72238 );
nand ( n72888 , n72886 , n72887 );
nand ( n72889 , n72888 , n53620 );
nand ( n72890 , n72883 , n72889 );
not ( n72891 , n72480 );
not ( n72892 , n72891 );
not ( n72893 , n70500 );
or ( n72894 , n72892 , n72893 );
not ( n72895 , n66140 );
not ( n72896 , n40855 );
and ( n72897 , n72895 , n72896 );
and ( n72898 , n66140 , n40855 );
nor ( n72899 , n72897 , n72898 );
not ( n72900 , n72899 );
nand ( n72901 , n72900 , n70930 );
nand ( n72902 , n72894 , n72901 );
not ( n72903 , n72902 );
xor ( n72904 , n72890 , n72903 );
not ( n72905 , n72142 );
not ( n72906 , n72548 );
or ( n72907 , n72905 , n72906 );
not ( n72908 , n40364 );
not ( n72909 , n54302 );
or ( n72910 , n72908 , n72909 );
nand ( n72911 , n54811 , n54725 );
nand ( n72912 , n72910 , n72911 );
nand ( n72913 , n72912 , n54327 );
nand ( n72914 , n72907 , n72913 );
xor ( n72915 , n72904 , n72914 );
not ( n72916 , n70193 );
not ( n72917 , n72560 );
or ( n72918 , n72916 , n72917 );
buf ( n72919 , n55582 );
not ( n72920 , n72919 );
not ( n72921 , n53289 );
or ( n72922 , n72920 , n72921 );
not ( n72923 , n55582 );
nand ( n72924 , n72923 , n54646 );
nand ( n72925 , n72922 , n72924 );
nand ( n72926 , n72925 , n70183 );
nand ( n72927 , n72918 , n72926 );
not ( n72928 , n67862 );
not ( n72929 , n72571 );
or ( n72930 , n72928 , n72929 );
not ( n72931 , n72288 );
not ( n72932 , n40627 );
or ( n72933 , n72931 , n72932 );
nand ( n72934 , n68049 , n55846 );
nand ( n72935 , n72933 , n72934 );
nand ( n72936 , n72935 , n59984 );
nand ( n72937 , n72930 , n72936 );
xor ( n72938 , n72927 , n72937 );
not ( n72939 , n56777 );
not ( n72940 , n72595 );
or ( n72941 , n72939 , n72940 );
not ( n72942 , n69820 );
not ( n72943 , n40528 );
or ( n72944 , n72942 , n72943 );
not ( n72945 , n40527 );
nand ( n72946 , n72945 , n56785 );
nand ( n72947 , n72944 , n72946 );
nand ( n72948 , n72947 , n72185 );
nand ( n72949 , n72941 , n72948 );
xor ( n72950 , n72938 , n72949 );
xor ( n72951 , n72915 , n72950 );
not ( n72952 , n67568 );
not ( n72953 , n70638 );
or ( n72954 , n72952 , n72953 );
not ( n72955 , n40733 );
nand ( n72956 , n72955 , n67890 );
nand ( n72957 , n72954 , n72956 );
not ( n72958 , n72957 );
not ( n72959 , n70604 );
or ( n72960 , n72958 , n72959 );
buf ( n72961 , n60482 );
not ( n72962 , n72961 );
or ( n72963 , n72716 , n72962 );
nand ( n72964 , n72960 , n72963 );
or ( n72965 , n72609 , n52124 );
not ( n72966 , n56455 );
not ( n72967 , n52487 );
and ( n72968 , n72966 , n72967 );
not ( n72969 , n67193 );
and ( n72970 , n72969 , n52113 );
nor ( n72971 , n72968 , n72970 );
or ( n72972 , n72971 , n62302 );
nand ( n72973 , n72965 , n72972 );
xor ( n72974 , n72964 , n72973 );
not ( n72975 , n72529 );
or ( n72976 , n72975 , n70585 );
not ( n72977 , n69458 );
not ( n72978 , n55630 );
or ( n72979 , n72977 , n72978 );
not ( n72980 , n52841 );
nand ( n72981 , n72980 , n72217 );
nand ( n72982 , n72979 , n72981 );
not ( n72983 , n72982 );
or ( n72984 , n72983 , n56861 );
nand ( n72985 , n72976 , n72984 );
xor ( n72986 , n72974 , n72985 );
xor ( n72987 , n72951 , n72986 );
xor ( n72988 , n72915 , n72950 );
and ( n72989 , n72988 , n72986 );
and ( n72990 , n72915 , n72950 );
or ( n72991 , n72989 , n72990 );
not ( n72992 , n59950 );
not ( n72993 , n72693 );
or ( n72994 , n72992 , n72993 );
not ( n72995 , n59345 );
not ( n72996 , n69961 );
or ( n72997 , n72995 , n72996 );
not ( n72998 , n72252 );
nand ( n72999 , n72998 , n65743 );
nand ( n73000 , n72997 , n72999 );
nand ( n73001 , n73000 , n56639 );
nand ( n73002 , n72994 , n73001 );
xor ( n73003 , n72473 , n73002 );
xor ( n73004 , n73003 , n72509 );
xor ( n73005 , n72796 , n73004 );
not ( n73006 , n62654 );
not ( n73007 , n61951 );
not ( n73008 , n69072 );
or ( n73009 , n73007 , n73008 );
nand ( n73010 , n71547 , n66690 );
nand ( n73011 , n73009 , n73010 );
not ( n73012 , n73011 );
or ( n73013 , n73006 , n73012 );
nand ( n73014 , n72634 , n66696 );
nand ( n73015 , n73013 , n73014 );
not ( n73016 , n52022 );
not ( n73017 , n72684 );
or ( n73018 , n73016 , n73017 );
nand ( n73019 , n54623 , n59174 );
nand ( n73020 , n73018 , n73019 );
xor ( n73021 , n73015 , n73020 );
or ( n73022 , n72658 , n59820 );
and ( n73023 , n64191 , n68206 );
not ( n73024 , n64191 );
and ( n73025 , n73024 , n39714 );
or ( n73026 , n73023 , n73025 );
or ( n73027 , n73026 , n59828 );
nand ( n73028 , n73022 , n73027 );
xor ( n73029 , n73021 , n73028 );
xor ( n73030 , n73005 , n73029 );
xor ( n73031 , n72796 , n73004 );
and ( n73032 , n73031 , n73029 );
and ( n73033 , n72796 , n73004 );
or ( n73034 , n73032 , n73033 );
not ( n73035 , n51533 );
not ( n73036 , n53931 );
not ( n73037 , n60167 );
or ( n73038 , n73036 , n73037 );
nand ( n73039 , n39847 , n71053 );
nand ( n73040 , n73038 , n73039 );
not ( n73041 , n73040 );
or ( n73042 , n73035 , n73041 );
nand ( n73043 , n72585 , n72198 );
nand ( n73044 , n73042 , n73043 );
not ( n73045 , n58977 );
and ( n73046 , n62577 , n67269 );
not ( n73047 , n62577 );
not ( n73048 , n66301 );
and ( n73049 , n73047 , n73048 );
or ( n73050 , n73046 , n73049 );
not ( n73051 , n73050 );
not ( n73052 , n73051 );
or ( n73053 , n73045 , n73052 );
not ( n73054 , n72646 );
nand ( n73055 , n73054 , n59633 );
nand ( n73056 , n73053 , n73055 );
xor ( n73057 , n73044 , n73056 );
not ( n73058 , n62085 );
not ( n73059 , n72624 );
not ( n73060 , n73059 );
or ( n73061 , n73058 , n73060 );
buf ( n73062 , n62960 );
and ( n73063 , n69893 , n73062 );
not ( n73064 , n69893 );
not ( n73065 , n73062 );
and ( n73066 , n73064 , n73065 );
or ( n73067 , n73063 , n73066 );
not ( n73068 , n73067 );
nand ( n73069 , n73068 , n52191 );
nand ( n73070 , n73061 , n73069 );
xor ( n73071 , n73057 , n73070 );
xor ( n73072 , n73071 , n72808 );
xor ( n73073 , n73072 , n72515 );
xor ( n73074 , n73071 , n72808 );
and ( n73075 , n73074 , n72515 );
and ( n73076 , n73071 , n72808 );
or ( n73077 , n73075 , n73076 );
not ( n73078 , n52151 );
not ( n73079 , n72674 );
or ( n73080 , n73078 , n73079 );
not ( n73081 , n57187 );
not ( n73082 , n67040 );
or ( n73083 , n73081 , n73082 );
nand ( n73084 , n71509 , n71042 );
nand ( n73085 , n73083 , n73084 );
nand ( n73086 , n73085 , n50922 );
nand ( n73087 , n73080 , n73086 );
xor ( n73088 , n73087 , n72870 );
xor ( n73089 , n73088 , n72841 );
xor ( n73090 , n73089 , n72521 );
xor ( n73091 , n73090 , n72618 );
xor ( n73092 , n73089 , n72521 );
and ( n73093 , n73092 , n72618 );
and ( n73094 , n73089 , n72521 );
or ( n73095 , n73093 , n73094 );
xor ( n73096 , n72762 , n72784 );
xor ( n73097 , n73096 , n72788 );
xor ( n73098 , n73097 , n72987 );
xor ( n73099 , n73098 , n72876 );
xor ( n73100 , n73097 , n72987 );
and ( n73101 , n73100 , n72876 );
and ( n73102 , n73097 , n72987 );
or ( n73103 , n73101 , n73102 );
xor ( n73104 , n72666 , n72728 );
xor ( n73105 , n73104 , n73030 );
xor ( n73106 , n72666 , n72728 );
and ( n73107 , n73106 , n73030 );
and ( n73108 , n72666 , n72728 );
or ( n73109 , n73107 , n73108 );
xor ( n73110 , n72734 , n73073 );
xor ( n73111 , n73110 , n73091 );
xor ( n73112 , n72734 , n73073 );
and ( n73113 , n73112 , n73091 );
and ( n73114 , n72734 , n73073 );
or ( n73115 , n73113 , n73114 );
xor ( n73116 , n72740 , n72746 );
xor ( n73117 , n73116 , n73099 );
xor ( n73118 , n72740 , n72746 );
and ( n73119 , n73118 , n73099 );
and ( n73120 , n72740 , n72746 );
or ( n73121 , n73119 , n73120 );
xor ( n73122 , n73105 , n73111 );
xor ( n73123 , n73122 , n72752 );
xor ( n73124 , n73105 , n73111 );
and ( n73125 , n73124 , n72752 );
and ( n73126 , n73105 , n73111 );
or ( n73127 , n73125 , n73126 );
xor ( n73128 , n72964 , n72973 );
and ( n73129 , n73128 , n72985 );
and ( n73130 , n72964 , n72973 );
or ( n73131 , n73129 , n73130 );
xor ( n73132 , n73117 , n72758 );
xor ( n73133 , n73132 , n72768 );
xor ( n73134 , n73117 , n72758 );
and ( n73135 , n73134 , n72768 );
and ( n73136 , n73117 , n72758 );
or ( n73137 , n73135 , n73136 );
xor ( n73138 , n73123 , n73133 );
xor ( n73139 , n73138 , n72774 );
xor ( n73140 , n73123 , n73133 );
and ( n73141 , n73140 , n72774 );
and ( n73142 , n73123 , n73133 );
or ( n73143 , n73141 , n73142 );
xor ( n73144 , n72890 , n72903 );
and ( n73145 , n73144 , n72914 );
and ( n73146 , n72890 , n72903 );
or ( n73147 , n73145 , n73146 );
xor ( n73148 , n72927 , n72937 );
and ( n73149 , n73148 , n72949 );
and ( n73150 , n72927 , n72937 );
or ( n73151 , n73149 , n73150 );
xor ( n73152 , n73044 , n73056 );
and ( n73153 , n73152 , n73070 );
and ( n73154 , n73044 , n73056 );
or ( n73155 , n73153 , n73154 );
xor ( n73156 , n73015 , n73020 );
and ( n73157 , n73156 , n73028 );
and ( n73158 , n73015 , n73020 );
or ( n73159 , n73157 , n73158 );
xor ( n73160 , n72473 , n73002 );
and ( n73161 , n73160 , n72509 );
and ( n73162 , n72473 , n73002 );
or ( n73163 , n73161 , n73162 );
xor ( n73164 , n73087 , n72870 );
and ( n73165 , n73164 , n72841 );
and ( n73166 , n73087 , n72870 );
or ( n73167 , n73165 , n73166 );
xor ( n73168 , n72762 , n72784 );
and ( n73169 , n73168 , n72788 );
and ( n73170 , n72762 , n72784 );
or ( n73171 , n73169 , n73170 );
not ( n73172 , n54622 );
not ( n73173 , n66735 );
or ( n73174 , n73172 , n73173 );
nand ( n73175 , n73174 , n59174 );
not ( n73176 , n72853 );
not ( n73177 , n70915 );
or ( n73178 , n73176 , n73177 );
not ( n73179 , n59340 );
not ( n73180 , n70889 );
or ( n73181 , n73179 , n73180 );
not ( n73182 , n52079 );
nand ( n73183 , n73182 , n62513 );
nand ( n73184 , n73181 , n73183 );
nand ( n73185 , n59575 , n73184 );
nand ( n73186 , n73178 , n73185 );
xor ( n73187 , n73175 , n73186 );
or ( n73188 , n60960 , n72899 );
not ( n73189 , n70930 );
not ( n73190 , n70506 );
and ( n73191 , n71691 , n73190 );
not ( n73192 , n71691 );
and ( n73193 , n73192 , n70506 );
nor ( n73194 , n73191 , n73193 );
or ( n73195 , n73189 , n73194 );
nand ( n73196 , n73188 , n73195 );
xor ( n73197 , n73187 , n73196 );
xor ( n73198 , n73175 , n73186 );
and ( n73199 , n73198 , n73196 );
and ( n73200 , n73175 , n73186 );
or ( n73201 , n73199 , n73200 );
not ( n73202 , n72818 );
not ( n73203 , n61550 );
or ( n73204 , n73202 , n73203 );
not ( n73205 , n53706 );
not ( n73206 , n61417 );
or ( n73207 , n73205 , n73206 );
nand ( n73208 , n61416 , n52796 );
nand ( n73209 , n73207 , n73208 );
nand ( n73210 , n61558 , n73209 );
nand ( n73211 , n73204 , n73210 );
not ( n73212 , n72828 );
not ( n73213 , n67061 );
or ( n73214 , n73212 , n73213 );
not ( n73215 , n67441 );
not ( n73216 , n64167 );
or ( n73217 , n73215 , n73216 );
nand ( n73218 , n62451 , n48679 );
nand ( n73219 , n73217 , n73218 );
nand ( n73220 , n67068 , n73219 );
nand ( n73221 , n73214 , n73220 );
xor ( n73222 , n73211 , n73221 );
or ( n73223 , n71959 , n72837 );
not ( n73224 , n62319 );
not ( n73225 , n63415 );
or ( n73226 , n73224 , n73225 );
nand ( n73227 , n67969 , n44112 );
nand ( n73228 , n73226 , n73227 );
not ( n73229 , n73228 );
or ( n73230 , n70965 , n73229 );
nand ( n73231 , n73223 , n73230 );
xor ( n73232 , n73222 , n73231 );
xor ( n73233 , n73211 , n73221 );
and ( n73234 , n73233 , n73231 );
and ( n73235 , n73211 , n73221 );
or ( n73236 , n73234 , n73235 );
xor ( n73237 , n73151 , n73159 );
xor ( n73238 , n73237 , n73163 );
xor ( n73239 , n73151 , n73159 );
and ( n73240 , n73239 , n73163 );
and ( n73241 , n73151 , n73159 );
or ( n73242 , n73240 , n73241 );
not ( n73243 , n59984 );
not ( n73244 , n72288 );
not ( n73245 , n54415 );
or ( n73246 , n73244 , n73245 );
nand ( n73247 , n59612 , n55846 );
nand ( n73248 , n73246 , n73247 );
not ( n73249 , n73248 );
or ( n73250 , n73243 , n73249 );
nand ( n73251 , n72935 , n71099 );
nand ( n73252 , n73250 , n73251 );
not ( n73253 , n56777 );
not ( n73254 , n72947 );
or ( n73255 , n73253 , n73254 );
not ( n73256 , n40592 );
not ( n73257 , n56785 );
or ( n73258 , n73256 , n73257 );
nand ( n73259 , n53730 , n56786 );
nand ( n73260 , n73258 , n73259 );
nand ( n73261 , n73260 , n60472 );
nand ( n73262 , n73255 , n73261 );
xor ( n73263 , n73252 , n73262 );
not ( n73264 , n56355 );
not ( n73265 , n73040 );
or ( n73266 , n73264 , n73265 );
not ( n73267 , n53931 );
not ( n73268 , n68510 );
not ( n73269 , n73268 );
or ( n73270 , n73267 , n73269 );
not ( n73271 , n68507 );
nand ( n73272 , n73271 , n71053 );
nand ( n73273 , n73270 , n73272 );
nand ( n73274 , n73273 , n51533 );
nand ( n73275 , n73266 , n73274 );
xor ( n73276 , n73263 , n73275 );
not ( n73277 , n54327 );
not ( n73278 , n71395 );
buf ( n73279 , n40148 );
not ( n73280 , n73279 );
or ( n73281 , n73278 , n73280 );
not ( n73282 , n70627 );
nand ( n73283 , n73282 , n71067 );
nand ( n73284 , n73281 , n73283 );
not ( n73285 , n73284 );
or ( n73286 , n73277 , n73285 );
nand ( n73287 , n72912 , n54316 );
nand ( n73288 , n73286 , n73287 );
not ( n73289 , n70183 );
not ( n73290 , n55120 );
not ( n73291 , n71073 );
not ( n73292 , n73291 );
or ( n73293 , n73290 , n73292 );
nand ( n73294 , n40226 , n71409 );
nand ( n73295 , n73293 , n73294 );
not ( n73296 , n73295 );
or ( n73297 , n73289 , n73296 );
nand ( n73298 , n55144 , n72925 );
nand ( n73299 , n73297 , n73298 );
xor ( n73300 , n73288 , n73299 );
xor ( n73301 , n73300 , n72902 );
xor ( n73302 , n73276 , n73301 );
not ( n73303 , n70604 );
not ( n73304 , n66963 );
not ( n73305 , n51601 );
or ( n73306 , n73304 , n73305 );
buf ( n73307 , n66963 );
or ( n73308 , n73307 , n52223 );
nand ( n73309 , n73306 , n73308 );
not ( n73310 , n73309 );
or ( n73311 , n73303 , n73310 );
nand ( n73312 , n72957 , n72182 );
nand ( n73313 , n73311 , n73312 );
not ( n73314 , n53571 );
not ( n73315 , n52841 );
not ( n73316 , n70290 );
or ( n73317 , n73315 , n73316 );
nand ( n73318 , n67721 , n55104 );
nand ( n73319 , n73317 , n73318 );
not ( n73320 , n73319 );
or ( n73321 , n73314 , n73320 );
nand ( n73322 , n72982 , n53182 );
nand ( n73323 , n73321 , n73322 );
xor ( n73324 , n73313 , n73323 );
not ( n73325 , n53620 );
not ( n73326 , n53596 );
not ( n73327 , n71052 );
not ( n73328 , n73327 );
or ( n73329 , n73326 , n73328 );
nand ( n73330 , n40382 , n71756 );
nand ( n73331 , n73329 , n73330 );
not ( n73332 , n73331 );
or ( n73333 , n73325 , n73332 );
nand ( n73334 , n72888 , n68603 );
nand ( n73335 , n73333 , n73334 );
xor ( n73336 , n73324 , n73335 );
xor ( n73337 , n73302 , n73336 );
xor ( n73338 , n73276 , n73301 );
and ( n73339 , n73338 , n73336 );
and ( n73340 , n73276 , n73301 );
or ( n73341 , n73339 , n73340 );
and ( n73342 , n72846 , n58458 );
and ( n73343 , n51574 , n62496 );
not ( n73344 , n51574 );
and ( n73345 , n73344 , n62497 );
or ( n73346 , n73343 , n73345 );
not ( n73347 , n73346 );
or ( n73348 , n73347 , n71467 );
not ( n73349 , n71689 );
nand ( n73350 , n73349 , n72865 );
nand ( n73351 , n73348 , n73350 );
xor ( n73352 , n73342 , n73351 );
not ( n73353 , n72220 );
not ( n73354 , n52114 );
not ( n73355 , n39963 );
or ( n73356 , n73354 , n73355 );
buf ( n73357 , n57801 );
nand ( n73358 , n73357 , n52130 );
nand ( n73359 , n73356 , n73358 );
not ( n73360 , n73359 );
or ( n73361 , n73353 , n73360 );
or ( n73362 , n72971 , n52481 );
nand ( n73363 , n73361 , n73362 );
xor ( n73364 , n73352 , n73363 );
xor ( n73365 , n73364 , n73155 );
or ( n73366 , n73050 , n59632 );
not ( n73367 , n66784 );
not ( n73368 , n73367 );
not ( n73369 , n52728 );
and ( n73370 , n73368 , n73369 );
not ( n73371 , n71162 );
not ( n73372 , n73371 );
and ( n73373 , n73372 , n52728 );
nor ( n73374 , n73370 , n73373 );
or ( n73375 , n73374 , n59630 );
nand ( n73376 , n73366 , n73375 );
not ( n73377 , n62085 );
or ( n73378 , n73067 , n73377 );
xor ( n73379 , n60289 , n69530 );
or ( n73380 , n73379 , n59811 );
nand ( n73381 , n73378 , n73380 );
xor ( n73382 , n73376 , n73381 );
not ( n73383 , n73011 );
or ( n73384 , n73383 , n72628 );
not ( n73385 , n61951 );
not ( n73386 , n62394 );
or ( n73387 , n73385 , n73386 );
nand ( n73388 , n67482 , n66690 );
nand ( n73389 , n73387 , n73388 );
not ( n73390 , n73389 );
or ( n73391 , n73390 , n72636 );
nand ( n73392 , n73384 , n73391 );
xor ( n73393 , n73382 , n73392 );
xor ( n73394 , n73365 , n73393 );
xor ( n73395 , n73364 , n73155 );
and ( n73396 , n73395 , n73393 );
and ( n73397 , n73364 , n73155 );
or ( n73398 , n73396 , n73397 );
or ( n73399 , n73026 , n59820 );
not ( n73400 , n39574 );
and ( n73401 , n66705 , n73400 );
not ( n73402 , n66705 );
and ( n73403 , n73402 , n68667 );
or ( n73404 , n73401 , n73403 );
or ( n73405 , n73404 , n59828 );
nand ( n73406 , n73399 , n73405 );
xor ( n73407 , n73406 , n72845 );
not ( n73408 , n73000 );
not ( n73409 , n59950 );
or ( n73410 , n73408 , n73409 );
and ( n73411 , n65743 , n68381 );
not ( n73412 , n65743 );
and ( n73413 , n73412 , n42399 );
nor ( n73414 , n73411 , n73413 );
or ( n73415 , n73414 , n68961 );
nand ( n73416 , n73410 , n73415 );
xor ( n73417 , n73407 , n73416 );
xor ( n73418 , n73167 , n73417 );
xor ( n73419 , n73418 , n73171 );
xor ( n73420 , n73167 , n73417 );
and ( n73421 , n73420 , n73171 );
and ( n73422 , n73167 , n73417 );
or ( n73423 , n73421 , n73422 );
not ( n73424 , n52151 );
not ( n73425 , n73085 );
or ( n73426 , n73424 , n73425 );
not ( n73427 , n51465 );
not ( n73428 , n66546 );
not ( n73429 , n73428 );
or ( n73430 , n73427 , n73429 );
nand ( n73431 , n66546 , n71042 );
nand ( n73432 , n73430 , n73431 );
nand ( n73433 , n73432 , n50922 );
nand ( n73434 , n73426 , n73433 );
xor ( n73435 , n73434 , n73232 );
xor ( n73436 , n73435 , n73197 );
xor ( n73437 , n73436 , n72880 );
xor ( n73438 , n73437 , n72991 );
xor ( n73439 , n73436 , n72880 );
and ( n73440 , n73439 , n72991 );
and ( n73441 , n73436 , n72880 );
or ( n73442 , n73440 , n73441 );
xor ( n73443 , n72874 , n73131 );
xor ( n73444 , n73443 , n73147 );
xor ( n73445 , n73444 , n73034 );
xor ( n73446 , n73445 , n73394 );
xor ( n73447 , n73444 , n73034 );
and ( n73448 , n73447 , n73394 );
and ( n73449 , n73444 , n73034 );
or ( n73450 , n73448 , n73449 );
xor ( n73451 , n73337 , n73238 );
xor ( n73452 , n73451 , n73077 );
xor ( n73453 , n73337 , n73238 );
and ( n73454 , n73453 , n73077 );
and ( n73455 , n73337 , n73238 );
or ( n73456 , n73454 , n73455 );
xor ( n73457 , n73419 , n73095 );
xor ( n73458 , n73457 , n73103 );
xor ( n73459 , n73419 , n73095 );
and ( n73460 , n73459 , n73103 );
and ( n73461 , n73419 , n73095 );
or ( n73462 , n73460 , n73461 );
xor ( n73463 , n73438 , n73109 );
xor ( n73464 , n73463 , n73452 );
xor ( n73465 , n73438 , n73109 );
and ( n73466 , n73465 , n73452 );
and ( n73467 , n73438 , n73109 );
or ( n73468 , n73466 , n73467 );
xor ( n73469 , n73446 , n73458 );
xor ( n73470 , n73469 , n73115 );
xor ( n73471 , n73446 , n73458 );
and ( n73472 , n73471 , n73115 );
and ( n73473 , n73446 , n73458 );
or ( n73474 , n73472 , n73473 );
xor ( n73475 , n73342 , n73351 );
and ( n73476 , n73475 , n73363 );
and ( n73477 , n73342 , n73351 );
or ( n73478 , n73476 , n73477 );
xor ( n73479 , n73121 , n73464 );
xor ( n73480 , n73479 , n73127 );
xor ( n73481 , n73121 , n73464 );
and ( n73482 , n73481 , n73127 );
and ( n73483 , n73121 , n73464 );
or ( n73484 , n73482 , n73483 );
xor ( n73485 , n73470 , n73480 );
xor ( n73486 , n73485 , n73137 );
xor ( n73487 , n73470 , n73480 );
and ( n73488 , n73487 , n73137 );
and ( n73489 , n73470 , n73480 );
or ( n73490 , n73488 , n73489 );
xor ( n73491 , n73313 , n73323 );
and ( n73492 , n73491 , n73335 );
and ( n73493 , n73313 , n73323 );
or ( n73494 , n73492 , n73493 );
xor ( n73495 , n73288 , n73299 );
and ( n73496 , n73495 , n72902 );
and ( n73497 , n73288 , n73299 );
or ( n73498 , n73496 , n73497 );
xor ( n73499 , n73252 , n73262 );
and ( n73500 , n73499 , n73275 );
and ( n73501 , n73252 , n73262 );
or ( n73502 , n73500 , n73501 );
xor ( n73503 , n73376 , n73381 );
and ( n73504 , n73503 , n73392 );
and ( n73505 , n73376 , n73381 );
or ( n73506 , n73504 , n73505 );
xor ( n73507 , n73406 , n72845 );
and ( n73508 , n73507 , n73416 );
and ( n73509 , n73406 , n72845 );
or ( n73510 , n73508 , n73509 );
xor ( n73511 , n73434 , n73232 );
and ( n73512 , n73511 , n73197 );
and ( n73513 , n73434 , n73232 );
or ( n73514 , n73512 , n73513 );
xor ( n73515 , n72874 , n73131 );
and ( n73516 , n73515 , n73147 );
and ( n73517 , n72874 , n73131 );
or ( n73518 , n73516 , n73517 );
not ( n73519 , n73209 );
not ( n73520 , n61548 );
or ( n73521 , n73519 , n73520 );
not ( n73522 , n50008 );
not ( n73523 , n61939 );
or ( n73524 , n73522 , n73523 );
nand ( n73525 , n64633 , n50004 );
nand ( n73526 , n73524 , n73525 );
nand ( n73527 , n73526 , n62428 );
nand ( n73528 , n73521 , n73527 );
not ( n73529 , n73228 );
not ( n73530 , n63410 );
or ( n73531 , n73529 , n73530 );
not ( n73532 , n48486 );
not ( n73533 , n63415 );
or ( n73534 , n73532 , n73533 );
nand ( n73535 , n63681 , n48951 );
nand ( n73536 , n73534 , n73535 );
nand ( n73537 , n63398 , n73536 );
nand ( n73538 , n73531 , n73537 );
xor ( n73539 , n73528 , n73538 );
not ( n73540 , n73219 );
not ( n73541 , n62463 );
or ( n73542 , n73540 , n73541 );
not ( n73543 , n64166 );
not ( n73544 , n52592 );
not ( n73545 , n66089 );
or ( n73546 , n73544 , n73545 );
not ( n73547 , n64687 );
nand ( n73548 , n73547 , n41287 );
nand ( n73549 , n73546 , n73548 );
nand ( n73550 , n73543 , n73549 );
nand ( n73551 , n73542 , n73550 );
xor ( n73552 , n73539 , n73551 );
xor ( n73553 , n73528 , n73538 );
and ( n73554 , n73553 , n73551 );
and ( n73555 , n73528 , n73538 );
or ( n73556 , n73554 , n73555 );
and ( n73557 , n72846 , n58915 );
not ( n73558 , n59575 );
not ( n73559 , n72464 );
not ( n73560 , n50654 );
or ( n73561 , n73559 , n73560 );
nand ( n73562 , n40692 , n59340 );
nand ( n73563 , n73561 , n73562 );
not ( n73564 , n73563 );
or ( n73565 , n73558 , n73564 );
not ( n73566 , n67584 );
nand ( n73567 , n73566 , n73184 );
nand ( n73568 , n73565 , n73567 );
xor ( n73569 , n73557 , n73568 );
not ( n73570 , n71466 );
not ( n73571 , n62496 );
not ( n73572 , n40733 );
or ( n73573 , n73571 , n73572 );
nand ( n73574 , n54032 , n66652 );
nand ( n73575 , n73573 , n73574 );
not ( n73576 , n73575 );
or ( n73577 , n73570 , n73576 );
nand ( n73578 , n73346 , n72106 );
nand ( n73579 , n73577 , n73578 );
xor ( n73580 , n73569 , n73579 );
xor ( n73581 , n73557 , n73568 );
and ( n73582 , n73581 , n73579 );
and ( n73583 , n73557 , n73568 );
or ( n73584 , n73582 , n73583 );
not ( n73585 , n56777 );
not ( n73586 , n73260 );
or ( n73587 , n73585 , n73586 );
not ( n73588 , n69820 );
not ( n73589 , n40627 );
or ( n73590 , n73588 , n73589 );
nand ( n73591 , n40626 , n67454 );
nand ( n73592 , n73590 , n73591 );
nand ( n73593 , n73592 , n60472 );
nand ( n73594 , n73587 , n73593 );
not ( n73595 , n73309 );
not ( n73596 , n72182 );
or ( n73597 , n73595 , n73596 );
not ( n73598 , n66642 );
not ( n73599 , n52570 );
or ( n73600 , n73598 , n73599 );
nand ( n73601 , n51916 , n66963 );
nand ( n73602 , n73600 , n73601 );
nand ( n73603 , n73602 , n72710 );
nand ( n73604 , n73597 , n73603 );
xor ( n73605 , n73594 , n73604 );
not ( n73606 , n51766 );
not ( n73607 , n52487 );
not ( n73608 , n73607 );
not ( n73609 , n62970 );
or ( n73610 , n73608 , n73609 );
nand ( n73611 , n66215 , n52130 );
nand ( n73612 , n73610 , n73611 );
not ( n73613 , n73612 );
or ( n73614 , n73606 , n73613 );
nand ( n73615 , n73359 , n52482 );
nand ( n73616 , n73614 , n73615 );
xor ( n73617 , n73605 , n73616 );
not ( n73618 , n52854 );
not ( n73619 , n73319 );
or ( n73620 , n73618 , n73619 );
not ( n73621 , n54283 );
not ( n73622 , n63180 );
or ( n73623 , n73621 , n73622 );
nand ( n73624 , n67196 , n55104 );
nand ( n73625 , n73623 , n73624 );
nand ( n73626 , n73625 , n53571 );
nand ( n73627 , n73620 , n73626 );
not ( n73628 , n53620 );
not ( n73629 , n55089 );
not ( n73630 , n70661 );
or ( n73631 , n73629 , n73630 );
nand ( n73632 , n68980 , n69444 );
nand ( n73633 , n73631 , n73632 );
not ( n73634 , n73633 );
or ( n73635 , n73628 , n73634 );
nand ( n73636 , n73331 , n68603 );
nand ( n73637 , n73635 , n73636 );
xor ( n73638 , n73627 , n73637 );
not ( n73639 , n54316 );
not ( n73640 , n73284 );
or ( n73641 , n73639 , n73640 );
not ( n73642 , n71395 );
not ( n73643 , n57390 );
or ( n73644 , n73642 , n73643 );
nand ( n73645 , n68990 , n55276 );
nand ( n73646 , n73644 , n73645 );
nand ( n73647 , n73646 , n54327 );
nand ( n73648 , n73641 , n73647 );
xor ( n73649 , n73638 , n73648 );
xor ( n73650 , n73617 , n73649 );
xor ( n73651 , n73650 , n73510 );
xor ( n73652 , n73617 , n73649 );
and ( n73653 , n73652 , n73510 );
and ( n73654 , n73617 , n73649 );
or ( n73655 , n73653 , n73654 );
xor ( n73656 , n73502 , n73506 );
or ( n73657 , n73379 , n73377 );
not ( n73658 , n66234 );
not ( n73659 , n66052 );
or ( n73660 , n73658 , n73659 );
nand ( n73661 , n66053 , n60289 );
nand ( n73662 , n73660 , n73661 );
not ( n73663 , n73662 );
or ( n73664 , n73663 , n59811 );
nand ( n73665 , n73657 , n73664 );
xor ( n73666 , n73236 , n73665 );
not ( n73667 , n72198 );
not ( n73668 , n73273 );
or ( n73669 , n73667 , n73668 );
not ( n73670 , n53931 );
not ( n73671 , n67040 );
or ( n73672 , n73670 , n73671 );
nand ( n73673 , n71509 , n71445 );
nand ( n73674 , n73672 , n73673 );
nand ( n73675 , n73674 , n51533 );
nand ( n73676 , n73669 , n73675 );
xor ( n73677 , n73666 , n73676 );
xor ( n73678 , n73656 , n73677 );
xor ( n73679 , n73502 , n73506 );
and ( n73680 , n73679 , n73677 );
and ( n73681 , n73502 , n73506 );
or ( n73682 , n73680 , n73681 );
or ( n73683 , n73414 , n73409 );
not ( n73684 , n73048 );
not ( n73685 , n65743 );
and ( n73686 , n73684 , n73685 );
and ( n73687 , n73048 , n65743 );
nor ( n73688 , n73686 , n73687 );
or ( n73689 , n68961 , n73688 );
nand ( n73690 , n73683 , n73689 );
not ( n73691 , n62654 );
not ( n73692 , n61951 );
not ( n73693 , n62959 );
or ( n73694 , n73692 , n73693 );
nand ( n73695 , n39332 , n61952 );
nand ( n73696 , n73694 , n73695 );
not ( n73697 , n73696 );
or ( n73698 , n73691 , n73697 );
nand ( n73699 , n73389 , n66696 );
nand ( n73700 , n73698 , n73699 );
xor ( n73701 , n73690 , n73700 );
or ( n73702 , n73404 , n59820 );
not ( n73703 , n64190 );
not ( n73704 , n69072 );
or ( n73705 , n73703 , n73704 );
nand ( n73706 , n39056 , n66705 );
nand ( n73707 , n73705 , n73706 );
not ( n73708 , n73707 );
or ( n73709 , n73708 , n59828 );
nand ( n73710 , n73702 , n73709 );
xor ( n73711 , n73701 , n73710 );
xor ( n73712 , n73711 , n73514 );
not ( n73713 , n58977 );
not ( n73714 , n58982 );
or ( n73715 , n73713 , n73714 );
or ( n73716 , n73374 , n49420 );
nand ( n73717 , n73715 , n73716 );
not ( n73718 , n52151 );
not ( n73719 , n73432 );
or ( n73720 , n73718 , n73719 );
not ( n73721 , n50895 );
not ( n73722 , n62931 );
or ( n73723 , n73721 , n73722 );
nand ( n73724 , n71567 , n50916 );
nand ( n73725 , n73723 , n73724 );
nand ( n73726 , n73725 , n50922 );
nand ( n73727 , n73720 , n73726 );
xor ( n73728 , n73717 , n73727 );
xor ( n73729 , n73728 , n73201 );
xor ( n73730 , n73712 , n73729 );
xor ( n73731 , n73711 , n73514 );
and ( n73732 , n73731 , n73729 );
and ( n73733 , n73711 , n73514 );
or ( n73734 , n73732 , n73733 );
xor ( n73735 , n73494 , n73498 );
not ( n73736 , n73194 );
not ( n73737 , n73736 );
not ( n73738 , n70500 );
or ( n73739 , n73737 , n73738 );
not ( n73740 , n51891 );
not ( n73741 , n66141 );
or ( n73742 , n73740 , n73741 );
nand ( n73743 , n68878 , n63930 );
nand ( n73744 , n73742 , n73743 );
nand ( n73745 , n70930 , n73744 );
nand ( n73746 , n73739 , n73745 );
not ( n73747 , n73746 );
not ( n73748 , n55144 );
not ( n73749 , n73295 );
or ( n73750 , n73748 , n73749 );
not ( n73751 , n55582 );
not ( n73752 , n63201 );
or ( n73753 , n73751 , n73752 );
nand ( n73754 , n59195 , n55148 );
nand ( n73755 , n73753 , n73754 );
nand ( n73756 , n73755 , n70183 );
nand ( n73757 , n73750 , n73756 );
xor ( n73758 , n73747 , n73757 );
not ( n73759 , n71099 );
not ( n73760 , n73248 );
or ( n73761 , n73759 , n73760 );
not ( n73762 , n55846 );
not ( n73763 , n40377 );
or ( n73764 , n73762 , n73763 );
not ( n73765 , n72148 );
nand ( n73766 , n73765 , n72288 );
nand ( n73767 , n73764 , n73766 );
nand ( n73768 , n73767 , n55458 );
nand ( n73769 , n73761 , n73768 );
xor ( n73770 , n73758 , n73769 );
xor ( n73771 , n73735 , n73770 );
xor ( n73772 , n73518 , n73771 );
xor ( n73773 , n73772 , n73341 );
xor ( n73774 , n73518 , n73771 );
and ( n73775 , n73774 , n73341 );
and ( n73776 , n73518 , n73771 );
or ( n73777 , n73775 , n73776 );
xor ( n73778 , n73552 , n73580 );
xor ( n73779 , n73778 , n73478 );
xor ( n73780 , n73242 , n73779 );
xor ( n73781 , n73780 , n73398 );
xor ( n73782 , n73242 , n73779 );
and ( n73783 , n73782 , n73398 );
and ( n73784 , n73242 , n73779 );
or ( n73785 , n73783 , n73784 );
xor ( n73786 , n73678 , n73651 );
xor ( n73787 , n73786 , n73730 );
xor ( n73788 , n73678 , n73651 );
and ( n73789 , n73788 , n73730 );
and ( n73790 , n73678 , n73651 );
or ( n73791 , n73789 , n73790 );
xor ( n73792 , n73423 , n73442 );
xor ( n73793 , n73792 , n73781 );
xor ( n73794 , n73423 , n73442 );
and ( n73795 , n73794 , n73781 );
and ( n73796 , n73423 , n73442 );
or ( n73797 , n73795 , n73796 );
xor ( n73798 , n73450 , n73773 );
xor ( n73799 , n73798 , n73787 );
xor ( n73800 , n73450 , n73773 );
and ( n73801 , n73800 , n73787 );
and ( n73802 , n73450 , n73773 );
or ( n73803 , n73801 , n73802 );
xor ( n73804 , n73456 , n73462 );
xor ( n73805 , n73804 , n73793 );
xor ( n73806 , n73456 , n73462 );
and ( n73807 , n73806 , n73793 );
and ( n73808 , n73456 , n73462 );
or ( n73809 , n73807 , n73808 );
xor ( n73810 , n73799 , n73468 );
xor ( n73811 , n73810 , n73474 );
xor ( n73812 , n73799 , n73468 );
and ( n73813 , n73812 , n73474 );
and ( n73814 , n73799 , n73468 );
or ( n73815 , n73813 , n73814 );
xor ( n73816 , n73627 , n73637 );
and ( n73817 , n73816 , n73648 );
and ( n73818 , n73627 , n73637 );
or ( n73819 , n73817 , n73818 );
xor ( n73820 , n73805 , n73811 );
xor ( n73821 , n73820 , n73484 );
xor ( n73822 , n73805 , n73811 );
and ( n73823 , n73822 , n73484 );
and ( n73824 , n73805 , n73811 );
or ( n73825 , n73823 , n73824 );
xor ( n73826 , n73747 , n73757 );
and ( n73827 , n73826 , n73769 );
and ( n73828 , n73747 , n73757 );
or ( n73829 , n73827 , n73828 );
xor ( n73830 , n73594 , n73604 );
and ( n73831 , n73830 , n73616 );
and ( n73832 , n73594 , n73604 );
or ( n73833 , n73831 , n73832 );
xor ( n73834 , n73690 , n73700 );
and ( n73835 , n73834 , n73710 );
and ( n73836 , n73690 , n73700 );
or ( n73837 , n73835 , n73836 );
xor ( n73838 , n73717 , n73727 );
and ( n73839 , n73838 , n73201 );
and ( n73840 , n73717 , n73727 );
or ( n73841 , n73839 , n73840 );
xor ( n73842 , n73236 , n73665 );
and ( n73843 , n73842 , n73676 );
and ( n73844 , n73236 , n73665 );
or ( n73845 , n73843 , n73844 );
xor ( n73846 , n73552 , n73580 );
and ( n73847 , n73846 , n73478 );
and ( n73848 , n73552 , n73580 );
or ( n73849 , n73847 , n73848 );
xor ( n73850 , n73494 , n73498 );
and ( n73851 , n73850 , n73770 );
and ( n73852 , n73494 , n73498 );
or ( n73853 , n73851 , n73852 );
not ( n73854 , n52722 );
not ( n73855 , n49420 );
or ( n73856 , n73854 , n73855 );
nand ( n73857 , n73856 , n58982 );
not ( n73858 , n73744 );
not ( n73859 , n65130 );
or ( n73860 , n73858 , n73859 );
not ( n73861 , n66140 );
not ( n73862 , n52076 );
or ( n73863 , n73861 , n73862 );
nand ( n73864 , n67084 , n41132 );
nand ( n73865 , n73863 , n73864 );
nand ( n73866 , n60427 , n73865 );
nand ( n73867 , n73860 , n73866 );
xor ( n73868 , n73857 , n73867 );
not ( n73869 , n73526 );
or ( n73870 , n69728 , n73869 );
and ( n73871 , n64452 , n61537 );
not ( n73872 , n64452 );
and ( n73873 , n73872 , n61540 );
nor ( n73874 , n73871 , n73873 );
or ( n73875 , n69731 , n73874 );
nand ( n73876 , n73870 , n73875 );
xor ( n73877 , n73868 , n73876 );
xor ( n73878 , n73857 , n73867 );
and ( n73879 , n73878 , n73876 );
and ( n73880 , n73857 , n73867 );
or ( n73881 , n73879 , n73880 );
not ( n73882 , n73549 );
not ( n73883 , n67061 );
or ( n73884 , n73882 , n73883 );
not ( n73885 , n62451 );
not ( n73886 , n49837 );
and ( n73887 , n73885 , n73886 );
and ( n73888 , n64170 , n49210 );
nor ( n73889 , n73887 , n73888 );
not ( n73890 , n73889 );
nand ( n73891 , n73890 , n67068 );
nand ( n73892 , n73884 , n73891 );
not ( n73893 , n73536 );
not ( n73894 , n66569 );
or ( n73895 , n73893 , n73894 );
not ( n73896 , n67441 );
not ( n73897 , n65094 );
or ( n73898 , n73896 , n73897 );
nand ( n73899 , n67072 , n49190 );
nand ( n73900 , n73898 , n73899 );
nand ( n73901 , n65092 , n73900 );
nand ( n73902 , n73895 , n73901 );
xor ( n73903 , n73892 , n73902 );
and ( n73904 , n72846 , n41532 );
xor ( n73905 , n73903 , n73904 );
xor ( n73906 , n73892 , n73902 );
and ( n73907 , n73906 , n73904 );
and ( n73908 , n73892 , n73902 );
or ( n73909 , n73907 , n73908 );
not ( n73910 , n53956 );
not ( n73911 , n73633 );
or ( n73912 , n73910 , n73911 );
not ( n73913 , n55089 );
not ( n73914 , n72606 );
or ( n73915 , n73913 , n73914 );
nand ( n73916 , n40514 , n55090 );
nand ( n73917 , n73915 , n73916 );
nand ( n73918 , n73917 , n54364 );
nand ( n73919 , n73912 , n73918 );
not ( n73920 , n54327 );
not ( n73921 , n70627 );
not ( n73922 , n59694 );
or ( n73923 , n73921 , n73922 );
nand ( n73924 , n71829 , n54322 );
nand ( n73925 , n73923 , n73924 );
not ( n73926 , n73925 );
or ( n73927 , n73920 , n73926 );
nand ( n73928 , n73646 , n54316 );
nand ( n73929 , n73927 , n73928 );
xor ( n73930 , n73919 , n73929 );
xor ( n73931 , n73930 , n73746 );
not ( n73932 , n59575 );
not ( n73933 , n72464 );
not ( n73934 , n51574 );
or ( n73935 , n73933 , n73934 );
nand ( n73936 , n40677 , n70920 );
nand ( n73937 , n73935 , n73936 );
not ( n73938 , n73937 );
or ( n73939 , n73932 , n73938 );
nand ( n73940 , n73563 , n70487 );
nand ( n73941 , n73939 , n73940 );
not ( n73942 , n53182 );
not ( n73943 , n73625 );
or ( n73944 , n73942 , n73943 );
not ( n73945 , n54283 );
not ( n73946 , n39963 );
or ( n73947 , n73945 , n73946 );
nand ( n73948 , n59654 , n53947 );
nand ( n73949 , n73947 , n73948 );
nand ( n73950 , n73949 , n53571 );
nand ( n73951 , n73944 , n73950 );
xor ( n73952 , n73941 , n73951 );
not ( n73953 , n71466 );
not ( n73954 , n62496 );
not ( n73955 , n51602 );
or ( n73956 , n73954 , n73955 );
nand ( n73957 , n51601 , n62497 );
nand ( n73958 , n73956 , n73957 );
not ( n73959 , n73958 );
or ( n73960 , n73953 , n73959 );
nand ( n73961 , n73575 , n72106 );
nand ( n73962 , n73960 , n73961 );
xor ( n73963 , n73952 , n73962 );
xor ( n73964 , n73931 , n73963 );
xor ( n73965 , n73964 , n73845 );
xor ( n73966 , n73931 , n73963 );
and ( n73967 , n73966 , n73845 );
and ( n73968 , n73931 , n73963 );
or ( n73969 , n73967 , n73968 );
xor ( n73970 , n73833 , n73837 );
xor ( n73971 , n73970 , n73841 );
xor ( n73972 , n73833 , n73837 );
and ( n73973 , n73972 , n73841 );
and ( n73974 , n73833 , n73837 );
or ( n73975 , n73973 , n73974 );
not ( n73976 , n70604 );
not ( n73977 , n73307 );
not ( n73978 , n73977 );
not ( n73979 , n66798 );
or ( n73980 , n73978 , n73979 );
nand ( n73981 , n40592 , n67890 );
nand ( n73982 , n73980 , n73981 );
not ( n73983 , n73982 );
or ( n73984 , n73976 , n73983 );
nand ( n73985 , n73602 , n60482 );
nand ( n73986 , n73984 , n73985 );
not ( n73987 , n53197 );
not ( n73988 , n73612 );
or ( n73989 , n73987 , n73988 );
not ( n73990 , n52490 );
not ( n73991 , n59414 );
or ( n73992 , n73990 , n73991 );
not ( n73993 , n39894 );
nand ( n73994 , n73993 , n52130 );
nand ( n73995 , n73992 , n73994 );
nand ( n73996 , n73995 , n72220 );
nand ( n73997 , n73989 , n73996 );
xor ( n73998 , n73986 , n73997 );
not ( n73999 , n56639 );
not ( n74000 , n59345 );
not ( n74001 , n71163 );
or ( n74002 , n74000 , n74001 );
nand ( n74003 , n42654 , n65743 );
nand ( n74004 , n74002 , n74003 );
not ( n74005 , n74004 );
or ( n74006 , n73999 , n74005 );
not ( n74007 , n73688 );
nand ( n74008 , n74007 , n59950 );
nand ( n74009 , n74006 , n74008 );
xor ( n74010 , n73998 , n74009 );
not ( n74011 , n60927 );
not ( n74012 , n66234 );
not ( n74013 , n42399 );
or ( n74014 , n74012 , n74013 );
nand ( n74015 , n65546 , n60289 );
nand ( n74016 , n74014 , n74015 );
not ( n74017 , n74016 );
or ( n74018 , n74011 , n74017 );
nand ( n74019 , n73662 , n58168 );
nand ( n74020 , n74018 , n74019 );
xor ( n74021 , n73556 , n74020 );
not ( n74022 , n51533 );
not ( n74023 , n53931 );
not ( n74024 , n58482 );
or ( n74025 , n74023 , n74024 );
nand ( n74026 , n60386 , n71445 );
nand ( n74027 , n74025 , n74026 );
not ( n74028 , n74027 );
or ( n74029 , n74022 , n74028 );
nand ( n74030 , n73674 , n56355 );
nand ( n74031 , n74029 , n74030 );
xor ( n74032 , n74021 , n74031 );
xor ( n74033 , n74010 , n74032 );
not ( n74034 , n62664 );
not ( n74035 , n73696 );
or ( n74036 , n74034 , n74035 );
not ( n74037 , n61951 );
not ( n74038 , n66500 );
or ( n74039 , n74037 , n74038 );
nand ( n74040 , n39253 , n61952 );
nand ( n74041 , n74039 , n74040 );
nand ( n74042 , n74041 , n62654 );
nand ( n74043 , n74036 , n74042 );
not ( n74044 , n63708 );
not ( n74045 , n73707 );
or ( n74046 , n74044 , n74045 );
not ( n74047 , n50306 );
not ( n74048 , n68652 );
or ( n74049 , n74047 , n74048 );
nand ( n74050 , n67482 , n66705 );
nand ( n74051 , n74049 , n74050 );
nand ( n74052 , n74051 , n52757 );
nand ( n74053 , n74046 , n74052 );
xor ( n74054 , n74043 , n74053 );
not ( n74055 , n52151 );
not ( n74056 , n73725 );
or ( n74057 , n74055 , n74056 );
not ( n74058 , n65773 );
not ( n74059 , n39575 );
not ( n74060 , n74059 );
or ( n74061 , n74058 , n74060 );
nand ( n74062 , n39575 , n71042 );
nand ( n74063 , n74061 , n74062 );
nand ( n74064 , n74063 , n50922 );
nand ( n74065 , n74057 , n74064 );
xor ( n74066 , n74054 , n74065 );
xor ( n74067 , n74033 , n74066 );
xor ( n74068 , n74010 , n74032 );
and ( n74069 , n74068 , n74066 );
and ( n74070 , n74010 , n74032 );
or ( n74071 , n74069 , n74070 );
xor ( n74072 , n73905 , n73877 );
xor ( n74073 , n74072 , n73584 );
xor ( n74074 , n73849 , n74073 );
xor ( n74075 , n74074 , n73655 );
xor ( n74076 , n73849 , n74073 );
and ( n74077 , n74076 , n73655 );
and ( n74078 , n73849 , n74073 );
or ( n74079 , n74077 , n74078 );
xor ( n74080 , n73819 , n73829 );
not ( n74081 , n70193 );
not ( n74082 , n73755 );
or ( n74083 , n74081 , n74082 );
and ( n74084 , n55124 , n40148 );
not ( n74085 , n55124 );
and ( n74086 , n74085 , n69409 );
or ( n74087 , n74084 , n74086 );
nand ( n74088 , n74087 , n70183 );
nand ( n74089 , n74083 , n74088 );
not ( n74090 , n59984 );
not ( n74091 , n72288 );
not ( n74092 , n55242 );
or ( n74093 , n74091 , n74092 );
not ( n74094 , n69695 );
nand ( n74095 , n53660 , n74094 );
nand ( n74096 , n74093 , n74095 );
not ( n74097 , n74096 );
or ( n74098 , n74090 , n74097 );
nand ( n74099 , n71099 , n73767 );
nand ( n74100 , n74098 , n74099 );
xor ( n74101 , n74089 , n74100 );
not ( n74102 , n72185 );
not ( n74103 , n56786 );
not ( n74104 , n54415 );
or ( n74105 , n74103 , n74104 );
nand ( n74106 , n59612 , n71362 );
nand ( n74107 , n74105 , n74106 );
not ( n74108 , n74107 );
or ( n74109 , n74102 , n74108 );
nand ( n74110 , n73592 , n56777 );
nand ( n74111 , n74109 , n74110 );
xor ( n74112 , n74101 , n74111 );
xor ( n74113 , n74080 , n74112 );
xor ( n74114 , n73853 , n74113 );
xor ( n74115 , n74114 , n73734 );
xor ( n74116 , n73853 , n74113 );
and ( n74117 , n74116 , n73734 );
and ( n74118 , n73853 , n74113 );
or ( n74119 , n74117 , n74118 );
xor ( n74120 , n73971 , n73682 );
xor ( n74121 , n74120 , n73965 );
xor ( n74122 , n73971 , n73682 );
and ( n74123 , n74122 , n73965 );
and ( n74124 , n73971 , n73682 );
or ( n74125 , n74123 , n74124 );
xor ( n74126 , n74067 , n73777 );
xor ( n74127 , n74126 , n74075 );
xor ( n74128 , n74067 , n73777 );
and ( n74129 , n74128 , n74075 );
and ( n74130 , n74067 , n73777 );
or ( n74131 , n74129 , n74130 );
xor ( n74132 , n73785 , n74115 );
xor ( n74133 , n74132 , n73791 );
xor ( n74134 , n73785 , n74115 );
and ( n74135 , n74134 , n73791 );
and ( n74136 , n73785 , n74115 );
or ( n74137 , n74135 , n74136 );
xor ( n74138 , n74121 , n73797 );
xor ( n74139 , n74138 , n74127 );
xor ( n74140 , n74121 , n73797 );
and ( n74141 , n74140 , n74127 );
and ( n74142 , n74121 , n73797 );
or ( n74143 , n74141 , n74142 );
xor ( n74144 , n74133 , n73803 );
xor ( n74145 , n74144 , n73809 );
xor ( n74146 , n74133 , n73803 );
and ( n74147 , n74146 , n73809 );
and ( n74148 , n74133 , n73803 );
or ( n74149 , n74147 , n74148 );
xor ( n74150 , n73941 , n73951 );
and ( n74151 , n74150 , n73962 );
and ( n74152 , n73941 , n73951 );
or ( n74153 , n74151 , n74152 );
xor ( n74154 , n74139 , n74145 );
xor ( n74155 , n74154 , n73815 );
xor ( n74156 , n74139 , n74145 );
and ( n74157 , n74156 , n73815 );
and ( n74158 , n74139 , n74145 );
or ( n74159 , n74157 , n74158 );
xor ( n74160 , n73919 , n73929 );
and ( n74161 , n74160 , n73746 );
and ( n74162 , n73919 , n73929 );
or ( n74163 , n74161 , n74162 );
xor ( n74164 , n74089 , n74100 );
and ( n74165 , n74164 , n74111 );
and ( n74166 , n74089 , n74100 );
or ( n74167 , n74165 , n74166 );
xor ( n74168 , n73986 , n73997 );
and ( n74169 , n74168 , n74009 );
and ( n74170 , n73986 , n73997 );
or ( n74171 , n74169 , n74170 );
xor ( n74172 , n74043 , n74053 );
and ( n74173 , n74172 , n74065 );
and ( n74174 , n74043 , n74053 );
or ( n74175 , n74173 , n74174 );
xor ( n74176 , n73556 , n74020 );
and ( n74177 , n74176 , n74031 );
and ( n74178 , n73556 , n74020 );
or ( n74179 , n74177 , n74178 );
xor ( n74180 , n73905 , n73877 );
and ( n74181 , n74180 , n73584 );
and ( n74182 , n73905 , n73877 );
or ( n74183 , n74181 , n74182 );
xor ( n74184 , n73819 , n73829 );
and ( n74185 , n74184 , n74112 );
and ( n74186 , n73819 , n73829 );
or ( n74187 , n74185 , n74186 );
or ( n74188 , n64684 , n73889 );
and ( n74189 , n62452 , n56239 );
and ( n74190 , n67555 , n62861 );
nor ( n74191 , n74189 , n74190 );
or ( n74192 , n74191 , n64166 );
nand ( n74193 , n74188 , n74192 );
and ( n74194 , n66155 , n65969 );
xor ( n74195 , n74193 , n74194 );
not ( n74196 , n73900 );
not ( n74197 , n65795 );
or ( n74198 , n74196 , n74197 );
and ( n74199 , n41288 , n64443 );
not ( n74200 , n41288 );
and ( n74201 , n74200 , n63922 );
or ( n74202 , n74199 , n74201 );
nand ( n74203 , n74202 , n65092 );
nand ( n74204 , n74198 , n74203 );
xor ( n74205 , n74195 , n74204 );
xor ( n74206 , n74193 , n74194 );
and ( n74207 , n74206 , n74204 );
and ( n74208 , n74193 , n74194 );
or ( n74209 , n74207 , n74208 );
not ( n74210 , n73865 );
not ( n74211 , n66136 );
or ( n74212 , n74210 , n74211 );
not ( n74213 , n70506 );
not ( n74214 , n50654 );
or ( n74215 , n74213 , n74214 );
nand ( n74216 , n71361 , n73190 );
nand ( n74217 , n74215 , n74216 );
nand ( n74218 , n74217 , n70930 );
nand ( n74219 , n74212 , n74218 );
not ( n74220 , n60542 );
and ( n74221 , n51929 , n59340 );
not ( n74222 , n51929 );
and ( n74223 , n74222 , n72464 );
or ( n74224 , n74221 , n74223 );
not ( n74225 , n74224 );
or ( n74226 , n74220 , n74225 );
nand ( n74227 , n73937 , n72131 );
nand ( n74228 , n74226 , n74227 );
xor ( n74229 , n74219 , n74228 );
not ( n74230 , n54364 );
not ( n74231 , n53596 );
not ( n74232 , n63180 );
or ( n74233 , n74231 , n74232 );
nand ( n74234 , n56455 , n71756 );
nand ( n74235 , n74233 , n74234 );
not ( n74236 , n74235 );
or ( n74237 , n74230 , n74236 );
nand ( n74238 , n73917 , n68603 );
nand ( n74239 , n74237 , n74238 );
xor ( n74240 , n74229 , n74239 );
xor ( n74241 , n74219 , n74228 );
and ( n74242 , n74241 , n74239 );
and ( n74243 , n74219 , n74228 );
or ( n74244 , n74242 , n74243 );
xor ( n74245 , n74175 , n74171 );
not ( n74246 , n54316 );
not ( n74247 , n73925 );
or ( n74248 , n74246 , n74247 );
not ( n74249 , n54725 );
not ( n74250 , n70661 );
or ( n74251 , n74249 , n74250 );
nand ( n74252 , n68980 , n54302 );
nand ( n74253 , n74251 , n74252 );
nand ( n74254 , n74253 , n54327 );
nand ( n74255 , n74248 , n74254 );
not ( n74256 , n55144 );
not ( n74257 , n74087 );
or ( n74258 , n74256 , n74257 );
not ( n74259 , n55582 );
not ( n74260 , n68073 );
or ( n74261 , n74259 , n74260 );
nand ( n74262 , n55642 , n55119 );
nand ( n74263 , n74261 , n74262 );
nand ( n74264 , n74263 , n70183 );
nand ( n74265 , n74258 , n74264 );
xor ( n74266 , n74255 , n74265 );
not ( n74267 , n73874 );
not ( n74268 , n74267 );
not ( n74269 , n64111 );
or ( n74270 , n74268 , n74269 );
not ( n74271 , n50021 );
not ( n74272 , n61537 );
or ( n74273 , n74271 , n74272 );
not ( n74274 , n51891 );
nand ( n74275 , n74274 , n61540 );
nand ( n74276 , n74273 , n74275 );
nand ( n74277 , n61558 , n74276 );
nand ( n74278 , n74270 , n74277 );
not ( n74279 , n74278 );
xor ( n74280 , n74266 , n74279 );
xor ( n74281 , n74245 , n74280 );
xor ( n74282 , n74175 , n74171 );
and ( n74283 , n74282 , n74280 );
and ( n74284 , n74175 , n74171 );
or ( n74285 , n74283 , n74284 );
not ( n74286 , n72106 );
not ( n74287 , n73958 );
or ( n74288 , n74286 , n74287 );
not ( n74289 , n66652 );
not ( n74290 , n74289 );
not ( n74291 , n40527 );
or ( n74292 , n74290 , n74291 );
nand ( n74293 , n72945 , n66652 );
nand ( n74294 , n74292 , n74293 );
nand ( n74295 , n74294 , n71466 );
nand ( n74296 , n74288 , n74295 );
not ( n74297 , n52469 );
not ( n74298 , n54283 );
not ( n74299 , n39846 );
or ( n74300 , n74298 , n74299 );
nand ( n74301 , n68145 , n52837 );
nand ( n74302 , n74300 , n74301 );
not ( n74303 , n74302 );
or ( n74304 , n74297 , n74303 );
nand ( n74305 , n73949 , n52854 );
nand ( n74306 , n74304 , n74305 );
xor ( n74307 , n74296 , n74306 );
not ( n74308 , n62085 );
not ( n74309 , n74016 );
or ( n74310 , n74308 , n74309 );
not ( n74311 , n60289 );
not ( n74312 , n71525 );
or ( n74313 , n74311 , n74312 );
nand ( n74314 , n66301 , n62077 );
nand ( n74315 , n74313 , n74314 );
nand ( n74316 , n74315 , n52191 );
nand ( n74317 , n74310 , n74316 );
xor ( n74318 , n74307 , n74317 );
not ( n74319 , n62654 );
not ( n74320 , n61951 );
not ( n74321 , n66052 );
or ( n74322 , n74320 , n74321 );
nand ( n74323 , n61907 , n61952 );
nand ( n74324 , n74322 , n74323 );
not ( n74325 , n74324 );
or ( n74326 , n74319 , n74325 );
nand ( n74327 , n74041 , n52058 );
nand ( n74328 , n74326 , n74327 );
not ( n74329 , n72220 );
not ( n74330 , n52114 );
not ( n74331 , n67040 );
or ( n74332 , n74330 , n74331 );
nand ( n74333 , n59913 , n52130 );
nand ( n74334 , n74332 , n74333 );
not ( n74335 , n74334 );
or ( n74336 , n74329 , n74335 );
nand ( n74337 , n53197 , n73995 );
nand ( n74338 , n74336 , n74337 );
xor ( n74339 , n74328 , n74338 );
xor ( n74340 , n74339 , n74205 );
xor ( n74341 , n74318 , n74340 );
not ( n74342 , n52749 );
not ( n74343 , n74051 );
or ( n74344 , n74342 , n74343 );
not ( n74345 , n50306 );
not ( n74346 , n39333 );
or ( n74347 , n74345 , n74346 );
nand ( n74348 , n62963 , n66705 );
nand ( n74349 , n74347 , n74348 );
nand ( n74350 , n74349 , n52757 );
nand ( n74351 , n74344 , n74350 );
not ( n74352 , n50922 );
not ( n74353 , n51465 );
not ( n74354 , n69072 );
or ( n74355 , n74353 , n74354 );
nand ( n74356 , n39056 , n71042 );
nand ( n74357 , n74355 , n74356 );
not ( n74358 , n74357 );
or ( n74359 , n74352 , n74358 );
nand ( n74360 , n74063 , n52151 );
nand ( n74361 , n74359 , n74360 );
xor ( n74362 , n74351 , n74361 );
not ( n74363 , n59950 );
not ( n74364 , n74004 );
or ( n74365 , n74363 , n74364 );
nand ( n74366 , n56639 , n59345 );
nand ( n74367 , n74365 , n74366 );
xor ( n74368 , n74362 , n74367 );
xor ( n74369 , n74341 , n74368 );
xor ( n74370 , n74318 , n74340 );
and ( n74371 , n74370 , n74368 );
and ( n74372 , n74318 , n74340 );
or ( n74373 , n74371 , n74372 );
not ( n74374 , n72198 );
not ( n74375 , n74027 );
or ( n74376 , n74374 , n74375 );
not ( n74377 , n53931 );
not ( n74378 , n68206 );
or ( n74379 , n74377 , n74378 );
nand ( n74380 , n39714 , n71053 );
nand ( n74381 , n74379 , n74380 );
nand ( n74382 , n74381 , n51533 );
nand ( n74383 , n74376 , n74382 );
xor ( n74384 , n73881 , n74383 );
xor ( n74385 , n74384 , n73909 );
xor ( n74386 , n74385 , n74183 );
xor ( n74387 , n74386 , n74187 );
xor ( n74388 , n74385 , n74183 );
and ( n74389 , n74388 , n74187 );
and ( n74390 , n74385 , n74183 );
or ( n74391 , n74389 , n74390 );
xor ( n74392 , n73975 , n73969 );
xor ( n74393 , n74153 , n74163 );
xor ( n74394 , n74393 , n74167 );
xor ( n74395 , n74392 , n74394 );
xor ( n74396 , n73975 , n73969 );
and ( n74397 , n74396 , n74394 );
and ( n74398 , n73975 , n73969 );
or ( n74399 , n74397 , n74398 );
xor ( n74400 , n74071 , n74281 );
not ( n74401 , n59984 );
not ( n74402 , n69237 );
not ( n74403 , n74402 );
not ( n74404 , n54811 );
or ( n74405 , n74403 , n74404 );
nand ( n74406 , n59195 , n74094 );
nand ( n74407 , n74405 , n74406 );
not ( n74408 , n74407 );
or ( n74409 , n74401 , n74408 );
nand ( n74410 , n74096 , n67862 );
nand ( n74411 , n74409 , n74410 );
not ( n74412 , n56777 );
not ( n74413 , n74107 );
or ( n74414 , n74412 , n74413 );
not ( n74415 , n56786 );
not ( n74416 , n56476 );
or ( n74417 , n74415 , n74416 );
nand ( n74418 , n54646 , n71362 );
nand ( n74419 , n74417 , n74418 );
nand ( n74420 , n74419 , n60472 );
nand ( n74421 , n74414 , n74420 );
xor ( n74422 , n74411 , n74421 );
not ( n74423 , n72961 );
not ( n74424 , n73982 );
or ( n74425 , n74423 , n74424 );
not ( n74426 , n73977 );
not ( n74427 , n52432 );
or ( n74428 , n74426 , n74427 );
nand ( n74429 , n68049 , n67890 );
nand ( n74430 , n74428 , n74429 );
nand ( n74431 , n74430 , n72710 );
nand ( n74432 , n74425 , n74431 );
xor ( n74433 , n74422 , n74432 );
xor ( n74434 , n74179 , n74433 );
xor ( n74435 , n74434 , n74240 );
xor ( n74436 , n74400 , n74435 );
xor ( n74437 , n74071 , n74281 );
and ( n74438 , n74437 , n74435 );
and ( n74439 , n74071 , n74281 );
or ( n74440 , n74438 , n74439 );
xor ( n74441 , n74369 , n74079 );
xor ( n74442 , n74441 , n74387 );
xor ( n74443 , n74369 , n74079 );
and ( n74444 , n74443 , n74387 );
and ( n74445 , n74369 , n74079 );
or ( n74446 , n74444 , n74445 );
xor ( n74447 , n74395 , n74125 );
xor ( n74448 , n74447 , n74119 );
xor ( n74449 , n74395 , n74125 );
and ( n74450 , n74449 , n74119 );
and ( n74451 , n74395 , n74125 );
or ( n74452 , n74450 , n74451 );
xor ( n74453 , n74436 , n74131 );
xor ( n74454 , n74453 , n74442 );
xor ( n74455 , n74436 , n74131 );
and ( n74456 , n74455 , n74442 );
and ( n74457 , n74436 , n74131 );
or ( n74458 , n74456 , n74457 );
xor ( n74459 , n74448 , n74137 );
xor ( n74460 , n74459 , n74143 );
xor ( n74461 , n74448 , n74137 );
and ( n74462 , n74461 , n74143 );
and ( n74463 , n74448 , n74137 );
or ( n74464 , n74462 , n74463 );
xor ( n74465 , n74454 , n74460 );
xor ( n74466 , n74465 , n74149 );
xor ( n74467 , n74454 , n74460 );
and ( n74468 , n74467 , n74149 );
and ( n74469 , n74454 , n74460 );
or ( n74470 , n74468 , n74469 );
xor ( n74471 , n74255 , n74265 );
and ( n74472 , n74471 , n74279 );
and ( n74473 , n74255 , n74265 );
or ( n74474 , n74472 , n74473 );
xor ( n74475 , n74411 , n74421 );
and ( n74476 , n74475 , n74432 );
and ( n74477 , n74411 , n74421 );
or ( n74478 , n74476 , n74477 );
xor ( n74479 , n74296 , n74306 );
and ( n74480 , n74479 , n74317 );
and ( n74481 , n74296 , n74306 );
or ( n74482 , n74480 , n74481 );
xor ( n74483 , n74351 , n74361 );
and ( n74484 , n74483 , n74367 );
and ( n74485 , n74351 , n74361 );
or ( n74486 , n74484 , n74485 );
xor ( n74487 , n73881 , n74383 );
and ( n74488 , n74487 , n73909 );
and ( n74489 , n73881 , n74383 );
or ( n74490 , n74488 , n74489 );
xor ( n74491 , n74328 , n74338 );
and ( n74492 , n74491 , n74205 );
and ( n74493 , n74328 , n74338 );
or ( n74494 , n74492 , n74493 );
xor ( n74495 , n74153 , n74163 );
and ( n74496 , n74495 , n74167 );
and ( n74497 , n74153 , n74163 );
or ( n74498 , n74496 , n74497 );
xor ( n74499 , n74179 , n74433 );
and ( n74500 , n74499 , n74240 );
and ( n74501 , n74179 , n74433 );
or ( n74502 , n74500 , n74501 );
not ( n74503 , n68961 );
not ( n74504 , n73409 );
or ( n74505 , n74503 , n74504 );
nand ( n74506 , n74505 , n59345 );
not ( n74507 , n74276 );
not ( n74508 , n72810 );
or ( n74509 , n74507 , n74508 );
not ( n74510 , n71307 );
not ( n74511 , n41132 );
or ( n74512 , n74510 , n74511 );
not ( n74513 , n70889 );
nand ( n74514 , n74513 , n71309 );
nand ( n74515 , n74512 , n74514 );
nand ( n74516 , n61558 , n74515 );
nand ( n74517 , n74509 , n74516 );
xor ( n74518 , n74506 , n74517 );
or ( n74519 , n64164 , n74191 );
and ( n74520 , n69704 , n71691 );
and ( n74521 , n64170 , n64451 );
nor ( n74522 , n74520 , n74521 );
or ( n74523 , n64166 , n74522 );
nand ( n74524 , n74519 , n74523 );
xor ( n74525 , n74518 , n74524 );
xor ( n74526 , n74506 , n74517 );
and ( n74527 , n74526 , n74524 );
and ( n74528 , n74506 , n74517 );
or ( n74529 , n74527 , n74528 );
not ( n74530 , n74202 );
not ( n74531 , n65795 );
or ( n74532 , n74530 , n74531 );
and ( n74533 , n70908 , n64443 );
not ( n74534 , n70908 );
and ( n74535 , n74534 , n66575 );
or ( n74536 , n74533 , n74535 );
nand ( n74537 , n70964 , n74536 );
nand ( n74538 , n74532 , n74537 );
and ( n74539 , n71971 , n67441 );
xor ( n74540 , n74538 , n74539 );
not ( n74541 , n70930 );
not ( n74542 , n70506 );
not ( n74543 , n51574 );
or ( n74544 , n74542 , n74543 );
nand ( n74545 , n68598 , n67084 );
nand ( n74546 , n74544 , n74545 );
not ( n74547 , n74546 );
or ( n74548 , n74541 , n74547 );
nand ( n74549 , n70500 , n74217 );
nand ( n74550 , n74548 , n74549 );
xor ( n74551 , n74540 , n74550 );
xor ( n74552 , n74538 , n74539 );
and ( n74553 , n74552 , n74550 );
and ( n74554 , n74538 , n74539 );
or ( n74555 , n74553 , n74554 );
not ( n74556 , n60472 );
not ( n74557 , n72589 );
not ( n74558 , n40225 );
or ( n74559 , n74557 , n74558 );
nand ( n74560 , n54433 , n56785 );
nand ( n74561 , n74559 , n74560 );
not ( n74562 , n74561 );
or ( n74563 , n74556 , n74562 );
nand ( n74564 , n56777 , n74419 );
nand ( n74565 , n74563 , n74564 );
not ( n74566 , n70604 );
not ( n74567 , n63656 );
not ( n74568 , n73977 );
or ( n74569 , n74567 , n74568 );
nand ( n74570 , n71770 , n67890 );
nand ( n74571 , n74569 , n74570 );
not ( n74572 , n74571 );
or ( n74573 , n74566 , n74572 );
nand ( n74574 , n74430 , n72182 );
nand ( n74575 , n74573 , n74574 );
xor ( n74576 , n74565 , n74575 );
not ( n74577 , n61465 );
not ( n74578 , n62496 );
not ( n74579 , n66798 );
or ( n74580 , n74578 , n74579 );
not ( n74581 , n66798 );
nand ( n74582 , n65183 , n74581 );
nand ( n74583 , n74580 , n74582 );
not ( n74584 , n74583 );
or ( n74585 , n74577 , n74584 );
nand ( n74586 , n74294 , n65646 );
nand ( n74587 , n74585 , n74586 );
xor ( n74588 , n74576 , n74587 );
not ( n74589 , n68603 );
not ( n74590 , n74235 );
or ( n74591 , n74589 , n74590 );
not ( n74592 , n53596 );
not ( n74593 , n68611 );
or ( n74594 , n74592 , n74593 );
nand ( n74595 , n39964 , n70991 );
nand ( n74596 , n74594 , n74595 );
nand ( n74597 , n74596 , n53620 );
nand ( n74598 , n74591 , n74597 );
not ( n74599 , n60542 );
not ( n74600 , n59341 );
not ( n74601 , n70278 );
or ( n74602 , n74600 , n74601 );
nand ( n74603 , n69442 , n59340 );
nand ( n74604 , n74602 , n74603 );
not ( n74605 , n74604 );
or ( n74606 , n74599 , n74605 );
nand ( n74607 , n74224 , n70487 );
nand ( n74608 , n74606 , n74607 );
xor ( n74609 , n74598 , n74608 );
not ( n74610 , n54327 );
not ( n74611 , n54725 );
not ( n74612 , n70290 );
or ( n74613 , n74611 , n74612 );
nand ( n74614 , n72607 , n54468 );
nand ( n74615 , n74613 , n74614 );
not ( n74616 , n74615 );
or ( n74617 , n74610 , n74616 );
nand ( n74618 , n74253 , n54316 );
nand ( n74619 , n74617 , n74618 );
xor ( n74620 , n74609 , n74619 );
xor ( n74621 , n74588 , n74620 );
xor ( n74622 , n74621 , n74490 );
xor ( n74623 , n74588 , n74620 );
and ( n74624 , n74623 , n74490 );
and ( n74625 , n74588 , n74620 );
or ( n74626 , n74624 , n74625 );
not ( n74627 , n53571 );
not ( n74628 , n52841 );
not ( n74629 , n59414 );
or ( n74630 , n74628 , n74629 );
nand ( n74631 , n65708 , n52837 );
nand ( n74632 , n74630 , n74631 );
not ( n74633 , n74632 );
or ( n74634 , n74627 , n74633 );
nand ( n74635 , n74302 , n53182 );
nand ( n74636 , n74634 , n74635 );
not ( n74637 , n60927 );
not ( n74638 , n62077 );
not ( n74639 , n42654 );
not ( n74640 , n74639 );
or ( n74641 , n74638 , n74640 );
nand ( n74642 , n71875 , n60289 );
nand ( n74643 , n74641 , n74642 );
not ( n74644 , n74643 );
or ( n74645 , n74637 , n74644 );
nand ( n74646 , n74315 , n58168 );
nand ( n74647 , n74645 , n74646 );
xor ( n74648 , n74636 , n74647 );
not ( n74649 , n52757 );
not ( n74650 , n50306 );
not ( n74651 , n71176 );
or ( n74652 , n74650 , n74651 );
nand ( n74653 , n69530 , n64191 );
nand ( n74654 , n74652 , n74653 );
not ( n74655 , n74654 );
or ( n74656 , n74649 , n74655 );
nand ( n74657 , n74349 , n63708 );
nand ( n74658 , n74656 , n74657 );
xor ( n74659 , n74648 , n74658 );
xor ( n74660 , n74486 , n74659 );
not ( n74661 , n62654 );
not ( n74662 , n61951 );
not ( n74663 , n71139 );
or ( n74664 , n74662 , n74663 );
nand ( n74665 , n42400 , n66690 );
nand ( n74666 , n74664 , n74665 );
not ( n74667 , n74666 );
or ( n74668 , n74661 , n74667 );
nand ( n74669 , n74324 , n66696 );
nand ( n74670 , n74668 , n74669 );
not ( n74671 , n72220 );
not ( n74672 , n52490 );
not ( n74673 , n66546 );
not ( n74674 , n74673 );
or ( n74675 , n74672 , n74674 );
nand ( n74676 , n58485 , n52130 );
nand ( n74677 , n74675 , n74676 );
not ( n74678 , n74677 );
or ( n74679 , n74671 , n74678 );
nand ( n74680 , n74334 , n53197 );
nand ( n74681 , n74679 , n74680 );
xor ( n74682 , n74670 , n74681 );
xor ( n74683 , n74682 , n74525 );
xor ( n74684 , n74660 , n74683 );
xor ( n74685 , n74486 , n74659 );
and ( n74686 , n74685 , n74683 );
and ( n74687 , n74486 , n74659 );
or ( n74688 , n74686 , n74687 );
not ( n74689 , n52151 );
not ( n74690 , n74357 );
or ( n74691 , n74689 , n74690 );
not ( n74692 , n57187 );
not ( n74693 , n62394 );
or ( n74694 , n74692 , n74693 );
nand ( n74695 , n67482 , n50946 );
nand ( n74696 , n74694 , n74695 );
nand ( n74697 , n74696 , n50922 );
nand ( n74698 , n74691 , n74697 );
xor ( n74699 , n74698 , n74209 );
not ( n74700 , n51533 );
not ( n74701 , n53931 );
not ( n74702 , n65532 );
or ( n74703 , n74701 , n74702 );
nand ( n74704 , n39575 , n71053 );
nand ( n74705 , n74703 , n74704 );
not ( n74706 , n74705 );
or ( n74707 , n74700 , n74706 );
nand ( n74708 , n74381 , n72198 );
nand ( n74709 , n74707 , n74708 );
xor ( n74710 , n74699 , n74709 );
xor ( n74711 , n74710 , n74494 );
xor ( n74712 , n74711 , n74498 );
xor ( n74713 , n74710 , n74494 );
and ( n74714 , n74713 , n74498 );
and ( n74715 , n74710 , n74494 );
or ( n74716 , n74714 , n74715 );
xor ( n74717 , n74502 , n74285 );
xor ( n74718 , n74551 , n74244 );
xor ( n74719 , n74718 , n74474 );
xor ( n74720 , n74717 , n74719 );
xor ( n74721 , n74502 , n74285 );
and ( n74722 , n74721 , n74719 );
and ( n74723 , n74502 , n74285 );
or ( n74724 , n74722 , n74723 );
xor ( n74725 , n74373 , n74622 );
xor ( n74726 , n74478 , n74482 );
not ( n74727 , n70183 );
not ( n74728 , n55124 );
not ( n74729 , n59694 );
or ( n74730 , n74728 , n74729 );
nand ( n74731 , n71052 , n71409 );
nand ( n74732 , n74730 , n74731 );
not ( n74733 , n74732 );
or ( n74734 , n74727 , n74733 );
nand ( n74735 , n74263 , n70193 );
nand ( n74736 , n74734 , n74735 );
xor ( n74737 , n74736 , n74278 );
not ( n74738 , n59984 );
not ( n74739 , n72288 );
not ( n74740 , n54402 );
or ( n74741 , n74739 , n74740 );
not ( n74742 , n69695 );
nand ( n74743 , n74742 , n40149 );
nand ( n74744 , n74741 , n74743 );
not ( n74745 , n74744 );
or ( n74746 , n74738 , n74745 );
nand ( n74747 , n74407 , n67862 );
nand ( n74748 , n74746 , n74747 );
xor ( n74749 , n74737 , n74748 );
xor ( n74750 , n74726 , n74749 );
xor ( n74751 , n74725 , n74750 );
xor ( n74752 , n74373 , n74622 );
and ( n74753 , n74752 , n74750 );
and ( n74754 , n74373 , n74622 );
or ( n74755 , n74753 , n74754 );
xor ( n74756 , n74712 , n74684 );
xor ( n74757 , n74756 , n74399 );
xor ( n74758 , n74712 , n74684 );
and ( n74759 , n74758 , n74399 );
and ( n74760 , n74712 , n74684 );
or ( n74761 , n74759 , n74760 );
xor ( n74762 , n74391 , n74720 );
xor ( n74763 , n74762 , n74440 );
xor ( n74764 , n74391 , n74720 );
and ( n74765 , n74764 , n74440 );
and ( n74766 , n74391 , n74720 );
or ( n74767 , n74765 , n74766 );
xor ( n74768 , n74751 , n74446 );
xor ( n74769 , n74768 , n74757 );
xor ( n74770 , n74751 , n74446 );
and ( n74771 , n74770 , n74757 );
and ( n74772 , n74751 , n74446 );
or ( n74773 , n74771 , n74772 );
xor ( n74774 , n74452 , n74763 );
xor ( n74775 , n74774 , n74769 );
xor ( n74776 , n74452 , n74763 );
and ( n74777 , n74776 , n74769 );
and ( n74778 , n74452 , n74763 );
or ( n74779 , n74777 , n74778 );
xor ( n74780 , n74458 , n74775 );
xor ( n74781 , n74780 , n74464 );
xor ( n74782 , n74458 , n74775 );
and ( n74783 , n74782 , n74464 );
and ( n74784 , n74458 , n74775 );
or ( n74785 , n74783 , n74784 );
xor ( n74786 , n74598 , n74608 );
and ( n74787 , n74786 , n74619 );
and ( n74788 , n74598 , n74608 );
or ( n74789 , n74787 , n74788 );
xor ( n74790 , n74736 , n74278 );
and ( n74791 , n74790 , n74748 );
and ( n74792 , n74736 , n74278 );
or ( n74793 , n74791 , n74792 );
xor ( n74794 , n74565 , n74575 );
and ( n74795 , n74794 , n74587 );
and ( n74796 , n74565 , n74575 );
or ( n74797 , n74795 , n74796 );
xor ( n74798 , n74636 , n74647 );
and ( n74799 , n74798 , n74658 );
and ( n74800 , n74636 , n74647 );
or ( n74801 , n74799 , n74800 );
xor ( n74802 , n74698 , n74209 );
and ( n74803 , n74802 , n74709 );
and ( n74804 , n74698 , n74209 );
or ( n74805 , n74803 , n74804 );
xor ( n74806 , n74670 , n74681 );
and ( n74807 , n74806 , n74525 );
and ( n74808 , n74670 , n74681 );
or ( n74809 , n74807 , n74808 );
xor ( n74810 , n74551 , n74244 );
and ( n74811 , n74810 , n74474 );
and ( n74812 , n74551 , n74244 );
or ( n74813 , n74811 , n74812 );
xor ( n74814 , n74478 , n74482 );
and ( n74815 , n74814 , n74749 );
and ( n74816 , n74478 , n74482 );
or ( n74817 , n74815 , n74816 );
not ( n74818 , n74536 );
not ( n74819 , n65795 );
or ( n74820 , n74818 , n74819 );
xor ( n74821 , n49549 , n67072 );
nand ( n74822 , n70964 , n74821 );
nand ( n74823 , n74820 , n74822 );
and ( n74824 , n64444 , n41288 );
xor ( n74825 , n74823 , n74824 );
not ( n74826 , n61558 );
and ( n74827 , n71361 , n71307 );
not ( n74828 , n71361 );
and ( n74829 , n74828 , n71309 );
or ( n74830 , n74827 , n74829 );
not ( n74831 , n74830 );
or ( n74832 , n74826 , n74831 );
nand ( n74833 , n72484 , n74515 );
nand ( n74834 , n74832 , n74833 );
xor ( n74835 , n74825 , n74834 );
xor ( n74836 , n74823 , n74824 );
and ( n74837 , n74836 , n74834 );
and ( n74838 , n74823 , n74824 );
or ( n74839 , n74837 , n74838 );
not ( n74840 , n70930 );
not ( n74841 , n68878 );
not ( n74842 , n51925 );
or ( n74843 , n74841 , n74842 );
nand ( n74844 , n53258 , n72477 );
nand ( n74845 , n74843 , n74844 );
not ( n74846 , n74845 );
or ( n74847 , n74840 , n74846 );
not ( n74848 , n60960 );
nand ( n74849 , n74848 , n74546 );
nand ( n74850 , n74847 , n74849 );
not ( n74851 , n54316 );
not ( n74852 , n74615 );
or ( n74853 , n74851 , n74852 );
not ( n74854 , n70627 );
not ( n74855 , n63180 );
or ( n74856 , n74854 , n74855 );
nand ( n74857 , n72969 , n54468 );
nand ( n74858 , n74856 , n74857 );
nand ( n74859 , n74858 , n54327 );
nand ( n74860 , n74853 , n74859 );
xor ( n74861 , n74850 , n74860 );
not ( n74862 , n55144 );
not ( n74863 , n74732 );
or ( n74864 , n74862 , n74863 );
not ( n74865 , n72919 );
not ( n74866 , n56407 );
or ( n74867 , n74865 , n74866 );
nand ( n74868 , n72217 , n71409 );
nand ( n74869 , n74867 , n74868 );
nand ( n74870 , n74869 , n70183 );
nand ( n74871 , n74864 , n74870 );
xor ( n74872 , n74861 , n74871 );
xor ( n74873 , n74850 , n74860 );
and ( n74874 , n74873 , n74871 );
and ( n74875 , n74850 , n74860 );
or ( n74876 , n74874 , n74875 );
not ( n74877 , n51766 );
not ( n74878 , n73607 );
not ( n74879 , n62931 );
or ( n74880 , n74878 , n74879 );
nand ( n74881 , n71567 , n52487 );
nand ( n74882 , n74880 , n74881 );
not ( n74883 , n74882 );
or ( n74884 , n74877 , n74883 );
nand ( n74885 , n74677 , n53197 );
nand ( n74886 , n74884 , n74885 );
not ( n74887 , n52757 );
not ( n74888 , n64190 );
not ( n74889 , n69961 );
or ( n74890 , n74888 , n74889 );
nand ( n74891 , n72998 , n64191 );
nand ( n74892 , n74890 , n74891 );
not ( n74893 , n74892 );
or ( n74894 , n74887 , n74893 );
nand ( n74895 , n74654 , n63708 );
nand ( n74896 , n74894 , n74895 );
xor ( n74897 , n74886 , n74896 );
not ( n74898 , n52469 );
not ( n74899 , n69458 );
not ( n74900 , n59913 );
not ( n74901 , n74900 );
or ( n74902 , n74899 , n74901 );
nand ( n74903 , n71509 , n55104 );
nand ( n74904 , n74902 , n74903 );
not ( n74905 , n74904 );
or ( n74906 , n74898 , n74905 );
nand ( n74907 , n74632 , n52854 );
nand ( n74908 , n74906 , n74907 );
xor ( n74909 , n74897 , n74908 );
xor ( n74910 , n74805 , n74909 );
xor ( n74911 , n74910 , n74809 );
xor ( n74912 , n74805 , n74909 );
and ( n74913 , n74912 , n74809 );
and ( n74914 , n74805 , n74909 );
or ( n74915 , n74913 , n74914 );
not ( n74916 , n51533 );
not ( n74917 , n53931 );
not ( n74918 , n59891 );
or ( n74919 , n74917 , n74918 );
nand ( n74920 , n39056 , n71053 );
nand ( n74921 , n74919 , n74920 );
not ( n74922 , n74921 );
or ( n74923 , n74916 , n74922 );
nand ( n74924 , n56355 , n74705 );
nand ( n74925 , n74923 , n74924 );
not ( n74926 , n62085 );
not ( n74927 , n74643 );
or ( n74928 , n74926 , n74927 );
nand ( n74929 , n52191 , n62077 );
nand ( n74930 , n74928 , n74929 );
xor ( n74931 , n74925 , n74930 );
xor ( n74932 , n74931 , n74529 );
not ( n74933 , n54364 );
not ( n74934 , n53596 );
not ( n74935 , n71418 );
or ( n74936 , n74934 , n74935 );
not ( n74937 , n68142 );
nand ( n74938 , n74937 , n71756 );
nand ( n74939 , n74936 , n74938 );
not ( n74940 , n74939 );
or ( n74941 , n74933 , n74940 );
nand ( n74942 , n74596 , n68603 );
nand ( n74943 , n74941 , n74942 );
not ( n74944 , n62654 );
not ( n74945 , n61951 );
not ( n74946 , n72307 );
or ( n74947 , n74945 , n74946 );
nand ( n74948 , n66304 , n66690 );
nand ( n74949 , n74947 , n74948 );
not ( n74950 , n74949 );
or ( n74951 , n74944 , n74950 );
nand ( n74952 , n74666 , n66696 );
nand ( n74953 , n74951 , n74952 );
xor ( n74954 , n74943 , n74953 );
not ( n74955 , n50922 );
not ( n74956 , n65773 );
not ( n74957 , n39333 );
or ( n74958 , n74956 , n74957 );
nand ( n74959 , n39332 , n71042 );
nand ( n74960 , n74958 , n74959 );
not ( n74961 , n74960 );
or ( n74962 , n74955 , n74961 );
nand ( n74963 , n74696 , n52151 );
nand ( n74964 , n74962 , n74963 );
xor ( n74965 , n74954 , n74964 );
xor ( n74966 , n74932 , n74965 );
xor ( n74967 , n74966 , n74813 );
xor ( n74968 , n74932 , n74965 );
and ( n74969 , n74968 , n74813 );
and ( n74970 , n74932 , n74965 );
or ( n74971 , n74969 , n74970 );
xor ( n74972 , n74793 , n74797 );
not ( n74973 , n74744 );
not ( n74974 , n71099 );
or ( n74975 , n74973 , n74974 );
not ( n74976 , n72288 );
not ( n74977 , n57390 );
or ( n74978 , n74976 , n74977 );
nand ( n74979 , n68990 , n74094 );
nand ( n74980 , n74978 , n74979 );
nand ( n74981 , n74980 , n59984 );
nand ( n74982 , n74975 , n74981 );
not ( n74983 , n64164 );
not ( n74984 , n74522 );
and ( n74985 , n74983 , n74984 );
and ( n74986 , n64170 , n71330 );
not ( n74987 , n64170 );
and ( n74988 , n74987 , n51891 );
or ( n74989 , n74986 , n74988 );
not ( n74990 , n74989 );
nor ( n74991 , n74990 , n69703 );
nor ( n74992 , n74985 , n74991 );
xor ( n74993 , n74982 , n74992 );
not ( n74994 , n56777 );
not ( n74995 , n74561 );
or ( n74996 , n74994 , n74995 );
not ( n74997 , n69820 );
not ( n74998 , n71476 );
or ( n74999 , n74997 , n74998 );
nand ( n75000 , n63204 , n56785 );
nand ( n75001 , n74999 , n75000 );
nand ( n75002 , n75001 , n60472 );
nand ( n75003 , n74996 , n75002 );
xor ( n75004 , n74993 , n75003 );
xor ( n75005 , n74972 , n75004 );
xor ( n75006 , n75005 , n74626 );
xor ( n75007 , n75006 , n74817 );
xor ( n75008 , n75005 , n74626 );
and ( n75009 , n75008 , n74817 );
and ( n75010 , n75005 , n74626 );
or ( n75011 , n75009 , n75010 );
xor ( n75012 , n74835 , n74555 );
xor ( n75013 , n75012 , n74789 );
xor ( n75014 , n75013 , n74688 );
not ( n75015 , n72961 );
not ( n75016 , n74571 );
or ( n75017 , n75015 , n75016 );
not ( n75018 , n67568 );
not ( n75019 , n53289 );
or ( n75020 , n75018 , n75019 );
nand ( n75021 , n54646 , n73307 );
nand ( n75022 , n75020 , n75021 );
nand ( n75023 , n75022 , n70604 );
nand ( n75024 , n75017 , n75023 );
buf ( n75025 , n65646 );
not ( n75026 , n75025 );
not ( n75027 , n74583 );
or ( n75028 , n75026 , n75027 );
not ( n75029 , n65184 );
not ( n75030 , n40627 );
or ( n75031 , n75029 , n75030 );
nand ( n75032 , n72160 , n65183 );
nand ( n75033 , n75031 , n75032 );
nand ( n75034 , n75033 , n71466 );
nand ( n75035 , n75028 , n75034 );
xor ( n75036 , n75024 , n75035 );
not ( n75037 , n70487 );
not ( n75038 , n74604 );
or ( n75039 , n75037 , n75038 );
and ( n75040 , n72464 , n51913 );
not ( n75041 , n72464 );
and ( n75042 , n75041 , n51916 );
or ( n75043 , n75040 , n75042 );
nand ( n75044 , n75043 , n60542 );
nand ( n75045 , n75039 , n75044 );
xor ( n75046 , n75036 , n75045 );
xor ( n75047 , n75046 , n74872 );
xor ( n75048 , n75047 , n74801 );
xor ( n75049 , n75014 , n75048 );
xor ( n75050 , n75013 , n74688 );
and ( n75051 , n75050 , n75048 );
and ( n75052 , n75013 , n74688 );
or ( n75053 , n75051 , n75052 );
xor ( n75054 , n74967 , n74911 );
xor ( n75055 , n75054 , n74716 );
xor ( n75056 , n74967 , n74911 );
and ( n75057 , n75056 , n74716 );
and ( n75058 , n74967 , n74911 );
or ( n75059 , n75057 , n75058 );
xor ( n75060 , n74724 , n74755 );
xor ( n75061 , n75060 , n75007 );
xor ( n75062 , n74724 , n74755 );
and ( n75063 , n75062 , n75007 );
and ( n75064 , n74724 , n74755 );
or ( n75065 , n75063 , n75064 );
xor ( n75066 , n75049 , n74761 );
xor ( n75067 , n75066 , n75055 );
xor ( n75068 , n75049 , n74761 );
and ( n75069 , n75068 , n75055 );
and ( n75070 , n75049 , n74761 );
or ( n75071 , n75069 , n75070 );
xor ( n75072 , n74767 , n75061 );
xor ( n75073 , n75072 , n74773 );
xor ( n75074 , n74767 , n75061 );
and ( n75075 , n75074 , n74773 );
and ( n75076 , n74767 , n75061 );
or ( n75077 , n75075 , n75076 );
xor ( n75078 , n75067 , n75073 );
xor ( n75079 , n75078 , n74779 );
xor ( n75080 , n75067 , n75073 );
and ( n75081 , n75080 , n74779 );
and ( n75082 , n75067 , n75073 );
or ( n75083 , n75081 , n75082 );
xor ( n75084 , n74982 , n74992 );
and ( n75085 , n75084 , n75003 );
and ( n75086 , n74982 , n74992 );
or ( n75087 , n75085 , n75086 );
xor ( n75088 , n75024 , n75035 );
and ( n75089 , n75088 , n75045 );
and ( n75090 , n75024 , n75035 );
or ( n75091 , n75089 , n75090 );
xor ( n75092 , n74943 , n74953 );
and ( n75093 , n75092 , n74964 );
and ( n75094 , n74943 , n74953 );
or ( n75095 , n75093 , n75094 );
xor ( n75096 , n74925 , n74930 );
and ( n75097 , n75096 , n74529 );
and ( n75098 , n74925 , n74930 );
or ( n75099 , n75097 , n75098 );
xor ( n75100 , n74886 , n74896 );
and ( n75101 , n75100 , n74908 );
and ( n75102 , n74886 , n74896 );
or ( n75103 , n75101 , n75102 );
xor ( n75104 , n74835 , n74555 );
and ( n75105 , n75104 , n74789 );
and ( n75106 , n74835 , n74555 );
or ( n75107 , n75105 , n75106 );
xor ( n75108 , n74793 , n74797 );
and ( n75109 , n75108 , n75004 );
and ( n75110 , n74793 , n74797 );
or ( n75111 , n75109 , n75110 );
xor ( n75112 , n75046 , n74872 );
and ( n75113 , n75112 , n74801 );
and ( n75114 , n75046 , n74872 );
or ( n75115 , n75113 , n75114 );
not ( n75116 , n59811 );
not ( n75117 , n58167 );
or ( n75118 , n75116 , n75117 );
nand ( n75119 , n75118 , n62077 );
not ( n75120 , n74989 );
not ( n75121 , n67061 );
or ( n75122 , n75120 , n75121 );
not ( n75123 , n69704 );
not ( n75124 , n70889 );
or ( n75125 , n75123 , n75124 );
not ( n75126 , n52079 );
nand ( n75127 , n75126 , n64170 );
nand ( n75128 , n75125 , n75127 );
nand ( n75129 , n67068 , n75128 );
nand ( n75130 , n75122 , n75129 );
xor ( n75131 , n75119 , n75130 );
not ( n75132 , n74821 );
or ( n75133 , n71959 , n75132 );
and ( n75134 , n64443 , n71691 );
and ( n75135 , n71971 , n64451 );
nor ( n75136 , n75134 , n75135 );
or ( n75137 , n75136 , n70965 );
nand ( n75138 , n75133 , n75137 );
xor ( n75139 , n75131 , n75138 );
xor ( n75140 , n75119 , n75130 );
and ( n75141 , n75140 , n75138 );
and ( n75142 , n75119 , n75130 );
or ( n75143 , n75141 , n75142 );
and ( n75144 , n71971 , n41217 );
not ( n75145 , n61558 );
not ( n75146 , n71309 );
not ( n75147 , n70186 );
or ( n75148 , n75146 , n75147 );
nand ( n75149 , n68598 , n69333 );
nand ( n75150 , n75148 , n75149 );
not ( n75151 , n75150 );
or ( n75152 , n75145 , n75151 );
not ( n75153 , n69728 );
nand ( n75154 , n75153 , n74830 );
nand ( n75155 , n75152 , n75154 );
xor ( n75156 , n75144 , n75155 );
not ( n75157 , n54316 );
not ( n75158 , n74858 );
or ( n75159 , n75157 , n75158 );
not ( n75160 , n71395 );
buf ( n75161 , n67702 );
not ( n75162 , n75161 );
not ( n75163 , n75162 );
or ( n75164 , n75160 , n75163 );
nand ( n75165 , n62618 , n54468 );
nand ( n75166 , n75164 , n75165 );
nand ( n75167 , n75166 , n54327 );
nand ( n75168 , n75159 , n75167 );
xor ( n75169 , n75156 , n75168 );
xor ( n75170 , n75144 , n75155 );
and ( n75171 , n75170 , n75168 );
and ( n75172 , n75144 , n75155 );
or ( n75173 , n75171 , n75172 );
xor ( n75174 , n75095 , n75103 );
not ( n75175 , n61465 );
and ( n75176 , n66652 , n71767 );
not ( n75177 , n66652 );
and ( n75178 , n75177 , n59612 );
nor ( n75179 , n75176 , n75178 );
not ( n75180 , n75179 );
or ( n75181 , n75175 , n75180 );
nand ( n75182 , n75033 , n75025 );
nand ( n75183 , n75181 , n75182 );
not ( n75184 , n75043 );
not ( n75185 , n70487 );
or ( n75186 , n75184 , n75185 );
not ( n75187 , n72464 );
not ( n75188 , n66798 );
or ( n75189 , n75187 , n75188 );
nand ( n75190 , n74581 , n66983 );
nand ( n75191 , n75189 , n75190 );
nand ( n75192 , n75191 , n60542 );
nand ( n75193 , n75186 , n75192 );
xor ( n75194 , n75183 , n75193 );
not ( n75195 , n68603 );
not ( n75196 , n74939 );
or ( n75197 , n75195 , n75196 );
not ( n75198 , n55089 );
not ( n75199 , n39894 );
or ( n75200 , n75198 , n75199 );
nand ( n75201 , n71863 , n72238 );
nand ( n75202 , n75200 , n75201 );
nand ( n75203 , n75202 , n53620 );
nand ( n75204 , n75197 , n75203 );
xor ( n75205 , n75194 , n75204 );
xor ( n75206 , n75174 , n75205 );
xor ( n75207 , n75095 , n75103 );
and ( n75208 , n75207 , n75205 );
and ( n75209 , n75095 , n75103 );
or ( n75210 , n75208 , n75209 );
not ( n75211 , n51766 );
not ( n75212 , n73607 );
not ( n75213 , n73400 );
or ( n75214 , n75212 , n75213 );
nand ( n75215 , n68667 , n52487 );
nand ( n75216 , n75214 , n75215 );
not ( n75217 , n75216 );
or ( n75218 , n75211 , n75217 );
nand ( n75219 , n74882 , n53197 );
nand ( n75220 , n75218 , n75219 );
not ( n75221 , n63708 );
not ( n75222 , n74892 );
or ( n75223 , n75221 , n75222 );
not ( n75224 , n50306 );
not ( n75225 , n42399 );
or ( n75226 , n75224 , n75225 );
nand ( n75227 , n68381 , n66705 );
nand ( n75228 , n75226 , n75227 );
nand ( n75229 , n75228 , n52757 );
nand ( n75230 , n75223 , n75229 );
xor ( n75231 , n75220 , n75230 );
not ( n75232 , n53571 );
not ( n75233 , n69458 );
not ( n75234 , n73428 );
or ( n75235 , n75233 , n75234 );
nand ( n75236 , n60386 , n55104 );
nand ( n75237 , n75235 , n75236 );
not ( n75238 , n75237 );
or ( n75239 , n75232 , n75238 );
nand ( n75240 , n74904 , n52854 );
nand ( n75241 , n75239 , n75240 );
xor ( n75242 , n75231 , n75241 );
not ( n75243 , n62654 );
not ( n75244 , n61951 );
not ( n75245 , n74639 );
or ( n75246 , n75244 , n75245 );
nand ( n75247 , n71875 , n66690 );
nand ( n75248 , n75246 , n75247 );
not ( n75249 , n75248 );
or ( n75250 , n75243 , n75249 );
nand ( n75251 , n74949 , n66696 );
nand ( n75252 , n75250 , n75251 );
not ( n75253 , n52151 );
not ( n75254 , n74960 );
or ( n75255 , n75253 , n75254 );
not ( n75256 , n65773 );
not ( n75257 , n39254 );
or ( n75258 , n75256 , n75257 );
nand ( n75259 , n69530 , n71042 );
nand ( n75260 , n75258 , n75259 );
nand ( n75261 , n75260 , n50922 );
nand ( n75262 , n75255 , n75261 );
xor ( n75263 , n75252 , n75262 );
not ( n75264 , n72198 );
not ( n75265 , n74921 );
or ( n75266 , n75264 , n75265 );
not ( n75267 , n53931 );
not ( n75268 , n62394 );
or ( n75269 , n75267 , n75268 );
nand ( n75270 , n38499 , n71053 );
nand ( n75271 , n75269 , n75270 );
nand ( n75272 , n75271 , n51533 );
nand ( n75273 , n75266 , n75272 );
xor ( n75274 , n75263 , n75273 );
xor ( n75275 , n75242 , n75274 );
xor ( n75276 , n75275 , n75107 );
xor ( n75277 , n75242 , n75274 );
and ( n75278 , n75277 , n75107 );
and ( n75279 , n75242 , n75274 );
or ( n75280 , n75278 , n75279 );
xor ( n75281 , n75139 , n74839 );
xor ( n75282 , n75281 , n74876 );
xor ( n75283 , n75282 , n75115 );
xor ( n75284 , n75087 , n75091 );
not ( n75285 , n70930 );
not ( n75286 , n72477 );
not ( n75287 , n75286 );
not ( n75288 , n70278 );
or ( n75289 , n75287 , n75288 );
nand ( n75290 , n69442 , n72477 );
nand ( n75291 , n75289 , n75290 );
not ( n75292 , n75291 );
or ( n75293 , n75285 , n75292 );
nand ( n75294 , n74845 , n66136 );
nand ( n75295 , n75293 , n75294 );
not ( n75296 , n70183 );
not ( n75297 , n55120 );
not ( n75298 , n70290 );
or ( n75299 , n75297 , n75298 );
nand ( n75300 , n72607 , n71409 );
nand ( n75301 , n75299 , n75300 );
not ( n75302 , n75301 );
or ( n75303 , n75296 , n75302 );
nand ( n75304 , n74869 , n55144 );
nand ( n75305 , n75303 , n75304 );
xor ( n75306 , n75295 , n75305 );
not ( n75307 , n74992 );
xor ( n75308 , n75306 , n75307 );
xor ( n75309 , n75284 , n75308 );
xor ( n75310 , n75283 , n75309 );
xor ( n75311 , n75282 , n75115 );
and ( n75312 , n75311 , n75309 );
and ( n75313 , n75282 , n75115 );
or ( n75314 , n75312 , n75313 );
xor ( n75315 , n75111 , n74915 );
xor ( n75316 , n75315 , n75206 );
xor ( n75317 , n75111 , n74915 );
and ( n75318 , n75317 , n75206 );
and ( n75319 , n75111 , n74915 );
or ( n75320 , n75318 , n75319 );
not ( n75321 , n59984 );
not ( n75322 , n74402 );
not ( n75323 , n73327 );
or ( n75324 , n75322 , n75323 );
nand ( n75325 , n40382 , n72289 );
nand ( n75326 , n75324 , n75325 );
not ( n75327 , n75326 );
or ( n75328 , n75321 , n75327 );
nand ( n75329 , n74980 , n67862 );
nand ( n75330 , n75328 , n75329 );
not ( n75331 , n60472 );
not ( n75332 , n69820 );
not ( n75333 , n54402 );
or ( n75334 , n75332 , n75333 );
nand ( n75335 , n69409 , n69819 );
nand ( n75336 , n75334 , n75335 );
not ( n75337 , n75336 );
or ( n75338 , n75331 , n75337 );
nand ( n75339 , n75001 , n56777 );
nand ( n75340 , n75338 , n75339 );
xor ( n75341 , n75330 , n75340 );
not ( n75342 , n72710 );
not ( n75343 , n66963 );
not ( n75344 , n75343 );
not ( n75345 , n53661 );
or ( n75346 , n75344 , n75345 );
nand ( n75347 , n59601 , n73307 );
nand ( n75348 , n75346 , n75347 );
not ( n75349 , n75348 );
or ( n75350 , n75342 , n75349 );
nand ( n75351 , n72961 , n75022 );
nand ( n75352 , n75350 , n75351 );
xor ( n75353 , n75341 , n75352 );
xor ( n75354 , n75353 , n75169 );
xor ( n75355 , n75354 , n75099 );
xor ( n75356 , n75355 , n75276 );
xor ( n75357 , n75356 , n74971 );
xor ( n75358 , n75355 , n75276 );
and ( n75359 , n75358 , n74971 );
and ( n75360 , n75355 , n75276 );
or ( n75361 , n75359 , n75360 );
xor ( n75362 , n75011 , n75310 );
xor ( n75363 , n75362 , n75053 );
xor ( n75364 , n75011 , n75310 );
and ( n75365 , n75364 , n75053 );
and ( n75366 , n75011 , n75310 );
or ( n75367 , n75365 , n75366 );
xor ( n75368 , n75316 , n75059 );
xor ( n75369 , n75368 , n75357 );
xor ( n75370 , n75316 , n75059 );
and ( n75371 , n75370 , n75357 );
and ( n75372 , n75316 , n75059 );
or ( n75373 , n75371 , n75372 );
xor ( n75374 , n75065 , n75363 );
xor ( n75375 , n75374 , n75071 );
xor ( n75376 , n75065 , n75363 );
and ( n75377 , n75376 , n75071 );
and ( n75378 , n75065 , n75363 );
or ( n75379 , n75377 , n75378 );
xor ( n75380 , n75369 , n75375 );
xor ( n75381 , n75380 , n75077 );
xor ( n75382 , n75369 , n75375 );
and ( n75383 , n75382 , n75077 );
and ( n75384 , n75369 , n75375 );
or ( n75385 , n75383 , n75384 );
xor ( n75386 , n75295 , n75305 );
and ( n75387 , n75386 , n75307 );
and ( n75388 , n75295 , n75305 );
or ( n75389 , n75387 , n75388 );
xor ( n75390 , n75330 , n75340 );
and ( n75391 , n75390 , n75352 );
and ( n75392 , n75330 , n75340 );
or ( n75393 , n75391 , n75392 );
xor ( n75394 , n75183 , n75193 );
and ( n75395 , n75394 , n75204 );
and ( n75396 , n75183 , n75193 );
or ( n75397 , n75395 , n75396 );
xor ( n75398 , n75252 , n75262 );
and ( n75399 , n75398 , n75273 );
and ( n75400 , n75252 , n75262 );
or ( n75401 , n75399 , n75400 );
xor ( n75402 , n75220 , n75230 );
and ( n75403 , n75402 , n75241 );
and ( n75404 , n75220 , n75230 );
or ( n75405 , n75403 , n75404 );
xor ( n75406 , n75139 , n74839 );
and ( n75407 , n75406 , n74876 );
and ( n75408 , n75139 , n74839 );
or ( n75409 , n75407 , n75408 );
xor ( n75410 , n75087 , n75091 );
and ( n75411 , n75410 , n75308 );
and ( n75412 , n75087 , n75091 );
or ( n75413 , n75411 , n75412 );
xor ( n75414 , n75353 , n75169 );
and ( n75415 , n75414 , n75099 );
and ( n75416 , n75353 , n75169 );
or ( n75417 , n75415 , n75416 );
and ( n75418 , n49549 , n67072 );
not ( n75419 , n75128 );
not ( n75420 , n67061 );
or ( n75421 , n75419 , n75420 );
not ( n75422 , n72083 );
not ( n75423 , n50654 );
or ( n75424 , n75422 , n75423 );
nand ( n75425 , n71361 , n69704 );
nand ( n75426 , n75424 , n75425 );
buf ( n75427 , n67068 );
nand ( n75428 , n75426 , n75427 );
nand ( n75429 , n75421 , n75428 );
xor ( n75430 , n75418 , n75429 );
not ( n75431 , n63411 );
not ( n75432 , n75136 );
and ( n75433 , n75431 , n75432 );
not ( n75434 , n71331 );
not ( n75435 , n64443 );
or ( n75436 , n75434 , n75435 );
nand ( n75437 , n67072 , n41037 );
nand ( n75438 , n75436 , n75437 );
not ( n75439 , n75438 );
nor ( n75440 , n75439 , n70965 );
nor ( n75441 , n75433 , n75440 );
xor ( n75442 , n75430 , n75441 );
xor ( n75443 , n75418 , n75429 );
and ( n75444 , n75443 , n75441 );
and ( n75445 , n75418 , n75429 );
or ( n75446 , n75444 , n75445 );
not ( n75447 , n61558 );
not ( n75448 , n61540 );
not ( n75449 , n51925 );
or ( n75450 , n75448 , n75449 );
nand ( n75451 , n53258 , n69333 );
nand ( n75452 , n75450 , n75451 );
not ( n75453 , n75452 );
or ( n75454 , n75447 , n75453 );
nand ( n75455 , n75150 , n72810 );
nand ( n75456 , n75454 , n75455 );
not ( n75457 , n70193 );
not ( n75458 , n75301 );
or ( n75459 , n75457 , n75458 );
not ( n75460 , n55120 );
not ( n75461 , n63180 );
or ( n75462 , n75460 , n75461 );
nand ( n75463 , n70653 , n71409 );
nand ( n75464 , n75462 , n75463 );
nand ( n75465 , n75464 , n70183 );
nand ( n75466 , n75459 , n75465 );
xor ( n75467 , n75456 , n75466 );
not ( n75468 , n67862 );
not ( n75469 , n75326 );
or ( n75470 , n75468 , n75469 );
not ( n75471 , n74402 );
not ( n75472 , n70661 );
or ( n75473 , n75471 , n75472 );
nand ( n75474 , n72217 , n55846 );
nand ( n75475 , n75473 , n75474 );
nand ( n75476 , n75475 , n59984 );
nand ( n75477 , n75470 , n75476 );
xor ( n75478 , n75467 , n75477 );
xor ( n75479 , n75456 , n75466 );
and ( n75480 , n75479 , n75477 );
and ( n75481 , n75456 , n75466 );
or ( n75482 , n75480 , n75481 );
not ( n75483 , n66696 );
not ( n75484 , n75248 );
or ( n75485 , n75483 , n75484 );
nand ( n75486 , n62654 , n61951 );
nand ( n75487 , n75485 , n75486 );
xor ( n75488 , n75143 , n75487 );
not ( n75489 , n52469 );
and ( n75490 , n52841 , n71567 );
not ( n75491 , n52841 );
and ( n75492 , n75491 , n68206 );
nor ( n75493 , n75490 , n75492 );
not ( n75494 , n75493 );
or ( n75495 , n75489 , n75494 );
nand ( n75496 , n75237 , n52854 );
nand ( n75497 , n75495 , n75496 );
xor ( n75498 , n75488 , n75497 );
not ( n75499 , n63708 );
not ( n75500 , n75228 );
or ( n75501 , n75499 , n75500 );
not ( n75502 , n50306 );
not ( n75503 , n67269 );
or ( n75504 , n75502 , n75503 );
nand ( n75505 , n73048 , n64191 );
nand ( n75506 , n75504 , n75505 );
nand ( n75507 , n75506 , n52757 );
nand ( n75508 , n75501 , n75507 );
not ( n75509 , n72198 );
not ( n75510 , n75271 );
or ( n75511 , n75509 , n75510 );
not ( n75512 , n53931 );
not ( n75513 , n60855 );
or ( n75514 , n75512 , n75513 );
nand ( n75515 , n69919 , n71053 );
nand ( n75516 , n75514 , n75515 );
nand ( n75517 , n75516 , n51533 );
nand ( n75518 , n75511 , n75517 );
xor ( n75519 , n75508 , n75518 );
not ( n75520 , n72220 );
not ( n75521 , n73607 );
not ( n75522 , n59891 );
or ( n75523 , n75521 , n75522 );
nand ( n75524 , n39056 , n52110 );
nand ( n75525 , n75523 , n75524 );
not ( n75526 , n75525 );
or ( n75527 , n75520 , n75526 );
nand ( n75528 , n75216 , n53197 );
nand ( n75529 , n75527 , n75528 );
xor ( n75530 , n75519 , n75529 );
xor ( n75531 , n75498 , n75530 );
not ( n75532 , n52151 );
not ( n75533 , n75260 );
or ( n75534 , n75532 , n75533 );
not ( n75535 , n57187 );
not ( n75536 , n72252 );
or ( n75537 , n75535 , n75536 );
nand ( n75538 , n71577 , n71042 );
nand ( n75539 , n75537 , n75538 );
nand ( n75540 , n75539 , n50922 );
nand ( n75541 , n75534 , n75540 );
not ( n75542 , n68603 );
not ( n75543 , n75202 );
or ( n75544 , n75542 , n75543 );
not ( n75545 , n55089 );
not ( n75546 , n67037 );
or ( n75547 , n75545 , n75546 );
not ( n75548 , n67040 );
nand ( n75549 , n75548 , n72238 );
nand ( n75550 , n75547 , n75549 );
nand ( n75551 , n75550 , n54364 );
nand ( n75552 , n75544 , n75551 );
xor ( n75553 , n75541 , n75552 );
xor ( n75554 , n75553 , n75442 );
xor ( n75555 , n75531 , n75554 );
xor ( n75556 , n75498 , n75530 );
and ( n75557 , n75556 , n75554 );
and ( n75558 , n75498 , n75530 );
or ( n75559 , n75557 , n75558 );
xor ( n75560 , n75409 , n75210 );
xor ( n75561 , n75173 , n75389 );
xor ( n75562 , n75561 , n75393 );
xor ( n75563 , n75560 , n75562 );
xor ( n75564 , n75409 , n75210 );
and ( n75565 , n75564 , n75562 );
and ( n75566 , n75409 , n75210 );
or ( n75567 , n75565 , n75566 );
xor ( n75568 , n75417 , n75413 );
xor ( n75569 , n75397 , n75401 );
not ( n75570 , n72131 );
not ( n75571 , n75191 );
or ( n75572 , n75570 , n75571 );
not ( n75573 , n72464 );
not ( n75574 , n52432 );
or ( n75575 , n75573 , n75574 );
nand ( n75576 , n72160 , n66983 );
nand ( n75577 , n75575 , n75576 );
buf ( n75578 , n60542 );
nand ( n75579 , n75577 , n75578 );
nand ( n75580 , n75572 , n75579 );
not ( n75581 , n70500 );
not ( n75582 , n75291 );
or ( n75583 , n75581 , n75582 );
not ( n75584 , n70506 );
not ( n75585 , n60138 );
or ( n75586 , n75584 , n75585 );
nand ( n75587 , n72945 , n67084 );
nand ( n75588 , n75586 , n75587 );
nand ( n75589 , n75588 , n70930 );
nand ( n75590 , n75583 , n75589 );
xor ( n75591 , n75580 , n75590 );
not ( n75592 , n54327 );
not ( n75593 , n70627 );
not ( n75594 , n66215 );
not ( n75595 , n75594 );
or ( n75596 , n75593 , n75595 );
nand ( n75597 , n66215 , n54468 );
nand ( n75598 , n75596 , n75597 );
not ( n75599 , n75598 );
or ( n75600 , n75592 , n75599 );
nand ( n75601 , n75166 , n72142 );
nand ( n75602 , n75600 , n75601 );
xor ( n75603 , n75591 , n75602 );
xor ( n75604 , n75569 , n75603 );
xor ( n75605 , n75568 , n75604 );
xor ( n75606 , n75417 , n75413 );
and ( n75607 , n75606 , n75604 );
and ( n75608 , n75417 , n75413 );
or ( n75609 , n75607 , n75608 );
not ( n75610 , n56777 );
not ( n75611 , n75336 );
or ( n75612 , n75610 , n75611 );
not ( n75613 , n72589 );
not ( n75614 , n57390 );
or ( n75615 , n75613 , n75614 );
nand ( n75616 , n68994 , n71362 );
nand ( n75617 , n75615 , n75616 );
nand ( n75618 , n75617 , n72185 );
nand ( n75619 , n75612 , n75618 );
not ( n75620 , n72182 );
not ( n75621 , n75348 );
or ( n75622 , n75620 , n75621 );
not ( n75623 , n73977 );
not ( n75624 , n66236 );
or ( n75625 , n75623 , n75624 );
nand ( n75626 , n40364 , n66963 );
nand ( n75627 , n75625 , n75626 );
nand ( n75628 , n75627 , n72710 );
nand ( n75629 , n75622 , n75628 );
xor ( n75630 , n75619 , n75629 );
not ( n75631 , n75025 );
not ( n75632 , n75179 );
or ( n75633 , n75631 , n75632 );
not ( n75634 , n58642 );
not ( n75635 , n54020 );
or ( n75636 , n75634 , n75635 );
nand ( n75637 , n54646 , n66652 );
nand ( n75638 , n75636 , n75637 );
nand ( n75639 , n75638 , n61465 );
nand ( n75640 , n75633 , n75639 );
xor ( n75641 , n75630 , n75640 );
xor ( n75642 , n75478 , n75641 );
xor ( n75643 , n75642 , n75405 );
xor ( n75644 , n75643 , n75280 );
xor ( n75645 , n75644 , n75555 );
xor ( n75646 , n75643 , n75280 );
and ( n75647 , n75646 , n75555 );
and ( n75648 , n75643 , n75280 );
or ( n75649 , n75647 , n75648 );
xor ( n75650 , n75314 , n75563 );
xor ( n75651 , n75650 , n75320 );
xor ( n75652 , n75314 , n75563 );
and ( n75653 , n75652 , n75320 );
and ( n75654 , n75314 , n75563 );
or ( n75655 , n75653 , n75654 );
xor ( n75656 , n75605 , n75361 );
xor ( n75657 , n75656 , n75645 );
xor ( n75658 , n75605 , n75361 );
and ( n75659 , n75658 , n75645 );
and ( n75660 , n75605 , n75361 );
or ( n75661 , n75659 , n75660 );
xor ( n75662 , n75367 , n75651 );
xor ( n75663 , n75662 , n75373 );
xor ( n75664 , n75367 , n75651 );
and ( n75665 , n75664 , n75373 );
and ( n75666 , n75367 , n75651 );
or ( n75667 , n75665 , n75666 );
xor ( n75668 , n75657 , n75663 );
xor ( n75669 , n75668 , n75379 );
xor ( n75670 , n75657 , n75663 );
and ( n75671 , n75670 , n75379 );
and ( n75672 , n75657 , n75663 );
or ( n75673 , n75671 , n75672 );
xor ( n75674 , n75619 , n75629 );
and ( n75675 , n75674 , n75640 );
and ( n75676 , n75619 , n75629 );
or ( n75677 , n75675 , n75676 );
xor ( n75678 , n75580 , n75590 );
and ( n75679 , n75678 , n75602 );
and ( n75680 , n75580 , n75590 );
or ( n75681 , n75679 , n75680 );
xor ( n75682 , n75508 , n75518 );
and ( n75683 , n75682 , n75529 );
and ( n75684 , n75508 , n75518 );
or ( n75685 , n75683 , n75684 );
xor ( n75686 , n75143 , n75487 );
and ( n75687 , n75686 , n75497 );
and ( n75688 , n75143 , n75487 );
or ( n75689 , n75687 , n75688 );
xor ( n75690 , n75541 , n75552 );
and ( n75691 , n75690 , n75442 );
and ( n75692 , n75541 , n75552 );
or ( n75693 , n75691 , n75692 );
xor ( n75694 , n75173 , n75389 );
and ( n75695 , n75694 , n75393 );
and ( n75696 , n75173 , n75389 );
or ( n75697 , n75695 , n75696 );
xor ( n75698 , n75478 , n75641 );
and ( n75699 , n75698 , n75405 );
and ( n75700 , n75478 , n75641 );
or ( n75701 , n75699 , n75700 );
xor ( n75702 , n75397 , n75401 );
and ( n75703 , n75702 , n75603 );
and ( n75704 , n75397 , n75401 );
or ( n75705 , n75703 , n75704 );
not ( n75706 , n72636 );
not ( n75707 , n62663 );
or ( n75708 , n75706 , n75707 );
nand ( n75709 , n75708 , n61951 );
not ( n75710 , n75438 );
not ( n75711 , n65089 );
or ( n75712 , n75710 , n75711 );
xor ( n75713 , n70889 , n66575 );
nand ( n75714 , n70964 , n75713 );
nand ( n75715 , n75712 , n75714 );
xor ( n75716 , n75709 , n75715 );
and ( n75717 , n67072 , n71691 );
xor ( n75718 , n75716 , n75717 );
xor ( n75719 , n75709 , n75715 );
and ( n75720 , n75719 , n75717 );
and ( n75721 , n75709 , n75715 );
or ( n75722 , n75720 , n75721 );
not ( n75723 , n75427 );
not ( n75724 , n64170 );
not ( n75725 , n52286 );
or ( n75726 , n75724 , n75725 );
nand ( n75727 , n71093 , n66089 );
nand ( n75728 , n75726 , n75727 );
not ( n75729 , n75728 );
or ( n75730 , n75723 , n75729 );
nand ( n75731 , n67061 , n75426 );
nand ( n75732 , n75730 , n75731 );
not ( n75733 , n55144 );
not ( n75734 , n75464 );
or ( n75735 , n75733 , n75734 );
not ( n75736 , n55120 );
not ( n75737 , n59651 );
or ( n75738 , n75736 , n75737 );
nand ( n75739 , n75161 , n71409 );
nand ( n75740 , n75738 , n75739 );
nand ( n75741 , n75740 , n70183 );
nand ( n75742 , n75735 , n75741 );
xor ( n75743 , n75732 , n75742 );
not ( n75744 , n61558 );
not ( n75745 , n61540 );
not ( n75746 , n51602 );
or ( n75747 , n75745 , n75746 );
not ( n75748 , n61540 );
nand ( n75749 , n69442 , n75748 );
nand ( n75750 , n75747 , n75749 );
not ( n75751 , n75750 );
or ( n75752 , n75744 , n75751 );
not ( n75753 , n69728 );
nand ( n75754 , n75452 , n75753 );
nand ( n75755 , n75752 , n75754 );
xor ( n75756 , n75743 , n75755 );
xor ( n75757 , n75732 , n75742 );
and ( n75758 , n75757 , n75755 );
and ( n75759 , n75732 , n75742 );
or ( n75760 , n75758 , n75759 );
not ( n75761 , n50922 );
and ( n75762 , n50895 , n68381 );
not ( n75763 , n50895 );
and ( n75764 , n75763 , n42399 );
nor ( n75765 , n75762 , n75764 );
not ( n75766 , n75765 );
or ( n75767 , n75761 , n75766 );
nand ( n75768 , n75539 , n52151 );
nand ( n75769 , n75767 , n75768 );
not ( n75770 , n53620 );
not ( n75771 , n55089 );
not ( n75772 , n71904 );
or ( n75773 , n75771 , n75772 );
nand ( n75774 , n72238 , n39681 );
nand ( n75775 , n75773 , n75774 );
not ( n75776 , n75775 );
or ( n75777 , n75770 , n75776 );
nand ( n75778 , n75550 , n68603 );
nand ( n75779 , n75777 , n75778 );
xor ( n75780 , n75769 , n75779 );
xor ( n75781 , n75780 , n75718 );
not ( n75782 , n51533 );
not ( n75783 , n53931 );
not ( n75784 , n71176 );
or ( n75785 , n75783 , n75784 );
nand ( n75786 , n69530 , n71053 );
nand ( n75787 , n75785 , n75786 );
not ( n75788 , n75787 );
or ( n75789 , n75782 , n75788 );
nand ( n75790 , n75516 , n56355 );
nand ( n75791 , n75789 , n75790 );
not ( n75792 , n53197 );
not ( n75793 , n75525 );
or ( n75794 , n75792 , n75793 );
not ( n75795 , n73607 );
not ( n75796 , n68652 );
or ( n75797 , n75795 , n75796 );
nand ( n75798 , n38499 , n52487 );
nand ( n75799 , n75797 , n75798 );
nand ( n75800 , n75799 , n72220 );
nand ( n75801 , n75794 , n75800 );
xor ( n75802 , n75791 , n75801 );
not ( n75803 , n52854 );
not ( n75804 , n75493 );
or ( n75805 , n75803 , n75804 );
not ( n75806 , n69458 );
not ( n75807 , n65532 );
or ( n75808 , n75806 , n75807 );
nand ( n75809 , n39575 , n53947 );
nand ( n75810 , n75808 , n75809 );
nand ( n75811 , n75810 , n53571 );
nand ( n75812 , n75805 , n75811 );
xor ( n75813 , n75802 , n75812 );
xor ( n75814 , n75781 , n75813 );
not ( n75815 , n66136 );
not ( n75816 , n75588 );
or ( n75817 , n75815 , n75816 );
not ( n75818 , n68878 );
not ( n75819 , n52208 );
or ( n75820 , n75818 , n75819 );
nand ( n75821 , n40592 , n67084 );
nand ( n75822 , n75820 , n75821 );
nand ( n75823 , n75822 , n70930 );
nand ( n75824 , n75817 , n75823 );
not ( n75825 , n54316 );
not ( n75826 , n75598 );
or ( n75827 , n75825 , n75826 );
not ( n75828 , n70627 );
not ( n75829 , n59414 );
or ( n75830 , n75828 , n75829 );
nand ( n75831 , n71013 , n54468 );
nand ( n75832 , n75830 , n75831 );
nand ( n75833 , n75832 , n54327 );
nand ( n75834 , n75827 , n75833 );
xor ( n75835 , n75824 , n75834 );
not ( n75836 , n52757 );
and ( n75837 , n64191 , n73371 );
not ( n75838 , n64191 );
and ( n75839 , n75838 , n71162 );
nor ( n75840 , n75837 , n75839 );
not ( n75841 , n75840 );
or ( n75842 , n75836 , n75841 );
nand ( n75843 , n75506 , n63708 );
nand ( n75844 , n75842 , n75843 );
xor ( n75845 , n75835 , n75844 );
xor ( n75846 , n75814 , n75845 );
xor ( n75847 , n75781 , n75813 );
and ( n75848 , n75847 , n75845 );
and ( n75849 , n75781 , n75813 );
or ( n75850 , n75848 , n75849 );
xor ( n75851 , n75697 , n75693 );
xor ( n75852 , n75851 , n75705 );
xor ( n75853 , n75697 , n75693 );
and ( n75854 , n75853 , n75705 );
and ( n75855 , n75697 , n75693 );
or ( n75856 , n75854 , n75855 );
xor ( n75857 , n75446 , n75482 );
xor ( n75858 , n75857 , n75677 );
xor ( n75859 , n75701 , n75858 );
not ( n75860 , n59984 );
not ( n75861 , n71371 );
not ( n75862 , n72606 );
or ( n75863 , n75861 , n75862 );
nand ( n75864 , n69237 , n40514 );
nand ( n75865 , n75863 , n75864 );
not ( n75866 , n75865 );
or ( n75867 , n75860 , n75866 );
nand ( n75868 , n75475 , n71099 );
nand ( n75869 , n75867 , n75868 );
not ( n75870 , n75441 );
xor ( n75871 , n75869 , n75870 );
not ( n75872 , n72185 );
not ( n75873 , n56786 );
not ( n75874 , n59694 );
or ( n75875 , n75873 , n75874 );
nand ( n75876 , n40382 , n56785 );
nand ( n75877 , n75875 , n75876 );
not ( n75878 , n75877 );
or ( n75879 , n75872 , n75878 );
nand ( n75880 , n75617 , n56777 );
nand ( n75881 , n75879 , n75880 );
xor ( n75882 , n75871 , n75881 );
xor ( n75883 , n75756 , n75882 );
xor ( n75884 , n75883 , n75681 );
xor ( n75885 , n75859 , n75884 );
xor ( n75886 , n75701 , n75858 );
and ( n75887 , n75886 , n75884 );
and ( n75888 , n75701 , n75858 );
or ( n75889 , n75887 , n75888 );
xor ( n75890 , n75685 , n75689 );
not ( n75891 , n72710 );
not ( n75892 , n73977 );
not ( n75893 , n54402 );
or ( n75894 , n75892 , n75893 );
nand ( n75895 , n40149 , n66963 );
nand ( n75896 , n75894 , n75895 );
not ( n75897 , n75896 );
or ( n75898 , n75891 , n75897 );
nand ( n75899 , n75627 , n72182 );
nand ( n75900 , n75898 , n75899 );
not ( n75901 , n61465 );
not ( n75902 , n58642 );
not ( n75903 , n40225 );
or ( n75904 , n75902 , n75903 );
nand ( n75905 , n53660 , n66652 );
nand ( n75906 , n75904 , n75905 );
not ( n75907 , n75906 );
or ( n75908 , n75901 , n75907 );
nand ( n75909 , n75025 , n75638 );
nand ( n75910 , n75908 , n75909 );
xor ( n75911 , n75900 , n75910 );
not ( n75912 , n60542 );
not ( n75913 , n59341 );
not ( n75914 , n54415 );
or ( n75915 , n75913 , n75914 );
nand ( n75916 , n66704 , n66983 );
nand ( n75917 , n75915 , n75916 );
not ( n75918 , n75917 );
or ( n75919 , n75912 , n75918 );
nand ( n75920 , n75577 , n70487 );
nand ( n75921 , n75919 , n75920 );
xor ( n75922 , n75911 , n75921 );
xor ( n75923 , n75890 , n75922 );
xor ( n75924 , n75923 , n75846 );
xor ( n75925 , n75924 , n75559 );
xor ( n75926 , n75923 , n75846 );
and ( n75927 , n75926 , n75559 );
and ( n75928 , n75923 , n75846 );
or ( n75929 , n75927 , n75928 );
xor ( n75930 , n75567 , n75852 );
xor ( n75931 , n75930 , n75609 );
xor ( n75932 , n75567 , n75852 );
and ( n75933 , n75932 , n75609 );
and ( n75934 , n75567 , n75852 );
or ( n75935 , n75933 , n75934 );
xor ( n75936 , n75885 , n75649 );
xor ( n75937 , n75936 , n75925 );
xor ( n75938 , n75885 , n75649 );
and ( n75939 , n75938 , n75925 );
and ( n75940 , n75885 , n75649 );
or ( n75941 , n75939 , n75940 );
xor ( n75942 , n75931 , n75655 );
xor ( n75943 , n75942 , n75661 );
xor ( n75944 , n75931 , n75655 );
and ( n75945 , n75944 , n75661 );
and ( n75946 , n75931 , n75655 );
or ( n75947 , n75945 , n75946 );
xor ( n75948 , n75937 , n75943 );
xor ( n75949 , n75948 , n75667 );
xor ( n75950 , n75937 , n75943 );
and ( n75951 , n75950 , n75667 );
and ( n75952 , n75937 , n75943 );
or ( n75953 , n75951 , n75952 );
xor ( n75954 , n75869 , n75870 );
and ( n75955 , n75954 , n75881 );
and ( n75956 , n75869 , n75870 );
or ( n75957 , n75955 , n75956 );
xor ( n75958 , n75900 , n75910 );
and ( n75959 , n75958 , n75921 );
and ( n75960 , n75900 , n75910 );
or ( n75961 , n75959 , n75960 );
xor ( n75962 , n75824 , n75834 );
and ( n75963 , n75962 , n75844 );
and ( n75964 , n75824 , n75834 );
or ( n75965 , n75963 , n75964 );
xor ( n75966 , n75791 , n75801 );
and ( n75967 , n75966 , n75812 );
and ( n75968 , n75791 , n75801 );
or ( n75969 , n75967 , n75968 );
xor ( n75970 , n75769 , n75779 );
and ( n75971 , n75970 , n75718 );
and ( n75972 , n75769 , n75779 );
or ( n75973 , n75971 , n75972 );
xor ( n75974 , n75446 , n75482 );
and ( n75975 , n75974 , n75677 );
and ( n75976 , n75446 , n75482 );
or ( n75977 , n75975 , n75976 );
xor ( n75978 , n75756 , n75882 );
and ( n75979 , n75978 , n75681 );
and ( n75980 , n75756 , n75882 );
or ( n75981 , n75979 , n75980 );
xor ( n75982 , n75685 , n75689 );
and ( n75983 , n75982 , n75922 );
and ( n75984 , n75685 , n75689 );
or ( n75985 , n75983 , n75984 );
not ( n75986 , n70964 );
not ( n75987 , n67072 );
not ( n75988 , n75987 );
not ( n75989 , n40691 );
or ( n75990 , n75988 , n75989 );
not ( n75991 , n71361 );
nand ( n75992 , n75991 , n71971 );
nand ( n75993 , n75990 , n75992 );
not ( n75994 , n75993 );
or ( n75995 , n75986 , n75994 );
nand ( n75996 , n65795 , n75713 );
nand ( n75997 , n75995 , n75996 );
not ( n75998 , n67061 );
not ( n75999 , n75728 );
or ( n76000 , n75998 , n75999 );
not ( n76001 , n64170 );
not ( n76002 , n70638 );
or ( n76003 , n76001 , n76002 );
not ( n76004 , n64170 );
nand ( n76005 , n53258 , n76004 );
nand ( n76006 , n76003 , n76005 );
nand ( n76007 , n76006 , n75427 );
nand ( n76008 , n76000 , n76007 );
xor ( n76009 , n75997 , n76008 );
not ( n76010 , n71099 );
not ( n76011 , n75865 );
or ( n76012 , n76010 , n76011 );
not ( n76013 , n55872 );
not ( n76014 , n63180 );
or ( n76015 , n76013 , n76014 );
not ( n76016 , n71371 );
nand ( n76017 , n70653 , n76016 );
nand ( n76018 , n76015 , n76017 );
nand ( n76019 , n76018 , n59984 );
nand ( n76020 , n76012 , n76019 );
xor ( n76021 , n76009 , n76020 );
xor ( n76022 , n75997 , n76008 );
and ( n76023 , n76022 , n76020 );
and ( n76024 , n75997 , n76008 );
or ( n76025 , n76023 , n76024 );
not ( n76026 , n56777 );
not ( n76027 , n75877 );
or ( n76028 , n76026 , n76027 );
not ( n76029 , n56786 );
not ( n76030 , n70661 );
or ( n76031 , n76029 , n76030 );
nand ( n76032 , n72217 , n69819 );
nand ( n76033 , n76031 , n76032 );
nand ( n76034 , n76033 , n60472 );
nand ( n76035 , n76028 , n76034 );
nand ( n76036 , n72846 , n41038 );
xor ( n76037 , n76035 , n76036 );
not ( n76038 , n72710 );
and ( n76039 , n73977 , n54791 );
not ( n76040 , n73977 );
and ( n76041 , n76040 , n57390 );
nor ( n76042 , n76039 , n76041 );
not ( n76043 , n76042 );
or ( n76044 , n76038 , n76043 );
nand ( n76045 , n75896 , n72961 );
nand ( n76046 , n76044 , n76045 );
xor ( n76047 , n76037 , n76046 );
xor ( n76048 , n76035 , n76036 );
and ( n76049 , n76048 , n76046 );
and ( n76050 , n76035 , n76036 );
or ( n76051 , n76049 , n76050 );
not ( n76052 , n53197 );
not ( n76053 , n75799 );
or ( n76054 , n76052 , n76053 );
not ( n76055 , n52114 );
not ( n76056 , n39333 );
or ( n76057 , n76055 , n76056 );
not ( n76058 , n73607 );
nand ( n76059 , n76058 , n69919 );
nand ( n76060 , n76057 , n76059 );
nand ( n76061 , n76060 , n51766 );
nand ( n76062 , n76054 , n76061 );
not ( n76063 , n52854 );
not ( n76064 , n75810 );
or ( n76065 , n76063 , n76064 );
not ( n76066 , n52841 );
not ( n76067 , n59891 );
or ( n76068 , n76066 , n76067 );
nand ( n76069 , n39056 , n53947 );
nand ( n76070 , n76068 , n76069 );
nand ( n76071 , n76070 , n53571 );
nand ( n76072 , n76065 , n76071 );
xor ( n76073 , n76062 , n76072 );
xor ( n76074 , n76073 , n75722 );
xor ( n76075 , n76074 , n75977 );
not ( n76076 , n72142 );
not ( n76077 , n75832 );
or ( n76078 , n76076 , n76077 );
not ( n76079 , n71395 );
not ( n76080 , n67040 );
or ( n76081 , n76079 , n76080 );
not ( n76082 , n74900 );
nand ( n76083 , n76082 , n54468 );
nand ( n76084 , n76081 , n76083 );
nand ( n76085 , n76084 , n54327 );
nand ( n76086 , n76078 , n76085 );
xor ( n76087 , n76086 , n75760 );
xor ( n76088 , n76087 , n75957 );
xor ( n76089 , n76075 , n76088 );
xor ( n76090 , n76074 , n75977 );
and ( n76091 , n76090 , n76088 );
and ( n76092 , n76074 , n75977 );
or ( n76093 , n76091 , n76092 );
xor ( n76094 , n75985 , n75981 );
xor ( n76095 , n76094 , n75850 );
xor ( n76096 , n75985 , n75981 );
and ( n76097 , n76096 , n75850 );
and ( n76098 , n75985 , n75981 );
or ( n76099 , n76097 , n76098 );
xor ( n76100 , n75961 , n76021 );
xor ( n76101 , n76100 , n76047 );
xor ( n76102 , n75965 , n75969 );
not ( n76103 , n61465 );
not ( n76104 , n58642 );
not ( n76105 , n71476 );
or ( n76106 , n76104 , n76105 );
nand ( n76107 , n59195 , n65183 );
nand ( n76108 , n76106 , n76107 );
not ( n76109 , n76108 );
or ( n76110 , n76103 , n76109 );
nand ( n76111 , n75906 , n75025 );
nand ( n76112 , n76110 , n76111 );
not ( n76113 , n70487 );
not ( n76114 , n75917 );
or ( n76115 , n76113 , n76114 );
and ( n76116 , n53289 , n59341 );
not ( n76117 , n53289 );
and ( n76118 , n76117 , n59340 );
or ( n76119 , n76116 , n76118 );
nand ( n76120 , n76119 , n75578 );
nand ( n76121 , n76115 , n76120 );
xor ( n76122 , n76112 , n76121 );
not ( n76123 , n70930 );
not ( n76124 , n70506 );
not ( n76125 , n52432 );
or ( n76126 , n76124 , n76125 );
nand ( n76127 , n72160 , n60286 );
nand ( n76128 , n76126 , n76127 );
not ( n76129 , n76128 );
or ( n76130 , n76123 , n76129 );
nand ( n76131 , n75822 , n70500 );
nand ( n76132 , n76130 , n76131 );
xor ( n76133 , n76122 , n76132 );
xor ( n76134 , n76102 , n76133 );
xor ( n76135 , n76101 , n76134 );
not ( n76136 , n52749 );
not ( n76137 , n75840 );
or ( n76138 , n76136 , n76137 );
nand ( n76139 , n52757 , n64190 );
nand ( n76140 , n76138 , n76139 );
not ( n76141 , n68603 );
not ( n76142 , n75775 );
or ( n76143 , n76141 , n76142 );
not ( n76144 , n55089 );
not ( n76145 , n67014 );
or ( n76146 , n76144 , n76145 );
not ( n76147 , n53596 );
not ( n76148 , n67014 );
nand ( n76149 , n76147 , n76148 );
nand ( n76150 , n76146 , n76149 );
nand ( n76151 , n76150 , n54364 );
nand ( n76152 , n76143 , n76151 );
xor ( n76153 , n76140 , n76152 );
not ( n76154 , n56355 );
not ( n76155 , n75787 );
or ( n76156 , n76154 , n76155 );
not ( n76157 , n53931 );
not ( n76158 , n69961 );
or ( n76159 , n76157 , n76158 );
nand ( n76160 , n69962 , n71053 );
nand ( n76161 , n76159 , n76160 );
nand ( n76162 , n76161 , n51533 );
nand ( n76163 , n76156 , n76162 );
xor ( n76164 , n76153 , n76163 );
xor ( n76165 , n76164 , n75973 );
not ( n76166 , n75753 );
not ( n76167 , n75750 );
or ( n76168 , n76166 , n76167 );
not ( n76169 , n61540 );
not ( n76170 , n52570 );
or ( n76171 , n76169 , n76170 );
nand ( n76172 , n51916 , n71307 );
nand ( n76173 , n76171 , n76172 );
nand ( n76174 , n76173 , n61558 );
nand ( n76175 , n76168 , n76174 );
not ( n76176 , n70183 );
and ( n76177 , n55120 , n68142 );
not ( n76178 , n55120 );
and ( n76179 , n76178 , n39847 );
or ( n76180 , n76177 , n76179 );
not ( n76181 , n76180 );
or ( n76182 , n76176 , n76181 );
nand ( n76183 , n75740 , n55144 );
nand ( n76184 , n76182 , n76183 );
xor ( n76185 , n76175 , n76184 );
not ( n76186 , n52151 );
not ( n76187 , n75765 );
or ( n76188 , n76186 , n76187 );
not ( n76189 , n57187 );
not ( n76190 , n72307 );
or ( n76191 , n76189 , n76190 );
nand ( n76192 , n71525 , n50946 );
nand ( n76193 , n76191 , n76192 );
nand ( n76194 , n76193 , n50922 );
nand ( n76195 , n76188 , n76194 );
xor ( n76196 , n76185 , n76195 );
xor ( n76197 , n76165 , n76196 );
xor ( n76198 , n76135 , n76197 );
xor ( n76199 , n76101 , n76134 );
and ( n76200 , n76199 , n76197 );
and ( n76201 , n76101 , n76134 );
or ( n76202 , n76200 , n76201 );
xor ( n76203 , n76089 , n75856 );
xor ( n76204 , n76203 , n75889 );
xor ( n76205 , n76089 , n75856 );
and ( n76206 , n76205 , n75889 );
and ( n76207 , n76089 , n75856 );
or ( n76208 , n76206 , n76207 );
xor ( n76209 , n76095 , n75929 );
xor ( n76210 , n76209 , n76198 );
xor ( n76211 , n76095 , n75929 );
and ( n76212 , n76211 , n76198 );
and ( n76213 , n76095 , n75929 );
or ( n76214 , n76212 , n76213 );
xor ( n76215 , n76204 , n75935 );
xor ( n76216 , n76215 , n75941 );
xor ( n76217 , n76204 , n75935 );
and ( n76218 , n76217 , n75941 );
and ( n76219 , n76204 , n75935 );
or ( n76220 , n76218 , n76219 );
xor ( n76221 , n76210 , n76216 );
xor ( n76222 , n76221 , n75947 );
xor ( n76223 , n76210 , n76216 );
and ( n76224 , n76223 , n75947 );
and ( n76225 , n76210 , n76216 );
or ( n76226 , n76224 , n76225 );
xor ( n76227 , n76112 , n76121 );
and ( n76228 , n76227 , n76132 );
and ( n76229 , n76112 , n76121 );
or ( n76230 , n76228 , n76229 );
xor ( n76231 , n76175 , n76184 );
and ( n76232 , n76231 , n76195 );
and ( n76233 , n76175 , n76184 );
or ( n76234 , n76232 , n76233 );
xor ( n76235 , n76062 , n76072 );
and ( n76236 , n76235 , n75722 );
and ( n76237 , n76062 , n76072 );
or ( n76238 , n76236 , n76237 );
xor ( n76239 , n76140 , n76152 );
and ( n76240 , n76239 , n76163 );
and ( n76241 , n76140 , n76152 );
or ( n76242 , n76240 , n76241 );
xor ( n76243 , n76086 , n75760 );
and ( n76244 , n76243 , n75957 );
and ( n76245 , n76086 , n75760 );
or ( n76246 , n76244 , n76245 );
xor ( n76247 , n75961 , n76021 );
and ( n76248 , n76247 , n76047 );
and ( n76249 , n75961 , n76021 );
or ( n76250 , n76248 , n76249 );
xor ( n76251 , n75965 , n75969 );
and ( n76252 , n76251 , n76133 );
and ( n76253 , n75965 , n75969 );
or ( n76254 , n76252 , n76253 );
xor ( n76255 , n76164 , n75973 );
and ( n76256 , n76255 , n76196 );
and ( n76257 , n76164 , n75973 );
or ( n76258 , n76256 , n76257 );
not ( n76259 , n59828 );
not ( n76260 , n59820 );
or ( n76261 , n76259 , n76260 );
nand ( n76262 , n76261 , n50306 );
and ( n76263 , n70889 , n66575 );
xor ( n76264 , n76262 , n76263 );
not ( n76265 , n71099 );
not ( n76266 , n76018 );
or ( n76267 , n76265 , n76266 );
not ( n76268 , n55872 );
not ( n76269 , n75162 );
or ( n76270 , n76268 , n76269 );
nand ( n76271 , n62618 , n71094 );
nand ( n76272 , n76270 , n76271 );
nand ( n76273 , n76272 , n59984 );
nand ( n76274 , n76267 , n76273 );
xor ( n76275 , n76264 , n76274 );
xor ( n76276 , n76262 , n76263 );
and ( n76277 , n76276 , n76274 );
and ( n76278 , n76262 , n76263 );
or ( n76279 , n76277 , n76278 );
not ( n76280 , n70964 );
not ( n76281 , n71971 );
not ( n76282 , n52286 );
or ( n76283 , n76281 , n76282 );
nand ( n76284 , n71093 , n64443 );
nand ( n76285 , n76283 , n76284 );
not ( n76286 , n76285 );
or ( n76287 , n76280 , n76286 );
nand ( n76288 , n75993 , n65795 );
nand ( n76289 , n76287 , n76288 );
not ( n76290 , n67068 );
not ( n76291 , n72083 );
not ( n76292 , n51602 );
or ( n76293 , n76291 , n76292 );
nand ( n76294 , n51601 , n76004 );
nand ( n76295 , n76293 , n76294 );
not ( n76296 , n76295 );
or ( n76297 , n76290 , n76296 );
nand ( n76298 , n76006 , n67061 );
nand ( n76299 , n76297 , n76298 );
xor ( n76300 , n76289 , n76299 );
not ( n76301 , n76036 );
xor ( n76302 , n76300 , n76301 );
xor ( n76303 , n76289 , n76299 );
and ( n76304 , n76303 , n76301 );
and ( n76305 , n76289 , n76299 );
or ( n76306 , n76304 , n76305 );
not ( n76307 , n70183 );
not ( n76308 , n55120 );
not ( n76309 , n65708 );
not ( n76310 , n76309 );
or ( n76311 , n76308 , n76310 );
nand ( n76312 , n71013 , n71409 );
nand ( n76313 , n76311 , n76312 );
not ( n76314 , n76313 );
or ( n76315 , n76307 , n76314 );
nand ( n76316 , n76180 , n55144 );
nand ( n76317 , n76315 , n76316 );
not ( n76318 , n52151 );
not ( n76319 , n76193 );
or ( n76320 , n76318 , n76319 );
not ( n76321 , n57187 );
not ( n76322 , n71876 );
or ( n76323 , n76321 , n76322 );
nand ( n76324 , n71875 , n67639 );
nand ( n76325 , n76323 , n76324 );
nand ( n76326 , n76325 , n50922 );
nand ( n76327 , n76320 , n76326 );
xor ( n76328 , n76317 , n76327 );
not ( n76329 , n72220 );
not ( n76330 , n52114 );
not ( n76331 , n71176 );
or ( n76332 , n76330 , n76331 );
nand ( n76333 , n39255 , n52113 );
nand ( n76334 , n76332 , n76333 );
not ( n76335 , n76334 );
or ( n76336 , n76329 , n76335 );
nand ( n76337 , n53197 , n76060 );
nand ( n76338 , n76336 , n76337 );
xor ( n76339 , n76328 , n76338 );
xor ( n76340 , n76339 , n76246 );
xor ( n76341 , n76340 , n76254 );
xor ( n76342 , n76339 , n76246 );
and ( n76343 , n76342 , n76254 );
and ( n76344 , n76339 , n76246 );
or ( n76345 , n76343 , n76344 );
xor ( n76346 , n76051 , n76230 );
xor ( n76347 , n76346 , n76302 );
xor ( n76348 , n76250 , n76347 );
not ( n76349 , n54327 );
and ( n76350 , n70627 , n39681 );
not ( n76351 , n70627 );
and ( n76352 , n76351 , n73428 );
nor ( n76353 , n76350 , n76352 );
not ( n76354 , n76353 );
or ( n76355 , n76349 , n76354 );
nand ( n76356 , n76084 , n72142 );
nand ( n76357 , n76355 , n76356 );
xor ( n76358 , n76357 , n76275 );
xor ( n76359 , n76358 , n76025 );
xor ( n76360 , n76348 , n76359 );
xor ( n76361 , n76250 , n76347 );
and ( n76362 , n76361 , n76359 );
and ( n76363 , n76250 , n76347 );
or ( n76364 , n76362 , n76363 );
not ( n76365 , n75578 );
not ( n76366 , n66985 );
not ( n76367 , n73291 );
or ( n76368 , n76366 , n76367 );
nand ( n76369 , n40226 , n59340 );
nand ( n76370 , n76368 , n76369 );
not ( n76371 , n76370 );
or ( n76372 , n76365 , n76371 );
nand ( n76373 , n70487 , n76119 );
nand ( n76374 , n76372 , n76373 );
not ( n76375 , n70930 );
not ( n76376 , n68878 );
not ( n76377 , n71767 );
or ( n76378 , n76376 , n76377 );
nand ( n76379 , n71770 , n60286 );
nand ( n76380 , n76378 , n76379 );
not ( n76381 , n76380 );
or ( n76382 , n76375 , n76381 );
nand ( n76383 , n76128 , n70500 );
nand ( n76384 , n76382 , n76383 );
xor ( n76385 , n76374 , n76384 );
not ( n76386 , n72484 );
not ( n76387 , n76173 );
or ( n76388 , n76386 , n76387 );
not ( n76389 , n61540 );
not ( n76390 , n66798 );
or ( n76391 , n76389 , n76390 );
nand ( n76392 , n40592 , n71307 );
nand ( n76393 , n76391 , n76392 );
nand ( n76394 , n76393 , n61558 );
nand ( n76395 , n76388 , n76394 );
xor ( n76396 , n76385 , n76395 );
not ( n76397 , n72185 );
not ( n76398 , n72589 );
not ( n76399 , n70290 );
or ( n76400 , n76398 , n76399 );
nand ( n76401 , n72607 , n72593 );
nand ( n76402 , n76400 , n76401 );
not ( n76403 , n76402 );
or ( n76404 , n76397 , n76403 );
nand ( n76405 , n76033 , n56777 );
nand ( n76406 , n76404 , n76405 );
not ( n76407 , n72182 );
not ( n76408 , n76042 );
or ( n76409 , n76407 , n76408 );
not ( n76410 , n67568 );
not ( n76411 , n73327 );
or ( n76412 , n76410 , n76411 );
nand ( n76413 , n71052 , n73307 );
nand ( n76414 , n76412 , n76413 );
nand ( n76415 , n76414 , n72710 );
nand ( n76416 , n76409 , n76415 );
xor ( n76417 , n76406 , n76416 );
not ( n76418 , n75025 );
not ( n76419 , n76108 );
or ( n76420 , n76418 , n76419 );
not ( n76421 , n65184 );
not ( n76422 , n62626 );
or ( n76423 , n76421 , n76422 );
buf ( n76424 , n69409 );
nand ( n76425 , n76424 , n62497 );
nand ( n76426 , n76423 , n76425 );
nand ( n76427 , n76426 , n71466 );
nand ( n76428 , n76420 , n76427 );
xor ( n76429 , n76417 , n76428 );
xor ( n76430 , n76396 , n76429 );
not ( n76431 , n52854 );
not ( n76432 , n76070 );
or ( n76433 , n76431 , n76432 );
not ( n76434 , n52841 );
not ( n76435 , n68652 );
or ( n76436 , n76434 , n76435 );
nand ( n76437 , n38499 , n53947 );
nand ( n76438 , n76436 , n76437 );
nand ( n76439 , n76438 , n52469 );
nand ( n76440 , n76433 , n76439 );
not ( n76441 , n53620 );
and ( n76442 , n55089 , n39575 );
not ( n76443 , n55089 );
not ( n76444 , n39575 );
and ( n76445 , n76443 , n76444 );
nor ( n76446 , n76442 , n76445 );
not ( n76447 , n76446 );
or ( n76448 , n76441 , n76447 );
nand ( n76449 , n76150 , n68603 );
nand ( n76450 , n76448 , n76449 );
xor ( n76451 , n76440 , n76450 );
not ( n76452 , n51533 );
not ( n76453 , n53931 );
buf ( n76454 , n68381 );
not ( n76455 , n76454 );
not ( n76456 , n76455 );
or ( n76457 , n76453 , n76456 );
nand ( n76458 , n76454 , n71053 );
nand ( n76459 , n76457 , n76458 );
not ( n76460 , n76459 );
or ( n76461 , n76452 , n76460 );
nand ( n76462 , n76161 , n72198 );
nand ( n76463 , n76461 , n76462 );
xor ( n76464 , n76451 , n76463 );
xor ( n76465 , n76430 , n76464 );
xor ( n76466 , n76258 , n76465 );
xor ( n76467 , n76234 , n76238 );
xor ( n76468 , n76467 , n76242 );
xor ( n76469 , n76466 , n76468 );
xor ( n76470 , n76258 , n76465 );
and ( n76471 , n76470 , n76468 );
and ( n76472 , n76258 , n76465 );
or ( n76473 , n76471 , n76472 );
xor ( n76474 , n76093 , n76341 );
xor ( n76475 , n76474 , n76360 );
xor ( n76476 , n76093 , n76341 );
and ( n76477 , n76476 , n76360 );
and ( n76478 , n76093 , n76341 );
or ( n76479 , n76477 , n76478 );
xor ( n76480 , n76099 , n76202 );
xor ( n76481 , n76480 , n76469 );
xor ( n76482 , n76099 , n76202 );
and ( n76483 , n76482 , n76469 );
and ( n76484 , n76099 , n76202 );
or ( n76485 , n76483 , n76484 );
xor ( n76486 , n76475 , n76208 );
xor ( n76487 , n76486 , n76214 );
xor ( n76488 , n76475 , n76208 );
and ( n76489 , n76488 , n76214 );
and ( n76490 , n76475 , n76208 );
or ( n76491 , n76489 , n76490 );
xor ( n76492 , n76481 , n76487 );
xor ( n76493 , n76492 , n76220 );
xor ( n76494 , n76481 , n76487 );
and ( n76495 , n76494 , n76220 );
and ( n76496 , n76481 , n76487 );
or ( n76497 , n76495 , n76496 );
xor ( n76498 , n76406 , n76416 );
and ( n76499 , n76498 , n76428 );
and ( n76500 , n76406 , n76416 );
or ( n76501 , n76499 , n76500 );
xor ( n76502 , n76374 , n76384 );
and ( n76503 , n76502 , n76395 );
and ( n76504 , n76374 , n76384 );
or ( n76505 , n76503 , n76504 );
xor ( n76506 , n76317 , n76327 );
and ( n76507 , n76506 , n76338 );
and ( n76508 , n76317 , n76327 );
or ( n76509 , n76507 , n76508 );
xor ( n76510 , n76440 , n76450 );
and ( n76511 , n76510 , n76463 );
and ( n76512 , n76440 , n76450 );
or ( n76513 , n76511 , n76512 );
xor ( n76514 , n76357 , n76275 );
and ( n76515 , n76514 , n76025 );
and ( n76516 , n76357 , n76275 );
or ( n76517 , n76515 , n76516 );
xor ( n76518 , n76051 , n76230 );
and ( n76519 , n76518 , n76302 );
and ( n76520 , n76051 , n76230 );
or ( n76521 , n76519 , n76520 );
xor ( n76522 , n76234 , n76238 );
and ( n76523 , n76522 , n76242 );
and ( n76524 , n76234 , n76238 );
or ( n76525 , n76523 , n76524 );
xor ( n76526 , n76396 , n76429 );
and ( n76527 , n76526 , n76464 );
and ( n76528 , n76396 , n76429 );
or ( n76529 , n76527 , n76528 );
not ( n76530 , n56777 );
not ( n76531 , n76402 );
or ( n76532 , n76530 , n76531 );
not ( n76533 , n56786 );
not ( n76534 , n63180 );
or ( n76535 , n76533 , n76534 );
nand ( n76536 , n72205 , n56785 );
nand ( n76537 , n76535 , n76536 );
nand ( n76538 , n76537 , n72185 );
nand ( n76539 , n76532 , n76538 );
not ( n76540 , n70964 );
xor ( n76541 , n66581 , n40736 );
not ( n76542 , n76541 );
or ( n76543 , n76540 , n76542 );
nand ( n76544 , n76285 , n65795 );
nand ( n76545 , n76543 , n76544 );
xor ( n76546 , n76539 , n76545 );
not ( n76547 , n72182 );
not ( n76548 , n76414 );
or ( n76549 , n76547 , n76548 );
not ( n76550 , n75343 );
not ( n76551 , n55630 );
or ( n76552 , n76550 , n76551 );
nand ( n76553 , n68980 , n73307 );
nand ( n76554 , n76552 , n76553 );
nand ( n76555 , n76554 , n72710 );
nand ( n76556 , n76549 , n76555 );
xor ( n76557 , n76546 , n76556 );
xor ( n76558 , n76539 , n76545 );
and ( n76559 , n76558 , n76556 );
and ( n76560 , n76539 , n76545 );
or ( n76561 , n76559 , n76560 );
not ( n76562 , n75025 );
not ( n76563 , n76426 );
or ( n76564 , n76562 , n76563 );
not ( n76565 , n65184 );
not ( n76566 , n68073 );
or ( n76567 , n76565 , n76566 );
nand ( n76568 , n68994 , n65187 );
nand ( n76569 , n76567 , n76568 );
nand ( n76570 , n76569 , n71466 );
nand ( n76571 , n76564 , n76570 );
not ( n76572 , n75578 );
not ( n76573 , n59341 );
not ( n76574 , n54811 );
or ( n76575 , n76573 , n76574 );
nand ( n76576 , n40364 , n70920 );
nand ( n76577 , n76575 , n76576 );
not ( n76578 , n76577 );
or ( n76579 , n76572 , n76578 );
nand ( n76580 , n76370 , n70487 );
nand ( n76581 , n76579 , n76580 );
xor ( n76582 , n76571 , n76581 );
not ( n76583 , n70500 );
not ( n76584 , n76380 );
or ( n76585 , n76583 , n76584 );
not ( n76586 , n66140 );
not ( n76587 , n53289 );
or ( n76588 , n76586 , n76587 );
nand ( n76589 , n54646 , n67084 );
nand ( n76590 , n76588 , n76589 );
nand ( n76591 , n76590 , n70930 );
nand ( n76592 , n76585 , n76591 );
xor ( n76593 , n76582 , n76592 );
xor ( n76594 , n76571 , n76581 );
and ( n76595 , n76594 , n76592 );
and ( n76596 , n76571 , n76581 );
or ( n76597 , n76595 , n76596 );
xor ( n76598 , n76306 , n76501 );
xor ( n76599 , n76598 , n76505 );
xor ( n76600 , n76521 , n76599 );
xor ( n76601 , n76600 , n76525 );
xor ( n76602 , n76521 , n76599 );
and ( n76603 , n76602 , n76525 );
and ( n76604 , n76521 , n76599 );
or ( n76605 , n76603 , n76604 );
not ( n76606 , n61558 );
not ( n76607 , n61540 );
not ( n76608 , n52432 );
or ( n76609 , n76607 , n76608 );
nand ( n76610 , n72160 , n61537 );
nand ( n76611 , n76609 , n76610 );
not ( n76612 , n76611 );
or ( n76613 , n76606 , n76612 );
nand ( n76614 , n76393 , n75753 );
nand ( n76615 , n76613 , n76614 );
not ( n76616 , n72083 );
not ( n76617 , n60138 );
or ( n76618 , n76616 , n76617 );
not ( n76619 , n40528 );
nand ( n76620 , n76619 , n76004 );
nand ( n76621 , n76618 , n76620 );
nand ( n76622 , n76621 , n75427 );
nand ( n76623 , n67061 , n76295 );
nand ( n76624 , n76622 , n76623 );
xor ( n76625 , n76615 , n76624 );
nand ( n76626 , n40691 , n71971 );
xor ( n76627 , n76625 , n76626 );
xor ( n76628 , n76627 , n76593 );
not ( n76629 , n68603 );
not ( n76630 , n76446 );
or ( n76631 , n76629 , n76630 );
not ( n76632 , n55089 );
not ( n76633 , n69072 );
or ( n76634 , n76632 , n76633 );
nand ( n76635 , n71547 , n72238 );
nand ( n76636 , n76634 , n76635 );
nand ( n76637 , n76636 , n53620 );
nand ( n76638 , n76631 , n76637 );
not ( n76639 , n52151 );
not ( n76640 , n76325 );
or ( n76641 , n76639 , n76640 );
nand ( n76642 , n50922 , n57187 );
nand ( n76643 , n76641 , n76642 );
xor ( n76644 , n76638 , n76643 );
not ( n76645 , n54316 );
not ( n76646 , n76353 );
or ( n76647 , n76645 , n76646 );
not ( n76648 , n70627 );
not ( n76649 , n67014 );
or ( n76650 , n76648 , n76649 );
nand ( n76651 , n76148 , n54302 );
nand ( n76652 , n76650 , n76651 );
nand ( n76653 , n76652 , n54327 );
nand ( n76654 , n76647 , n76653 );
xor ( n76655 , n76644 , n76654 );
xor ( n76656 , n76628 , n76655 );
xor ( n76657 , n76656 , n76529 );
xor ( n76658 , n76557 , n76509 );
xor ( n76659 , n76658 , n76513 );
xor ( n76660 , n76657 , n76659 );
xor ( n76661 , n76656 , n76529 );
and ( n76662 , n76661 , n76659 );
and ( n76663 , n76656 , n76529 );
or ( n76664 , n76662 , n76663 );
xor ( n76665 , n76364 , n76345 );
not ( n76666 , n59984 );
not ( n76667 , n71371 );
not ( n76668 , n71418 );
or ( n76669 , n76667 , n76668 );
nand ( n76670 , n39847 , n76016 );
nand ( n76671 , n76669 , n76670 );
not ( n76672 , n76671 );
or ( n76673 , n76666 , n76672 );
nand ( n76674 , n76272 , n71099 );
nand ( n76675 , n76673 , n76674 );
not ( n76676 , n72198 );
not ( n76677 , n76459 );
or ( n76678 , n76676 , n76677 );
not ( n76679 , n53931 );
not ( n76680 , n72307 );
or ( n76681 , n76679 , n76680 );
nand ( n76682 , n42556 , n71053 );
nand ( n76683 , n76681 , n76682 );
nand ( n76684 , n76683 , n51533 );
nand ( n76685 , n76678 , n76684 );
xor ( n76686 , n76675 , n76685 );
not ( n76687 , n52469 );
not ( n76688 , n69458 );
not ( n76689 , n60855 );
or ( n76690 , n76688 , n76689 );
nand ( n76691 , n39332 , n55104 );
nand ( n76692 , n76690 , n76691 );
not ( n76693 , n76692 );
or ( n76694 , n76687 , n76693 );
nand ( n76695 , n76438 , n52854 );
nand ( n76696 , n76694 , n76695 );
xor ( n76697 , n76686 , n76696 );
not ( n76698 , n53197 );
not ( n76699 , n76334 );
or ( n76700 , n76698 , n76699 );
not ( n76701 , n73607 );
not ( n76702 , n69961 );
or ( n76703 , n76701 , n76702 );
nand ( n76704 , n72998 , n52110 );
nand ( n76705 , n76703 , n76704 );
nand ( n76706 , n76705 , n72220 );
nand ( n76707 , n76700 , n76706 );
not ( n76708 , n70193 );
not ( n76709 , n76313 );
or ( n76710 , n76708 , n76709 );
not ( n76711 , n55120 );
not ( n76712 , n74900 );
or ( n76713 , n76711 , n76712 );
not ( n76714 , n72919 );
nand ( n76715 , n75548 , n76714 );
nand ( n76716 , n76713 , n76715 );
nand ( n76717 , n76716 , n70183 );
nand ( n76718 , n76710 , n76717 );
xor ( n76719 , n76707 , n76718 );
xor ( n76720 , n76719 , n76279 );
xor ( n76721 , n76697 , n76720 );
xor ( n76722 , n76721 , n76517 );
xor ( n76723 , n76665 , n76722 );
xor ( n76724 , n76364 , n76345 );
and ( n76725 , n76724 , n76722 );
and ( n76726 , n76364 , n76345 );
or ( n76727 , n76725 , n76726 );
xor ( n76728 , n76601 , n76473 );
xor ( n76729 , n76728 , n76660 );
xor ( n76730 , n76601 , n76473 );
and ( n76731 , n76730 , n76660 );
and ( n76732 , n76601 , n76473 );
or ( n76733 , n76731 , n76732 );
xor ( n76734 , n76723 , n76479 );
xor ( n76735 , n76734 , n76729 );
xor ( n76736 , n76723 , n76479 );
and ( n76737 , n76736 , n76729 );
and ( n76738 , n76723 , n76479 );
or ( n76739 , n76737 , n76738 );
xor ( n76740 , n76485 , n76735 );
xor ( n76741 , n76740 , n76491 );
xor ( n76742 , n76485 , n76735 );
and ( n76743 , n76742 , n76491 );
and ( n76744 , n76485 , n76735 );
or ( n76745 , n76743 , n76744 );
xor ( n76746 , n76615 , n76624 );
and ( n76747 , n76746 , n76626 );
and ( n76748 , n76615 , n76624 );
or ( n76749 , n76747 , n76748 );
xor ( n76750 , n76675 , n76685 );
and ( n76751 , n76750 , n76696 );
and ( n76752 , n76675 , n76685 );
or ( n76753 , n76751 , n76752 );
xor ( n76754 , n76638 , n76643 );
and ( n76755 , n76754 , n76654 );
and ( n76756 , n76638 , n76643 );
or ( n76757 , n76755 , n76756 );
xor ( n76758 , n76707 , n76718 );
and ( n76759 , n76758 , n76279 );
and ( n76760 , n76707 , n76718 );
or ( n76761 , n76759 , n76760 );
xor ( n76762 , n76306 , n76501 );
and ( n76763 , n76762 , n76505 );
and ( n76764 , n76306 , n76501 );
or ( n76765 , n76763 , n76764 );
xor ( n76766 , n76557 , n76509 );
and ( n76767 , n76766 , n76513 );
and ( n76768 , n76557 , n76509 );
or ( n76769 , n76767 , n76768 );
xor ( n76770 , n76627 , n76593 );
and ( n76771 , n76770 , n76655 );
and ( n76772 , n76627 , n76593 );
or ( n76773 , n76771 , n76772 );
xor ( n76774 , n76697 , n76720 );
and ( n76775 , n76774 , n76517 );
and ( n76776 , n76697 , n76720 );
or ( n76777 , n76775 , n76776 );
not ( n76778 , n50922 );
not ( n76779 , n76778 );
not ( n76780 , n54692 );
or ( n76781 , n76779 , n76780 );
nand ( n76782 , n76781 , n57187 );
not ( n76783 , n56777 );
not ( n76784 , n76537 );
or ( n76785 , n76783 , n76784 );
not ( n76786 , n72593 );
not ( n76787 , n76786 );
not ( n76788 , n59651 );
or ( n76789 , n76787 , n76788 );
nand ( n76790 , n75161 , n72593 );
nand ( n76791 , n76789 , n76790 );
nand ( n76792 , n76791 , n60472 );
nand ( n76793 , n76785 , n76792 );
xor ( n76794 , n76782 , n76793 );
not ( n76795 , n70964 );
xor ( n76796 , n66155 , n69442 );
not ( n76797 , n76796 );
or ( n76798 , n76795 , n76797 );
nand ( n76799 , n76541 , n71960 );
nand ( n76800 , n76798 , n76799 );
xor ( n76801 , n76794 , n76800 );
xor ( n76802 , n76782 , n76793 );
and ( n76803 , n76802 , n76800 );
and ( n76804 , n76782 , n76793 );
or ( n76805 , n76803 , n76804 );
and ( n76806 , n71093 , n66581 );
not ( n76807 , n72710 );
not ( n76808 , n67568 );
not ( n76809 , n70290 );
or ( n76810 , n76808 , n76809 );
not ( n76811 , n67568 );
nand ( n76812 , n67721 , n76811 );
nand ( n76813 , n76810 , n76812 );
not ( n76814 , n76813 );
or ( n76815 , n76807 , n76814 );
nand ( n76816 , n76554 , n72182 );
nand ( n76817 , n76815 , n76816 );
xor ( n76818 , n76806 , n76817 );
not ( n76819 , n71466 );
not ( n76820 , n65184 );
not ( n76821 , n40382 );
not ( n76822 , n76821 );
or ( n76823 , n76820 , n76822 );
nand ( n76824 , n71052 , n62497 );
nand ( n76825 , n76823 , n76824 );
not ( n76826 , n76825 );
or ( n76827 , n76819 , n76826 );
not ( n76828 , n71689 );
nand ( n76829 , n76569 , n76828 );
nand ( n76830 , n76827 , n76829 );
xor ( n76831 , n76818 , n76830 );
xor ( n76832 , n76806 , n76817 );
and ( n76833 , n76832 , n76830 );
and ( n76834 , n76806 , n76817 );
or ( n76835 , n76833 , n76834 );
xor ( n76836 , n76761 , n76769 );
xor ( n76837 , n76561 , n76597 );
xor ( n76838 , n76837 , n76801 );
xor ( n76839 , n76836 , n76838 );
xor ( n76840 , n76761 , n76769 );
and ( n76841 , n76840 , n76838 );
and ( n76842 , n76761 , n76769 );
or ( n76843 , n76841 , n76842 );
not ( n76844 , n60542 );
and ( n76845 , n66983 , n54402 );
not ( n76846 , n66983 );
and ( n76847 , n76846 , n69409 );
nor ( n76848 , n76845 , n76847 );
not ( n76849 , n76848 );
or ( n76850 , n76844 , n76849 );
nand ( n76851 , n76577 , n72131 );
nand ( n76852 , n76850 , n76851 );
not ( n76853 , n70930 );
not ( n76854 , n68878 );
not ( n76855 , n53661 );
or ( n76856 , n76854 , n76855 );
nand ( n76857 , n40226 , n67084 );
nand ( n76858 , n76856 , n76857 );
not ( n76859 , n76858 );
or ( n76860 , n76853 , n76859 );
nand ( n76861 , n66136 , n76590 );
nand ( n76862 , n76860 , n76861 );
xor ( n76863 , n76852 , n76862 );
not ( n76864 , n61558 );
not ( n76865 , n71309 );
not ( n76866 , n54415 );
or ( n76867 , n76865 , n76866 );
nand ( n76868 , n66704 , n75748 );
nand ( n76869 , n76867 , n76868 );
not ( n76870 , n76869 );
or ( n76871 , n76864 , n76870 );
nand ( n76872 , n76611 , n75753 );
nand ( n76873 , n76871 , n76872 );
xor ( n76874 , n76863 , n76873 );
xor ( n76875 , n76874 , n76831 );
not ( n76876 , n76652 );
not ( n76877 , n54316 );
or ( n76878 , n76876 , n76877 );
and ( n76879 , n54468 , n68667 );
not ( n76880 , n54468 );
and ( n76881 , n76880 , n74059 );
or ( n76882 , n76879 , n76881 );
nand ( n76883 , n76882 , n54327 );
nand ( n76884 , n76878 , n76883 );
not ( n76885 , n53197 );
not ( n76886 , n76705 );
or ( n76887 , n76885 , n76886 );
and ( n76888 , n73607 , n76454 );
not ( n76889 , n73607 );
and ( n76890 , n76889 , n42399 );
nor ( n76891 , n76888 , n76890 );
nand ( n76892 , n76891 , n72220 );
nand ( n76893 , n76887 , n76892 );
xor ( n76894 , n76884 , n76893 );
not ( n76895 , n70193 );
not ( n76896 , n76716 );
or ( n76897 , n76895 , n76896 );
not ( n76898 , n72919 );
not ( n76899 , n74673 );
or ( n76900 , n76898 , n76899 );
nand ( n76901 , n58485 , n71409 );
nand ( n76902 , n76900 , n76901 );
nand ( n76903 , n76902 , n70183 );
nand ( n76904 , n76897 , n76903 );
xor ( n76905 , n76894 , n76904 );
xor ( n76906 , n76875 , n76905 );
xor ( n76907 , n76773 , n76906 );
xor ( n76908 , n76749 , n76753 );
xor ( n76909 , n76908 , n76757 );
xor ( n76910 , n76907 , n76909 );
xor ( n76911 , n76773 , n76906 );
and ( n76912 , n76911 , n76909 );
and ( n76913 , n76773 , n76906 );
or ( n76914 , n76912 , n76913 );
not ( n76915 , n75427 );
not ( n76916 , n72083 );
not ( n76917 , n66798 );
or ( n76918 , n76916 , n76917 );
nand ( n76919 , n40592 , n76004 );
nand ( n76920 , n76918 , n76919 );
not ( n76921 , n76920 );
or ( n76922 , n76915 , n76921 );
nand ( n76923 , n76621 , n67061 );
nand ( n76924 , n76922 , n76923 );
not ( n76925 , n71099 );
not ( n76926 , n76671 );
or ( n76927 , n76925 , n76926 );
nand ( n76928 , n71863 , n76016 );
not ( n76929 , n76928 );
not ( n76930 , n73271 );
nand ( n76931 , n76930 , n55872 );
not ( n76932 , n76931 );
or ( n76933 , n76929 , n76932 );
nand ( n76934 , n76933 , n59984 );
nand ( n76935 , n76927 , n76934 );
xor ( n76936 , n76924 , n76935 );
not ( n76937 , n72198 );
not ( n76938 , n76683 );
or ( n76939 , n76937 , n76938 );
and ( n76940 , n71053 , n71875 );
not ( n76941 , n71053 );
and ( n76942 , n76941 , n71876 );
nor ( n76943 , n76940 , n76942 );
not ( n76944 , n76943 );
nand ( n76945 , n76944 , n51533 );
nand ( n76946 , n76939 , n76945 );
xor ( n76947 , n76936 , n76946 );
not ( n76948 , n52854 );
not ( n76949 , n76692 );
or ( n76950 , n76948 , n76949 );
not ( n76951 , n69458 );
not ( n76952 , n71176 );
or ( n76953 , n76951 , n76952 );
nand ( n76954 , n69530 , n55104 );
nand ( n76955 , n76953 , n76954 );
nand ( n76956 , n76955 , n53571 );
nand ( n76957 , n76950 , n76956 );
not ( n76958 , n76626 );
xor ( n76959 , n76957 , n76958 );
not ( n76960 , n54364 );
not ( n76961 , n53596 );
not ( n76962 , n62394 );
or ( n76963 , n76961 , n76962 );
nand ( n76964 , n38499 , n72238 );
nand ( n76965 , n76963 , n76964 );
not ( n76966 , n76965 );
or ( n76967 , n76960 , n76966 );
nand ( n76968 , n76636 , n68603 );
nand ( n76969 , n76967 , n76968 );
xor ( n76970 , n76959 , n76969 );
xor ( n76971 , n76947 , n76970 );
xor ( n76972 , n76971 , n76765 );
xor ( n76973 , n76972 , n76777 );
xor ( n76974 , n76973 , n76605 );
xor ( n76975 , n76972 , n76777 );
and ( n76976 , n76975 , n76605 );
and ( n76977 , n76972 , n76777 );
or ( n76978 , n76976 , n76977 );
xor ( n76979 , n76839 , n76664 );
xor ( n76980 , n76979 , n76910 );
xor ( n76981 , n76839 , n76664 );
and ( n76982 , n76981 , n76910 );
and ( n76983 , n76839 , n76664 );
or ( n76984 , n76982 , n76983 );
xor ( n76985 , n76727 , n76974 );
xor ( n76986 , n76985 , n76980 );
xor ( n76987 , n76727 , n76974 );
and ( n76988 , n76987 , n76980 );
and ( n76989 , n76727 , n76974 );
or ( n76990 , n76988 , n76989 );
xor ( n76991 , n76733 , n76986 );
xor ( n76992 , n76991 , n76739 );
xor ( n76993 , n76733 , n76986 );
and ( n76994 , n76993 , n76739 );
and ( n76995 , n76733 , n76986 );
or ( n76996 , n76994 , n76995 );
xor ( n76997 , n76852 , n76862 );
and ( n76998 , n76997 , n76873 );
and ( n76999 , n76852 , n76862 );
or ( n77000 , n76998 , n76999 );
xor ( n77001 , n76924 , n76935 );
and ( n77002 , n77001 , n76946 );
and ( n77003 , n76924 , n76935 );
or ( n77004 , n77002 , n77003 );
xor ( n77005 , n76957 , n76958 );
and ( n77006 , n77005 , n76969 );
and ( n77007 , n76957 , n76958 );
or ( n77008 , n77006 , n77007 );
xor ( n77009 , n76884 , n76893 );
and ( n77010 , n77009 , n76904 );
and ( n77011 , n76884 , n76893 );
or ( n77012 , n77010 , n77011 );
xor ( n77013 , n76561 , n76597 );
and ( n77014 , n77013 , n76801 );
and ( n77015 , n76561 , n76597 );
or ( n77016 , n77014 , n77015 );
xor ( n77017 , n76749 , n76753 );
and ( n77018 , n77017 , n76757 );
and ( n77019 , n76749 , n76753 );
or ( n77020 , n77018 , n77019 );
xor ( n77021 , n76874 , n76831 );
and ( n77022 , n77021 , n76905 );
and ( n77023 , n76874 , n76831 );
or ( n77024 , n77022 , n77023 );
xor ( n77025 , n76947 , n76970 );
and ( n77026 , n77025 , n76765 );
and ( n77027 , n76947 , n76970 );
or ( n77028 , n77026 , n77027 );
not ( n77029 , n76828 );
not ( n77030 , n76825 );
or ( n77031 , n77029 , n77030 );
not ( n77032 , n62496 );
not ( n77033 , n71442 );
or ( n77034 , n77032 , n77033 );
nand ( n77035 , n72217 , n66652 );
nand ( n77036 , n77034 , n77035 );
nand ( n77037 , n77036 , n71466 );
nand ( n77038 , n77031 , n77037 );
and ( n77039 , n66581 , n40736 );
xor ( n77040 , n77038 , n77039 );
not ( n77041 , n70487 );
not ( n77042 , n76848 );
or ( n77043 , n77041 , n77042 );
not ( n77044 , n72464 );
not ( n77045 , n68991 );
or ( n77046 , n77044 , n77045 );
nand ( n77047 , n68994 , n66983 );
nand ( n77048 , n77046 , n77047 );
nand ( n77049 , n77048 , n75578 );
nand ( n77050 , n77043 , n77049 );
xor ( n77051 , n77040 , n77050 );
xor ( n77052 , n77038 , n77039 );
and ( n77053 , n77052 , n77050 );
and ( n77054 , n77038 , n77039 );
or ( n77055 , n77053 , n77054 );
not ( n77056 , n66136 );
not ( n77057 , n76858 );
or ( n77058 , n77056 , n77057 );
not ( n77059 , n68878 );
not ( n77060 , n59194 );
or ( n77061 , n77059 , n77060 );
nand ( n77062 , n63204 , n72477 );
nand ( n77063 , n77061 , n77062 );
nand ( n77064 , n70930 , n77063 );
nand ( n77065 , n77058 , n77064 );
not ( n77066 , n72484 );
not ( n77067 , n76869 );
or ( n77068 , n77066 , n77067 );
not ( n77069 , n61540 );
not ( n77070 , n56476 );
or ( n77071 , n77069 , n77070 );
nand ( n77072 , n54646 , n75748 );
nand ( n77073 , n77071 , n77072 );
nand ( n77074 , n61558 , n77073 );
nand ( n77075 , n77068 , n77074 );
xor ( n77076 , n77065 , n77075 );
buf ( n77077 , n67061 );
not ( n77078 , n77077 );
not ( n77079 , n76920 );
or ( n77080 , n77078 , n77079 );
not ( n77081 , n64170 );
not ( n77082 , n52432 );
or ( n77083 , n77081 , n77082 );
nand ( n77084 , n72160 , n66089 );
nand ( n77085 , n77083 , n77084 );
nand ( n77086 , n77085 , n67068 );
nand ( n77087 , n77080 , n77086 );
xor ( n77088 , n77076 , n77087 );
xor ( n77089 , n77065 , n77075 );
and ( n77090 , n77089 , n77087 );
and ( n77091 , n77065 , n77075 );
or ( n77092 , n77090 , n77091 );
xor ( n77093 , n77000 , n77004 );
xor ( n77094 , n77093 , n77008 );
xor ( n77095 , n77012 , n77088 );
xor ( n77096 , n77095 , n77051 );
xor ( n77097 , n77094 , n77096 );
xor ( n77098 , n77097 , n77024 );
xor ( n77099 , n77094 , n77096 );
and ( n77100 , n77099 , n77024 );
and ( n77101 , n77094 , n77096 );
or ( n77102 , n77100 , n77101 );
not ( n77103 , n55144 );
not ( n77104 , n76902 );
or ( n77105 , n77103 , n77104 );
not ( n77106 , n55120 );
not ( n77107 , n67014 );
or ( n77108 , n77106 , n77107 );
nand ( n77109 , n71567 , n71409 );
nand ( n77110 , n77108 , n77109 );
nand ( n77111 , n77110 , n70183 );
nand ( n77112 , n77105 , n77111 );
not ( n77113 , n52854 );
not ( n77114 , n76955 );
or ( n77115 , n77113 , n77114 );
not ( n77116 , n69458 );
not ( n77117 , n69961 );
or ( n77118 , n77116 , n77117 );
nand ( n77119 , n69962 , n55104 );
nand ( n77120 , n77118 , n77119 );
nand ( n77121 , n52469 , n77120 );
nand ( n77122 , n77115 , n77121 );
xor ( n77123 , n77112 , n77122 );
not ( n77124 , n71099 );
nand ( n77125 , n76928 , n76931 );
not ( n77126 , n77125 );
or ( n77127 , n77124 , n77126 );
not ( n77128 , n69695 );
not ( n77129 , n59914 );
or ( n77130 , n77128 , n77129 );
nand ( n77131 , n59913 , n76016 );
nand ( n77132 , n77130 , n77131 );
nand ( n77133 , n77132 , n55458 );
nand ( n77134 , n77127 , n77133 );
xor ( n77135 , n77123 , n77134 );
not ( n77136 , n71960 );
not ( n77137 , n76796 );
or ( n77138 , n77136 , n77137 );
xor ( n77139 , n72846 , n40529 );
nand ( n77140 , n70964 , n77139 );
nand ( n77141 , n77138 , n77140 );
not ( n77142 , n72185 );
not ( n77143 , n72589 );
not ( n77144 , n71418 );
or ( n77145 , n77143 , n77144 );
nand ( n77146 , n72298 , n72593 );
nand ( n77147 , n77145 , n77146 );
not ( n77148 , n77147 );
or ( n77149 , n77142 , n77148 );
nand ( n77150 , n76791 , n56777 );
nand ( n77151 , n77149 , n77150 );
xor ( n77152 , n77141 , n77151 );
not ( n77153 , n53197 );
not ( n77154 , n76891 );
or ( n77155 , n77153 , n77154 );
not ( n77156 , n68931 );
not ( n77157 , n67269 );
or ( n77158 , n77156 , n77157 );
nand ( n77159 , n42555 , n52110 );
nand ( n77160 , n77158 , n77159 );
nand ( n77161 , n77160 , n72220 );
nand ( n77162 , n77155 , n77161 );
xor ( n77163 , n77152 , n77162 );
xor ( n77164 , n77135 , n77163 );
not ( n77165 , n68603 );
not ( n77166 , n76965 );
or ( n77167 , n77165 , n77166 );
not ( n77168 , n55089 );
not ( n77169 , n39333 );
or ( n77170 , n77168 , n77169 );
not ( n77171 , n39331 );
nand ( n77172 , n77171 , n72238 );
nand ( n77173 , n77170 , n77172 );
nand ( n77174 , n77173 , n53620 );
nand ( n77175 , n77167 , n77174 );
not ( n77176 , n54327 );
not ( n77177 , n54298 );
not ( n77178 , n69072 );
or ( n77179 , n77177 , n77178 );
nand ( n77180 , n39056 , n54302 );
nand ( n77181 , n77179 , n77180 );
not ( n77182 , n77181 );
or ( n77183 , n77176 , n77182 );
nand ( n77184 , n76882 , n54316 );
nand ( n77185 , n77183 , n77184 );
xor ( n77186 , n77175 , n77185 );
or ( n77187 , n76943 , n72197 );
or ( n77188 , n53927 , n71053 );
nand ( n77189 , n77187 , n77188 );
xor ( n77190 , n77186 , n77189 );
xor ( n77191 , n77164 , n77190 );
xor ( n77192 , n77028 , n77191 );
xor ( n77193 , n77192 , n76843 );
xor ( n77194 , n77028 , n77191 );
and ( n77195 , n77194 , n76843 );
and ( n77196 , n77028 , n77191 );
or ( n77197 , n77195 , n77196 );
not ( n77198 , n72182 );
not ( n77199 , n76813 );
or ( n77200 , n77198 , n77199 );
not ( n77201 , n73977 );
not ( n77202 , n67193 );
or ( n77203 , n77201 , n77202 );
nand ( n77204 , n67196 , n66963 );
nand ( n77205 , n77203 , n77204 );
nand ( n77206 , n77205 , n72710 );
nand ( n77207 , n77200 , n77206 );
not ( n77208 , n77207 );
xor ( n77209 , n77208 , n76805 );
xor ( n77210 , n77209 , n76835 );
xor ( n77211 , n77020 , n77210 );
xor ( n77212 , n77211 , n77016 );
xor ( n77213 , n76914 , n77212 );
xor ( n77214 , n77213 , n77098 );
xor ( n77215 , n76914 , n77212 );
and ( n77216 , n77215 , n77098 );
and ( n77217 , n76914 , n77212 );
or ( n77218 , n77216 , n77217 );
xor ( n77219 , n77193 , n76978 );
xor ( n77220 , n77219 , n76984 );
xor ( n77221 , n77193 , n76978 );
and ( n77222 , n77221 , n76984 );
and ( n77223 , n77193 , n76978 );
or ( n77224 , n77222 , n77223 );
xor ( n77225 , n77214 , n77220 );
xor ( n77226 , n77225 , n76990 );
xor ( n77227 , n77214 , n77220 );
and ( n77228 , n77227 , n76990 );
and ( n77229 , n77214 , n77220 );
or ( n77230 , n77228 , n77229 );
xor ( n77231 , n77141 , n77151 );
and ( n77232 , n77231 , n77162 );
and ( n77233 , n77141 , n77151 );
or ( n77234 , n77232 , n77233 );
xor ( n77235 , n77175 , n77185 );
and ( n77236 , n77235 , n77189 );
and ( n77237 , n77175 , n77185 );
or ( n77238 , n77236 , n77237 );
xor ( n77239 , n77112 , n77122 );
and ( n77240 , n77239 , n77134 );
and ( n77241 , n77112 , n77122 );
or ( n77242 , n77240 , n77241 );
xor ( n77243 , n77208 , n76805 );
and ( n77244 , n77243 , n76835 );
and ( n77245 , n77208 , n76805 );
or ( n77246 , n77244 , n77245 );
xor ( n77247 , n77000 , n77004 );
and ( n77248 , n77247 , n77008 );
and ( n77249 , n77000 , n77004 );
or ( n77250 , n77248 , n77249 );
xor ( n77251 , n77012 , n77088 );
and ( n77252 , n77251 , n77051 );
and ( n77253 , n77012 , n77088 );
or ( n77254 , n77252 , n77253 );
xor ( n77255 , n77135 , n77163 );
and ( n77256 , n77255 , n77190 );
and ( n77257 , n77135 , n77163 );
or ( n77258 , n77256 , n77257 );
xor ( n77259 , n77020 , n77210 );
and ( n77260 , n77259 , n77016 );
and ( n77261 , n77020 , n77210 );
or ( n77262 , n77260 , n77261 );
not ( n77263 , n53927 );
not ( n77264 , n65111 );
or ( n77265 , n77263 , n77264 );
nand ( n77266 , n77265 , n53931 );
not ( n77267 , n72961 );
not ( n77268 , n77205 );
or ( n77269 , n77267 , n77268 );
not ( n77270 , n75343 );
not ( n77271 , n59651 );
or ( n77272 , n77270 , n77271 );
nand ( n77273 , n59654 , n76811 );
nand ( n77274 , n77272 , n77273 );
nand ( n77275 , n77274 , n72710 );
nand ( n77276 , n77269 , n77275 );
xor ( n77277 , n77266 , n77276 );
and ( n77278 , n66155 , n69442 );
xor ( n77279 , n77277 , n77278 );
xor ( n77280 , n77266 , n77276 );
and ( n77281 , n77280 , n77278 );
and ( n77282 , n77266 , n77276 );
or ( n77283 , n77281 , n77282 );
not ( n77284 , n61465 );
not ( n77285 , n58642 );
not ( n77286 , n70290 );
or ( n77287 , n77285 , n77286 );
nand ( n77288 , n40514 , n66652 );
nand ( n77289 , n77287 , n77288 );
not ( n77290 , n77289 );
or ( n77291 , n77284 , n77290 );
nand ( n77292 , n77036 , n76828 );
nand ( n77293 , n77291 , n77292 );
not ( n77294 , n75578 );
not ( n77295 , n72464 );
not ( n77296 , n76821 );
or ( n77297 , n77295 , n77296 );
nand ( n77298 , n71829 , n66983 );
nand ( n77299 , n77297 , n77298 );
not ( n77300 , n77299 );
or ( n77301 , n77294 , n77300 );
nand ( n77302 , n77048 , n70487 );
nand ( n77303 , n77301 , n77302 );
xor ( n77304 , n77293 , n77303 );
not ( n77305 , n70930 );
not ( n77306 , n68878 );
not ( n77307 , n54402 );
or ( n77308 , n77306 , n77307 );
nand ( n77309 , n71067 , n72477 );
nand ( n77310 , n77308 , n77309 );
not ( n77311 , n77310 );
or ( n77312 , n77305 , n77311 );
nand ( n77313 , n77063 , n70500 );
nand ( n77314 , n77312 , n77313 );
xor ( n77315 , n77304 , n77314 );
xor ( n77316 , n77293 , n77303 );
and ( n77317 , n77316 , n77314 );
and ( n77318 , n77293 , n77303 );
or ( n77319 , n77317 , n77318 );
xor ( n77320 , n77250 , n77258 );
xor ( n77321 , n77092 , n77279 );
xor ( n77322 , n77321 , n77234 );
xor ( n77323 , n77320 , n77322 );
xor ( n77324 , n77250 , n77258 );
and ( n77325 , n77324 , n77322 );
and ( n77326 , n77250 , n77258 );
or ( n77327 , n77325 , n77326 );
xor ( n77328 , n77238 , n77242 );
not ( n77329 , n61558 );
not ( n77330 , n61540 );
not ( n77331 , n72544 );
or ( n77332 , n77330 , n77331 );
not ( n77333 , n71309 );
nand ( n77334 , n40226 , n77333 );
nand ( n77335 , n77332 , n77334 );
not ( n77336 , n77335 );
or ( n77337 , n77329 , n77336 );
nand ( n77338 , n72810 , n77073 );
nand ( n77339 , n77337 , n77338 );
not ( n77340 , n67068 );
not ( n77341 , n72083 );
not ( n77342 , n71767 );
or ( n77343 , n77341 , n77342 );
not ( n77344 , n72083 );
nand ( n77345 , n71770 , n77344 );
nand ( n77346 , n77343 , n77345 );
not ( n77347 , n77346 );
or ( n77348 , n77340 , n77347 );
nand ( n77349 , n77085 , n67061 );
nand ( n77350 , n77348 , n77349 );
xor ( n77351 , n77339 , n77350 );
not ( n77352 , n71960 );
not ( n77353 , n77139 );
or ( n77354 , n77352 , n77353 );
xor ( n77355 , n66155 , n74581 );
nand ( n77356 , n77355 , n70964 );
nand ( n77357 , n77354 , n77356 );
xor ( n77358 , n77351 , n77357 );
xor ( n77359 , n77328 , n77358 );
not ( n77360 , n77181 );
not ( n77361 , n54316 );
or ( n77362 , n77360 , n77361 );
not ( n77363 , n54298 );
not ( n77364 , n68652 );
or ( n77365 , n77363 , n77364 );
nand ( n77366 , n38499 , n54302 );
nand ( n77367 , n77365 , n77366 );
nand ( n77368 , n77367 , n54327 );
nand ( n77369 , n77362 , n77368 );
not ( n77370 , n70183 );
and ( n77371 , n71409 , n76444 );
not ( n77372 , n71409 );
and ( n77373 , n77372 , n39575 );
nor ( n77374 , n77371 , n77373 );
not ( n77375 , n77374 );
or ( n77376 , n77370 , n77375 );
nand ( n77377 , n77110 , n70193 );
nand ( n77378 , n77376 , n77377 );
xor ( n77379 , n77369 , n77378 );
not ( n77380 , n52854 );
not ( n77381 , n77120 );
or ( n77382 , n77380 , n77381 );
not ( n77383 , n54283 );
not ( n77384 , n42399 );
or ( n77385 , n77383 , n77384 );
nand ( n77386 , n42400 , n55104 );
nand ( n77387 , n77385 , n77386 );
nand ( n77388 , n77387 , n52469 );
nand ( n77389 , n77382 , n77388 );
xor ( n77390 , n77379 , n77389 );
xor ( n77391 , n77315 , n77390 );
not ( n77392 , n51766 );
not ( n77393 , n68931 );
not ( n77394 , n66784 );
or ( n77395 , n77393 , n77394 );
nand ( n77396 , n42654 , n52110 );
nand ( n77397 , n77395 , n77396 );
not ( n77398 , n77397 );
or ( n77399 , n77392 , n77398 );
nand ( n77400 , n77160 , n53197 );
nand ( n77401 , n77399 , n77400 );
not ( n77402 , n56777 );
not ( n77403 , n77147 );
or ( n77404 , n77402 , n77403 );
and ( n77405 , n65708 , n72593 );
not ( n77406 , n65708 );
and ( n77407 , n77406 , n56786 );
or ( n77408 , n77405 , n77407 );
nand ( n77409 , n77408 , n60472 );
nand ( n77410 , n77404 , n77409 );
xor ( n77411 , n77401 , n77410 );
not ( n77412 , n53620 );
and ( n77413 , n69530 , n71756 );
not ( n77414 , n69530 );
and ( n77415 , n77414 , n53596 );
or ( n77416 , n77413 , n77415 );
not ( n77417 , n77416 );
or ( n77418 , n77412 , n77417 );
nand ( n77419 , n77173 , n68603 );
nand ( n77420 , n77418 , n77419 );
xor ( n77421 , n77411 , n77420 );
xor ( n77422 , n77391 , n77421 );
xor ( n77423 , n77359 , n77422 );
not ( n77424 , n55458 );
not ( n77425 , n71371 );
not ( n77426 , n43513 );
or ( n77427 , n77425 , n77426 );
nand ( n77428 , n60386 , n69237 );
nand ( n77429 , n77427 , n77428 );
not ( n77430 , n77429 );
or ( n77431 , n77424 , n77430 );
nand ( n77432 , n77132 , n71099 );
nand ( n77433 , n77431 , n77432 );
xor ( n77434 , n77433 , n77207 );
xor ( n77435 , n77434 , n77055 );
xor ( n77436 , n77435 , n77246 );
xor ( n77437 , n77436 , n77254 );
xor ( n77438 , n77423 , n77437 );
xor ( n77439 , n77359 , n77422 );
and ( n77440 , n77439 , n77437 );
and ( n77441 , n77359 , n77422 );
or ( n77442 , n77440 , n77441 );
xor ( n77443 , n77262 , n77102 );
xor ( n77444 , n77443 , n77323 );
xor ( n77445 , n77262 , n77102 );
and ( n77446 , n77445 , n77323 );
and ( n77447 , n77262 , n77102 );
or ( n77448 , n77446 , n77447 );
xor ( n77449 , n77438 , n77197 );
xor ( n77450 , n77449 , n77218 );
xor ( n77451 , n77438 , n77197 );
and ( n77452 , n77451 , n77218 );
and ( n77453 , n77438 , n77197 );
or ( n77454 , n77452 , n77453 );
xor ( n77455 , n77444 , n77450 );
xor ( n77456 , n77455 , n77224 );
xor ( n77457 , n77444 , n77450 );
and ( n77458 , n77457 , n77224 );
and ( n77459 , n77444 , n77450 );
or ( n77460 , n77458 , n77459 );
xor ( n77461 , n77339 , n77350 );
and ( n77462 , n77461 , n77357 );
and ( n77463 , n77339 , n77350 );
or ( n77464 , n77462 , n77463 );
xor ( n77465 , n77401 , n77410 );
and ( n77466 , n77465 , n77420 );
and ( n77467 , n77401 , n77410 );
or ( n77468 , n77466 , n77467 );
xor ( n77469 , n77369 , n77378 );
and ( n77470 , n77469 , n77389 );
and ( n77471 , n77369 , n77378 );
or ( n77472 , n77470 , n77471 );
xor ( n77473 , n77433 , n77207 );
and ( n77474 , n77473 , n77055 );
and ( n77475 , n77433 , n77207 );
or ( n77476 , n77474 , n77475 );
xor ( n77477 , n77092 , n77279 );
and ( n77478 , n77477 , n77234 );
and ( n77479 , n77092 , n77279 );
or ( n77480 , n77478 , n77479 );
xor ( n77481 , n77238 , n77242 );
and ( n77482 , n77481 , n77358 );
and ( n77483 , n77238 , n77242 );
or ( n77484 , n77482 , n77483 );
xor ( n77485 , n77315 , n77390 );
and ( n77486 , n77485 , n77421 );
and ( n77487 , n77315 , n77390 );
or ( n77488 , n77486 , n77487 );
xor ( n77489 , n77435 , n77246 );
and ( n77490 , n77489 , n77254 );
and ( n77491 , n77435 , n77246 );
or ( n77492 , n77490 , n77491 );
not ( n77493 , n70487 );
not ( n77494 , n77299 );
or ( n77495 , n77493 , n77494 );
not ( n77496 , n59341 );
not ( n77497 , n71442 );
or ( n77498 , n77496 , n77497 );
nand ( n77499 , n72217 , n59340 );
nand ( n77500 , n77498 , n77499 );
nand ( n77501 , n77500 , n60542 );
nand ( n77502 , n77495 , n77501 );
not ( n77503 , n70500 );
not ( n77504 , n77310 );
or ( n77505 , n77503 , n77504 );
not ( n77506 , n68878 );
not ( n77507 , n68991 );
or ( n77508 , n77506 , n77507 );
nand ( n77509 , n68994 , n72477 );
nand ( n77510 , n77508 , n77509 );
nand ( n77511 , n77510 , n70930 );
nand ( n77512 , n77505 , n77511 );
xor ( n77513 , n77502 , n77512 );
not ( n77514 , n72484 );
not ( n77515 , n77335 );
or ( n77516 , n77514 , n77515 );
not ( n77517 , n71307 );
not ( n77518 , n77517 );
not ( n77519 , n66236 );
or ( n77520 , n77518 , n77519 );
nand ( n77521 , n71479 , n77333 );
nand ( n77522 , n77520 , n77521 );
nand ( n77523 , n77522 , n61558 );
nand ( n77524 , n77516 , n77523 );
xor ( n77525 , n77513 , n77524 );
xor ( n77526 , n77502 , n77512 );
and ( n77527 , n77526 , n77524 );
and ( n77528 , n77502 , n77512 );
or ( n77529 , n77527 , n77528 );
not ( n77530 , n77077 );
not ( n77531 , n77346 );
or ( n77532 , n77530 , n77531 );
and ( n77533 , n72148 , n76004 );
not ( n77534 , n72148 );
and ( n77535 , n77534 , n64170 );
or ( n77536 , n77533 , n77535 );
nand ( n77537 , n77536 , n67068 );
nand ( n77538 , n77532 , n77537 );
not ( n77539 , n70964 );
xor ( n77540 , n66155 , n72160 );
not ( n77541 , n77540 );
or ( n77542 , n77539 , n77541 );
nand ( n77543 , n77355 , n71960 );
nand ( n77544 , n77542 , n77543 );
xor ( n77545 , n77538 , n77544 );
and ( n77546 , n72846 , n40529 );
xor ( n77547 , n77545 , n77546 );
xor ( n77548 , n77538 , n77544 );
and ( n77549 , n77548 , n77546 );
and ( n77550 , n77538 , n77544 );
or ( n77551 , n77549 , n77550 );
not ( n77552 , n68603 );
not ( n77553 , n77416 );
or ( n77554 , n77552 , n77553 );
not ( n77555 , n53596 );
not ( n77556 , n69961 );
or ( n77557 , n77555 , n77556 );
nand ( n77558 , n69962 , n71756 );
nand ( n77559 , n77557 , n77558 );
nand ( n77560 , n77559 , n54364 );
nand ( n77561 , n77554 , n77560 );
not ( n77562 , n72185 );
not ( n77563 , n76786 );
not ( n77564 , n67040 );
or ( n77565 , n77563 , n77564 );
nand ( n77566 , n59913 , n72593 );
nand ( n77567 , n77565 , n77566 );
not ( n77568 , n77567 );
or ( n77569 , n77562 , n77568 );
nand ( n77570 , n77408 , n56777 );
nand ( n77571 , n77569 , n77570 );
xor ( n77572 , n77561 , n77571 );
and ( n77573 , n77289 , n75025 );
not ( n77574 , n74289 );
not ( n77575 , n70653 );
not ( n77576 , n77575 );
or ( n77577 , n77574 , n77576 );
nand ( n77578 , n70653 , n65187 );
nand ( n77579 , n77577 , n77578 );
and ( n77580 , n77579 , n61465 );
nor ( n77581 , n77573 , n77580 );
xor ( n77582 , n77572 , n77581 );
xor ( n77583 , n77525 , n77582 );
not ( n77584 , n70193 );
not ( n77585 , n77374 );
or ( n77586 , n77584 , n77585 );
not ( n77587 , n55120 );
not ( n77588 , n69072 );
or ( n77589 , n77587 , n77588 );
nand ( n77590 , n39056 , n71409 );
nand ( n77591 , n77589 , n77590 );
nand ( n77592 , n77591 , n70183 );
nand ( n77593 , n77586 , n77592 );
not ( n77594 , n53197 );
not ( n77595 , n77397 );
or ( n77596 , n77594 , n77595 );
not ( n77597 , n52113 );
nand ( n77598 , n77597 , n72220 );
nand ( n77599 , n77596 , n77598 );
xor ( n77600 , n77593 , n77599 );
not ( n77601 , n71099 );
not ( n77602 , n77429 );
or ( n77603 , n77601 , n77602 );
not ( n77604 , n74402 );
not ( n77605 , n62931 );
or ( n77606 , n77604 , n77605 );
nand ( n77607 , n39714 , n76016 );
nand ( n77608 , n77606 , n77607 );
nand ( n77609 , n77608 , n55458 );
nand ( n77610 , n77603 , n77609 );
xor ( n77611 , n77600 , n77610 );
xor ( n77612 , n77583 , n77611 );
xor ( n77613 , n77488 , n77612 );
xor ( n77614 , n77613 , n77492 );
xor ( n77615 , n77488 , n77612 );
and ( n77616 , n77615 , n77492 );
and ( n77617 , n77488 , n77612 );
or ( n77618 , n77616 , n77617 );
not ( n77619 , n52469 );
not ( n77620 , n54283 );
not ( n77621 , n67269 );
or ( n77622 , n77620 , n77621 );
nand ( n77623 , n73048 , n55104 );
nand ( n77624 , n77622 , n77623 );
not ( n77625 , n77624 );
or ( n77626 , n77619 , n77625 );
nand ( n77627 , n77387 , n52854 );
nand ( n77628 , n77626 , n77627 );
not ( n77629 , n72710 );
and ( n77630 , n73307 , n68142 );
not ( n77631 , n73307 );
and ( n77632 , n77631 , n66215 );
nor ( n77633 , n77630 , n77632 );
not ( n77634 , n77633 );
or ( n77635 , n77629 , n77634 );
nand ( n77636 , n77274 , n72961 );
nand ( n77637 , n77635 , n77636 );
xor ( n77638 , n77628 , n77637 );
not ( n77639 , n72142 );
not ( n77640 , n77367 );
or ( n77641 , n77639 , n77640 );
not ( n77642 , n70627 );
not ( n77643 , n73062 );
or ( n77644 , n77642 , n77643 );
or ( n77645 , n73062 , n70627 );
nand ( n77646 , n77644 , n77645 );
nand ( n77647 , n77646 , n54327 );
nand ( n77648 , n77641 , n77647 );
xor ( n77649 , n77638 , n77648 );
xor ( n77650 , n77649 , n77476 );
xor ( n77651 , n77650 , n77484 );
xor ( n77652 , n77651 , n77327 );
xor ( n77653 , n77283 , n77319 );
xor ( n77654 , n77653 , n77464 );
xor ( n77655 , n77654 , n77480 );
xor ( n77656 , n77468 , n77472 );
xor ( n77657 , n77656 , n77547 );
xor ( n77658 , n77655 , n77657 );
xor ( n77659 , n77652 , n77658 );
xor ( n77660 , n77651 , n77327 );
and ( n77661 , n77660 , n77658 );
and ( n77662 , n77651 , n77327 );
or ( n77663 , n77661 , n77662 );
xor ( n77664 , n77442 , n77614 );
xor ( n77665 , n77664 , n77659 );
xor ( n77666 , n77442 , n77614 );
and ( n77667 , n77666 , n77659 );
and ( n77668 , n77442 , n77614 );
or ( n77669 , n77667 , n77668 );
xor ( n77670 , n77448 , n77665 );
xor ( n77671 , n77670 , n77454 );
xor ( n77672 , n77448 , n77665 );
and ( n77673 , n77672 , n77454 );
and ( n77674 , n77448 , n77665 );
or ( n77675 , n77673 , n77674 );
xor ( n77676 , n77628 , n77637 );
and ( n77677 , n77676 , n77648 );
and ( n77678 , n77628 , n77637 );
or ( n77679 , n77677 , n77678 );
xor ( n77680 , n77593 , n77599 );
and ( n77681 , n77680 , n77610 );
and ( n77682 , n77593 , n77599 );
or ( n77683 , n77681 , n77682 );
xor ( n77684 , n77561 , n77571 );
and ( n77685 , n77684 , n77581 );
and ( n77686 , n77561 , n77571 );
or ( n77687 , n77685 , n77686 );
xor ( n77688 , n77283 , n77319 );
and ( n77689 , n77688 , n77464 );
and ( n77690 , n77283 , n77319 );
or ( n77691 , n77689 , n77690 );
xor ( n77692 , n77468 , n77472 );
and ( n77693 , n77692 , n77547 );
and ( n77694 , n77468 , n77472 );
or ( n77695 , n77693 , n77694 );
xor ( n77696 , n77525 , n77582 );
and ( n77697 , n77696 , n77611 );
and ( n77698 , n77525 , n77582 );
or ( n77699 , n77697 , n77698 );
xor ( n77700 , n77649 , n77476 );
and ( n77701 , n77700 , n77484 );
and ( n77702 , n77649 , n77476 );
or ( n77703 , n77701 , n77702 );
xor ( n77704 , n77654 , n77480 );
and ( n77705 , n77704 , n77657 );
and ( n77706 , n77654 , n77480 );
or ( n77707 , n77705 , n77706 );
not ( n77708 , n62302 );
not ( n77709 , n52481 );
or ( n77710 , n77708 , n77709 );
nand ( n77711 , n77710 , n52490 );
not ( n77712 , n75025 );
not ( n77713 , n77579 );
or ( n77714 , n77712 , n77713 );
not ( n77715 , n74289 );
not ( n77716 , n75162 );
or ( n77717 , n77715 , n77716 );
nand ( n77718 , n75161 , n65187 );
nand ( n77719 , n77717 , n77718 );
nand ( n77720 , n77719 , n71466 );
nand ( n77721 , n77714 , n77720 );
xor ( n77722 , n77711 , n77721 );
not ( n77723 , n75578 );
not ( n77724 , n66985 );
not ( n77725 , n70290 );
or ( n77726 , n77724 , n77725 );
nand ( n77727 , n40514 , n59340 );
nand ( n77728 , n77726 , n77727 );
not ( n77729 , n77728 );
or ( n77730 , n77723 , n77729 );
nand ( n77731 , n77500 , n70487 );
nand ( n77732 , n77730 , n77731 );
xor ( n77733 , n77722 , n77732 );
xor ( n77734 , n77711 , n77721 );
and ( n77735 , n77734 , n77732 );
and ( n77736 , n77711 , n77721 );
or ( n77737 , n77735 , n77736 );
not ( n77738 , n70500 );
not ( n77739 , n77510 );
or ( n77740 , n77738 , n77739 );
not ( n77741 , n68878 );
not ( n77742 , n73327 );
or ( n77743 , n77741 , n77742 );
nand ( n77744 , n40382 , n72477 );
nand ( n77745 , n77743 , n77744 );
nand ( n77746 , n77745 , n70930 );
nand ( n77747 , n77740 , n77746 );
not ( n77748 , n61558 );
and ( n77749 , n77333 , n54402 );
not ( n77750 , n77333 );
and ( n77751 , n77750 , n40149 );
nor ( n77752 , n77749 , n77751 );
not ( n77753 , n77752 );
or ( n77754 , n77748 , n77753 );
nand ( n77755 , n77522 , n75753 );
nand ( n77756 , n77754 , n77755 );
xor ( n77757 , n77747 , n77756 );
not ( n77758 , n75427 );
not ( n77759 , n72083 );
not ( n77760 , n40225 );
or ( n77761 , n77759 , n77760 );
nand ( n77762 , n40226 , n77344 );
nand ( n77763 , n77761 , n77762 );
not ( n77764 , n77763 );
or ( n77765 , n77758 , n77764 );
nand ( n77766 , n77077 , n77536 );
nand ( n77767 , n77765 , n77766 );
xor ( n77768 , n77757 , n77767 );
xor ( n77769 , n77747 , n77756 );
and ( n77770 , n77769 , n77767 );
and ( n77771 , n77747 , n77756 );
or ( n77772 , n77770 , n77771 );
not ( n77773 , n70964 );
not ( n77774 , n54415 );
xor ( n77775 , n72846 , n77774 );
not ( n77776 , n77775 );
or ( n77777 , n77773 , n77776 );
nand ( n77778 , n77540 , n71960 );
nand ( n77779 , n77777 , n77778 );
and ( n77780 , n66155 , n74581 );
xor ( n77781 , n77779 , n77780 );
not ( n77782 , n52469 );
buf ( n77783 , n70333 );
and ( n77784 , n54283 , n77783 );
not ( n77785 , n54283 );
and ( n77786 , n77785 , n71876 );
nor ( n77787 , n77784 , n77786 );
not ( n77788 , n77787 );
or ( n77789 , n77782 , n77788 );
nand ( n77790 , n77624 , n52854 );
nand ( n77791 , n77789 , n77790 );
xor ( n77792 , n77781 , n77791 );
xor ( n77793 , n77679 , n77792 );
xor ( n77794 , n77793 , n77683 );
xor ( n77795 , n77733 , n77768 );
not ( n77796 , n59984 );
and ( n77797 , n76016 , n76444 );
not ( n77798 , n76016 );
and ( n77799 , n77798 , n68667 );
nor ( n77800 , n77797 , n77799 );
not ( n77801 , n77800 );
or ( n77802 , n77796 , n77801 );
nand ( n77803 , n77608 , n71099 );
nand ( n77804 , n77802 , n77803 );
not ( n77805 , n53620 );
not ( n77806 , n55089 );
not ( n77807 , n72642 );
or ( n77808 , n77806 , n77807 );
nand ( n77809 , n76454 , n72238 );
nand ( n77810 , n77808 , n77809 );
not ( n77811 , n77810 );
or ( n77812 , n77805 , n77811 );
nand ( n77813 , n77559 , n68603 );
nand ( n77814 , n77812 , n77813 );
xor ( n77815 , n77804 , n77814 );
not ( n77816 , n72185 );
not ( n77817 , n76786 );
not ( n77818 , n73428 );
or ( n77819 , n77817 , n77818 );
nand ( n77820 , n60386 , n72593 );
nand ( n77821 , n77819 , n77820 );
not ( n77822 , n77821 );
or ( n77823 , n77816 , n77822 );
nand ( n77824 , n77567 , n56777 );
nand ( n77825 , n77823 , n77824 );
xor ( n77826 , n77815 , n77825 );
xor ( n77827 , n77795 , n77826 );
xor ( n77828 , n77794 , n77827 );
not ( n77829 , n59414 );
nand ( n77830 , n77829 , n75343 );
not ( n77831 , n77830 );
not ( n77832 , n75343 );
not ( n77833 , n73271 );
and ( n77834 , n77832 , n77833 );
nor ( n77835 , n77834 , n69648 );
not ( n77836 , n77835 );
or ( n77837 , n77831 , n77836 );
nand ( n77838 , n77633 , n72182 );
nand ( n77839 , n77837 , n77838 );
not ( n77840 , n77646 );
not ( n77841 , n54316 );
or ( n77842 , n77840 , n77841 );
not ( n77843 , n70627 );
not ( n77844 , n71176 );
or ( n77845 , n77843 , n77844 );
nand ( n77846 , n69530 , n54302 );
nand ( n77847 , n77845 , n77846 );
nand ( n77848 , n77847 , n54327 );
nand ( n77849 , n77842 , n77848 );
xor ( n77850 , n77839 , n77849 );
not ( n77851 , n70183 );
not ( n77852 , n55120 );
not ( n77853 , n68652 );
or ( n77854 , n77852 , n77853 );
nand ( n77855 , n38499 , n76714 );
nand ( n77856 , n77854 , n77855 );
not ( n77857 , n77856 );
or ( n77858 , n77851 , n77857 );
nand ( n77859 , n77591 , n55144 );
nand ( n77860 , n77858 , n77859 );
xor ( n77861 , n77850 , n77860 );
xor ( n77862 , n77861 , n77687 );
xor ( n77863 , n77862 , n77691 );
xor ( n77864 , n77828 , n77863 );
xor ( n77865 , n77794 , n77827 );
and ( n77866 , n77865 , n77863 );
and ( n77867 , n77794 , n77827 );
or ( n77868 , n77866 , n77867 );
xor ( n77869 , n77703 , n77707 );
not ( n77870 , n77581 );
xor ( n77871 , n77870 , n77529 );
xor ( n77872 , n77871 , n77551 );
xor ( n77873 , n77695 , n77872 );
xor ( n77874 , n77873 , n77699 );
xor ( n77875 , n77869 , n77874 );
xor ( n77876 , n77703 , n77707 );
and ( n77877 , n77876 , n77874 );
and ( n77878 , n77703 , n77707 );
or ( n77879 , n77877 , n77878 );
xor ( n77880 , n77864 , n77618 );
xor ( n77881 , n77880 , n77663 );
xor ( n77882 , n77864 , n77618 );
and ( n77883 , n77882 , n77663 );
and ( n77884 , n77864 , n77618 );
or ( n77885 , n77883 , n77884 );
xor ( n77886 , n77875 , n77881 );
xor ( n77887 , n77886 , n77669 );
xor ( n77888 , n77875 , n77881 );
and ( n77889 , n77888 , n77669 );
and ( n77890 , n77875 , n77881 );
or ( n77891 , n77889 , n77890 );
xor ( n77892 , n77779 , n77780 );
and ( n77893 , n77892 , n77791 );
and ( n77894 , n77779 , n77780 );
or ( n77895 , n77893 , n77894 );
xor ( n77896 , n77839 , n77849 );
and ( n77897 , n77896 , n77860 );
and ( n77898 , n77839 , n77849 );
or ( n77899 , n77897 , n77898 );
xor ( n77900 , n77804 , n77814 );
and ( n77901 , n77900 , n77825 );
and ( n77902 , n77804 , n77814 );
or ( n77903 , n77901 , n77902 );
xor ( n77904 , n77870 , n77529 );
and ( n77905 , n77904 , n77551 );
and ( n77906 , n77870 , n77529 );
or ( n77907 , n77905 , n77906 );
xor ( n77908 , n77679 , n77792 );
and ( n77909 , n77908 , n77683 );
and ( n77910 , n77679 , n77792 );
or ( n77911 , n77909 , n77910 );
xor ( n77912 , n77733 , n77768 );
and ( n77913 , n77912 , n77826 );
and ( n77914 , n77733 , n77768 );
or ( n77915 , n77913 , n77914 );
xor ( n77916 , n77861 , n77687 );
and ( n77917 , n77916 , n77691 );
and ( n77918 , n77861 , n77687 );
or ( n77919 , n77917 , n77918 );
xor ( n77920 , n77695 , n77872 );
and ( n77921 , n77920 , n77699 );
and ( n77922 , n77695 , n77872 );
or ( n77923 , n77921 , n77922 );
not ( n77924 , n72484 );
not ( n77925 , n77752 );
or ( n77926 , n77924 , n77925 );
not ( n77927 , n77517 );
not ( n77928 , n57390 );
or ( n77929 , n77927 , n77928 );
not ( n77930 , n68991 );
nand ( n77931 , n77930 , n71307 );
nand ( n77932 , n77929 , n77931 );
nand ( n77933 , n77932 , n61558 );
nand ( n77934 , n77926 , n77933 );
not ( n77935 , n70487 );
not ( n77936 , n77728 );
or ( n77937 , n77935 , n77936 );
not ( n77938 , n72464 );
not ( n77939 , n77575 );
or ( n77940 , n77938 , n77939 );
nand ( n77941 , n70653 , n70920 );
nand ( n77942 , n77940 , n77941 );
nand ( n77943 , n77942 , n75578 );
nand ( n77944 , n77937 , n77943 );
xor ( n77945 , n77934 , n77944 );
not ( n77946 , n71960 );
not ( n77947 , n77775 );
or ( n77948 , n77946 , n77947 );
xor ( n77949 , n72148 , n71971 );
nand ( n77950 , n77949 , n70964 );
nand ( n77951 , n77948 , n77950 );
xor ( n77952 , n77945 , n77951 );
xor ( n77953 , n77934 , n77944 );
and ( n77954 , n77953 , n77951 );
and ( n77955 , n77934 , n77944 );
or ( n77956 , n77954 , n77955 );
not ( n77957 , n77077 );
not ( n77958 , n77763 );
or ( n77959 , n77957 , n77958 );
not ( n77960 , n72083 );
not ( n77961 , n63201 );
or ( n77962 , n77960 , n77961 );
buf ( n77963 , n59195 );
nand ( n77964 , n77963 , n77344 );
nand ( n77965 , n77962 , n77964 );
nand ( n77966 , n77965 , n75427 );
nand ( n77967 , n77959 , n77966 );
and ( n77968 , n66155 , n72160 );
xor ( n77969 , n77967 , n77968 );
not ( n77970 , n54364 );
not ( n77971 , n55089 );
not ( n77972 , n42556 );
not ( n77973 , n77972 );
or ( n77974 , n77971 , n77973 );
nand ( n77975 , n42556 , n72238 );
nand ( n77976 , n77974 , n77975 );
not ( n77977 , n77976 );
or ( n77978 , n77970 , n77977 );
nand ( n77979 , n77810 , n68603 );
nand ( n77980 , n77978 , n77979 );
xor ( n77981 , n77969 , n77980 );
xor ( n77982 , n77967 , n77968 );
and ( n77983 , n77982 , n77980 );
and ( n77984 , n77967 , n77968 );
or ( n77985 , n77983 , n77984 );
not ( n77986 , n52854 );
not ( n77987 , n77787 );
or ( n77988 , n77986 , n77987 );
nand ( n77989 , n53571 , n69458 );
nand ( n77990 , n77988 , n77989 );
not ( n77991 , n56777 );
not ( n77992 , n77821 );
or ( n77993 , n77991 , n77992 );
not ( n77994 , n72589 );
not ( n77995 , n68206 );
or ( n77996 , n77994 , n77995 );
nand ( n77997 , n39714 , n71362 );
nand ( n77998 , n77996 , n77997 );
nand ( n77999 , n77998 , n72185 );
nand ( n78000 , n77993 , n77999 );
xor ( n78001 , n77990 , n78000 );
not ( n78002 , n54327 );
not ( n78003 , n70627 );
not ( n78004 , n69961 );
or ( n78005 , n78003 , n78004 );
nand ( n78006 , n69962 , n54468 );
nand ( n78007 , n78005 , n78006 );
not ( n78008 , n78007 );
or ( n78009 , n78002 , n78008 );
nand ( n78010 , n77847 , n72142 );
nand ( n78011 , n78009 , n78010 );
xor ( n78012 , n78001 , n78011 );
not ( n78013 , n71466 );
not ( n78014 , n65184 );
not ( n78015 , n75594 );
or ( n78016 , n78014 , n78015 );
nand ( n78017 , n39847 , n65183 );
nand ( n78018 , n78016 , n78017 );
not ( n78019 , n78018 );
or ( n78020 , n78013 , n78019 );
nand ( n78021 , n77719 , n75025 );
nand ( n78022 , n78020 , n78021 );
not ( n78023 , n55144 );
not ( n78024 , n77856 );
or ( n78025 , n78023 , n78024 );
not ( n78026 , n72919 );
not ( n78027 , n73062 );
or ( n78028 , n78026 , n78027 );
nand ( n78029 , n73065 , n76714 );
nand ( n78030 , n78028 , n78029 );
nand ( n78031 , n78030 , n70183 );
nand ( n78032 , n78025 , n78031 );
xor ( n78033 , n78022 , n78032 );
not ( n78034 , n77800 );
not ( n78035 , n71099 );
or ( n78036 , n78034 , n78035 );
not ( n78037 , n74402 );
not ( n78038 , n59891 );
or ( n78039 , n78037 , n78038 );
nand ( n78040 , n71547 , n69237 );
nand ( n78041 , n78039 , n78040 );
nand ( n78042 , n78041 , n59984 );
nand ( n78043 , n78036 , n78042 );
xor ( n78044 , n78033 , n78043 );
xor ( n78045 , n78012 , n78044 );
and ( n78046 , n75343 , n71863 );
not ( n78047 , n75343 );
and ( n78048 , n78047 , n76930 );
nor ( n78049 , n78046 , n78048 );
nand ( n78050 , n78049 , n72182 );
and ( n78051 , n67568 , n74900 );
not ( n78052 , n67568 );
and ( n78053 , n78052 , n75548 );
or ( n78054 , n78051 , n78053 );
nand ( n78055 , n78054 , n72710 );
nand ( n78056 , n78050 , n78055 );
not ( n78057 , n70500 );
not ( n78058 , n77745 );
or ( n78059 , n78057 , n78058 );
not ( n78060 , n75286 );
not ( n78061 , n71442 );
or ( n78062 , n78060 , n78061 );
nand ( n78063 , n72217 , n73190 );
nand ( n78064 , n78062 , n78063 );
nand ( n78065 , n78064 , n70930 );
nand ( n78066 , n78059 , n78065 );
not ( n78067 , n78066 );
xor ( n78068 , n78056 , n78067 );
xor ( n78069 , n78068 , n77737 );
xor ( n78070 , n78045 , n78069 );
xor ( n78071 , n78070 , n77923 );
xor ( n78072 , n77907 , n77911 );
xor ( n78073 , n77772 , n77899 );
xor ( n78074 , n78073 , n77895 );
xor ( n78075 , n78072 , n78074 );
xor ( n78076 , n78071 , n78075 );
xor ( n78077 , n78070 , n77923 );
and ( n78078 , n78077 , n78075 );
and ( n78079 , n78070 , n77923 );
or ( n78080 , n78078 , n78079 );
xor ( n78081 , n77903 , n77981 );
xor ( n78082 , n78081 , n77952 );
xor ( n78083 , n78082 , n77915 );
xor ( n78084 , n78083 , n77919 );
xor ( n78085 , n77868 , n78084 );
xor ( n78086 , n78085 , n77879 );
xor ( n78087 , n77868 , n78084 );
and ( n78088 , n78087 , n77879 );
and ( n78089 , n77868 , n78084 );
or ( n78090 , n78088 , n78089 );
xor ( n78091 , n78076 , n78086 );
xor ( n78092 , n78091 , n77885 );
xor ( n78093 , n78076 , n78086 );
and ( n78094 , n78093 , n77885 );
and ( n78095 , n78076 , n78086 );
or ( n78096 , n78094 , n78095 );
xor ( n78097 , n78022 , n78032 );
and ( n78098 , n78097 , n78043 );
and ( n78099 , n78022 , n78032 );
or ( n78100 , n78098 , n78099 );
xor ( n78101 , n77990 , n78000 );
and ( n78102 , n78101 , n78011 );
and ( n78103 , n77990 , n78000 );
or ( n78104 , n78102 , n78103 );
xor ( n78105 , n78056 , n78067 );
and ( n78106 , n78105 , n77737 );
and ( n78107 , n78056 , n78067 );
or ( n78108 , n78106 , n78107 );
xor ( n78109 , n77772 , n77899 );
and ( n78110 , n78109 , n77895 );
and ( n78111 , n77772 , n77899 );
or ( n78112 , n78110 , n78111 );
xor ( n78113 , n77903 , n77981 );
and ( n78114 , n78113 , n77952 );
and ( n78115 , n77903 , n77981 );
or ( n78116 , n78114 , n78115 );
xor ( n78117 , n78012 , n78044 );
and ( n78118 , n78117 , n78069 );
and ( n78119 , n78012 , n78044 );
or ( n78120 , n78118 , n78119 );
xor ( n78121 , n77907 , n77911 );
and ( n78122 , n78121 , n78074 );
and ( n78123 , n77907 , n77911 );
or ( n78124 , n78122 , n78123 );
xor ( n78125 , n78082 , n77915 );
and ( n78126 , n78125 , n77919 );
and ( n78127 , n78082 , n77915 );
or ( n78128 , n78126 , n78127 );
not ( n78129 , n56861 );
not ( n78130 , n70585 );
or ( n78131 , n78129 , n78130 );
nand ( n78132 , n78131 , n69458 );
not ( n78133 , n72131 );
not ( n78134 , n77942 );
or ( n78135 , n78133 , n78134 );
not ( n78136 , n59341 );
not ( n78137 , n75162 );
or ( n78138 , n78136 , n78137 );
nand ( n78139 , n75161 , n70920 );
nand ( n78140 , n78138 , n78139 );
nand ( n78141 , n78140 , n75578 );
nand ( n78142 , n78135 , n78141 );
xor ( n78143 , n78132 , n78142 );
not ( n78144 , n70930 );
not ( n78145 , n75286 );
not ( n78146 , n70290 );
or ( n78147 , n78145 , n78146 );
not ( n78148 , n70506 );
nand ( n78149 , n67721 , n78148 );
nand ( n78150 , n78147 , n78149 );
not ( n78151 , n78150 );
or ( n78152 , n78144 , n78151 );
nand ( n78153 , n78064 , n70500 );
nand ( n78154 , n78152 , n78153 );
xor ( n78155 , n78143 , n78154 );
xor ( n78156 , n78132 , n78142 );
and ( n78157 , n78156 , n78154 );
and ( n78158 , n78132 , n78142 );
or ( n78159 , n78157 , n78158 );
not ( n78160 , n75753 );
not ( n78161 , n77932 );
or ( n78162 , n78160 , n78161 );
not ( n78163 , n71309 );
not ( n78164 , n76821 );
or ( n78165 , n78163 , n78164 );
nand ( n78166 , n40382 , n64630 );
nand ( n78167 , n78165 , n78166 );
nand ( n78168 , n78167 , n61558 );
nand ( n78169 , n78162 , n78168 );
not ( n78170 , n77077 );
not ( n78171 , n77965 );
or ( n78172 , n78170 , n78171 );
not ( n78173 , n64170 );
not ( n78174 , n73279 );
or ( n78175 , n78173 , n78174 );
nand ( n78176 , n69409 , n76004 );
nand ( n78177 , n78175 , n78176 );
nand ( n78178 , n78177 , n75427 );
nand ( n78179 , n78172 , n78178 );
xor ( n78180 , n78169 , n78179 );
not ( n78181 , n70964 );
xor ( n78182 , n67072 , n40226 );
not ( n78183 , n78182 );
or ( n78184 , n78181 , n78183 );
nand ( n78185 , n71960 , n77949 );
nand ( n78186 , n78184 , n78185 );
xor ( n78187 , n78180 , n78186 );
xor ( n78188 , n78169 , n78179 );
and ( n78189 , n78188 , n78186 );
and ( n78190 , n78169 , n78179 );
or ( n78191 , n78189 , n78190 );
not ( n78192 , n54327 );
not ( n78193 , n70627 );
not ( n78194 , n71139 );
or ( n78195 , n78193 , n78194 );
nand ( n78196 , n42400 , n54468 );
nand ( n78197 , n78195 , n78196 );
not ( n78198 , n78197 );
or ( n78199 , n78192 , n78198 );
nand ( n78200 , n78007 , n72142 );
nand ( n78201 , n78199 , n78200 );
not ( n78202 , n72710 );
not ( n78203 , n67568 );
not ( n78204 , n43513 );
or ( n78205 , n78203 , n78204 );
nand ( n78206 , n60386 , n76811 );
nand ( n78207 , n78205 , n78206 );
not ( n78208 , n78207 );
or ( n78209 , n78202 , n78208 );
nand ( n78210 , n78054 , n72961 );
nand ( n78211 , n78209 , n78210 );
xor ( n78212 , n78201 , n78211 );
xor ( n78213 , n78212 , n78066 );
and ( n78214 , n72846 , n77774 );
not ( n78215 , n54364 );
not ( n78216 , n55089 );
not ( n78217 , n42655 );
or ( n78218 , n78216 , n78217 );
not ( n78219 , n42655 );
nand ( n78220 , n78219 , n72238 );
nand ( n78221 , n78218 , n78220 );
not ( n78222 , n78221 );
or ( n78223 , n78215 , n78222 );
nand ( n78224 , n77976 , n68603 );
nand ( n78225 , n78223 , n78224 );
xor ( n78226 , n78214 , n78225 );
not ( n78227 , n76828 );
not ( n78228 , n78018 );
or ( n78229 , n78227 , n78228 );
not ( n78230 , n65184 );
not ( n78231 , n39895 );
or ( n78232 , n78230 , n78231 );
nand ( n78233 , n39896 , n65183 );
nand ( n78234 , n78232 , n78233 );
nand ( n78235 , n78234 , n71466 );
nand ( n78236 , n78229 , n78235 );
xor ( n78237 , n78226 , n78236 );
xor ( n78238 , n78213 , n78237 );
not ( n78239 , n70183 );
not ( n78240 , n72919 );
not ( n78241 , n71176 );
or ( n78242 , n78240 , n78241 );
nand ( n78243 , n39255 , n76714 );
nand ( n78244 , n78242 , n78243 );
not ( n78245 , n78244 );
or ( n78246 , n78239 , n78245 );
nand ( n78247 , n78030 , n70193 );
nand ( n78248 , n78246 , n78247 );
not ( n78249 , n59984 );
not ( n78250 , n68652 );
not ( n78251 , n71371 );
or ( n78252 , n78250 , n78251 );
nand ( n78253 , n38499 , n69237 );
nand ( n78254 , n78252 , n78253 );
not ( n78255 , n78254 );
or ( n78256 , n78249 , n78255 );
nand ( n78257 , n78041 , n71099 );
nand ( n78258 , n78256 , n78257 );
xor ( n78259 , n78248 , n78258 );
not ( n78260 , n72185 );
not ( n78261 , n76786 );
not ( n78262 , n76444 );
or ( n78263 , n78261 , n78262 );
nand ( n78264 , n39575 , n71362 );
nand ( n78265 , n78263 , n78264 );
not ( n78266 , n78265 );
or ( n78267 , n78260 , n78266 );
nand ( n78268 , n77998 , n56777 );
nand ( n78269 , n78267 , n78268 );
xor ( n78270 , n78259 , n78269 );
xor ( n78271 , n78238 , n78270 );
xor ( n78272 , n78271 , n78124 );
xor ( n78273 , n78108 , n78116 );
xor ( n78274 , n78273 , n78112 );
xor ( n78275 , n78272 , n78274 );
xor ( n78276 , n78271 , n78124 );
and ( n78277 , n78276 , n78274 );
and ( n78278 , n78271 , n78124 );
or ( n78279 , n78277 , n78278 );
xor ( n78280 , n77956 , n78100 );
xor ( n78281 , n78280 , n77985 );
xor ( n78282 , n78187 , n78104 );
xor ( n78283 , n78282 , n78155 );
xor ( n78284 , n78281 , n78283 );
xor ( n78285 , n78284 , n78120 );
xor ( n78286 , n78285 , n78128 );
xor ( n78287 , n78286 , n78080 );
xor ( n78288 , n78285 , n78128 );
and ( n78289 , n78288 , n78080 );
and ( n78290 , n78285 , n78128 );
or ( n78291 , n78289 , n78290 );
xor ( n78292 , n78275 , n78287 );
xor ( n78293 , n78292 , n78090 );
xor ( n78294 , n78275 , n78287 );
and ( n78295 , n78294 , n78090 );
and ( n78296 , n78275 , n78287 );
or ( n78297 , n78295 , n78296 );
xor ( n78298 , n78214 , n78225 );
and ( n78299 , n78298 , n78236 );
and ( n78300 , n78214 , n78225 );
or ( n78301 , n78299 , n78300 );
xor ( n78302 , n78248 , n78258 );
and ( n78303 , n78302 , n78269 );
and ( n78304 , n78248 , n78258 );
or ( n78305 , n78303 , n78304 );
xor ( n78306 , n78201 , n78211 );
and ( n78307 , n78306 , n78066 );
and ( n78308 , n78201 , n78211 );
or ( n78309 , n78307 , n78308 );
xor ( n78310 , n77956 , n78100 );
and ( n78311 , n78310 , n77985 );
and ( n78312 , n77956 , n78100 );
or ( n78313 , n78311 , n78312 );
xor ( n78314 , n78187 , n78104 );
and ( n78315 , n78314 , n78155 );
and ( n78316 , n78187 , n78104 );
or ( n78317 , n78315 , n78316 );
xor ( n78318 , n78213 , n78237 );
and ( n78319 , n78318 , n78270 );
and ( n78320 , n78213 , n78237 );
or ( n78321 , n78319 , n78320 );
xor ( n78322 , n78108 , n78116 );
and ( n78323 , n78322 , n78112 );
and ( n78324 , n78108 , n78116 );
or ( n78325 , n78323 , n78324 );
xor ( n78326 , n78281 , n78283 );
and ( n78327 , n78326 , n78120 );
and ( n78328 , n78281 , n78283 );
or ( n78329 , n78327 , n78328 );
not ( n78330 , n77077 );
not ( n78331 , n78177 );
or ( n78332 , n78330 , n78331 );
not ( n78333 , n76004 );
not ( n78334 , n54791 );
or ( n78335 , n78333 , n78334 );
nand ( n78336 , n64170 , n68073 );
nand ( n78337 , n78335 , n78336 );
nand ( n78338 , n78337 , n67068 );
nand ( n78339 , n78332 , n78338 );
not ( n78340 , n70500 );
not ( n78341 , n78150 );
or ( n78342 , n78340 , n78341 );
not ( n78343 , n75286 );
not ( n78344 , n77575 );
or ( n78345 , n78343 , n78344 );
nand ( n78346 , n70653 , n73190 );
nand ( n78347 , n78345 , n78346 );
nand ( n78348 , n78347 , n70930 );
nand ( n78349 , n78342 , n78348 );
xor ( n78350 , n78339 , n78349 );
and ( n78351 , n72148 , n71971 );
xor ( n78352 , n78350 , n78351 );
xor ( n78353 , n78339 , n78349 );
and ( n78354 , n78353 , n78351 );
and ( n78355 , n78339 , n78349 );
or ( n78356 , n78354 , n78355 );
not ( n78357 , n71960 );
not ( n78358 , n78182 );
or ( n78359 , n78357 , n78358 );
xor ( n78360 , n69305 , n59195 );
nand ( n78361 , n78360 , n70964 );
nand ( n78362 , n78359 , n78361 );
not ( n78363 , n54327 );
and ( n78364 , n54725 , n42555 );
not ( n78365 , n54725 );
and ( n78366 , n78365 , n72307 );
nor ( n78367 , n78364 , n78366 );
not ( n78368 , n78367 );
or ( n78369 , n78363 , n78368 );
nand ( n78370 , n78197 , n72142 );
nand ( n78371 , n78369 , n78370 );
xor ( n78372 , n78362 , n78371 );
not ( n78373 , n75578 );
not ( n78374 , n59341 );
not ( n78375 , n75594 );
or ( n78376 , n78374 , n78375 );
nand ( n78377 , n39847 , n70920 );
nand ( n78378 , n78376 , n78377 );
not ( n78379 , n78378 );
or ( n78380 , n78373 , n78379 );
nand ( n78381 , n78140 , n72131 );
nand ( n78382 , n78380 , n78381 );
xor ( n78383 , n78372 , n78382 );
xor ( n78384 , n78362 , n78371 );
and ( n78385 , n78384 , n78382 );
and ( n78386 , n78362 , n78371 );
or ( n78387 , n78385 , n78386 );
xor ( n78388 , n78313 , n78321 );
xor ( n78389 , n78301 , n78352 );
xor ( n78390 , n78389 , n78305 );
xor ( n78391 , n78388 , n78390 );
xor ( n78392 , n78329 , n78391 );
not ( n78393 , n72961 );
not ( n78394 , n78207 );
or ( n78395 , n78393 , n78394 );
not ( n78396 , n67568 );
not ( n78397 , n39715 );
or ( n78398 , n78396 , n78397 );
nand ( n78399 , n71567 , n76811 );
nand ( n78400 , n78398 , n78399 );
nand ( n78401 , n78400 , n72710 );
nand ( n78402 , n78395 , n78401 );
not ( n78403 , n55144 );
not ( n78404 , n78244 );
or ( n78405 , n78403 , n78404 );
not ( n78406 , n72919 );
not ( n78407 , n69961 );
or ( n78408 , n78406 , n78407 );
nand ( n78409 , n69962 , n76714 );
nand ( n78410 , n78408 , n78409 );
nand ( n78411 , n78410 , n70183 );
nand ( n78412 , n78405 , n78411 );
xor ( n78413 , n78402 , n78412 );
not ( n78414 , n76828 );
not ( n78415 , n78234 );
or ( n78416 , n78414 , n78415 );
not ( n78417 , n65184 );
not ( n78418 , n74900 );
or ( n78419 , n78417 , n78418 );
nand ( n78420 , n75548 , n65183 );
nand ( n78421 , n78419 , n78420 );
nand ( n78422 , n78421 , n71466 );
nand ( n78423 , n78416 , n78422 );
xor ( n78424 , n78413 , n78423 );
xor ( n78425 , n78424 , n78383 );
not ( n78426 , n55872 );
not ( n78427 , n73062 );
or ( n78428 , n78426 , n78427 );
nand ( n78429 , n73065 , n76016 );
nand ( n78430 , n78428 , n78429 );
not ( n78431 , n78430 );
not ( n78432 , n59984 );
or ( n78433 , n78431 , n78432 );
nand ( n78434 , n78254 , n71099 );
nand ( n78435 , n78433 , n78434 );
not ( n78436 , n56777 );
not ( n78437 , n78265 );
or ( n78438 , n78436 , n78437 );
not ( n78439 , n72589 );
not ( n78440 , n59891 );
or ( n78441 , n78439 , n78440 );
nand ( n78442 , n71547 , n71362 );
nand ( n78443 , n78441 , n78442 );
nand ( n78444 , n78443 , n72185 );
nand ( n78445 , n78438 , n78444 );
xor ( n78446 , n78435 , n78445 );
not ( n78447 , n54364 );
not ( n78448 , n55089 );
or ( n78449 , n78447 , n78448 );
not ( n78450 , n78221 );
not ( n78451 , n68603 );
or ( n78452 , n78450 , n78451 );
nand ( n78453 , n78449 , n78452 );
xor ( n78454 , n78446 , n78453 );
xor ( n78455 , n78425 , n78454 );
xor ( n78456 , n78455 , n78325 );
not ( n78457 , n61558 );
xnor ( n78458 , n71309 , n71442 );
not ( n78459 , n78458 );
or ( n78460 , n78457 , n78459 );
nand ( n78461 , n78167 , n72484 );
nand ( n78462 , n78460 , n78461 );
not ( n78463 , n78462 );
xor ( n78464 , n78463 , n78191 );
xor ( n78465 , n78464 , n78159 );
xor ( n78466 , n78309 , n78465 );
xor ( n78467 , n78466 , n78317 );
xor ( n78468 , n78456 , n78467 );
xor ( n78469 , n78392 , n78468 );
xor ( n78470 , n78329 , n78391 );
and ( n78471 , n78470 , n78468 );
and ( n78472 , n78329 , n78391 );
or ( n78473 , n78471 , n78472 );
xor ( n78474 , n78279 , n78469 );
xor ( n78475 , n78474 , n78291 );
xor ( n78476 , n78279 , n78469 );
and ( n78477 , n78476 , n78291 );
and ( n78478 , n78279 , n78469 );
or ( n78479 , n78477 , n78478 );
xor ( n78480 , n78435 , n78445 );
and ( n78481 , n78480 , n78453 );
and ( n78482 , n78435 , n78445 );
or ( n78483 , n78481 , n78482 );
xor ( n78484 , n78402 , n78412 );
and ( n78485 , n78484 , n78423 );
and ( n78486 , n78402 , n78412 );
or ( n78487 , n78485 , n78486 );
xor ( n78488 , n78463 , n78191 );
and ( n78489 , n78488 , n78159 );
and ( n78490 , n78463 , n78191 );
or ( n78491 , n78489 , n78490 );
xor ( n78492 , n78301 , n78352 );
and ( n78493 , n78492 , n78305 );
and ( n78494 , n78301 , n78352 );
or ( n78495 , n78493 , n78494 );
xor ( n78496 , n78424 , n78383 );
and ( n78497 , n78496 , n78454 );
and ( n78498 , n78424 , n78383 );
or ( n78499 , n78497 , n78498 );
xor ( n78500 , n78309 , n78465 );
and ( n78501 , n78500 , n78317 );
and ( n78502 , n78309 , n78465 );
or ( n78503 , n78501 , n78502 );
xor ( n78504 , n78313 , n78321 );
and ( n78505 , n78504 , n78390 );
and ( n78506 , n78313 , n78321 );
or ( n78507 , n78505 , n78506 );
xor ( n78508 , n78455 , n78325 );
and ( n78509 , n78508 , n78467 );
and ( n78510 , n78455 , n78325 );
or ( n78511 , n78509 , n78510 );
not ( n78512 , n53620 );
not ( n78513 , n78512 );
not ( n78514 , n78451 );
or ( n78515 , n78513 , n78514 );
nand ( n78516 , n78515 , n55089 );
not ( n78517 , n70500 );
not ( n78518 , n78347 );
or ( n78519 , n78517 , n78518 );
and ( n78520 , n70506 , n59651 );
not ( n78521 , n70506 );
and ( n78522 , n78521 , n75161 );
or ( n78523 , n78520 , n78522 );
nand ( n78524 , n78523 , n70930 );
nand ( n78525 , n78519 , n78524 );
xor ( n78526 , n78516 , n78525 );
not ( n78527 , n61558 );
not ( n78528 , n61540 );
not ( n78529 , n70290 );
or ( n78530 , n78528 , n78529 );
not ( n78531 , n71309 );
nand ( n78532 , n78531 , n67721 );
nand ( n78533 , n78530 , n78532 );
not ( n78534 , n78533 );
or ( n78535 , n78527 , n78534 );
nand ( n78536 , n78458 , n75753 );
nand ( n78537 , n78535 , n78536 );
xor ( n78538 , n78526 , n78537 );
xor ( n78539 , n78516 , n78525 );
and ( n78540 , n78539 , n78537 );
and ( n78541 , n78516 , n78525 );
or ( n78542 , n78540 , n78541 );
not ( n78543 , n75427 );
not ( n78544 , n72083 );
not ( n78545 , n76821 );
or ( n78546 , n78544 , n78545 );
nand ( n78547 , n71829 , n77344 );
nand ( n78548 , n78546 , n78547 );
not ( n78549 , n78548 );
or ( n78550 , n78543 , n78549 );
nand ( n78551 , n78337 , n77077 );
nand ( n78552 , n78550 , n78551 );
not ( n78553 , n71960 );
not ( n78554 , n78360 );
or ( n78555 , n78553 , n78554 );
xor ( n78556 , n66155 , n69409 );
nand ( n78557 , n78556 , n70964 );
nand ( n78558 , n78555 , n78557 );
xor ( n78559 , n78552 , n78558 );
and ( n78560 , n67072 , n40226 );
xor ( n78561 , n78559 , n78560 );
xor ( n78562 , n78552 , n78558 );
and ( n78563 , n78562 , n78560 );
and ( n78564 , n78552 , n78558 );
or ( n78565 , n78563 , n78564 );
xor ( n78566 , n78495 , n78499 );
xor ( n78567 , n78561 , n78538 );
not ( n78568 , n54316 );
not ( n78569 , n78367 );
or ( n78570 , n78568 , n78569 );
and ( n78571 , n54302 , n71876 );
not ( n78572 , n54302 );
and ( n78573 , n78572 , n77783 );
nor ( n78574 , n78571 , n78573 );
nand ( n78575 , n78574 , n54327 );
nand ( n78576 , n78570 , n78575 );
not ( n78577 , n72131 );
not ( n78578 , n78378 );
or ( n78579 , n78577 , n78578 );
and ( n78580 , n59413 , n59340 );
not ( n78581 , n59413 );
and ( n78582 , n78581 , n59341 );
or ( n78583 , n78580 , n78582 );
nand ( n78584 , n78583 , n75578 );
nand ( n78585 , n78579 , n78584 );
xor ( n78586 , n78576 , n78585 );
not ( n78587 , n59984 );
not ( n78588 , n55872 );
not ( n78589 , n71176 );
or ( n78590 , n78588 , n78589 );
nand ( n78591 , n69530 , n76016 );
nand ( n78592 , n78590 , n78591 );
not ( n78593 , n78592 );
or ( n78594 , n78587 , n78593 );
nand ( n78595 , n78430 , n71099 );
nand ( n78596 , n78594 , n78595 );
xor ( n78597 , n78586 , n78596 );
xor ( n78598 , n78567 , n78597 );
xor ( n78599 , n78566 , n78598 );
xor ( n78600 , n78507 , n78599 );
xor ( n78601 , n78387 , n78483 );
xor ( n78602 , n78601 , n78487 );
xor ( n78603 , n78602 , n78503 );
not ( n78604 , n72185 );
not ( n78605 , n72589 );
not ( n78606 , n68652 );
or ( n78607 , n78605 , n78606 );
nand ( n78608 , n72622 , n72593 );
nand ( n78609 , n78607 , n78608 );
not ( n78610 , n78609 );
or ( n78611 , n78604 , n78610 );
nand ( n78612 , n78443 , n56777 );
nand ( n78613 , n78611 , n78612 );
not ( n78614 , n72710 );
and ( n78615 , n76811 , n73400 );
not ( n78616 , n76811 );
and ( n78617 , n78616 , n68667 );
nor ( n78618 , n78615 , n78617 );
not ( n78619 , n78618 );
or ( n78620 , n78614 , n78619 );
nand ( n78621 , n78400 , n72961 );
nand ( n78622 , n78620 , n78621 );
xor ( n78623 , n78613 , n78622 );
not ( n78624 , n70193 );
not ( n78625 , n78410 );
or ( n78626 , n78624 , n78625 );
not ( n78627 , n55120 );
not ( n78628 , n76455 );
or ( n78629 , n78627 , n78628 );
nand ( n78630 , n76454 , n71409 );
nand ( n78631 , n78629 , n78630 );
nand ( n78632 , n78631 , n70183 );
nand ( n78633 , n78626 , n78632 );
xor ( n78634 , n78623 , n78633 );
not ( n78635 , n71466 );
and ( n78636 , n74289 , n60386 );
not ( n78637 , n74289 );
and ( n78638 , n78637 , n71904 );
nor ( n78639 , n78636 , n78638 );
not ( n78640 , n78639 );
or ( n78641 , n78635 , n78640 );
nand ( n78642 , n78421 , n76828 );
nand ( n78643 , n78641 , n78642 );
xor ( n78644 , n78643 , n78462 );
xor ( n78645 , n78644 , n78356 );
xor ( n78646 , n78634 , n78645 );
xor ( n78647 , n78646 , n78491 );
xor ( n78648 , n78603 , n78647 );
xor ( n78649 , n78600 , n78648 );
xor ( n78650 , n78507 , n78599 );
and ( n78651 , n78650 , n78648 );
and ( n78652 , n78507 , n78599 );
or ( n78653 , n78651 , n78652 );
xor ( n78654 , n78511 , n78649 );
xor ( n78655 , n78654 , n78473 );
xor ( n78656 , n78511 , n78649 );
and ( n78657 , n78656 , n78473 );
and ( n78658 , n78511 , n78649 );
or ( n78659 , n78657 , n78658 );
xor ( n78660 , n78576 , n78585 );
and ( n78661 , n78660 , n78596 );
and ( n78662 , n78576 , n78585 );
or ( n78663 , n78661 , n78662 );
xor ( n78664 , n78613 , n78622 );
and ( n78665 , n78664 , n78633 );
and ( n78666 , n78613 , n78622 );
or ( n78667 , n78665 , n78666 );
xor ( n78668 , n78643 , n78462 );
and ( n78669 , n78668 , n78356 );
and ( n78670 , n78643 , n78462 );
or ( n78671 , n78669 , n78670 );
xor ( n78672 , n78387 , n78483 );
and ( n78673 , n78672 , n78487 );
and ( n78674 , n78387 , n78483 );
or ( n78675 , n78673 , n78674 );
xor ( n78676 , n78561 , n78538 );
and ( n78677 , n78676 , n78597 );
and ( n78678 , n78561 , n78538 );
or ( n78679 , n78677 , n78678 );
xor ( n78680 , n78634 , n78645 );
and ( n78681 , n78680 , n78491 );
and ( n78682 , n78634 , n78645 );
or ( n78683 , n78681 , n78682 );
xor ( n78684 , n78495 , n78499 );
and ( n78685 , n78684 , n78598 );
and ( n78686 , n78495 , n78499 );
or ( n78687 , n78685 , n78686 );
xor ( n78688 , n78602 , n78503 );
and ( n78689 , n78688 , n78647 );
and ( n78690 , n78602 , n78503 );
or ( n78691 , n78689 , n78690 );
not ( n78692 , n71960 );
not ( n78693 , n78556 );
or ( n78694 , n78692 , n78693 );
xor ( n78695 , n66155 , n68990 );
nand ( n78696 , n78695 , n70964 );
nand ( n78697 , n78694 , n78696 );
not ( n78698 , n72484 );
not ( n78699 , n78533 );
or ( n78700 , n78698 , n78699 );
not ( n78701 , n71309 );
not ( n78702 , n63180 );
or ( n78703 , n78701 , n78702 );
nand ( n78704 , n70653 , n75748 );
nand ( n78705 , n78703 , n78704 );
nand ( n78706 , n78705 , n61558 );
nand ( n78707 , n78700 , n78706 );
xor ( n78708 , n78697 , n78707 );
and ( n78709 , n69305 , n59195 );
xor ( n78710 , n78708 , n78709 );
xor ( n78711 , n78697 , n78707 );
and ( n78712 , n78711 , n78709 );
and ( n78713 , n78697 , n78707 );
or ( n78714 , n78712 , n78713 );
not ( n78715 , n55144 );
not ( n78716 , n78631 );
or ( n78717 , n78715 , n78716 );
not ( n78718 , n55120 );
not ( n78719 , n72307 );
or ( n78720 , n78718 , n78719 );
nand ( n78721 , n42556 , n71409 );
nand ( n78722 , n78720 , n78721 );
nand ( n78723 , n78722 , n70183 );
nand ( n78724 , n78717 , n78723 );
not ( n78725 , n70930 );
not ( n78726 , n75286 );
not ( n78727 , n75594 );
or ( n78728 , n78726 , n78727 );
nand ( n78729 , n39847 , n72477 );
nand ( n78730 , n78728 , n78729 );
not ( n78731 , n78730 );
or ( n78732 , n78725 , n78731 );
nand ( n78733 , n78523 , n70500 );
nand ( n78734 , n78732 , n78733 );
xor ( n78735 , n78724 , n78734 );
not ( n78736 , n56777 );
not ( n78737 , n78609 );
or ( n78738 , n78736 , n78737 );
not ( n78739 , n76786 );
not ( n78740 , n73062 );
or ( n78741 , n78739 , n78740 );
nand ( n78742 , n73065 , n72593 );
nand ( n78743 , n78741 , n78742 );
nand ( n78744 , n78743 , n72185 );
nand ( n78745 , n78738 , n78744 );
xor ( n78746 , n78735 , n78745 );
xor ( n78747 , n78724 , n78734 );
and ( n78748 , n78747 , n78745 );
and ( n78749 , n78724 , n78734 );
or ( n78750 , n78748 , n78749 );
xor ( n78751 , n78542 , n78565 );
xor ( n78752 , n78751 , n78710 );
xor ( n78753 , n78675 , n78752 );
xor ( n78754 , n78753 , n78679 );
xor ( n78755 , n78754 , n78687 );
xor ( n78756 , n78663 , n78667 );
not ( n78757 , n72961 );
not ( n78758 , n78618 );
or ( n78759 , n78757 , n78758 );
not ( n78760 , n75343 );
not ( n78761 , n69072 );
or ( n78762 , n78760 , n78761 );
nand ( n78763 , n39056 , n66963 );
nand ( n78764 , n78762 , n78763 );
nand ( n78765 , n78764 , n72710 );
nand ( n78766 , n78759 , n78765 );
not ( n78767 , n72142 );
not ( n78768 , n78574 );
or ( n78769 , n78767 , n78768 );
not ( n78770 , n54302 );
nand ( n78771 , n78770 , n54327 );
nand ( n78772 , n78769 , n78771 );
xor ( n78773 , n78766 , n78772 );
not ( n78774 , n76828 );
not ( n78775 , n78639 );
or ( n78776 , n78774 , n78775 );
not ( n78777 , n74289 );
not ( n78778 , n39715 );
or ( n78779 , n78777 , n78778 );
nand ( n78780 , n39714 , n66652 );
nand ( n78781 , n78779 , n78780 );
nand ( n78782 , n78781 , n71466 );
nand ( n78783 , n78776 , n78782 );
xor ( n78784 , n78773 , n78783 );
xor ( n78785 , n78756 , n78784 );
not ( n78786 , n71099 );
not ( n78787 , n78592 );
or ( n78788 , n78786 , n78787 );
not ( n78789 , n69695 );
not ( n78790 , n69961 );
or ( n78791 , n78789 , n78790 );
nand ( n78792 , n71577 , n76016 );
nand ( n78793 , n78791 , n78792 );
nand ( n78794 , n78793 , n59984 );
nand ( n78795 , n78788 , n78794 );
not ( n78796 , n72131 );
not ( n78797 , n78583 );
or ( n78798 , n78796 , n78797 );
not ( n78799 , n59341 );
not ( n78800 , n59914 );
or ( n78801 , n78799 , n78800 );
nand ( n78802 , n75548 , n66983 );
nand ( n78803 , n78801 , n78802 );
nand ( n78804 , n78803 , n75578 );
nand ( n78805 , n78798 , n78804 );
xor ( n78806 , n78795 , n78805 );
not ( n78807 , n77077 );
not ( n78808 , n78548 );
or ( n78809 , n78807 , n78808 );
not ( n78810 , n72083 );
not ( n78811 , n55630 );
or ( n78812 , n78810 , n78811 );
nand ( n78813 , n68980 , n76004 );
nand ( n78814 , n78812 , n78813 );
nand ( n78815 , n78814 , n67068 );
nand ( n78816 , n78809 , n78815 );
not ( n78817 , n78816 );
xor ( n78818 , n78806 , n78817 );
xor ( n78819 , n78746 , n78818 );
xor ( n78820 , n78819 , n78671 );
xor ( n78821 , n78785 , n78820 );
xor ( n78822 , n78821 , n78683 );
xor ( n78823 , n78755 , n78822 );
xor ( n78824 , n78691 , n78823 );
xor ( n78825 , n78824 , n78653 );
xor ( n78826 , n78691 , n78823 );
and ( n78827 , n78826 , n78653 );
and ( n78828 , n78691 , n78823 );
or ( n78829 , n78827 , n78828 );
xor ( n78830 , n78766 , n78772 );
and ( n78831 , n78830 , n78783 );
and ( n78832 , n78766 , n78772 );
or ( n78833 , n78831 , n78832 );
xor ( n78834 , n78795 , n78805 );
and ( n78835 , n78834 , n78817 );
and ( n78836 , n78795 , n78805 );
or ( n78837 , n78835 , n78836 );
xor ( n78838 , n78542 , n78565 );
and ( n78839 , n78838 , n78710 );
and ( n78840 , n78542 , n78565 );
or ( n78841 , n78839 , n78840 );
xor ( n78842 , n78663 , n78667 );
and ( n78843 , n78842 , n78784 );
and ( n78844 , n78663 , n78667 );
or ( n78845 , n78843 , n78844 );
xor ( n78846 , n78746 , n78818 );
and ( n78847 , n78846 , n78671 );
and ( n78848 , n78746 , n78818 );
or ( n78849 , n78847 , n78848 );
xor ( n78850 , n78675 , n78752 );
and ( n78851 , n78850 , n78679 );
and ( n78852 , n78675 , n78752 );
or ( n78853 , n78851 , n78852 );
xor ( n78854 , n78785 , n78820 );
and ( n78855 , n78854 , n78683 );
and ( n78856 , n78785 , n78820 );
or ( n78857 , n78855 , n78856 );
xor ( n78858 , n78754 , n78687 );
and ( n78859 , n78858 , n78822 );
and ( n78860 , n78754 , n78687 );
or ( n78861 , n78859 , n78860 );
not ( n78862 , n54326 );
not ( n78863 , n55161 );
or ( n78864 , n78862 , n78863 );
nand ( n78865 , n78864 , n71395 );
not ( n78866 , n72484 );
not ( n78867 , n78705 );
or ( n78868 , n78866 , n78867 );
not ( n78869 , n61540 );
not ( n78870 , n59651 );
or ( n78871 , n78869 , n78870 );
not ( n78872 , n71309 );
nand ( n78873 , n78872 , n75161 );
nand ( n78874 , n78871 , n78873 );
nand ( n78875 , n78874 , n61558 );
nand ( n78876 , n78868 , n78875 );
xor ( n78877 , n78865 , n78876 );
not ( n78878 , n75427 );
not ( n78879 , n72083 );
not ( n78880 , n70290 );
or ( n78881 , n78879 , n78880 );
nand ( n78882 , n67721 , n77344 );
nand ( n78883 , n78881 , n78882 );
not ( n78884 , n78883 );
or ( n78885 , n78878 , n78884 );
nand ( n78886 , n78814 , n77077 );
nand ( n78887 , n78885 , n78886 );
xor ( n78888 , n78877 , n78887 );
xor ( n78889 , n78865 , n78876 );
and ( n78890 , n78889 , n78887 );
and ( n78891 , n78865 , n78876 );
or ( n78892 , n78890 , n78891 );
not ( n78893 , n70964 );
xor ( n78894 , n67072 , n71829 );
not ( n78895 , n78894 );
or ( n78896 , n78893 , n78895 );
nand ( n78897 , n78695 , n65795 );
nand ( n78898 , n78896 , n78897 );
and ( n78899 , n66155 , n69409 );
xor ( n78900 , n78898 , n78899 );
not ( n78901 , n70183 );
not ( n78902 , n55120 );
not ( n78903 , n71876 );
or ( n78904 , n78902 , n78903 );
nand ( n78905 , n77783 , n71409 );
nand ( n78906 , n78904 , n78905 );
not ( n78907 , n78906 );
or ( n78908 , n78901 , n78907 );
nand ( n78909 , n78722 , n70193 );
nand ( n78910 , n78908 , n78909 );
xor ( n78911 , n78900 , n78910 );
xor ( n78912 , n78898 , n78899 );
and ( n78913 , n78912 , n78910 );
and ( n78914 , n78898 , n78899 );
or ( n78915 , n78913 , n78914 );
xor ( n78916 , n78911 , n78888 );
xor ( n78917 , n78916 , n78750 );
xor ( n78918 , n78917 , n78849 );
not ( n78919 , n55458 );
and ( n78920 , n71371 , n42400 );
not ( n78921 , n71371 );
and ( n78922 , n78921 , n71139 );
nor ( n78923 , n78920 , n78922 );
not ( n78924 , n78923 );
or ( n78925 , n78919 , n78924 );
nand ( n78926 , n78793 , n71099 );
nand ( n78927 , n78925 , n78926 );
not ( n78928 , n71466 );
and ( n78929 , n66652 , n76444 );
not ( n78930 , n66652 );
and ( n78931 , n78930 , n68667 );
nor ( n78932 , n78929 , n78931 );
not ( n78933 , n78932 );
or ( n78934 , n78928 , n78933 );
nand ( n78935 , n78781 , n75025 );
nand ( n78936 , n78934 , n78935 );
xor ( n78937 , n78927 , n78936 );
not ( n78938 , n75578 );
not ( n78939 , n72464 );
not ( n78940 , n43513 );
or ( n78941 , n78939 , n78940 );
nand ( n78942 , n60386 , n70920 );
nand ( n78943 , n78941 , n78942 );
not ( n78944 , n78943 );
or ( n78945 , n78938 , n78944 );
nand ( n78946 , n78803 , n72131 );
nand ( n78947 , n78945 , n78946 );
xor ( n78948 , n78937 , n78947 );
xor ( n78949 , n78837 , n78948 );
not ( n78950 , n70500 );
not ( n78951 , n78730 );
or ( n78952 , n78950 , n78951 );
and ( n78953 , n72477 , n59413 );
not ( n78954 , n72477 );
and ( n78955 , n78954 , n73268 );
or ( n78956 , n78953 , n78955 );
nand ( n78957 , n78956 , n70930 );
nand ( n78958 , n78952 , n78957 );
not ( n78959 , n56777 );
not ( n78960 , n78743 );
or ( n78961 , n78959 , n78960 );
not ( n78962 , n72589 );
not ( n78963 , n71176 );
or ( n78964 , n78962 , n78963 );
not ( n78965 , n76786 );
nand ( n78966 , n78965 , n39255 );
nand ( n78967 , n78964 , n78966 );
nand ( n78968 , n78967 , n72185 );
nand ( n78969 , n78961 , n78968 );
xor ( n78970 , n78958 , n78969 );
not ( n78971 , n72710 );
not ( n78972 , n67568 );
not ( n78973 , n62394 );
or ( n78974 , n78972 , n78973 );
nand ( n78975 , n72622 , n70608 );
nand ( n78976 , n78974 , n78975 );
not ( n78977 , n78976 );
or ( n78978 , n78971 , n78977 );
nand ( n78979 , n78764 , n72182 );
nand ( n78980 , n78978 , n78979 );
xor ( n78981 , n78970 , n78980 );
xor ( n78982 , n78949 , n78981 );
xor ( n78983 , n78918 , n78982 );
xor ( n78984 , n78816 , n78714 );
xor ( n78985 , n78984 , n78833 );
xor ( n78986 , n78985 , n78841 );
xor ( n78987 , n78986 , n78845 );
xor ( n78988 , n78987 , n78853 );
xor ( n78989 , n78988 , n78857 );
xor ( n78990 , n78983 , n78989 );
xor ( n78991 , n78990 , n78861 );
xor ( n78992 , n78983 , n78989 );
and ( n78993 , n78992 , n78861 );
and ( n78994 , n78983 , n78989 );
or ( n78995 , n78993 , n78994 );
xor ( n78996 , n78958 , n78969 );
and ( n78997 , n78996 , n78980 );
and ( n78998 , n78958 , n78969 );
or ( n78999 , n78997 , n78998 );
xor ( n79000 , n78927 , n78936 );
and ( n79001 , n79000 , n78947 );
and ( n79002 , n78927 , n78936 );
or ( n79003 , n79001 , n79002 );
xor ( n79004 , n78816 , n78714 );
and ( n79005 , n79004 , n78833 );
and ( n79006 , n78816 , n78714 );
or ( n79007 , n79005 , n79006 );
xor ( n79008 , n78911 , n78888 );
and ( n79009 , n79008 , n78750 );
and ( n79010 , n78911 , n78888 );
or ( n79011 , n79009 , n79010 );
xor ( n79012 , n78837 , n78948 );
and ( n79013 , n79012 , n78981 );
and ( n79014 , n78837 , n78948 );
or ( n79015 , n79013 , n79014 );
xor ( n79016 , n78985 , n78841 );
and ( n79017 , n79016 , n78845 );
and ( n79018 , n78985 , n78841 );
or ( n79019 , n79017 , n79018 );
xor ( n79020 , n78917 , n78849 );
and ( n79021 , n79020 , n78982 );
and ( n79022 , n78917 , n78849 );
or ( n79023 , n79021 , n79022 );
xor ( n79024 , n78987 , n78853 );
and ( n79025 , n79024 , n78857 );
and ( n79026 , n78987 , n78853 );
or ( n79027 , n79025 , n79026 );
and ( n79028 , n66155 , n68990 );
and ( n79029 , n63180 , n72083 );
not ( n79030 , n63180 );
and ( n79031 , n79030 , n77344 );
or ( n79032 , n79029 , n79031 );
not ( n79033 , n79032 );
not ( n79034 , n75427 );
or ( n79035 , n79033 , n79034 );
nand ( n79036 , n77077 , n78883 );
nand ( n79037 , n79035 , n79036 );
xor ( n79038 , n79028 , n79037 );
not ( n79039 , n71099 );
not ( n79040 , n78923 );
or ( n79041 , n79039 , n79040 );
not ( n79042 , n69695 );
not ( n79043 , n77972 );
or ( n79044 , n79042 , n79043 );
nand ( n79045 , n42556 , n69237 );
nand ( n79046 , n79044 , n79045 );
nand ( n79047 , n79046 , n59984 );
nand ( n79048 , n79041 , n79047 );
xor ( n79049 , n79038 , n79048 );
xor ( n79050 , n79028 , n79037 );
and ( n79051 , n79050 , n79048 );
and ( n79052 , n79028 , n79037 );
or ( n79053 , n79051 , n79052 );
not ( n79054 , n61558 );
not ( n79055 , n71309 );
not ( n79056 , n75594 );
or ( n79057 , n79055 , n79056 );
nand ( n79058 , n66215 , n77333 );
nand ( n79059 , n79057 , n79058 );
not ( n79060 , n79059 );
or ( n79061 , n79054 , n79060 );
nand ( n79062 , n78874 , n75753 );
nand ( n79063 , n79061 , n79062 );
not ( n79064 , n72710 );
and ( n79065 , n76811 , n39334 );
not ( n79066 , n76811 );
not ( n79067 , n39334 );
and ( n79068 , n79066 , n79067 );
nor ( n79069 , n79065 , n79068 );
not ( n79070 , n79069 );
or ( n79071 , n79064 , n79070 );
nand ( n79072 , n78976 , n72182 );
nand ( n79073 , n79071 , n79072 );
xor ( n79074 , n79063 , n79073 );
not ( n79075 , n76828 );
not ( n79076 , n78932 );
or ( n79077 , n79075 , n79076 );
not ( n79078 , n65184 );
not ( n79079 , n59891 );
or ( n79080 , n79078 , n79079 );
nand ( n79081 , n71547 , n65183 );
nand ( n79082 , n79080 , n79081 );
nand ( n79083 , n79082 , n71466 );
nand ( n79084 , n79077 , n79083 );
xor ( n79085 , n79074 , n79084 );
xor ( n79086 , n79063 , n79073 );
and ( n79087 , n79086 , n79084 );
and ( n79088 , n79063 , n79073 );
or ( n79089 , n79087 , n79088 );
not ( n79090 , n55144 );
not ( n79091 , n78906 );
or ( n79092 , n79090 , n79091 );
nand ( n79093 , n70183 , n72919 );
nand ( n79094 , n79092 , n79093 );
not ( n79095 , n56777 );
not ( n79096 , n78967 );
or ( n79097 , n79095 , n79096 );
not ( n79098 , n72589 );
not ( n79099 , n69961 );
or ( n79100 , n79098 , n79099 );
nand ( n79101 , n69962 , n71362 );
nand ( n79102 , n79100 , n79101 );
nand ( n79103 , n79102 , n72185 );
nand ( n79104 , n79097 , n79103 );
xor ( n79105 , n79094 , n79104 );
not ( n79106 , n75578 );
not ( n79107 , n70920 );
not ( n79108 , n79107 );
not ( n79109 , n58933 );
or ( n79110 , n79108 , n79109 );
nand ( n79111 , n39714 , n70920 );
nand ( n79112 , n79110 , n79111 );
not ( n79113 , n79112 );
or ( n79114 , n79106 , n79113 );
nand ( n79115 , n78943 , n72131 );
nand ( n79116 , n79114 , n79115 );
xor ( n79117 , n79105 , n79116 );
xor ( n79118 , n79094 , n79104 );
and ( n79119 , n79118 , n79116 );
and ( n79120 , n79094 , n79104 );
or ( n79121 , n79119 , n79120 );
not ( n79122 , n70500 );
not ( n79123 , n78956 );
or ( n79124 , n79122 , n79123 );
not ( n79125 , n70506 );
not ( n79126 , n67040 );
or ( n79127 , n79125 , n79126 );
nand ( n79128 , n76082 , n78148 );
nand ( n79129 , n79127 , n79128 );
nand ( n79130 , n79129 , n70930 );
nand ( n79131 , n79124 , n79130 );
not ( n79132 , n71960 );
not ( n79133 , n78894 );
or ( n79134 , n79132 , n79133 );
xor ( n79135 , n71971 , n72217 );
nand ( n79136 , n79135 , n70964 );
nand ( n79137 , n79134 , n79136 );
not ( n79138 , n79137 );
xor ( n79139 , n79131 , n79138 );
xor ( n79140 , n79139 , n78892 );
xor ( n79141 , n79131 , n79138 );
and ( n79142 , n79141 , n78892 );
and ( n79143 , n79131 , n79138 );
or ( n79144 , n79142 , n79143 );
xor ( n79145 , n79003 , n79049 );
xor ( n79146 , n79145 , n78999 );
xor ( n79147 , n79003 , n79049 );
and ( n79148 , n79147 , n78999 );
and ( n79149 , n79003 , n79049 );
or ( n79150 , n79148 , n79149 );
xor ( n79151 , n78915 , n79085 );
xor ( n79152 , n79151 , n79117 );
xor ( n79153 , n78915 , n79085 );
and ( n79154 , n79153 , n79117 );
and ( n79155 , n78915 , n79085 );
or ( n79156 , n79154 , n79155 );
xor ( n79157 , n79140 , n79007 );
xor ( n79158 , n79157 , n79011 );
xor ( n79159 , n79140 , n79007 );
and ( n79160 , n79159 , n79011 );
and ( n79161 , n79140 , n79007 );
or ( n79162 , n79160 , n79161 );
xor ( n79163 , n79015 , n79146 );
xor ( n79164 , n79163 , n79152 );
xor ( n79165 , n79015 , n79146 );
and ( n79166 , n79165 , n79152 );
and ( n79167 , n79015 , n79146 );
or ( n79168 , n79166 , n79167 );
xor ( n79169 , n79019 , n79158 );
xor ( n79170 , n79169 , n79023 );
xor ( n79171 , n79019 , n79158 );
and ( n79172 , n79171 , n79023 );
and ( n79173 , n79019 , n79158 );
or ( n79174 , n79172 , n79173 );
xor ( n79175 , n79164 , n79170 );
xor ( n79176 , n79175 , n79027 );
xor ( n79177 , n79164 , n79170 );
and ( n79178 , n79177 , n79027 );
and ( n79179 , n79164 , n79170 );
or ( n79180 , n79178 , n79179 );
not ( n79181 , n72562 );
not ( n79182 , n68334 );
or ( n79183 , n79181 , n79182 );
nand ( n79184 , n79183 , n72919 );
not ( n79185 , n77077 );
not ( n79186 , n79032 );
or ( n79187 , n79185 , n79186 );
not ( n79188 , n72083 );
not ( n79189 , n59651 );
or ( n79190 , n79188 , n79189 );
nand ( n79191 , n75161 , n77344 );
nand ( n79192 , n79190 , n79191 );
nand ( n79193 , n79192 , n75427 );
nand ( n79194 , n79187 , n79193 );
xor ( n79195 , n79184 , n79194 );
not ( n79196 , n70964 );
xor ( n79197 , n66155 , n67721 );
not ( n79198 , n79197 );
or ( n79199 , n79196 , n79198 );
nand ( n79200 , n79135 , n71960 );
nand ( n79201 , n79199 , n79200 );
xor ( n79202 , n79195 , n79201 );
xor ( n79203 , n79184 , n79194 );
and ( n79204 , n79203 , n79201 );
and ( n79205 , n79184 , n79194 );
or ( n79206 , n79204 , n79205 );
and ( n79207 , n67072 , n71829 );
not ( n79208 , n59984 );
not ( n79209 , n69695 );
not ( n79210 , n78219 );
not ( n79211 , n79210 );
or ( n79212 , n79209 , n79211 );
nand ( n79213 , n42656 , n74094 );
nand ( n79214 , n79212 , n79213 );
not ( n79215 , n79214 );
or ( n79216 , n79208 , n79215 );
nand ( n79217 , n79046 , n71099 );
nand ( n79218 , n79216 , n79217 );
xor ( n79219 , n79207 , n79218 );
not ( n79220 , n72484 );
not ( n79221 , n79059 );
or ( n79222 , n79220 , n79221 );
not ( n79223 , n71309 );
not ( n79224 , n39895 );
or ( n79225 , n79223 , n79224 );
nand ( n79226 , n39896 , n77333 );
nand ( n79227 , n79225 , n79226 );
nand ( n79228 , n79227 , n61558 );
nand ( n79229 , n79222 , n79228 );
xor ( n79230 , n79219 , n79229 );
xor ( n79231 , n79207 , n79218 );
and ( n79232 , n79231 , n79229 );
and ( n79233 , n79207 , n79218 );
or ( n79234 , n79232 , n79233 );
not ( n79235 , n72961 );
not ( n79236 , n79069 );
or ( n79237 , n79235 , n79236 );
not ( n79238 , n67568 );
not ( n79239 , n71176 );
or ( n79240 , n79238 , n79239 );
nand ( n79241 , n39255 , n76811 );
nand ( n79242 , n79240 , n79241 );
nand ( n79243 , n79242 , n72710 );
nand ( n79244 , n79237 , n79243 );
not ( n79245 , n71466 );
not ( n79246 , n72622 );
and ( n79247 , n65183 , n79246 );
not ( n79248 , n65183 );
and ( n79249 , n79248 , n72622 );
nor ( n79250 , n79247 , n79249 );
not ( n79251 , n79250 );
or ( n79252 , n79245 , n79251 );
nand ( n79253 , n79082 , n75025 );
nand ( n79254 , n79252 , n79253 );
xor ( n79255 , n79244 , n79254 );
not ( n79256 , n72185 );
not ( n79257 , n72589 );
not ( n79258 , n76455 );
or ( n79259 , n79257 , n79258 );
nand ( n79260 , n76454 , n71362 );
nand ( n79261 , n79259 , n79260 );
not ( n79262 , n79261 );
or ( n79263 , n79256 , n79262 );
nand ( n79264 , n79102 , n56777 );
nand ( n79265 , n79263 , n79264 );
xor ( n79266 , n79255 , n79265 );
xor ( n79267 , n79244 , n79254 );
and ( n79268 , n79267 , n79265 );
and ( n79269 , n79244 , n79254 );
or ( n79270 , n79268 , n79269 );
not ( n79271 , n75578 );
and ( n79272 , n70920 , n76444 );
not ( n79273 , n70920 );
and ( n79274 , n79273 , n39575 );
nor ( n79275 , n79272 , n79274 );
not ( n79276 , n79275 );
or ( n79277 , n79271 , n79276 );
nand ( n79278 , n79112 , n72131 );
nand ( n79279 , n79277 , n79278 );
buf ( n79280 , n70930 );
not ( n79281 , n79280 );
not ( n79282 , n70506 );
not ( n79283 , n43513 );
or ( n79284 , n79282 , n79283 );
nand ( n79285 , n72477 , n39681 );
nand ( n79286 , n79284 , n79285 );
not ( n79287 , n79286 );
or ( n79288 , n79281 , n79287 );
nand ( n79289 , n79129 , n70500 );
nand ( n79290 , n79288 , n79289 );
xor ( n79291 , n79279 , n79290 );
xor ( n79292 , n79291 , n79137 );
xor ( n79293 , n79279 , n79290 );
and ( n79294 , n79293 , n79137 );
and ( n79295 , n79279 , n79290 );
or ( n79296 , n79294 , n79295 );
xor ( n79297 , n79202 , n79121 );
xor ( n79298 , n79297 , n79053 );
xor ( n79299 , n79202 , n79121 );
and ( n79300 , n79299 , n79053 );
and ( n79301 , n79202 , n79121 );
or ( n79302 , n79300 , n79301 );
xor ( n79303 , n79089 , n79230 );
xor ( n79304 , n79303 , n79266 );
xor ( n79305 , n79089 , n79230 );
and ( n79306 , n79305 , n79266 );
and ( n79307 , n79089 , n79230 );
or ( n79308 , n79306 , n79307 );
xor ( n79309 , n79292 , n79144 );
xor ( n79310 , n79309 , n79150 );
xor ( n79311 , n79292 , n79144 );
and ( n79312 , n79311 , n79150 );
and ( n79313 , n79292 , n79144 );
or ( n79314 , n79312 , n79313 );
xor ( n79315 , n79156 , n79298 );
xor ( n79316 , n79315 , n79304 );
xor ( n79317 , n79156 , n79298 );
and ( n79318 , n79317 , n79304 );
and ( n79319 , n79156 , n79298 );
or ( n79320 , n79318 , n79319 );
xor ( n79321 , n79162 , n79310 );
xor ( n79322 , n79321 , n79168 );
xor ( n79323 , n79162 , n79310 );
and ( n79324 , n79323 , n79168 );
and ( n79325 , n79162 , n79310 );
or ( n79326 , n79324 , n79325 );
xor ( n79327 , n79316 , n79322 );
xor ( n79328 , n79327 , n79174 );
xor ( n79329 , n79316 , n79322 );
and ( n79330 , n79329 , n79174 );
and ( n79331 , n79316 , n79322 );
or ( n79332 , n79330 , n79331 );
and ( n79333 , n71971 , n72217 );
not ( n79334 , n56777 );
not ( n79335 , n79261 );
or ( n79336 , n79334 , n79335 );
not ( n79337 , n72589 );
not ( n79338 , n77972 );
or ( n79339 , n79337 , n79338 );
nand ( n79340 , n42556 , n71362 );
nand ( n79341 , n79339 , n79340 );
nand ( n79342 , n79341 , n72185 );
nand ( n79343 , n79336 , n79342 );
xor ( n79344 , n79333 , n79343 );
not ( n79345 , n75427 );
not ( n79346 , n72083 );
not ( n79347 , n39846 );
or ( n79348 , n79346 , n79347 );
nand ( n79349 , n39847 , n77344 );
nand ( n79350 , n79348 , n79349 );
not ( n79351 , n79350 );
or ( n79352 , n79345 , n79351 );
nand ( n79353 , n79192 , n77077 );
nand ( n79354 , n79352 , n79353 );
xor ( n79355 , n79344 , n79354 );
xor ( n79356 , n79333 , n79343 );
and ( n79357 , n79356 , n79354 );
and ( n79358 , n79333 , n79343 );
or ( n79359 , n79357 , n79358 );
not ( n79360 , n75025 );
not ( n79361 , n79250 );
or ( n79362 , n79360 , n79361 );
not ( n79363 , n65184 );
not ( n79364 , n39334 );
or ( n79365 , n79363 , n79364 );
nand ( n79366 , n79067 , n65183 );
nand ( n79367 , n79365 , n79366 );
nand ( n79368 , n79367 , n71466 );
nand ( n79369 , n79362 , n79368 );
not ( n79370 , n72131 );
not ( n79371 , n79275 );
or ( n79372 , n79370 , n79371 );
and ( n79373 , n59891 , n79107 );
not ( n79374 , n59891 );
and ( n79375 , n79374 , n70920 );
or ( n79376 , n79373 , n79375 );
nand ( n79377 , n79376 , n75578 );
nand ( n79378 , n79372 , n79377 );
xor ( n79379 , n79369 , n79378 );
not ( n79380 , n71099 );
not ( n79381 , n79214 );
or ( n79382 , n79380 , n79381 );
nand ( n79383 , n59984 , n69695 );
nand ( n79384 , n79382 , n79383 );
xor ( n79385 , n79379 , n79384 );
xor ( n79386 , n79369 , n79378 );
and ( n79387 , n79386 , n79384 );
and ( n79388 , n79369 , n79378 );
or ( n79389 , n79387 , n79388 );
not ( n79390 , n72961 );
not ( n79391 , n79242 );
or ( n79392 , n79390 , n79391 );
not ( n79393 , n67568 );
not ( n79394 , n69961 );
or ( n79395 , n79393 , n79394 );
nand ( n79396 , n69962 , n70608 );
nand ( n79397 , n79395 , n79396 );
nand ( n79398 , n79397 , n72710 );
nand ( n79399 , n79392 , n79398 );
not ( n79400 , n70500 );
not ( n79401 , n79286 );
or ( n79402 , n79400 , n79401 );
not ( n79403 , n75286 );
not ( n79404 , n39715 );
or ( n79405 , n79403 , n79404 );
not ( n79406 , n58933 );
nand ( n79407 , n79406 , n78148 );
nand ( n79408 , n79405 , n79407 );
nand ( n79409 , n79408 , n79280 );
nand ( n79410 , n79402 , n79409 );
xor ( n79411 , n79399 , n79410 );
not ( n79412 , n72484 );
not ( n79413 , n79227 );
or ( n79414 , n79412 , n79413 );
not ( n79415 , n71309 );
not ( n79416 , n74900 );
or ( n79417 , n79415 , n79416 );
nand ( n79418 , n76082 , n77333 );
nand ( n79419 , n79417 , n79418 );
nand ( n79420 , n79419 , n61558 );
nand ( n79421 , n79414 , n79420 );
xor ( n79422 , n79411 , n79421 );
xor ( n79423 , n79399 , n79410 );
and ( n79424 , n79423 , n79421 );
and ( n79425 , n79399 , n79410 );
or ( n79426 , n79424 , n79425 );
not ( n79427 , n71960 );
not ( n79428 , n79197 );
or ( n79429 , n79427 , n79428 );
and ( n79430 , n71971 , n77575 );
not ( n79431 , n71971 );
and ( n79432 , n79431 , n70653 );
or ( n79433 , n79430 , n79432 );
nand ( n79434 , n79433 , n70964 );
nand ( n79435 , n79429 , n79434 );
not ( n79436 , n79435 );
xor ( n79437 , n79436 , n79206 );
xor ( n79438 , n79437 , n79234 );
xor ( n79439 , n79436 , n79206 );
and ( n79440 , n79439 , n79234 );
and ( n79441 , n79436 , n79206 );
or ( n79442 , n79440 , n79441 );
xor ( n79443 , n79270 , n79355 );
xor ( n79444 , n79443 , n79385 );
xor ( n79445 , n79270 , n79355 );
and ( n79446 , n79445 , n79385 );
and ( n79447 , n79270 , n79355 );
or ( n79448 , n79446 , n79447 );
xor ( n79449 , n79422 , n79296 );
xor ( n79450 , n79449 , n79302 );
xor ( n79451 , n79422 , n79296 );
and ( n79452 , n79451 , n79302 );
and ( n79453 , n79422 , n79296 );
or ( n79454 , n79452 , n79453 );
xor ( n79455 , n79438 , n79308 );
xor ( n79456 , n79455 , n79444 );
xor ( n79457 , n79438 , n79308 );
and ( n79458 , n79457 , n79444 );
and ( n79459 , n79438 , n79308 );
or ( n79460 , n79458 , n79459 );
xor ( n79461 , n79450 , n79314 );
xor ( n79462 , n79461 , n79320 );
xor ( n79463 , n79450 , n79314 );
and ( n79464 , n79463 , n79320 );
and ( n79465 , n79450 , n79314 );
or ( n79466 , n79464 , n79465 );
xor ( n79467 , n79456 , n79462 );
xor ( n79468 , n79467 , n79326 );
xor ( n79469 , n79456 , n79462 );
and ( n79470 , n79469 , n79326 );
and ( n79471 , n79456 , n79462 );
or ( n79472 , n79470 , n79471 );
not ( n79473 , n58066 );
not ( n79474 , n69028 );
or ( n79475 , n79473 , n79474 );
nand ( n79476 , n79475 , n69695 );
not ( n79477 , n71960 );
not ( n79478 , n79433 );
or ( n79479 , n79477 , n79478 );
xor ( n79480 , n72846 , n62618 );
nand ( n79481 , n79480 , n70964 );
nand ( n79482 , n79479 , n79481 );
xor ( n79483 , n79476 , n79482 );
and ( n79484 , n66155 , n67721 );
xor ( n79485 , n79483 , n79484 );
xor ( n79486 , n79476 , n79482 );
and ( n79487 , n79486 , n79484 );
and ( n79488 , n79476 , n79482 );
or ( n79489 , n79487 , n79488 );
not ( n79490 , n72185 );
not ( n79491 , n72589 );
not ( n79492 , n79210 );
or ( n79493 , n79491 , n79492 );
buf ( n79494 , n77783 );
nand ( n79495 , n79494 , n71362 );
nand ( n79496 , n79493 , n79495 );
not ( n79497 , n79496 );
or ( n79498 , n79490 , n79497 );
nand ( n79499 , n79341 , n56777 );
nand ( n79500 , n79498 , n79499 );
not ( n79501 , n77077 );
not ( n79502 , n79350 );
or ( n79503 , n79501 , n79502 );
and ( n79504 , n72083 , n39895 );
not ( n79505 , n72083 );
and ( n79506 , n79505 , n39896 );
or ( n79507 , n79504 , n79506 );
nand ( n79508 , n79507 , n75427 );
nand ( n79509 , n79503 , n79508 );
xor ( n79510 , n79500 , n79509 );
not ( n79511 , n71466 );
not ( n79512 , n65184 );
not ( n79513 , n39254 );
or ( n79514 , n79512 , n79513 );
nand ( n79515 , n39255 , n65183 );
nand ( n79516 , n79514 , n79515 );
not ( n79517 , n79516 );
or ( n79518 , n79511 , n79517 );
nand ( n79519 , n79367 , n75025 );
nand ( n79520 , n79518 , n79519 );
xor ( n79521 , n79510 , n79520 );
xor ( n79522 , n79500 , n79509 );
and ( n79523 , n79522 , n79520 );
and ( n79524 , n79500 , n79509 );
or ( n79525 , n79523 , n79524 );
not ( n79526 , n75578 );
and ( n79527 , n70920 , n79246 );
not ( n79528 , n70920 );
and ( n79529 , n79528 , n72622 );
nor ( n79530 , n79527 , n79529 );
not ( n79531 , n79530 );
or ( n79532 , n79526 , n79531 );
nand ( n79533 , n79376 , n72131 );
nand ( n79534 , n79532 , n79533 );
not ( n79535 , n72710 );
and ( n79536 , n70608 , n76455 );
not ( n79537 , n70608 );
and ( n79538 , n79537 , n76454 );
nor ( n79539 , n79536 , n79538 );
not ( n79540 , n79539 );
or ( n79541 , n79535 , n79540 );
nand ( n79542 , n79397 , n72961 );
nand ( n79543 , n79541 , n79542 );
xor ( n79544 , n79534 , n79543 );
not ( n79545 , n79280 );
not ( n79546 , n70506 );
not ( n79547 , n39575 );
not ( n79548 , n79547 );
or ( n79549 , n79546 , n79548 );
nand ( n79550 , n39575 , n78148 );
nand ( n79551 , n79549 , n79550 );
not ( n79552 , n79551 );
or ( n79553 , n79545 , n79552 );
nand ( n79554 , n79408 , n70500 );
nand ( n79555 , n79553 , n79554 );
xor ( n79556 , n79544 , n79555 );
xor ( n79557 , n79534 , n79543 );
and ( n79558 , n79557 , n79555 );
and ( n79559 , n79534 , n79543 );
or ( n79560 , n79558 , n79559 );
not ( n79561 , n61558 );
and ( n79562 , n71309 , n39681 );
not ( n79563 , n71309 );
and ( n79564 , n79563 , n43513 );
nor ( n79565 , n79562 , n79564 );
not ( n79566 , n79565 );
or ( n79567 , n79561 , n79566 );
nand ( n79568 , n79419 , n72484 );
nand ( n79569 , n79567 , n79568 );
xor ( n79570 , n79569 , n79435 );
xor ( n79571 , n79570 , n79485 );
xor ( n79572 , n79569 , n79435 );
and ( n79573 , n79572 , n79485 );
and ( n79574 , n79569 , n79435 );
or ( n79575 , n79573 , n79574 );
xor ( n79576 , n79359 , n79389 );
xor ( n79577 , n79576 , n79426 );
xor ( n79578 , n79359 , n79389 );
and ( n79579 , n79578 , n79426 );
and ( n79580 , n79359 , n79389 );
or ( n79581 , n79579 , n79580 );
xor ( n79582 , n79556 , n79521 );
xor ( n79583 , n79582 , n79442 );
xor ( n79584 , n79556 , n79521 );
and ( n79585 , n79584 , n79442 );
and ( n79586 , n79556 , n79521 );
or ( n79587 , n79585 , n79586 );
xor ( n79588 , n79571 , n79577 );
xor ( n79589 , n79588 , n79448 );
xor ( n79590 , n79571 , n79577 );
and ( n79591 , n79590 , n79448 );
and ( n79592 , n79571 , n79577 );
or ( n79593 , n79591 , n79592 );
xor ( n79594 , n79583 , n79454 );
xor ( n79595 , n79594 , n79460 );
xor ( n79596 , n79583 , n79454 );
and ( n79597 , n79596 , n79460 );
and ( n79598 , n79583 , n79454 );
or ( n79599 , n79597 , n79598 );
xor ( n79600 , n79589 , n79595 );
xor ( n79601 , n79600 , n79466 );
xor ( n79602 , n79589 , n79595 );
and ( n79603 , n79602 , n79466 );
and ( n79604 , n79589 , n79595 );
or ( n79605 , n79603 , n79604 );
not ( n79606 , n72961 );
not ( n79607 , n79539 );
or ( n79608 , n79606 , n79607 );
not ( n79609 , n67568 );
not ( n79610 , n77972 );
or ( n79611 , n79609 , n79610 );
not ( n79612 , n77972 );
nand ( n79613 , n79612 , n70608 );
nand ( n79614 , n79611 , n79613 );
nand ( n79615 , n79614 , n72710 );
nand ( n79616 , n79608 , n79615 );
not ( n79617 , n70964 );
xor ( n79618 , n66581 , n39847 );
not ( n79619 , n79618 );
or ( n79620 , n79617 , n79619 );
nand ( n79621 , n79480 , n71960 );
nand ( n79622 , n79620 , n79621 );
xor ( n79623 , n79616 , n79622 );
not ( n79624 , n72131 );
not ( n79625 , n79530 );
or ( n79626 , n79624 , n79625 );
not ( n79627 , n79107 );
not ( n79628 , n39334 );
or ( n79629 , n79627 , n79628 );
nand ( n79630 , n79067 , n70920 );
nand ( n79631 , n79629 , n79630 );
nand ( n79632 , n79631 , n75578 );
nand ( n79633 , n79626 , n79632 );
xor ( n79634 , n79623 , n79633 );
xor ( n79635 , n79616 , n79622 );
and ( n79636 , n79635 , n79633 );
and ( n79637 , n79616 , n79622 );
or ( n79638 , n79636 , n79637 );
not ( n79639 , n56777 );
not ( n79640 , n79496 );
or ( n79641 , n79639 , n79640 );
nand ( n79642 , n72185 , n72589 );
nand ( n79643 , n79641 , n79642 );
not ( n79644 , n70500 );
not ( n79645 , n79551 );
or ( n79646 , n79644 , n79645 );
and ( n79647 , n75286 , n71547 );
not ( n79648 , n75286 );
and ( n79649 , n79648 , n59891 );
nor ( n79650 , n79647 , n79649 );
nand ( n79651 , n79650 , n79280 );
nand ( n79652 , n79646 , n79651 );
xor ( n79653 , n79643 , n79652 );
not ( n79654 , n75025 );
not ( n79655 , n79516 );
or ( n79656 , n79654 , n79655 );
not ( n79657 , n65184 );
not ( n79658 , n69961 );
or ( n79659 , n79657 , n79658 );
nand ( n79660 , n69962 , n65183 );
nand ( n79661 , n79659 , n79660 );
not ( n79662 , n79661 );
or ( n79663 , n79662 , n71467 );
nand ( n79664 , n79656 , n79663 );
xor ( n79665 , n79653 , n79664 );
xor ( n79666 , n79643 , n79652 );
and ( n79667 , n79666 , n79664 );
and ( n79668 , n79643 , n79652 );
or ( n79669 , n79667 , n79668 );
not ( n79670 , n72484 );
not ( n79671 , n79565 );
or ( n79672 , n79670 , n79671 );
not ( n79673 , n71309 );
not ( n79674 , n39715 );
or ( n79675 , n79673 , n79674 );
nand ( n79676 , n39716 , n77333 );
nand ( n79677 , n79675 , n79676 );
nand ( n79678 , n79677 , n61558 );
nand ( n79679 , n79672 , n79678 );
not ( n79680 , n77077 );
not ( n79681 , n79507 );
or ( n79682 , n79680 , n79681 );
and ( n79683 , n72083 , n76082 );
not ( n79684 , n72083 );
and ( n79685 , n79684 , n74900 );
nor ( n79686 , n79683 , n79685 );
nand ( n79687 , n79686 , n75427 );
nand ( n79688 , n79682 , n79687 );
xor ( n79689 , n79679 , n79688 );
nand ( n79690 , n70653 , n67072 );
xor ( n79691 , n79689 , n79690 );
xor ( n79692 , n79679 , n79688 );
and ( n79693 , n79692 , n79690 );
and ( n79694 , n79679 , n79688 );
or ( n79695 , n79693 , n79694 );
xor ( n79696 , n79489 , n79525 );
xor ( n79697 , n79696 , n79560 );
xor ( n79698 , n79489 , n79525 );
and ( n79699 , n79698 , n79560 );
and ( n79700 , n79489 , n79525 );
or ( n79701 , n79699 , n79700 );
xor ( n79702 , n79634 , n79691 );
xor ( n79703 , n79702 , n79665 );
xor ( n79704 , n79634 , n79691 );
and ( n79705 , n79704 , n79665 );
and ( n79706 , n79634 , n79691 );
or ( n79707 , n79705 , n79706 );
xor ( n79708 , n79581 , n79575 );
xor ( n79709 , n79708 , n79697 );
xor ( n79710 , n79581 , n79575 );
and ( n79711 , n79710 , n79697 );
and ( n79712 , n79581 , n79575 );
or ( n79713 , n79711 , n79712 );
xor ( n79714 , n79703 , n79587 );
xor ( n79715 , n79714 , n79593 );
xor ( n79716 , n79703 , n79587 );
and ( n79717 , n79716 , n79593 );
and ( n79718 , n79703 , n79587 );
or ( n79719 , n79717 , n79718 );
xor ( n79720 , n79709 , n79715 );
xor ( n79721 , n79720 , n79599 );
xor ( n79722 , n79709 , n79715 );
and ( n79723 , n79722 , n79599 );
and ( n79724 , n79709 , n79715 );
or ( n79725 , n79723 , n79724 );
or ( n79726 , n72185 , n56777 );
nand ( n79727 , n79726 , n72589 );
and ( n79728 , n72846 , n62618 );
xor ( n79729 , n79727 , n79728 );
not ( n79730 , n72710 );
not ( n79731 , n67568 );
not ( n79732 , n79210 );
or ( n79733 , n79731 , n79732 );
nand ( n79734 , n79494 , n70608 );
nand ( n79735 , n79733 , n79734 );
not ( n79736 , n79735 );
or ( n79737 , n79730 , n79736 );
nand ( n79738 , n79614 , n72961 );
nand ( n79739 , n79737 , n79738 );
xor ( n79740 , n79729 , n79739 );
xor ( n79741 , n79727 , n79728 );
and ( n79742 , n79741 , n79739 );
and ( n79743 , n79727 , n79728 );
or ( n79744 , n79742 , n79743 );
not ( n79745 , n71960 );
not ( n79746 , n79618 );
or ( n79747 , n79745 , n79746 );
xor ( n79748 , n66581 , n43609 );
nand ( n79749 , n79748 , n70964 );
nand ( n79750 , n79747 , n79749 );
not ( n79751 , n72131 );
not ( n79752 , n79631 );
or ( n79753 , n79751 , n79752 );
not ( n79754 , n79107 );
not ( n79755 , n39254 );
or ( n79756 , n79754 , n79755 );
nand ( n79757 , n70920 , n39255 );
nand ( n79758 , n79756 , n79757 );
nand ( n79759 , n79758 , n75578 );
nand ( n79760 , n79753 , n79759 );
xor ( n79761 , n79750 , n79760 );
not ( n79762 , n70500 );
not ( n79763 , n79650 );
or ( n79764 , n79762 , n79763 );
and ( n79765 , n72477 , n72622 );
not ( n79766 , n72477 );
and ( n79767 , n79766 , n79246 );
nor ( n79768 , n79765 , n79767 );
not ( n79769 , n79280 );
or ( n79770 , n79768 , n79769 );
nand ( n79771 , n79764 , n79770 );
xor ( n79772 , n79761 , n79771 );
xor ( n79773 , n79750 , n79760 );
and ( n79774 , n79773 , n79771 );
and ( n79775 , n79750 , n79760 );
or ( n79776 , n79774 , n79775 );
not ( n79777 , n71466 );
not ( n79778 , n65184 );
not ( n79779 , n76455 );
or ( n79780 , n79778 , n79779 );
nand ( n79781 , n76454 , n65183 );
nand ( n79782 , n79780 , n79781 );
not ( n79783 , n79782 );
or ( n79784 , n79777 , n79783 );
nand ( n79785 , n79661 , n75025 );
nand ( n79786 , n79784 , n79785 );
not ( n79787 , n72484 );
not ( n79788 , n79677 );
or ( n79789 , n79787 , n79788 );
not ( n79790 , n71309 );
not ( n79791 , n79547 );
or ( n79792 , n79790 , n79791 );
nand ( n79793 , n77333 , n39575 );
nand ( n79794 , n79792 , n79793 );
nand ( n79795 , n79794 , n61558 );
nand ( n79796 , n79789 , n79795 );
xor ( n79797 , n79786 , n79796 );
not ( n79798 , n77077 );
not ( n79799 , n79686 );
or ( n79800 , n79798 , n79799 );
and ( n79801 , n72083 , n43513 );
not ( n79802 , n72083 );
and ( n79803 , n79802 , n39681 );
nor ( n79804 , n79801 , n79803 );
not ( n79805 , n79804 );
nand ( n79806 , n79805 , n75427 );
nand ( n79807 , n79800 , n79806 );
xor ( n79808 , n79797 , n79807 );
xor ( n79809 , n79786 , n79796 );
and ( n79810 , n79809 , n79807 );
and ( n79811 , n79786 , n79796 );
or ( n79812 , n79810 , n79811 );
not ( n79813 , n79690 );
xor ( n79814 , n79813 , n79740 );
xor ( n79815 , n79814 , n79638 );
xor ( n79816 , n79813 , n79740 );
and ( n79817 , n79816 , n79638 );
and ( n79818 , n79813 , n79740 );
or ( n79819 , n79817 , n79818 );
xor ( n79820 , n79669 , n79808 );
xor ( n79821 , n79820 , n79695 );
xor ( n79822 , n79669 , n79808 );
and ( n79823 , n79822 , n79695 );
and ( n79824 , n79669 , n79808 );
or ( n79825 , n79823 , n79824 );
xor ( n79826 , n79772 , n79701 );
xor ( n79827 , n79826 , n79815 );
xor ( n79828 , n79772 , n79701 );
and ( n79829 , n79828 , n79815 );
and ( n79830 , n79772 , n79701 );
or ( n79831 , n79829 , n79830 );
xor ( n79832 , n79707 , n79821 );
xor ( n79833 , n79832 , n79827 );
xor ( n79834 , n79707 , n79821 );
and ( n79835 , n79834 , n79827 );
and ( n79836 , n79707 , n79821 );
or ( n79837 , n79835 , n79836 );
xor ( n79838 , n79713 , n79833 );
xor ( n79839 , n79838 , n79719 );
xor ( n79840 , n79713 , n79833 );
and ( n79841 , n79840 , n79719 );
and ( n79842 , n79713 , n79833 );
or ( n79843 , n79841 , n79842 );
not ( n79844 , n75025 );
not ( n79845 , n79782 );
or ( n79846 , n79844 , n79845 );
not ( n79847 , n65184 );
not ( n79848 , n77972 );
or ( n79849 , n79847 , n79848 );
nand ( n79850 , n79612 , n65183 );
nand ( n79851 , n79849 , n79850 );
nand ( n79852 , n79851 , n71466 );
nand ( n79853 , n79846 , n79852 );
and ( n79854 , n66581 , n39847 );
xor ( n79855 , n79853 , n79854 );
not ( n79856 , n79280 );
and ( n79857 , n75286 , n79067 );
not ( n79858 , n75286 );
and ( n79859 , n79858 , n39334 );
nor ( n79860 , n79857 , n79859 );
not ( n79861 , n79860 );
or ( n79862 , n79856 , n79861 );
not ( n79863 , n79768 );
nand ( n79864 , n79863 , n70500 );
nand ( n79865 , n79862 , n79864 );
xor ( n79866 , n79855 , n79865 );
xor ( n79867 , n79853 , n79854 );
and ( n79868 , n79867 , n79865 );
and ( n79869 , n79853 , n79854 );
or ( n79870 , n79868 , n79869 );
not ( n79871 , n72484 );
not ( n79872 , n79794 );
or ( n79873 , n79871 , n79872 );
not ( n79874 , n71309 );
not ( n79875 , n59891 );
or ( n79876 , n79874 , n79875 );
nand ( n79877 , n71547 , n77333 );
nand ( n79878 , n79876 , n79877 );
nand ( n79879 , n79878 , n61558 );
nand ( n79880 , n79873 , n79879 );
not ( n79881 , n72131 );
not ( n79882 , n79758 );
or ( n79883 , n79881 , n79882 );
not ( n79884 , n79107 );
not ( n79885 , n69961 );
or ( n79886 , n79884 , n79885 );
nand ( n79887 , n69962 , n70920 );
nand ( n79888 , n79886 , n79887 );
nand ( n79889 , n79888 , n75578 );
nand ( n79890 , n79883 , n79889 );
xor ( n79891 , n79880 , n79890 );
not ( n79892 , n75427 );
not ( n79893 , n72083 );
not ( n79894 , n39715 );
or ( n79895 , n79893 , n79894 );
nand ( n79896 , n39716 , n77344 );
nand ( n79897 , n79895 , n79896 );
not ( n79898 , n79897 );
or ( n79899 , n79892 , n79898 );
buf ( n79900 , n72495 );
or ( n79901 , n79804 , n79900 );
nand ( n79902 , n79899 , n79901 );
xor ( n79903 , n79891 , n79902 );
xor ( n79904 , n79880 , n79890 );
and ( n79905 , n79904 , n79902 );
and ( n79906 , n79880 , n79890 );
or ( n79907 , n79905 , n79906 );
not ( n79908 , n71960 );
not ( n79909 , n79748 );
or ( n79910 , n79908 , n79909 );
xor ( n79911 , n66581 , n76082 );
nand ( n79912 , n79911 , n70964 );
nand ( n79913 , n79910 , n79912 );
not ( n79914 , n69648 );
not ( n79915 , n70608 );
and ( n79916 , n79914 , n79915 );
and ( n79917 , n79735 , n72961 );
nor ( n79918 , n79916 , n79917 );
xor ( n79919 , n79913 , n79918 );
xor ( n79920 , n79919 , n79744 );
xor ( n79921 , n79913 , n79918 );
and ( n79922 , n79921 , n79744 );
and ( n79923 , n79913 , n79918 );
or ( n79924 , n79922 , n79923 );
xor ( n79925 , n79776 , n79812 );
xor ( n79926 , n79925 , n79903 );
xor ( n79927 , n79776 , n79812 );
and ( n79928 , n79927 , n79903 );
and ( n79929 , n79776 , n79812 );
or ( n79930 , n79928 , n79929 );
xor ( n79931 , n79866 , n79920 );
xor ( n79932 , n79931 , n79819 );
xor ( n79933 , n79866 , n79920 );
and ( n79934 , n79933 , n79819 );
and ( n79935 , n79866 , n79920 );
or ( n79936 , n79934 , n79935 );
xor ( n79937 , n79926 , n79825 );
xor ( n79938 , n79937 , n79932 );
xor ( n79939 , n79926 , n79825 );
and ( n79940 , n79939 , n79932 );
and ( n79941 , n79926 , n79825 );
or ( n79942 , n79940 , n79941 );
xor ( n79943 , n79831 , n79938 );
xor ( n79944 , n79943 , n79837 );
xor ( n79945 , n79831 , n79938 );
and ( n79946 , n79945 , n79837 );
and ( n79947 , n79831 , n79938 );
or ( n79948 , n79946 , n79947 );
not ( n79949 , n69648 );
not ( n79950 , n72962 );
or ( n79951 , n79949 , n79950 );
nand ( n79952 , n79951 , n67568 );
not ( n79953 , n71466 );
not ( n79954 , n79494 );
and ( n79955 , n65184 , n79954 );
not ( n79956 , n65184 );
and ( n79957 , n79956 , n42657 );
nor ( n79958 , n79955 , n79957 );
not ( n79959 , n79958 );
not ( n79960 , n79959 );
or ( n79961 , n79953 , n79960 );
nand ( n79962 , n79851 , n75025 );
nand ( n79963 , n79961 , n79962 );
xor ( n79964 , n79952 , n79963 );
not ( n79965 , n79280 );
not ( n79966 , n75286 );
not ( n79967 , n39254 );
or ( n79968 , n79966 , n79967 );
nand ( n79969 , n39255 , n72477 );
nand ( n79970 , n79968 , n79969 );
not ( n79971 , n79970 );
or ( n79972 , n79965 , n79971 );
nand ( n79973 , n79860 , n70500 );
nand ( n79974 , n79972 , n79973 );
xor ( n79975 , n79964 , n79974 );
xor ( n79976 , n79952 , n79963 );
and ( n79977 , n79976 , n79974 );
and ( n79978 , n79952 , n79963 );
or ( n79979 , n79977 , n79978 );
and ( n79980 , n66581 , n43609 );
not ( n79981 , n61558 );
and ( n79982 , n77333 , n79246 );
not ( n79983 , n77333 );
and ( n79984 , n79983 , n72622 );
nor ( n79985 , n79982 , n79984 );
not ( n79986 , n79985 );
or ( n79987 , n79981 , n79986 );
nand ( n79988 , n79878 , n72484 );
nand ( n79989 , n79987 , n79988 );
xor ( n79990 , n79980 , n79989 );
not ( n79991 , n75578 );
and ( n79992 , n79107 , n76454 );
not ( n79993 , n79107 );
and ( n79994 , n79993 , n76455 );
nor ( n79995 , n79992 , n79994 );
not ( n79996 , n79995 );
or ( n79997 , n79991 , n79996 );
not ( n79998 , n79888 );
not ( n79999 , n72131 );
or ( n80000 , n79998 , n79999 );
nand ( n80001 , n79997 , n80000 );
xor ( n80002 , n79990 , n80001 );
xor ( n80003 , n79980 , n79989 );
and ( n80004 , n80003 , n80001 );
and ( n80005 , n79980 , n79989 );
or ( n80006 , n80004 , n80005 );
not ( n80007 , n75427 );
buf ( n80008 , n72083 );
and ( n80009 , n80008 , n39575 );
not ( n80010 , n80008 );
and ( n80011 , n80010 , n79547 );
nor ( n80012 , n80009 , n80011 );
not ( n80013 , n80012 );
or ( n80014 , n80007 , n80013 );
nand ( n80015 , n79897 , n77077 );
nand ( n80016 , n80014 , n80015 );
not ( n80017 , n70964 );
xor ( n80018 , n66581 , n39681 );
not ( n80019 , n80018 );
or ( n80020 , n80017 , n80019 );
nand ( n80021 , n79911 , n71960 );
nand ( n80022 , n80020 , n80021 );
xor ( n80023 , n80016 , n80022 );
not ( n80024 , n79918 );
xor ( n80025 , n80023 , n80024 );
xor ( n80026 , n80016 , n80022 );
and ( n80027 , n80026 , n80024 );
and ( n80028 , n80016 , n80022 );
or ( n80029 , n80027 , n80028 );
xor ( n80030 , n79907 , n79870 );
xor ( n80031 , n80030 , n79975 );
xor ( n80032 , n79907 , n79870 );
and ( n80033 , n80032 , n79975 );
and ( n80034 , n79907 , n79870 );
or ( n80035 , n80033 , n80034 );
xor ( n80036 , n80002 , n80025 );
xor ( n80037 , n80036 , n79924 );
xor ( n80038 , n80002 , n80025 );
and ( n80039 , n80038 , n79924 );
and ( n80040 , n80002 , n80025 );
or ( n80041 , n80039 , n80040 );
xor ( n80042 , n80031 , n79930 );
xor ( n80043 , n80042 , n79936 );
xor ( n80044 , n80031 , n79930 );
and ( n80045 , n80044 , n79936 );
and ( n80046 , n80031 , n79930 );
or ( n80047 , n80045 , n80046 );
xor ( n80048 , n80037 , n80043 );
xor ( n80049 , n80048 , n79942 );
xor ( n80050 , n80037 , n80043 );
and ( n80051 , n80050 , n79942 );
and ( n80052 , n80037 , n80043 );
or ( n80053 , n80051 , n80052 );
not ( n80054 , n72131 );
not ( n80055 , n79995 );
or ( n80056 , n80054 , n80055 );
and ( n80057 , n70920 , n79612 );
not ( n80058 , n70920 );
and ( n80059 , n80058 , n77972 );
nor ( n80060 , n80057 , n80059 );
not ( n80061 , n80060 );
nand ( n80062 , n80061 , n75578 );
nand ( n80063 , n80056 , n80062 );
not ( n80064 , n61558 );
and ( n80065 , n71309 , n79067 );
not ( n80066 , n71309 );
and ( n80067 , n80066 , n39334 );
nor ( n80068 , n80065 , n80067 );
not ( n80069 , n80068 );
or ( n80070 , n80064 , n80069 );
nand ( n80071 , n79985 , n72484 );
nand ( n80072 , n80070 , n80071 );
xor ( n80073 , n80063 , n80072 );
not ( n80074 , n80012 );
or ( n80075 , n80074 , n79900 );
and ( n80076 , n77344 , n71547 );
not ( n80077 , n77344 );
and ( n80078 , n80077 , n59891 );
nor ( n80079 , n80076 , n80078 );
or ( n80080 , n80079 , n69703 );
nand ( n80081 , n80075 , n80080 );
xor ( n80082 , n80073 , n80081 );
xor ( n80083 , n80063 , n80072 );
and ( n80084 , n80083 , n80081 );
and ( n80085 , n80063 , n80072 );
or ( n80086 , n80084 , n80085 );
not ( n80087 , n70500 );
not ( n80088 , n79970 );
or ( n80089 , n80087 , n80088 );
not ( n80090 , n75286 );
not ( n80091 , n69961 );
or ( n80092 , n80090 , n80091 );
nand ( n80093 , n69962 , n78148 );
nand ( n80094 , n80092 , n80093 );
nand ( n80095 , n80094 , n79280 );
nand ( n80096 , n80089 , n80095 );
not ( n80097 , n71960 );
not ( n80098 , n80018 );
or ( n80099 , n80097 , n80098 );
xor ( n80100 , n67072 , n79406 );
nand ( n80101 , n80100 , n70964 );
nand ( n80102 , n80099 , n80101 );
xor ( n80103 , n80096 , n80102 );
and ( n80104 , n66581 , n76082 );
xor ( n80105 , n80103 , n80104 );
xor ( n80106 , n80096 , n80102 );
and ( n80107 , n80106 , n80104 );
and ( n80108 , n80096 , n80102 );
or ( n80109 , n80107 , n80108 );
not ( n80110 , n79958 );
not ( n80111 , n75025 );
not ( n80112 , n80111 );
and ( n80113 , n80110 , n80112 );
and ( n80114 , n71466 , n65184 );
nor ( n80115 , n80113 , n80114 );
xor ( n80116 , n80115 , n79979 );
xor ( n80117 , n80116 , n80006 );
xor ( n80118 , n80115 , n79979 );
and ( n80119 , n80118 , n80006 );
and ( n80120 , n80115 , n79979 );
or ( n80121 , n80119 , n80120 );
xor ( n80122 , n80105 , n80082 );
xor ( n80123 , n80122 , n80029 );
xor ( n80124 , n80105 , n80082 );
and ( n80125 , n80124 , n80029 );
and ( n80126 , n80105 , n80082 );
or ( n80127 , n80125 , n80126 );
xor ( n80128 , n80117 , n80035 );
xor ( n80129 , n80128 , n80123 );
xor ( n80130 , n80117 , n80035 );
and ( n80131 , n80130 , n80123 );
and ( n80132 , n80117 , n80035 );
or ( n80133 , n80131 , n80132 );
xor ( n80134 , n80041 , n80129 );
xor ( n80135 , n80134 , n80047 );
xor ( n80136 , n80041 , n80129 );
and ( n80137 , n80136 , n80047 );
and ( n80138 , n80041 , n80129 );
or ( n80139 , n80137 , n80138 );
or ( n80140 , n75025 , n71466 );
nand ( n80141 , n80140 , n65184 );
or ( n80142 , n80060 , n79999 );
and ( n80143 , n79107 , n79954 );
not ( n80144 , n79107 );
not ( n80145 , n79954 );
and ( n80146 , n80144 , n80145 );
nor ( n80147 , n80143 , n80146 );
not ( n80148 , n75578 );
or ( n80149 , n80147 , n80148 );
nand ( n80150 , n80142 , n80149 );
xor ( n80151 , n80141 , n80150 );
not ( n80152 , n72484 );
not ( n80153 , n80068 );
or ( n80154 , n80152 , n80153 );
and ( n80155 , n77333 , n39255 );
and ( n80156 , n39254 , n71309 );
nor ( n80157 , n80155 , n80156 );
or ( n80158 , n80157 , n69731 );
nand ( n80159 , n80154 , n80158 );
xor ( n80160 , n80151 , n80159 );
xor ( n80161 , n80141 , n80150 );
and ( n80162 , n80161 , n80159 );
and ( n80163 , n80141 , n80150 );
or ( n80164 , n80162 , n80163 );
not ( n80165 , n77077 );
not ( n80166 , n80079 );
not ( n80167 , n80166 );
or ( n80168 , n80165 , n80167 );
and ( n80169 , n72622 , n77344 );
and ( n80170 , n79246 , n80008 );
nor ( n80171 , n80169 , n80170 );
or ( n80172 , n80171 , n69703 );
nand ( n80173 , n80168 , n80172 );
not ( n80174 , n79280 );
and ( n80175 , n78148 , n76454 );
not ( n80176 , n78148 );
and ( n80177 , n80176 , n76455 );
nor ( n80178 , n80175 , n80177 );
not ( n80179 , n80178 );
not ( n80180 , n80179 );
or ( n80181 , n80174 , n80180 );
not ( n80182 , n80094 );
or ( n80183 , n80182 , n72474 );
nand ( n80184 , n80181 , n80183 );
xor ( n80185 , n80173 , n80184 );
not ( n80186 , n80100 );
not ( n80187 , n71960 );
or ( n80188 , n80186 , n80187 );
and ( n80189 , n39575 , n75987 );
and ( n80190 , n79547 , n67072 );
nor ( n80191 , n80189 , n80190 );
or ( n80192 , n80191 , n72838 );
nand ( n80193 , n80188 , n80192 );
xor ( n80194 , n80185 , n80193 );
xor ( n80195 , n80173 , n80184 );
and ( n80196 , n80195 , n80193 );
and ( n80197 , n80173 , n80184 );
or ( n80198 , n80196 , n80197 );
and ( n80199 , n66581 , n39681 );
not ( n80200 , n80115 );
xor ( n80201 , n80199 , n80200 );
xor ( n80202 , n80201 , n80086 );
xor ( n80203 , n80199 , n80200 );
and ( n80204 , n80203 , n80086 );
and ( n80205 , n80199 , n80200 );
or ( n80206 , n80204 , n80205 );
xor ( n80207 , n80109 , n80194 );
xor ( n80208 , n80207 , n80160 );
xor ( n80209 , n80109 , n80194 );
and ( n80210 , n80209 , n80160 );
and ( n80211 , n80109 , n80194 );
or ( n80212 , n80210 , n80211 );
xor ( n80213 , n80202 , n80121 );
xor ( n80214 , n80213 , n80127 );
xor ( n80215 , n80202 , n80121 );
and ( n80216 , n80215 , n80127 );
and ( n80217 , n80202 , n80121 );
or ( n80218 , n80216 , n80217 );
xor ( n80219 , n80208 , n80214 );
xor ( n80220 , n80219 , n80133 );
xor ( n80221 , n80208 , n80214 );
and ( n80222 , n80221 , n80133 );
and ( n80223 , n80208 , n80214 );
or ( n80224 , n80222 , n80223 );
or ( n80225 , n80171 , n79900 );
and ( n80226 , n79067 , n77344 );
not ( n80227 , n79067 );
and ( n80228 , n80227 , n72083 );
nor ( n80229 , n80226 , n80228 );
or ( n80230 , n80229 , n69703 );
nand ( n80231 , n80225 , n80230 );
or ( n80232 , n80191 , n80187 );
and ( n80233 , n67072 , n59891 );
not ( n80234 , n67072 );
and ( n80235 , n80234 , n71547 );
nor ( n80236 , n80233 , n80235 );
or ( n80237 , n80236 , n72838 );
nand ( n80238 , n80232 , n80237 );
xor ( n80239 , n80231 , n80238 );
or ( n80240 , n80147 , n79999 );
or ( n80241 , n80148 , n70920 );
nand ( n80242 , n80240 , n80241 );
xor ( n80243 , n80239 , n80242 );
xor ( n80244 , n80231 , n80238 );
and ( n80245 , n80244 , n80242 );
and ( n80246 , n80231 , n80238 );
or ( n80247 , n80245 , n80246 );
and ( n80248 , n67072 , n79406 );
not ( n80249 , n72484 );
or ( n80250 , n80157 , n80249 );
and ( n80251 , n69961 , n71309 );
not ( n80252 , n69961 );
and ( n80253 , n80252 , n77333 );
nor ( n80254 , n80251 , n80253 );
or ( n80255 , n80254 , n69731 );
nand ( n80256 , n80250 , n80255 );
xor ( n80257 , n80248 , n80256 );
or ( n80258 , n80178 , n72474 );
and ( n80259 , n42556 , n72477 );
and ( n80260 , n77972 , n75286 );
nor ( n80261 , n80259 , n80260 );
or ( n80262 , n80261 , n79769 );
nand ( n80263 , n80258 , n80262 );
not ( n80264 , n80263 );
xor ( n80265 , n80257 , n80264 );
xor ( n80266 , n80248 , n80256 );
and ( n80267 , n80266 , n80264 );
and ( n80268 , n80248 , n80256 );
or ( n80269 , n80267 , n80268 );
xor ( n80270 , n80198 , n80164 );
xor ( n80271 , n80270 , n80243 );
xor ( n80272 , n80198 , n80164 );
and ( n80273 , n80272 , n80243 );
and ( n80274 , n80198 , n80164 );
or ( n80275 , n80273 , n80274 );
xor ( n80276 , n80265 , n80206 );
xor ( n80277 , n80276 , n80212 );
xor ( n80278 , n80265 , n80206 );
and ( n80279 , n80278 , n80212 );
and ( n80280 , n80265 , n80206 );
or ( n80281 , n80279 , n80280 );
xor ( n80282 , n80271 , n80277 );
xor ( n80283 , n80282 , n80218 );
xor ( n80284 , n80271 , n80277 );
and ( n80285 , n80284 , n80218 );
and ( n80286 , n80271 , n80277 );
or ( n80287 , n80285 , n80286 );
or ( n80288 , n72131 , n75578 );
nand ( n80289 , n80288 , n79107 );
or ( n80290 , n80261 , n72474 );
and ( n80291 , n75286 , n42658 );
not ( n80292 , n75286 );
and ( n80293 , n80292 , n80145 );
nor ( n80294 , n80291 , n80293 );
or ( n80295 , n80294 , n79769 );
nand ( n80296 , n80290 , n80295 );
xor ( n80297 , n80289 , n80296 );
or ( n80298 , n80229 , n79900 );
and ( n80299 , n39255 , n77344 );
and ( n80300 , n39254 , n80008 );
nor ( n80301 , n80299 , n80300 );
or ( n80302 , n80301 , n69703 );
nand ( n80303 , n80298 , n80302 );
xor ( n80304 , n80297 , n80303 );
xor ( n80305 , n80289 , n80296 );
and ( n80306 , n80305 , n80303 );
and ( n80307 , n80289 , n80296 );
or ( n80308 , n80306 , n80307 );
and ( n80309 , n67072 , n79246 );
not ( n80310 , n67072 );
and ( n80311 , n80310 , n72622 );
nor ( n80312 , n80309 , n80311 );
not ( n80313 , n80312 );
not ( n80314 , n80313 );
not ( n80315 , n70964 );
or ( n80316 , n80314 , n80315 );
or ( n80317 , n80236 , n80187 );
nand ( n80318 , n80316 , n80317 );
or ( n80319 , n80254 , n80249 );
and ( n80320 , n76454 , n77333 );
and ( n80321 , n76455 , n71309 );
nor ( n80322 , n80320 , n80321 );
or ( n80323 , n80322 , n69731 );
nand ( n80324 , n80319 , n80323 );
xor ( n80325 , n80318 , n80324 );
nor ( n80326 , n76444 , n75987 );
xor ( n80327 , n80325 , n80326 );
xor ( n80328 , n80318 , n80324 );
and ( n80329 , n80328 , n80326 );
and ( n80330 , n80318 , n80324 );
or ( n80331 , n80329 , n80330 );
xor ( n80332 , n80263 , n80247 );
xor ( n80333 , n80332 , n80327 );
xor ( n80334 , n80263 , n80247 );
and ( n80335 , n80334 , n80327 );
and ( n80336 , n80263 , n80247 );
or ( n80337 , n80335 , n80336 );
xor ( n80338 , n80304 , n80269 );
xor ( n80339 , n80338 , n80333 );
xor ( n80340 , n80304 , n80269 );
and ( n80341 , n80340 , n80333 );
and ( n80342 , n80304 , n80269 );
or ( n80343 , n80341 , n80342 );
xor ( n80344 , n80275 , n80339 );
xor ( n80345 , n80344 , n80281 );
xor ( n80346 , n80275 , n80339 );
and ( n80347 , n80346 , n80281 );
and ( n80348 , n80275 , n80339 );
or ( n80349 , n80347 , n80348 );
or ( n80350 , n80312 , n71959 );
and ( n80351 , n39335 , n75987 );
and ( n80352 , n39334 , n67072 );
nor ( n80353 , n80351 , n80352 );
or ( n80354 , n80353 , n72838 );
nand ( n80355 , n80350 , n80354 );
not ( n80356 , n75987 );
and ( n80357 , n71547 , n80356 );
xor ( n80358 , n80355 , n80357 );
not ( n80359 , n75286 );
not ( n80360 , n79280 );
or ( n80361 , n80359 , n80360 );
or ( n80362 , n80294 , n72474 );
nand ( n80363 , n80361 , n80362 );
xor ( n80364 , n80358 , n80363 );
xor ( n80365 , n80355 , n80357 );
and ( n80366 , n80365 , n80363 );
and ( n80367 , n80355 , n80357 );
or ( n80368 , n80366 , n80367 );
or ( n80369 , n80301 , n79900 );
not ( n80370 , n69961 );
and ( n80371 , n80370 , n77344 );
and ( n80372 , n69961 , n80008 );
nor ( n80373 , n80371 , n80372 );
or ( n80374 , n80373 , n69703 );
nand ( n80375 , n80369 , n80374 );
or ( n80376 , n80322 , n80249 );
and ( n80377 , n71309 , n77972 );
not ( n80378 , n71309 );
and ( n80379 , n80378 , n79612 );
nor ( n80380 , n80377 , n80379 );
or ( n80381 , n80380 , n69731 );
nand ( n80382 , n80376 , n80381 );
not ( n80383 , n80382 );
xor ( n80384 , n80375 , n80383 );
xor ( n80385 , n80384 , n80331 );
xor ( n80386 , n80375 , n80383 );
and ( n80387 , n80386 , n80331 );
and ( n80388 , n80375 , n80383 );
or ( n80389 , n80387 , n80388 );
xor ( n80390 , n80308 , n80364 );
xor ( n80391 , n80390 , n80385 );
xor ( n80392 , n80308 , n80364 );
and ( n80393 , n80392 , n80385 );
and ( n80394 , n80308 , n80364 );
or ( n80395 , n80393 , n80394 );
xor ( n80396 , n80337 , n80391 );
xor ( n80397 , n80396 , n80343 );
xor ( n80398 , n80337 , n80391 );
and ( n80399 , n80398 , n80343 );
and ( n80400 , n80337 , n80391 );
or ( n80401 , n80399 , n80400 );
or ( n80402 , n70500 , n79280 );
nand ( n80403 , n80402 , n75286 );
not ( n80404 , n72484 );
not ( n80405 , n80380 );
not ( n80406 , n80405 );
or ( n80407 , n80404 , n80406 );
not ( n80408 , n42659 );
and ( n80409 , n80408 , n77333 );
and ( n80410 , n42659 , n71309 );
nor ( n80411 , n80409 , n80410 );
or ( n80412 , n80411 , n69731 );
nand ( n80413 , n80407 , n80412 );
xor ( n80414 , n80403 , n80413 );
or ( n80415 , n80353 , n71959 );
and ( n80416 , n39255 , n75987 );
and ( n80417 , n39254 , n67072 );
nor ( n80418 , n80416 , n80417 );
or ( n80419 , n80418 , n72838 );
nand ( n80420 , n80415 , n80419 );
xor ( n80421 , n80414 , n80420 );
xor ( n80422 , n80403 , n80413 );
and ( n80423 , n80422 , n80420 );
and ( n80424 , n80403 , n80413 );
or ( n80425 , n80423 , n80424 );
not ( n80426 , n72622 );
nor ( n80427 , n80426 , n75987 );
or ( n80428 , n80373 , n79900 );
and ( n80429 , n80008 , n76455 );
not ( n80430 , n80008 );
and ( n80431 , n80430 , n76454 );
nor ( n80432 , n80429 , n80431 );
or ( n80433 , n80432 , n69703 );
nand ( n80434 , n80428 , n80433 );
xor ( n80435 , n80427 , n80434 );
xor ( n80436 , n80435 , n80382 );
xor ( n80437 , n80427 , n80434 );
and ( n80438 , n80437 , n80382 );
and ( n80439 , n80427 , n80434 );
or ( n80440 , n80438 , n80439 );
xor ( n80441 , n80368 , n80421 );
xor ( n80442 , n80441 , n80436 );
xor ( n80443 , n80368 , n80421 );
and ( n80444 , n80443 , n80436 );
and ( n80445 , n80368 , n80421 );
or ( n80446 , n80444 , n80445 );
xor ( n80447 , n80389 , n80442 );
xor ( n80448 , n80447 , n80395 );
xor ( n80449 , n80389 , n80442 );
and ( n80450 , n80449 , n80395 );
and ( n80451 , n80389 , n80442 );
or ( n80452 , n80450 , n80451 );
nor ( n80453 , n39334 , n75987 );
or ( n80454 , n80432 , n79900 );
and ( n80455 , n42556 , n77344 );
and ( n80456 , n77972 , n80008 );
nor ( n80457 , n80455 , n80456 );
or ( n80458 , n80457 , n69703 );
nand ( n80459 , n80454 , n80458 );
xor ( n80460 , n80453 , n80459 );
or ( n80461 , n80418 , n80187 );
and ( n80462 , n80370 , n75987 );
and ( n80463 , n69961 , n80356 );
nor ( n80464 , n80462 , n80463 );
or ( n80465 , n80464 , n72838 );
nand ( n80466 , n80461 , n80465 );
xor ( n80467 , n80460 , n80466 );
xor ( n80468 , n80453 , n80459 );
and ( n80469 , n80468 , n80466 );
and ( n80470 , n80453 , n80459 );
or ( n80471 , n80469 , n80470 );
or ( n80472 , n80411 , n80249 );
or ( n80473 , n69731 , n77333 );
nand ( n80474 , n80472 , n80473 );
not ( n80475 , n80474 );
xor ( n80476 , n80475 , n80425 );
xor ( n80477 , n80476 , n80467 );
xor ( n80478 , n80475 , n80425 );
and ( n80479 , n80478 , n80467 );
and ( n80480 , n80475 , n80425 );
or ( n80481 , n80479 , n80480 );
xor ( n80482 , n80440 , n80477 );
xor ( n80483 , n80482 , n80446 );
xor ( n80484 , n80440 , n80477 );
and ( n80485 , n80484 , n80446 );
and ( n80486 , n80440 , n80477 );
or ( n80487 , n80485 , n80486 );
or ( n80488 , n72484 , n61558 );
nand ( n80489 , n80488 , n71309 );
not ( n80490 , n75427 );
or ( n80491 , n42660 , n72083 );
not ( n80492 , n42660 );
or ( n80493 , n80492 , n77344 );
nand ( n80494 , n80491 , n80493 );
not ( n80495 , n80494 );
or ( n80496 , n80490 , n80495 );
or ( n80497 , n80457 , n79900 );
nand ( n80498 , n80496 , n80497 );
xor ( n80499 , n80489 , n80498 );
nor ( n80500 , n39254 , n75987 );
xor ( n80501 , n80499 , n80500 );
xor ( n80502 , n80489 , n80498 );
and ( n80503 , n80502 , n80500 );
and ( n80504 , n80489 , n80498 );
or ( n80505 , n80503 , n80504 );
or ( n80506 , n80464 , n80187 );
and ( n80507 , n76454 , n75987 );
and ( n80508 , n76455 , n67072 );
nor ( n80509 , n80507 , n80508 );
or ( n80510 , n80509 , n72838 );
nand ( n80511 , n80506 , n80510 );
xor ( n80512 , n80511 , n80474 );
xor ( n80513 , n80512 , n80471 );
xor ( n80514 , n80511 , n80474 );
and ( n80515 , n80514 , n80471 );
and ( n80516 , n80511 , n80474 );
or ( n80517 , n80515 , n80516 );
xor ( n80518 , n80501 , n80513 );
xor ( n80519 , n80518 , n80481 );
xor ( n80520 , n80501 , n80513 );
and ( n80521 , n80520 , n80481 );
and ( n80522 , n80501 , n80513 );
or ( n80523 , n80521 , n80522 );
or ( n80524 , n80509 , n80187 );
and ( n80525 , n42557 , n75987 );
not ( n80526 , n42557 );
and ( n80527 , n80526 , n80356 );
nor ( n80528 , n80525 , n80527 );
or ( n80529 , n80528 , n72838 );
nand ( n80530 , n80524 , n80529 );
not ( n80531 , n80370 );
nor ( n80532 , n80531 , n75987 );
xor ( n80533 , n80530 , n80532 );
and ( n80534 , n80494 , n77077 );
and ( n80535 , n75427 , n72083 );
nor ( n80536 , n80534 , n80535 );
xor ( n80537 , n80533 , n80536 );
xor ( n80538 , n80530 , n80532 );
and ( n80539 , n80538 , n80536 );
and ( n80540 , n80530 , n80532 );
or ( n80541 , n80539 , n80540 );
xor ( n80542 , n80505 , n80537 );
xor ( n80543 , n80542 , n80517 );
xor ( n80544 , n80505 , n80537 );
and ( n80545 , n80544 , n80517 );
and ( n80546 , n80505 , n80537 );
or ( n80547 , n80545 , n80546 );
or ( n80548 , n77077 , n75427 );
nand ( n80549 , n80548 , n72083 );
or ( n80550 , n80528 , n80187 );
xnor ( n80551 , n42661 , n75987 );
or ( n80552 , n80551 , n72838 );
nand ( n80553 , n80550 , n80552 );
xor ( n80554 , n80549 , n80553 );
nor ( n80555 , n76455 , n75987 );
xor ( n80556 , n80554 , n80555 );
xor ( n80557 , n80549 , n80553 );
and ( n80558 , n80557 , n80555 );
and ( n80559 , n80549 , n80553 );
or ( n80560 , n80558 , n80559 );
not ( n80561 , n80536 );
xor ( n80562 , n80561 , n80556 );
xor ( n80563 , n80562 , n80541 );
xor ( n80564 , n80561 , n80556 );
and ( n80565 , n80564 , n80541 );
and ( n80566 , n80561 , n80556 );
or ( n80567 , n80565 , n80566 );
or ( n80568 , n80551 , n80187 );
nand ( n80569 , n70964 , n80356 );
nand ( n80570 , n80568 , n80569 );
nand ( n80571 , n42557 , n80356 );
xor ( n80572 , n80570 , n80571 );
xor ( n80573 , n80572 , n80560 );
xor ( n80574 , n80570 , n80571 );
and ( n80575 , n80574 , n80560 );
and ( n80576 , n80570 , n80571 );
or ( n80577 , n80575 , n80576 );
or ( n80578 , n80452 , n80483 );
not ( n80579 , n80578 );
nor ( n80580 , n77887 , n77675 );
nor ( n80581 , n78092 , n77891 );
nor ( n80582 , n80580 , n80581 );
not ( n80583 , n78293 );
not ( n80584 , n78096 );
nand ( n80585 , n80583 , n80584 );
buf ( n80586 , n80585 );
or ( n80587 , n78297 , n78475 );
and ( n80588 , n80582 , n80586 , n80587 );
not ( n80589 , n80588 );
nor ( n80590 , n78659 , n78825 );
not ( n80591 , n80590 );
or ( n80592 , n78829 , n78991 );
nand ( n80593 , n80591 , n80592 );
nor ( n80594 , n78479 , n78655 );
nor ( n80595 , n80593 , n80594 );
buf ( n80596 , n80595 );
nor ( n80597 , n79176 , n78995 );
nor ( n80598 , n79180 , n79328 );
nor ( n80599 , n80597 , n80598 );
or ( n80600 , n79332 , n79468 );
not ( n80601 , n80600 );
nor ( n80602 , n79472 , n79601 );
nor ( n80603 , n80601 , n80602 );
nand ( n80604 , n80599 , n80603 );
not ( n80605 , n79725 );
not ( n80606 , n79839 );
and ( n80607 , n80605 , n80606 );
nor ( n80608 , n79721 , n79605 );
nor ( n80609 , n80607 , n80608 );
or ( n80610 , n80053 , n80135 );
not ( n80611 , n80610 );
nor ( n80612 , n80049 , n79948 );
nor ( n80613 , n79843 , n79944 );
nor ( n80614 , n80611 , n80612 , n80613 );
nand ( n80615 , n80609 , n80614 );
nor ( n80616 , n80604 , n80615 );
nand ( n80617 , n80596 , n80616 );
nor ( n80618 , n80589 , n80617 );
or ( n80619 , n80220 , n80139 );
nor ( n80620 , n80283 , n80224 );
not ( n80621 , n80620 );
nand ( n80622 , n80619 , n80621 );
or ( n80623 , n80349 , n80397 );
or ( n80624 , n80287 , n80345 );
or ( n80625 , n80401 , n80448 );
nand ( n80626 , n80623 , n80624 , n80625 );
nor ( n80627 , n80622 , n80626 );
and ( n80628 , n80618 , n80627 );
not ( n80629 , n80628 );
or ( n80630 , n71253 , n70850 );
buf ( n80631 , n71257 );
buf ( n80632 , n71645 );
nor ( n80633 , n80631 , n80632 );
not ( n80634 , n80633 );
not ( n80635 , n72033 );
not ( n80636 , n72412 );
nand ( n80637 , n80635 , n80636 );
not ( n80638 , n71649 );
not ( n80639 , n72029 );
nand ( n80640 , n80638 , n80639 );
buf ( n80641 , n80640 );
nand ( n80642 , n80630 , n80634 , n80637 , n80641 );
nor ( n80643 , n73490 , n73821 );
nor ( n80644 , n74155 , n73825 );
nor ( n80645 , n80643 , n80644 );
nor ( n80646 , n74466 , n74159 );
nor ( n80647 , n74470 , n74781 );
nor ( n80648 , n80646 , n80647 );
and ( n80649 , n80645 , n80648 );
not ( n80650 , n73486 );
not ( n80651 , n73143 );
nand ( n80652 , n80650 , n80651 );
not ( n80653 , n72776 );
not ( n80654 , n72416 );
nand ( n80655 , n80653 , n80654 );
not ( n80656 , n72780 );
not ( n80657 , n73139 );
nand ( n80658 , n80656 , n80657 );
and ( n80659 , n80652 , n80655 , n80658 );
nand ( n80660 , n80649 , n80659 );
nor ( n80661 , n80642 , n80660 );
buf ( n80662 , n75381 );
buf ( n80663 , n75083 );
nor ( n80664 , n80662 , n80663 );
not ( n80665 , n80664 );
not ( n80666 , n75385 );
not ( n80667 , n75669 );
nand ( n80668 , n80666 , n80667 );
buf ( n80669 , n80668 );
or ( n80670 , n75079 , n74785 );
not ( n80671 , n75949 );
not ( n80672 , n75673 );
nand ( n80673 , n80671 , n80672 );
and ( n80674 , n80665 , n80669 , n80670 , n80673 );
nor ( n80675 , n76992 , n76745 );
nor ( n80676 , n77226 , n76996 );
nor ( n80677 , n80675 , n80676 );
nor ( n80678 , n77456 , n77230 );
nor ( n80679 , n77460 , n77671 );
nor ( n80680 , n80678 , n80679 );
nand ( n80681 , n80677 , n80680 );
not ( n80682 , n76493 );
not ( n80683 , n76226 );
nand ( n80684 , n80682 , n80683 );
not ( n80685 , n75953 );
not ( n80686 , n76222 );
nand ( n80687 , n80685 , n80686 );
not ( n80688 , n76741 );
not ( n80689 , n76497 );
nand ( n80690 , n80688 , n80689 );
nand ( n80691 , n80684 , n80687 , n80690 );
nor ( n80692 , n80681 , n80691 );
nand ( n80693 , n80674 , n80692 );
not ( n80694 , n80693 );
and ( n80695 , n80661 , n80694 );
not ( n80696 , n80695 );
not ( n80697 , n70029 );
not ( n80698 , n69618 );
nand ( n80699 , n80697 , n80698 );
not ( n80700 , n70033 );
not ( n80701 , n70446 );
nand ( n80702 , n80700 , n80701 );
not ( n80703 , n69189 );
not ( n80704 , n69614 );
nand ( n80705 , n80703 , n80704 );
and ( n80706 , n80699 , n80702 , n80705 );
buf ( n80707 , n66889 );
buf ( n80708 , n66403 );
nor ( n80709 , n80707 , n80708 );
nor ( n80710 , n66399 , n65920 );
nor ( n80711 , n80709 , n80710 );
not ( n80712 , n67829 );
not ( n80713 , n67370 );
and ( n80714 , n80712 , n80713 );
not ( n80715 , n67366 );
not ( n80716 , n66893 );
nand ( n80717 , n80715 , n80716 );
not ( n80718 , n80717 );
nor ( n80719 , n80714 , n80718 );
nand ( n80720 , n80711 , n80719 );
not ( n80721 , n80720 );
nor ( n80722 , n68738 , n68283 );
nor ( n80723 , n68742 , n69185 );
nor ( n80724 , n68279 , n67833 );
nor ( n80725 , n80722 , n80723 , n80724 );
or ( n80726 , n70846 , n70450 );
and ( n80727 , n80706 , n80721 , n80725 , n80726 );
not ( n80728 , n80727 );
nor ( n80729 , n62794 , n63326 );
nor ( n80730 , n63888 , n63330 );
nor ( n80731 , n80729 , n80730 );
buf ( n80732 , n64404 );
not ( n80733 , n80732 );
not ( n80734 , n63892 );
nand ( n80735 , n80733 , n80734 );
or ( n80736 , n64910 , n64408 );
nand ( n80737 , n80731 , n80735 , n80736 );
or ( n80738 , n65417 , n64914 );
or ( n80739 , n65916 , n65421 );
nand ( n80740 , n80738 , n80739 );
nor ( n80741 , n80737 , n80740 );
not ( n80742 , n80741 );
or ( n80743 , n61753 , n62246 );
not ( n80744 , n80743 );
nor ( n80745 , n61749 , n61243 );
not ( n80746 , n80745 );
not ( n80747 , n80746 );
not ( n80748 , n61239 );
not ( n80749 , n60745 );
nand ( n80750 , n80748 , n80749 );
not ( n80751 , n80750 );
nor ( n80752 , n60741 , n60241 );
nand ( n80753 , n60237 , n59780 );
or ( n80754 , n80752 , n80753 );
nand ( n80755 , n60741 , n60241 );
nand ( n80756 , n80754 , n80755 );
not ( n80757 , n80756 );
or ( n80758 , n80751 , n80757 );
nand ( n80759 , n61239 , n60745 );
nand ( n80760 , n80758 , n80759 );
not ( n80761 , n80760 );
or ( n80762 , n80747 , n80761 );
nand ( n80763 , n61749 , n61243 );
nand ( n80764 , n80762 , n80763 );
not ( n80765 , n80764 );
or ( n80766 , n80744 , n80765 );
nand ( n80767 , n61753 , n62246 );
nand ( n80768 , n80766 , n80767 );
nor ( n80769 , n62790 , n62250 );
not ( n80770 , n80769 );
nand ( n80771 , n80768 , n80770 );
nor ( n80772 , n57934 , n57468 );
not ( n80773 , n80772 );
or ( n80774 , n57938 , n58362 );
or ( n80775 , n58820 , n58366 );
nand ( n80776 , n80773 , n80774 , n80775 );
or ( n80777 , n59776 , n59274 );
or ( n80778 , n59270 , n58824 );
nand ( n80779 , n80777 , n80778 );
nor ( n80780 , n80776 , n80779 );
not ( n80781 , n80780 );
nor ( n80782 , n56157 , n56574 );
nor ( n80783 , n56153 , n55730 );
nor ( n80784 , n80782 , n80783 );
not ( n80785 , n57464 );
not ( n80786 , n57034 );
nand ( n80787 , n80785 , n80786 );
or ( n80788 , n57030 , n56578 );
and ( n80789 , n80784 , n80787 , n80788 );
not ( n80790 , n80789 );
nor ( n80791 , n55338 , n54919 );
nor ( n80792 , n55342 , n55726 );
nor ( n80793 , n54915 , n54524 );
nor ( n80794 , n80791 , n80792 , n80793 );
not ( n80795 , n80794 );
nor ( n80796 , n54520 , n54127 );
nor ( n80797 , n53775 , n54123 );
nor ( n80798 , n53771 , n53383 );
nor ( n80799 , n80796 , n80797 , n80798 );
not ( n80800 , n80799 );
not ( n80801 , n53379 );
not ( n80802 , n53026 );
and ( n80803 , n80801 , n80802 );
not ( n80804 , n53022 );
not ( n80805 , n52654 );
and ( n80806 , n80804 , n80805 );
nor ( n80807 , n80803 , n80806 );
not ( n80808 , n80807 );
nor ( n80809 , n51630 , n51303 );
nor ( n80810 , n51299 , n51010 );
nor ( n80811 , n51006 , n50704 );
nor ( n80812 , n80809 , n80810 , n80811 );
not ( n80813 , n80812 );
nor ( n80814 , n50700 , n50425 );
nor ( n80815 , n50421 , n50117 );
nor ( n80816 , n80814 , n80815 );
not ( n80817 , n80816 );
nor ( n80818 , n50113 , n49859 );
nor ( n80819 , n49855 , n49567 );
nor ( n80820 , n80818 , n80819 );
not ( n80821 , n80820 );
nor ( n80822 , n49563 , n49332 );
nor ( n80823 , n49328 , n49047 );
nor ( n80824 , n80822 , n80823 );
not ( n80825 , n80824 );
not ( n80826 , n48369 );
not ( n80827 , n48156 );
and ( n80828 , n80826 , n80827 );
nor ( n80829 , n48152 , n47954 );
nor ( n80830 , n80828 , n80829 );
not ( n80831 , n80830 );
nor ( n80832 , n47950 , n47738 );
nor ( n80833 , n47734 , n47556 );
nor ( n80834 , n80832 , n80833 );
not ( n80835 , n80834 );
or ( n80836 , n47552 , n47361 );
not ( n80837 , n80836 );
nor ( n80838 , n47357 , n47204 );
not ( n80839 , n80838 );
not ( n80840 , n80839 );
nor ( n80841 , n47200 , n47033 );
not ( n80842 , n80841 );
not ( n80843 , n80842 );
nor ( n80844 , n47029 , n46906 );
nor ( n80845 , n46902 , n46743 );
nor ( n80846 , n80844 , n80845 );
not ( n80847 , n80846 );
or ( n80848 , n46739 , n46626 );
not ( n80849 , n80848 );
or ( n80850 , n46622 , n46487 );
not ( n80851 , n80850 );
or ( n80852 , n46483 , n46372 );
not ( n80853 , n80852 );
or ( n80854 , n46368 , n46259 );
not ( n80855 , n80854 );
nor ( n80856 , n46173 , n46088 );
or ( n80857 , n46084 , n46024 );
xor ( n80858 , n45870 , n45929 );
xor ( n80859 , n45780 , n45787 );
not ( n80860 , n44004 );
and ( n80861 , n45777 , n45834 );
not ( n80862 , n45777 );
and ( n80863 , n80862 , n46111 );
or ( n80864 , n80861 , n80863 );
not ( n80865 , n80864 );
or ( n80866 , n80860 , n80865 );
and ( n80867 , n45777 , n30633 );
not ( n80868 , n45777 );
and ( n80869 , n80868 , n45752 );
or ( n80870 , n80867 , n80869 );
or ( n80871 , n80870 , n45862 );
nand ( n80872 , n80866 , n80871 );
xor ( n80873 , n80859 , n80872 );
nor ( n80874 , n45747 , n45794 );
xnor ( n80875 , n1212 , n37651 );
not ( n80876 , n80875 );
not ( n80877 , n45861 );
and ( n80878 , n80876 , n80877 );
and ( n80879 , n45776 , n42065 );
nor ( n80880 , n80879 , n45774 );
nor ( n80881 , n80880 , n45862 );
nor ( n80882 , n80878 , n80881 );
nor ( n80883 , n45774 , n45861 );
not ( n80884 , n80883 );
nand ( n80885 , n80884 , n45777 );
nor ( n80886 , n80882 , n80885 );
xor ( n80887 , n80874 , n80886 );
or ( n80888 , n80870 , n45861 );
or ( n80889 , n80875 , n45862 );
nand ( n80890 , n80888 , n80889 );
and ( n80891 , n80887 , n80890 );
or ( n80892 , n80891 , C0 );
and ( n80893 , n80873 , n80892 );
and ( n80894 , n80859 , n80872 );
or ( n80895 , n80893 , n80894 );
not ( n80896 , n80895 );
not ( n80897 , n45789 );
and ( n80898 , n45860 , n44004 );
not ( n80899 , n80864 );
nor ( n80900 , n80899 , n45862 );
nor ( n80901 , n80898 , n80900 );
nand ( n80902 , n80897 , n80901 );
not ( n80903 , n80902 );
or ( n80904 , n80896 , n80903 );
not ( n80905 , n80897 );
not ( n80906 , n80901 );
nand ( n80907 , n80905 , n80906 );
nand ( n80908 , n80904 , n80907 );
xor ( n80909 , n45793 , n80908 );
and ( n80910 , n80909 , n45866 );
and ( n80911 , n45793 , n80908 );
or ( n80912 , n80910 , n80911 );
and ( n80913 , n80858 , n80912 );
and ( n80914 , n45870 , n45929 );
or ( n80915 , n80913 , n80914 );
not ( n80916 , n80915 );
or ( n80917 , n46020 , n45933 );
not ( n80918 , n80917 );
or ( n80919 , n80916 , n80918 );
nand ( n80920 , n45933 , n46020 );
nand ( n80921 , n80919 , n80920 );
and ( n80922 , n80857 , n80921 );
and ( n80923 , n46084 , n46024 );
nor ( n80924 , n80922 , n80923 );
or ( n80925 , n80856 , n80924 );
nand ( n80926 , n46173 , n46088 );
nand ( n80927 , n80925 , n80926 );
not ( n80928 , n80927 );
or ( n80929 , n46255 , n46177 );
not ( n80930 , n80929 );
or ( n80931 , n80928 , n80930 );
nand ( n80932 , n46255 , n46177 );
nand ( n80933 , n80931 , n80932 );
not ( n80934 , n80933 );
or ( n80935 , n80855 , n80934 );
nand ( n80936 , n46368 , n46259 );
nand ( n80937 , n80935 , n80936 );
not ( n80938 , n80937 );
or ( n80939 , n80853 , n80938 );
nand ( n80940 , n46483 , n46372 );
nand ( n80941 , n80939 , n80940 );
not ( n80942 , n80941 );
or ( n80943 , n80851 , n80942 );
nand ( n80944 , n46622 , n46487 );
nand ( n80945 , n80943 , n80944 );
not ( n80946 , n80945 );
or ( n80947 , n80849 , n80946 );
nand ( n80948 , n46739 , n46626 );
nand ( n80949 , n80947 , n80948 );
not ( n80950 , n80949 );
or ( n80951 , n80847 , n80950 );
nand ( n80952 , n46902 , n46743 );
not ( n80953 , n80952 );
nand ( n80954 , n47029 , n46906 );
not ( n80955 , n80954 );
or ( n80956 , n80953 , n80955 );
not ( n80957 , n80844 );
nand ( n80958 , n80956 , n80957 );
nand ( n80959 , n80951 , n80958 );
not ( n80960 , n80959 );
or ( n80961 , n80843 , n80960 );
nand ( n80962 , n47200 , n47033 );
nand ( n80963 , n80961 , n80962 );
not ( n80964 , n80963 );
or ( n80965 , n80840 , n80964 );
nand ( n80966 , n47357 , n47204 );
nand ( n80967 , n80965 , n80966 );
not ( n80968 , n80967 );
or ( n80969 , n80837 , n80968 );
nand ( n80970 , n47552 , n47361 );
nand ( n80971 , n80969 , n80970 );
not ( n80972 , n80971 );
or ( n80973 , n80835 , n80972 );
not ( n80974 , n80832 );
and ( n80975 , n47734 , n47556 );
and ( n80976 , n80974 , n80975 );
nand ( n80977 , n47950 , n47738 );
not ( n80978 , n80977 );
nor ( n80979 , n80976 , n80978 );
nand ( n80980 , n80973 , n80979 );
not ( n80981 , n80980 );
or ( n80982 , n80831 , n80981 );
or ( n80983 , n48369 , n48156 );
and ( n80984 , n48152 , n47954 );
and ( n80985 , n80983 , n80984 );
and ( n80986 , n48369 , n48156 );
nor ( n80987 , n80985 , n80986 );
nand ( n80988 , n80982 , n80987 );
nor ( n80989 , n48791 , n48550 );
nor ( n80990 , n48546 , n48373 );
nor ( n80991 , n80989 , n80990 );
nor ( n80992 , n49043 , n48795 );
not ( n80993 , n80992 );
nand ( n80994 , n80988 , n80991 , n80993 );
nand ( n80995 , n48791 , n48550 );
nand ( n80996 , n48546 , n48373 );
and ( n80997 , n80995 , n80996 );
nor ( n80998 , n80997 , n80989 );
nand ( n80999 , n80993 , n80998 );
nand ( n81000 , n48795 , n49043 );
nand ( n81001 , n80994 , n80999 , n81000 );
not ( n81002 , n81001 );
or ( n81003 , n80825 , n81002 );
not ( n81004 , n80822 );
nand ( n81005 , n49328 , n49047 );
not ( n81006 , n81005 );
and ( n81007 , n81004 , n81006 );
nand ( n81008 , n49563 , n49332 );
not ( n81009 , n81008 );
nor ( n81010 , n81007 , n81009 );
nand ( n81011 , n81003 , n81010 );
not ( n81012 , n81011 );
or ( n81013 , n80821 , n81012 );
not ( n81014 , n80818 );
nand ( n81015 , n49855 , n49567 );
not ( n81016 , n81015 );
and ( n81017 , n81014 , n81016 );
and ( n81018 , n50113 , n49859 );
nor ( n81019 , n81017 , n81018 );
nand ( n81020 , n81013 , n81019 );
not ( n81021 , n81020 );
or ( n81022 , n80817 , n81021 );
not ( n81023 , n80814 );
nand ( n81024 , n50421 , n50117 );
not ( n81025 , n81024 );
and ( n81026 , n81023 , n81025 );
nand ( n81027 , n50700 , n50425 );
not ( n81028 , n81027 );
nor ( n81029 , n81026 , n81028 );
nand ( n81030 , n81022 , n81029 );
not ( n81031 , n81030 );
or ( n81032 , n80813 , n81031 );
nand ( n81033 , n51006 , n50704 );
nor ( n81034 , n80810 , n81033 );
not ( n81035 , n51303 );
not ( n81036 , n51630 );
or ( n81037 , n81035 , n81036 );
nand ( n81038 , n51299 , n51010 );
nand ( n81039 , n81037 , n81038 );
or ( n81040 , n81034 , n81039 );
or ( n81041 , n51630 , n51303 );
nand ( n81042 , n81040 , n81041 );
nand ( n81043 , n81032 , n81042 );
not ( n81044 , n81043 );
nor ( n81045 , n52316 , n51960 );
nor ( n81046 , n51956 , n51634 );
nor ( n81047 , n81045 , n81046 );
not ( n81048 , n52650 );
not ( n81049 , n52320 );
nand ( n81050 , n81048 , n81049 );
nand ( n81051 , n81047 , n81050 );
not ( n81052 , n81051 );
not ( n81053 , n81052 );
or ( n81054 , n81044 , n81053 );
nand ( n81055 , n51956 , n51634 );
or ( n81056 , n81045 , n81055 );
nand ( n81057 , n52316 , n51960 );
nand ( n81058 , n81056 , n81057 );
not ( n81059 , n52650 );
nand ( n81060 , n81059 , n81049 );
and ( n81061 , n81058 , n81060 );
and ( n81062 , n52650 , n52320 );
nor ( n81063 , n81061 , n81062 );
nand ( n81064 , n81054 , n81063 );
not ( n81065 , n81064 );
or ( n81066 , n80808 , n81065 );
nor ( n81067 , n53379 , n53026 );
not ( n81068 , n81067 );
nand ( n81069 , n53022 , n52654 );
not ( n81070 , n81069 );
and ( n81071 , n81068 , n81070 );
and ( n81072 , n53379 , n53026 );
nor ( n81073 , n81071 , n81072 );
nand ( n81074 , n81066 , n81073 );
not ( n81075 , n81074 );
or ( n81076 , n80800 , n81075 );
nor ( n81077 , n54123 , n53775 );
nand ( n81078 , n53771 , n53383 );
or ( n81079 , n81077 , n81078 );
nand ( n81080 , n54123 , n53775 );
nand ( n81081 , n81079 , n81080 );
or ( n81082 , n54520 , n54127 );
and ( n81083 , n81081 , n81082 );
and ( n81084 , n54520 , n54127 );
nor ( n81085 , n81083 , n81084 );
nand ( n81086 , n81076 , n81085 );
not ( n81087 , n81086 );
or ( n81088 , n80795 , n81087 );
nor ( n81089 , n55338 , n54919 );
nand ( n81090 , n54915 , n54524 );
or ( n81091 , n81089 , n81090 );
nand ( n81092 , n54919 , n55338 );
nand ( n81093 , n81091 , n81092 );
or ( n81094 , n55342 , n55726 );
and ( n81095 , n81093 , n81094 );
nand ( n81096 , n55342 , n55726 );
not ( n81097 , n81096 );
nor ( n81098 , n81095 , n81097 );
nand ( n81099 , n81088 , n81098 );
not ( n81100 , n81099 );
or ( n81101 , n80790 , n81100 );
nand ( n81102 , n57030 , n56578 );
not ( n81103 , n81102 );
and ( n81104 , n57464 , n57034 );
nor ( n81105 , n81103 , n81104 );
not ( n81106 , n81105 );
nand ( n81107 , n56153 , n55730 );
or ( n81108 , n80782 , n81107 );
nand ( n81109 , n56574 , n56157 );
nand ( n81110 , n81108 , n81109 );
nand ( n81111 , n80788 , n81110 );
not ( n81112 , n81111 );
or ( n81113 , n81106 , n81112 );
not ( n81114 , n57464 );
nand ( n81115 , n81114 , n80786 );
nand ( n81116 , n81113 , n81115 );
nand ( n81117 , n81101 , n81116 );
not ( n81118 , n81117 );
or ( n81119 , n80781 , n81118 );
nand ( n81120 , n59776 , n59274 );
not ( n81121 , n81120 );
not ( n81122 , n81121 );
not ( n81123 , n81122 );
nor ( n81124 , n59776 , n59274 );
not ( n81125 , n81124 );
or ( n81126 , n81123 , n81125 );
not ( n81127 , n58820 );
not ( n81128 , n58366 );
nand ( n81129 , n81127 , n81128 );
not ( n81130 , n81129 );
nor ( n81131 , n58362 , n57938 );
nand ( n81132 , n57468 , n57934 );
or ( n81133 , n81131 , n81132 );
nand ( n81134 , n57938 , n58362 );
nand ( n81135 , n81133 , n81134 );
not ( n81136 , n81135 );
or ( n81137 , n81130 , n81136 );
nand ( n81138 , n58820 , n58366 );
nand ( n81139 , n81137 , n81138 );
or ( n81140 , n59270 , n58824 );
nand ( n81141 , n81139 , n81140 );
nand ( n81142 , n59270 , n58824 );
nand ( n81143 , n81141 , n81122 , n81142 );
nand ( n81144 , n81126 , n81143 );
nand ( n81145 , n81119 , n81144 );
nor ( n81146 , n61749 , n61243 );
not ( n81147 , n81146 );
buf ( n81148 , n60237 );
buf ( n81149 , n59780 );
nor ( n81150 , n81148 , n81149 );
buf ( n81151 , n80752 );
nor ( n81152 , n81150 , n81151 );
not ( n81153 , n61239 );
nand ( n81154 , n81153 , n80749 );
nand ( n81155 , n81147 , n81152 , n81154 );
not ( n81156 , n80769 );
nand ( n81157 , n81156 , n80743 );
nor ( n81158 , n81155 , n81157 );
nand ( n81159 , n81145 , n81158 );
nand ( n81160 , n62790 , n62250 );
nand ( n81161 , n80771 , n81159 , n81160 );
not ( n81162 , n81161 );
or ( n81163 , n80742 , n81162 );
buf ( n81164 , n65417 );
not ( n81165 , n81164 );
not ( n81166 , n64914 );
and ( n81167 , n81165 , n81166 );
buf ( n81168 , n65421 );
nor ( n81169 , n81168 , n65916 );
nor ( n81170 , n81167 , n81169 );
nand ( n81171 , n65916 , n81168 );
not ( n81172 , n81171 );
or ( n81173 , n81170 , n81172 );
not ( n81174 , n64408 );
not ( n81175 , n81174 );
not ( n81176 , n64910 );
not ( n81177 , n81176 );
or ( n81178 , n81175 , n81177 );
not ( n81179 , n64404 );
nand ( n81180 , n81179 , n80734 );
not ( n81181 , n81180 );
nor ( n81182 , n63888 , n63330 );
nand ( n81183 , n63326 , n62794 );
or ( n81184 , n81182 , n81183 );
nand ( n81185 , n63888 , n63330 );
nand ( n81186 , n81184 , n81185 );
not ( n81187 , n81186 );
or ( n81188 , n81181 , n81187 );
nand ( n81189 , n80732 , n63892 );
nand ( n81190 , n81188 , n81189 );
nand ( n81191 , n81178 , n81190 );
nand ( n81192 , n81164 , n64914 );
nand ( n81193 , n64910 , n64408 );
nand ( n81194 , n81191 , n81192 , n81171 , n81193 );
nand ( n81195 , n81173 , n81194 );
nand ( n81196 , n81163 , n81195 );
not ( n81197 , n81196 );
or ( n81198 , n80728 , n81197 );
not ( n81199 , n80725 );
not ( n81200 , n67829 );
not ( n81201 , n67370 );
nand ( n81202 , n81200 , n81201 );
not ( n81203 , n81202 );
not ( n81204 , n67366 );
nand ( n81205 , n81204 , n80716 );
not ( n81206 , n81205 );
nor ( n81207 , n66889 , n66403 );
nand ( n81208 , n66399 , n65920 );
or ( n81209 , n81207 , n81208 );
nand ( n81210 , n66889 , n66403 );
nand ( n81211 , n81209 , n81210 );
not ( n81212 , n81211 );
or ( n81213 , n81206 , n81212 );
buf ( n81214 , n67366 );
nand ( n81215 , n81214 , n66893 );
nand ( n81216 , n81213 , n81215 );
not ( n81217 , n81216 );
or ( n81218 , n81203 , n81217 );
or ( n81219 , n81200 , n81201 );
nand ( n81220 , n81218 , n81219 );
not ( n81221 , n81220 );
or ( n81222 , n81199 , n81221 );
nor ( n81223 , n68283 , n68738 );
nand ( n81224 , n68279 , n67833 );
or ( n81225 , n81223 , n81224 );
nand ( n81226 , n68738 , n68283 );
nand ( n81227 , n81225 , n81226 );
or ( n81228 , n68742 , n69185 );
and ( n81229 , n81227 , n81228 );
nand ( n81230 , n69185 , n68742 );
not ( n81231 , n81230 );
nor ( n81232 , n81229 , n81231 );
nand ( n81233 , n81222 , n81232 );
nand ( n81234 , n80703 , n80704 );
and ( n81235 , n80699 , n80702 , n80726 , n81234 );
and ( n81236 , n81233 , n81235 );
not ( n81237 , n80701 );
nand ( n81238 , n81237 , n70033 );
not ( n81239 , n81238 );
nand ( n81240 , n81239 , n80726 );
nor ( n81241 , n80703 , n80704 );
not ( n81242 , n81241 );
not ( n81243 , n80699 );
or ( n81244 , n81242 , n81243 );
or ( n81245 , n80697 , n80698 );
nand ( n81246 , n81244 , n81245 );
nand ( n81247 , n80726 , n81246 , n80702 );
nand ( n81248 , n70846 , n70450 );
nand ( n81249 , n81240 , n81247 , n81248 );
nor ( n81250 , n81236 , n81249 );
nand ( n81251 , n81198 , n81250 );
not ( n81252 , n81251 );
or ( n81253 , n80696 , n81252 );
not ( n81254 , n80649 );
and ( n81255 , n80652 , n80655 , n80658 );
not ( n81256 , n81255 );
not ( n81257 , n80637 );
not ( n81258 , n80640 );
nor ( n81259 , n71257 , n71645 );
nand ( n81260 , n71253 , n70850 );
or ( n81261 , n81259 , n81260 );
nand ( n81262 , n71257 , n71645 );
nand ( n81263 , n81261 , n81262 );
not ( n81264 , n81263 );
or ( n81265 , n81258 , n81264 );
not ( n81266 , n80639 );
nand ( n81267 , n81266 , n71649 );
nand ( n81268 , n81265 , n81267 );
not ( n81269 , n81268 );
or ( n81270 , n81257 , n81269 );
not ( n81271 , n80636 );
nand ( n81272 , n81271 , n72033 );
nand ( n81273 , n81270 , n81272 );
not ( n81274 , n81273 );
or ( n81275 , n81256 , n81274 );
nand ( n81276 , n72776 , n72416 );
nor ( n81277 , n73139 , n72780 );
or ( n81278 , n81276 , n81277 );
nand ( n81279 , n73139 , n72780 );
nand ( n81280 , n81278 , n81279 );
nand ( n81281 , n80650 , n80651 );
and ( n81282 , n81280 , n81281 );
nor ( n81283 , n80650 , n80651 );
nor ( n81284 , n81282 , n81283 );
nand ( n81285 , n81275 , n81284 );
not ( n81286 , n81285 );
or ( n81287 , n81254 , n81286 );
not ( n81288 , n80646 );
not ( n81289 , n81288 );
nand ( n81290 , n73490 , n73821 );
or ( n81291 , n81290 , n80644 );
nand ( n81292 , n74155 , n73825 );
nand ( n81293 , n81291 , n81292 );
not ( n81294 , n81293 );
or ( n81295 , n81289 , n81294 );
nand ( n81296 , n74466 , n74159 );
nand ( n81297 , n81295 , n81296 );
not ( n81298 , n80647 );
and ( n81299 , n81297 , n81298 );
and ( n81300 , n74470 , n74781 );
nor ( n81301 , n81299 , n81300 );
nand ( n81302 , n81287 , n81301 );
and ( n81303 , n81302 , n80694 );
not ( n81304 , n80681 );
not ( n81305 , n81304 );
not ( n81306 , n80691 );
not ( n81307 , n81306 );
not ( n81308 , n80673 );
not ( n81309 , n80668 );
nor ( n81310 , n75381 , n75083 );
nand ( n81311 , n75079 , n74785 );
or ( n81312 , n81310 , n81311 );
nand ( n81313 , n75381 , n75083 );
nand ( n81314 , n81312 , n81313 );
not ( n81315 , n81314 );
or ( n81316 , n81309 , n81315 );
not ( n81317 , n80667 );
nand ( n81318 , n81317 , n75385 );
nand ( n81319 , n81316 , n81318 );
not ( n81320 , n81319 );
or ( n81321 , n81308 , n81320 );
nand ( n81322 , n75949 , n75673 );
nand ( n81323 , n81321 , n81322 );
not ( n81324 , n81323 );
or ( n81325 , n81307 , n81324 );
nor ( n81326 , n76493 , n76226 );
nand ( n81327 , n75953 , n76222 );
or ( n81328 , n81326 , n81327 );
nand ( n81329 , n76493 , n76226 );
nand ( n81330 , n81328 , n81329 );
buf ( n81331 , n80690 );
and ( n81332 , n81330 , n81331 );
nor ( n81333 , n80688 , n80689 );
nor ( n81334 , n81332 , n81333 );
nand ( n81335 , n81325 , n81334 );
not ( n81336 , n81335 );
or ( n81337 , n81305 , n81336 );
not ( n81338 , n80678 );
not ( n81339 , n81338 );
nor ( n81340 , n77226 , n76996 );
nand ( n81341 , n76992 , n76745 );
or ( n81342 , n81340 , n81341 );
nand ( n81343 , n76996 , n77226 );
nand ( n81344 , n81342 , n81343 );
not ( n81345 , n81344 );
or ( n81346 , n81339 , n81345 );
nand ( n81347 , n77456 , n77230 );
nand ( n81348 , n81346 , n81347 );
not ( n81349 , n80679 );
buf ( n81350 , n81349 );
and ( n81351 , n81348 , n81350 );
and ( n81352 , n77460 , n77671 );
nor ( n81353 , n81351 , n81352 );
nand ( n81354 , n81337 , n81353 );
nor ( n81355 , n81303 , n81354 );
nand ( n81356 , n81253 , n81355 );
not ( n81357 , n81356 );
or ( n81358 , n80629 , n81357 );
not ( n81359 , n80627 );
not ( n81360 , n80616 );
not ( n81361 , n80595 );
not ( n81362 , n80587 );
not ( n81363 , n80585 );
nand ( n81364 , n77887 , n77675 );
or ( n81365 , n80581 , n81364 );
nand ( n81366 , n78092 , n77891 );
nand ( n81367 , n81365 , n81366 );
not ( n81368 , n81367 );
or ( n81369 , n81363 , n81368 );
nand ( n81370 , n78293 , n78096 );
nand ( n81371 , n81369 , n81370 );
not ( n81372 , n81371 );
or ( n81373 , n81362 , n81372 );
nand ( n81374 , n78297 , n78475 );
nand ( n81375 , n81373 , n81374 );
not ( n81376 , n81375 );
or ( n81377 , n81361 , n81376 );
not ( n81378 , n80592 );
nand ( n81379 , n78479 , n78655 );
or ( n81380 , n81379 , n80590 );
nand ( n81381 , n78659 , n78825 );
nand ( n81382 , n81380 , n81381 );
not ( n81383 , n81382 );
or ( n81384 , n81378 , n81383 );
nand ( n81385 , n78829 , n78991 );
nand ( n81386 , n81384 , n81385 );
not ( n81387 , n81386 );
nand ( n81388 , n81377 , n81387 );
not ( n81389 , n81388 );
or ( n81390 , n81360 , n81389 );
not ( n81391 , n80609 );
not ( n81392 , n80602 );
not ( n81393 , n81392 );
not ( n81394 , n80600 );
nand ( n81395 , n79176 , n78995 );
or ( n81396 , n80598 , n81395 );
nand ( n81397 , n79180 , n79328 );
nand ( n81398 , n81396 , n81397 );
not ( n81399 , n81398 );
or ( n81400 , n81394 , n81399 );
nand ( n81401 , n79332 , n79468 );
nand ( n81402 , n81400 , n81401 );
not ( n81403 , n81402 );
or ( n81404 , n81393 , n81403 );
nand ( n81405 , n79472 , n79601 );
nand ( n81406 , n81404 , n81405 );
not ( n81407 , n81406 );
or ( n81408 , n81391 , n81407 );
or ( n81409 , n79839 , n79725 );
and ( n81410 , n79605 , n79721 );
and ( n81411 , n81409 , n81410 );
nand ( n81412 , n79839 , n79725 );
not ( n81413 , n81412 );
nor ( n81414 , n81411 , n81413 );
nand ( n81415 , n81408 , n81414 );
and ( n81416 , n81415 , n80614 );
not ( n81417 , n80610 );
nand ( n81418 , n79843 , n79944 );
or ( n81419 , n81418 , n80612 );
nand ( n81420 , n80049 , n79948 );
nand ( n81421 , n81419 , n81420 );
not ( n81422 , n81421 );
or ( n81423 , n81417 , n81422 );
nand ( n81424 , n80053 , n80135 );
nand ( n81425 , n81423 , n81424 );
nor ( n81426 , n81416 , n81425 );
nand ( n81427 , n81390 , n81426 );
not ( n81428 , n81427 );
or ( n81429 , n81359 , n81428 );
nand ( n81430 , n80220 , n80139 );
or ( n81431 , n81430 , n80620 );
nand ( n81432 , n80283 , n80224 );
nand ( n81433 , n81431 , n81432 );
not ( n81434 , n80626 );
and ( n81435 , n81433 , n81434 );
not ( n81436 , n80625 );
nor ( n81437 , n80349 , n80397 );
nand ( n81438 , n80287 , n80345 );
or ( n81439 , n81437 , n81438 );
nand ( n81440 , n80349 , n80397 );
nand ( n81441 , n81439 , n81440 );
not ( n81442 , n81441 );
or ( n81443 , n81436 , n81442 );
nand ( n81444 , n80401 , n80448 );
nand ( n81445 , n81443 , n81444 );
nor ( n81446 , n81435 , n81445 );
nand ( n81447 , n81429 , n81446 );
buf ( n81448 , n81447 );
not ( n81449 , n81448 );
nand ( n81450 , n81358 , n81449 );
not ( n81451 , n81450 );
or ( n81452 , n80579 , n81451 );
nand ( n81453 , n80452 , n80483 );
nand ( n81454 , n81452 , n81453 );
nor ( n81455 , n80487 , n80519 );
not ( n81456 , n81455 );
nand ( n81457 , n80487 , n80519 );
nand ( n81458 , n81456 , n81457 );
not ( n81459 , n81458 );
and ( n81460 , n81454 , n81459 );
not ( n81461 , n81454 );
and ( n81462 , n81461 , n81458 );
nor ( n81463 , n81460 , n81462 );
not ( n81464 , n80586 );
not ( n81465 , n80582 );
not ( n81466 , n81356 );
or ( n81467 , n81465 , n81466 );
not ( n81468 , n81367 );
nand ( n81469 , n81467 , n81468 );
not ( n81470 , n81469 );
or ( n81471 , n81464 , n81470 );
nand ( n81472 , n81471 , n81370 );
nand ( n81473 , n80587 , n81374 );
not ( n81474 , n81473 );
and ( n81475 , n81472 , n81474 );
not ( n81476 , n81472 );
and ( n81477 , n81476 , n81473 );
nor ( n81478 , n81475 , n81477 );
not ( n81479 , n81288 );
buf ( n81480 , n80659 );
buf ( n81481 , n80645 );
and ( n81482 , n81480 , n81481 );
not ( n81483 , n81482 );
not ( n81484 , n80642 );
not ( n81485 , n81484 );
not ( n81486 , n81251 );
or ( n81487 , n81485 , n81486 );
buf ( n81488 , n81273 );
not ( n81489 , n81488 );
nand ( n81490 , n81487 , n81489 );
not ( n81491 , n81490 );
or ( n81492 , n81483 , n81491 );
buf ( n81493 , n81284 );
not ( n81494 , n81493 );
and ( n81495 , n81494 , n81481 );
buf ( n81496 , n81293 );
nor ( n81497 , n81495 , n81496 );
nand ( n81498 , n81492 , n81497 );
not ( n81499 , n81498 );
or ( n81500 , n81479 , n81499 );
nand ( n81501 , n81500 , n81296 );
not ( n81502 , n81300 );
nand ( n81503 , n81502 , n81298 );
not ( n81504 , n81503 );
and ( n81505 , n81501 , n81504 );
not ( n81506 , n81501 );
and ( n81507 , n81506 , n81503 );
nor ( n81508 , n81505 , n81507 );
not ( n81509 , n80619 );
buf ( n81510 , n80694 );
not ( n81511 , n80588 );
nor ( n81512 , n81511 , n80617 );
nand ( n81513 , n81510 , n81512 );
not ( n81514 , n81513 );
not ( n81515 , n81514 );
buf ( n81516 , n80661 );
not ( n81517 , n81516 );
not ( n81518 , n80727 );
not ( n81519 , n81196 );
or ( n81520 , n81518 , n81519 );
and ( n81521 , n81233 , n81235 );
nor ( n81522 , n81521 , n81249 );
nand ( n81523 , n81520 , n81522 );
not ( n81524 , n81523 );
or ( n81525 , n81517 , n81524 );
not ( n81526 , n81302 );
nand ( n81527 , n81525 , n81526 );
not ( n81528 , n81527 );
or ( n81529 , n81515 , n81528 );
not ( n81530 , n81512 );
not ( n81531 , n81354 );
or ( n81532 , n81530 , n81531 );
not ( n81533 , n81427 );
nand ( n81534 , n81532 , n81533 );
not ( n81535 , n81534 );
nand ( n81536 , n81529 , n81535 );
not ( n81537 , n81536 );
or ( n81538 , n81509 , n81537 );
nand ( n81539 , n81538 , n81430 );
nand ( n81540 , n80621 , n81432 );
not ( n81541 , n81540 );
and ( n81542 , n81539 , n81541 );
not ( n81543 , n81539 );
and ( n81544 , n81543 , n81540 );
nor ( n81545 , n81542 , n81544 );
not ( n81546 , n80604 );
and ( n81547 , n80596 , n81546 );
not ( n81548 , n81547 );
nor ( n81549 , n81548 , n80608 );
not ( n81550 , n81549 );
buf ( n81551 , n81523 );
buf ( n81552 , n80588 );
nand ( n81553 , n80695 , n81552 );
not ( n81554 , n81553 );
nand ( n81555 , n81551 , n81554 );
and ( n81556 , n80694 , n80588 );
and ( n81557 , n81556 , n81302 );
not ( n81558 , n81304 );
not ( n81559 , n81335 );
or ( n81560 , n81558 , n81559 );
nand ( n81561 , n81560 , n81353 );
nand ( n81562 , n81561 , n80588 );
buf ( n81563 , n81375 );
not ( n81564 , n81563 );
nand ( n81565 , n81562 , n81564 );
nor ( n81566 , n81557 , n81565 );
nand ( n81567 , n81555 , n81566 );
not ( n81568 , n81567 );
or ( n81569 , n81550 , n81568 );
not ( n81570 , n81546 );
not ( n81571 , n81386 );
or ( n81572 , n81570 , n81571 );
not ( n81573 , n81406 );
nand ( n81574 , n81572 , n81573 );
not ( n81575 , n80608 );
and ( n81576 , n81574 , n81575 );
nor ( n81577 , n81576 , n81410 );
nand ( n81578 , n81569 , n81577 );
nand ( n81579 , n81409 , n81412 );
not ( n81580 , n81579 );
and ( n81581 , n81578 , n81580 );
not ( n81582 , n81578 );
and ( n81583 , n81582 , n81579 );
nor ( n81584 , n81581 , n81583 );
not ( n81585 , n80594 );
not ( n81586 , n81585 );
not ( n81587 , n81567 );
or ( n81588 , n81586 , n81587 );
nand ( n81589 , n81588 , n81379 );
nand ( n81590 , n80591 , n81381 );
not ( n81591 , n81590 );
and ( n81592 , n81589 , n81591 );
not ( n81593 , n81589 );
and ( n81594 , n81593 , n81590 );
nor ( n81595 , n81592 , n81594 );
nand ( n81596 , n80596 , n80599 );
nor ( n81597 , n81596 , n80601 );
not ( n81598 , n81597 );
not ( n81599 , n81567 );
or ( n81600 , n81598 , n81599 );
not ( n81601 , n80599 );
not ( n81602 , n81386 );
or ( n81603 , n81601 , n81602 );
not ( n81604 , n81398 );
nand ( n81605 , n81603 , n81604 );
or ( n81606 , n79332 , n79468 );
and ( n81607 , n81605 , n81606 );
not ( n81608 , n81401 );
nor ( n81609 , n81607 , n81608 );
nand ( n81610 , n81600 , n81609 );
nand ( n81611 , n81392 , n81405 );
not ( n81612 , n81611 );
and ( n81613 , n81610 , n81612 );
not ( n81614 , n81610 );
and ( n81615 , n81614 , n81611 );
nor ( n81616 , n81613 , n81615 );
not ( n81617 , n80596 );
not ( n81618 , n81567 );
or ( n81619 , n81617 , n81618 );
nand ( n81620 , n81619 , n81387 );
not ( n81621 , n80597 );
nand ( n81622 , n81621 , n81395 );
not ( n81623 , n81622 );
and ( n81624 , n81620 , n81623 );
not ( n81625 , n81620 );
and ( n81626 , n81625 , n81622 );
nor ( n81627 , n81624 , n81626 );
not ( n81628 , n80677 );
and ( n81629 , n80674 , n81306 );
nand ( n81630 , n81551 , n81516 , n81629 );
not ( n81631 , n81526 );
and ( n81632 , n81631 , n81629 );
buf ( n81633 , n81335 );
nor ( n81634 , n81632 , n81633 );
nand ( n81635 , n81630 , n81634 );
not ( n81636 , n81635 );
or ( n81637 , n81628 , n81636 );
not ( n81638 , n81344 );
nand ( n81639 , n81637 , n81638 );
nand ( n81640 , n81338 , n81347 );
not ( n81641 , n81640 );
and ( n81642 , n81639 , n81641 );
not ( n81643 , n81639 );
and ( n81644 , n81643 , n81640 );
nor ( n81645 , n81642 , n81644 );
not ( n81646 , n80675 );
not ( n81647 , n81646 );
not ( n81648 , n81635 );
or ( n81649 , n81647 , n81648 );
nand ( n81650 , n81649 , n81341 );
not ( n81651 , n81340 );
nand ( n81652 , n81651 , n81343 );
not ( n81653 , n81652 );
and ( n81654 , n81650 , n81653 );
not ( n81655 , n81650 );
and ( n81656 , n81655 , n81652 );
nor ( n81657 , n81654 , n81656 );
not ( n81658 , n81484 );
not ( n81659 , n81251 );
or ( n81660 , n81658 , n81659 );
not ( n81661 , n81488 );
nand ( n81662 , n81660 , n81661 );
nand ( n81663 , n81662 , n81480 );
buf ( n81664 , n80643 );
or ( n81665 , n81663 , n81664 );
not ( n81666 , n81664 );
and ( n81667 , n81494 , n81666 );
not ( n81668 , n81290 );
nor ( n81669 , n81667 , n81668 );
nand ( n81670 , n81665 , n81669 );
or ( n81671 , n74155 , n73825 );
nand ( n81672 , n81671 , n81292 );
not ( n81673 , n81672 );
and ( n81674 , n81670 , n81673 );
not ( n81675 , n81670 );
and ( n81676 , n81675 , n81672 );
nor ( n81677 , n81674 , n81676 );
not ( n81678 , n80655 );
nor ( n81679 , n81678 , n81277 );
not ( n81680 , n81679 );
not ( n81681 , n81662 );
or ( n81682 , n81680 , n81681 );
not ( n81683 , n81280 );
nand ( n81684 , n81682 , n81683 );
not ( n81685 , n81283 );
nand ( n81686 , n81685 , n81281 );
not ( n81687 , n81686 );
and ( n81688 , n81684 , n81687 );
not ( n81689 , n81684 );
and ( n81690 , n81689 , n81686 );
nor ( n81691 , n81688 , n81690 );
not ( n81692 , n80578 );
nor ( n81693 , n81692 , n81455 );
nand ( n81694 , n80627 , n81693 );
nor ( n81695 , n81513 , n81694 );
not ( n81696 , n81695 );
not ( n81697 , n81527 );
or ( n81698 , n81696 , n81697 );
not ( n81699 , n81694 );
and ( n81700 , n81699 , n81534 );
not ( n81701 , n81446 );
and ( n81702 , n81701 , n80578 );
not ( n81703 , n81453 );
nor ( n81704 , n81702 , n81703 );
or ( n81705 , n81704 , n81455 );
nand ( n81706 , n81705 , n81457 );
nor ( n81707 , n81700 , n81706 );
nand ( n81708 , n81698 , n81707 );
nor ( n81709 , n80523 , n80543 );
not ( n81710 , n81709 );
nand ( n81711 , n80523 , n80543 );
nand ( n81712 , n81710 , n81711 );
not ( n81713 , n81712 );
and ( n81714 , n81708 , n81713 );
not ( n81715 , n81708 );
and ( n81716 , n81715 , n81712 );
nor ( n81717 , n81714 , n81716 );
nor ( n81718 , n80613 , n80612 );
nand ( n81719 , n80609 , n81718 );
nor ( n81720 , n81548 , n81719 );
not ( n81721 , n81720 );
not ( n81722 , n81567 );
or ( n81723 , n81721 , n81722 );
not ( n81724 , n81719 );
and ( n81725 , n81574 , n81724 );
not ( n81726 , n81414 );
not ( n81727 , n80613 );
and ( n81728 , n81726 , n81727 );
not ( n81729 , n81418 );
nor ( n81730 , n81728 , n81729 );
or ( n81731 , n81730 , n80612 );
nand ( n81732 , n81731 , n81420 );
nor ( n81733 , n81725 , n81732 );
nand ( n81734 , n81723 , n81733 );
nand ( n81735 , n80610 , n81424 );
not ( n81736 , n81735 );
and ( n81737 , n81734 , n81736 );
not ( n81738 , n81734 );
and ( n81739 , n81738 , n81735 );
nor ( n81740 , n81737 , n81739 );
and ( n81741 , n80665 , n80673 , n80669 , n80670 );
nand ( n81742 , n81741 , n80687 );
not ( n81743 , n81742 );
not ( n81744 , n81743 );
buf ( n81745 , n81527 );
not ( n81746 , n81745 );
or ( n81747 , n81744 , n81746 );
not ( n81748 , n80687 );
not ( n81749 , n81323 );
or ( n81750 , n81748 , n81749 );
nand ( n81751 , n81750 , n81327 );
not ( n81752 , n81751 );
nand ( n81753 , n81747 , n81752 );
nand ( n81754 , n80684 , n81329 );
not ( n81755 , n81754 );
and ( n81756 , n81753 , n81755 );
not ( n81757 , n81753 );
and ( n81758 , n81757 , n81754 );
nor ( n81759 , n81756 , n81758 );
nor ( n81760 , n81742 , n81326 );
not ( n81761 , n81760 );
not ( n81762 , n81745 );
or ( n81763 , n81761 , n81762 );
nand ( n81764 , n81751 , n80684 );
and ( n81765 , n81764 , n81329 );
nand ( n81766 , n81763 , n81765 );
not ( n81767 , n81333 );
nand ( n81768 , n81767 , n80690 );
not ( n81769 , n81768 );
and ( n81770 , n81766 , n81769 );
not ( n81771 , n81766 );
and ( n81772 , n81771 , n81768 );
nor ( n81773 , n81770 , n81772 );
not ( n81774 , n80580 );
not ( n81775 , n81774 );
buf ( n81776 , n81356 );
not ( n81777 , n81776 );
or ( n81778 , n81775 , n81777 );
nand ( n81779 , n81778 , n81364 );
not ( n81780 , n80581 );
nand ( n81781 , n81780 , n81366 );
not ( n81782 , n81781 );
and ( n81783 , n81779 , n81782 );
not ( n81784 , n81779 );
and ( n81785 , n81784 , n81781 );
nor ( n81786 , n81783 , n81785 );
not ( n81787 , n81552 );
nand ( n81788 , n81585 , n80591 );
nor ( n81789 , n81787 , n81788 );
not ( n81790 , n81789 );
not ( n81791 , n81776 );
or ( n81792 , n81790 , n81791 );
not ( n81793 , n81585 );
not ( n81794 , n81563 );
or ( n81795 , n81793 , n81794 );
nand ( n81796 , n81795 , n81379 );
and ( n81797 , n81796 , n80591 );
not ( n81798 , n81381 );
nor ( n81799 , n81797 , n81798 );
nand ( n81800 , n81792 , n81799 );
nand ( n81801 , n80592 , n81385 );
not ( n81802 , n81801 );
and ( n81803 , n81800 , n81802 );
not ( n81804 , n81800 );
and ( n81805 , n81804 , n81801 );
nor ( n81806 , n81803 , n81805 );
nor ( n81807 , n81787 , n81596 );
not ( n81808 , n81807 );
not ( n81809 , n81776 );
or ( n81810 , n81808 , n81809 );
buf ( n81811 , n81388 );
and ( n81812 , n81811 , n80599 );
buf ( n81813 , n81398 );
nor ( n81814 , n81812 , n81813 );
nand ( n81815 , n81810 , n81814 );
nand ( n81816 , n81606 , n81401 );
not ( n81817 , n81816 );
and ( n81818 , n81815 , n81817 );
not ( n81819 , n81815 );
and ( n81820 , n81819 , n81816 );
nor ( n81821 , n81818 , n81820 );
nand ( n81822 , n80596 , n81621 );
nor ( n81823 , n81787 , n81822 );
not ( n81824 , n81823 );
not ( n81825 , n81776 );
or ( n81826 , n81824 , n81825 );
and ( n81827 , n81811 , n81621 );
not ( n81828 , n81395 );
nor ( n81829 , n81827 , n81828 );
nand ( n81830 , n81826 , n81829 );
not ( n81831 , n80598 );
nand ( n81832 , n81831 , n81397 );
not ( n81833 , n81832 );
and ( n81834 , n81830 , n81833 );
not ( n81835 , n81830 );
and ( n81836 , n81835 , n81832 );
nor ( n81837 , n81834 , n81836 );
nand ( n81838 , n80609 , n81727 );
nor ( n81839 , n80604 , n81838 );
nand ( n81840 , n80596 , n81839 );
nor ( n81841 , n81787 , n81840 );
not ( n81842 , n81841 );
not ( n81843 , n81776 );
or ( n81844 , n81842 , n81843 );
and ( n81845 , n81811 , n81839 );
not ( n81846 , n81727 );
not ( n81847 , n81415 );
or ( n81848 , n81846 , n81847 );
nand ( n81849 , n81848 , n81418 );
nor ( n81850 , n81845 , n81849 );
nand ( n81851 , n81844 , n81850 );
not ( n81852 , n80612 );
nand ( n81853 , n81852 , n81420 );
not ( n81854 , n81853 );
and ( n81855 , n81851 , n81854 );
not ( n81856 , n81851 );
and ( n81857 , n81856 , n81853 );
nor ( n81858 , n81855 , n81857 );
nand ( n81859 , n81547 , n81552 );
not ( n81860 , n81859 );
not ( n81861 , n81860 );
not ( n81862 , n81776 );
or ( n81863 , n81861 , n81862 );
and ( n81864 , n81563 , n81547 );
nor ( n81865 , n81864 , n81574 );
nand ( n81866 , n81863 , n81865 );
nor ( n81867 , n81410 , n80608 );
and ( n81868 , n81866 , n81867 );
not ( n81869 , n81866 );
not ( n81870 , n81867 );
and ( n81871 , n81869 , n81870 );
nor ( n81872 , n81868 , n81871 );
not ( n81873 , n81512 );
not ( n81874 , n81776 );
or ( n81875 , n81873 , n81874 );
nand ( n81876 , n81875 , n81533 );
nand ( n81877 , n80619 , n81430 );
not ( n81878 , n81877 );
and ( n81879 , n81876 , n81878 );
not ( n81880 , n81876 );
and ( n81881 , n81880 , n81877 );
nor ( n81882 , n81879 , n81881 );
not ( n81883 , n80669 );
not ( n81884 , n80670 );
nor ( n81885 , n81883 , n80664 , n81884 );
not ( n81886 , n81885 );
not ( n81887 , n81745 );
or ( n81888 , n81886 , n81887 );
not ( n81889 , n80668 );
buf ( n81890 , n81314 );
not ( n81891 , n81890 );
or ( n81892 , n81889 , n81891 );
nand ( n81893 , n81892 , n81318 );
not ( n81894 , n81893 );
nand ( n81895 , n81888 , n81894 );
nand ( n81896 , n80673 , n81322 );
not ( n81897 , n81896 );
and ( n81898 , n81895 , n81897 );
not ( n81899 , n81895 );
and ( n81900 , n81899 , n81896 );
nor ( n81901 , n81898 , n81900 );
nor ( n81902 , n80664 , n81884 );
not ( n81903 , n81902 );
not ( n81904 , n81745 );
or ( n81905 , n81903 , n81904 );
not ( n81906 , n81890 );
nand ( n81907 , n81905 , n81906 );
nand ( n81908 , n80669 , n81318 );
not ( n81909 , n81908 );
and ( n81910 , n81907 , n81909 );
not ( n81911 , n81907 );
and ( n81912 , n81911 , n81908 );
nor ( n81913 , n81910 , n81912 );
not ( n81914 , n80670 );
not ( n81915 , n81745 );
or ( n81916 , n81914 , n81915 );
buf ( n81917 , n81311 );
nand ( n81918 , n81916 , n81917 );
nand ( n81919 , n80665 , n81313 );
not ( n81920 , n81919 );
and ( n81921 , n81918 , n81920 );
not ( n81922 , n81918 );
and ( n81923 , n81922 , n81919 );
nor ( n81924 , n81921 , n81923 );
nand ( n81925 , n81288 , n81296 );
not ( n81926 , n81925 );
and ( n81927 , n81498 , n81926 );
not ( n81928 , n81498 );
and ( n81929 , n81928 , n81925 );
nor ( n81930 , n81927 , n81929 );
not ( n81931 , n81480 );
not ( n81932 , n81490 );
or ( n81933 , n81931 , n81932 );
nand ( n81934 , n81933 , n81493 );
nand ( n81935 , n81666 , n81290 );
not ( n81936 , n81935 );
and ( n81937 , n81934 , n81936 );
not ( n81938 , n81934 );
and ( n81939 , n81938 , n81935 );
nor ( n81940 , n81937 , n81939 );
not ( n81941 , n80655 );
not ( n81942 , n81490 );
or ( n81943 , n81941 , n81942 );
nand ( n81944 , n81943 , n81276 );
nand ( n81945 , n80658 , n81279 );
not ( n81946 , n81945 );
and ( n81947 , n81944 , n81946 );
not ( n81948 , n81944 );
and ( n81949 , n81948 , n81945 );
nor ( n81950 , n81947 , n81949 );
not ( n81951 , n80641 );
not ( n81952 , n80630 );
nor ( n81953 , n81952 , n80633 );
not ( n81954 , n81953 );
not ( n81955 , n81251 );
or ( n81956 , n81954 , n81955 );
buf ( n81957 , n81263 );
not ( n81958 , n81957 );
nand ( n81959 , n81956 , n81958 );
not ( n81960 , n81959 );
or ( n81961 , n81951 , n81960 );
buf ( n81962 , n81267 );
nand ( n81963 , n81961 , n81962 );
nand ( n81964 , n80637 , n81272 );
not ( n81965 , n81964 );
and ( n81966 , n81963 , n81965 );
not ( n81967 , n81963 );
and ( n81968 , n81967 , n81964 );
nor ( n81969 , n81966 , n81968 );
not ( n81970 , n81234 );
buf ( n81971 , n80725 );
not ( n81972 , n81971 );
not ( n81973 , n80721 );
not ( n81974 , n81196 );
or ( n81975 , n81973 , n81974 );
buf ( n81976 , n81220 );
not ( n81977 , n81976 );
nand ( n81978 , n81975 , n81977 );
not ( n81979 , n81978 );
or ( n81980 , n81972 , n81979 );
and ( n81981 , n81227 , n81228 );
nor ( n81982 , n81981 , n81231 );
not ( n81983 , n81982 );
not ( n81984 , n81983 );
nand ( n81985 , n81980 , n81984 );
not ( n81986 , n81985 );
or ( n81987 , n81970 , n81986 );
not ( n81988 , n80704 );
nand ( n81989 , n81988 , n69189 );
nand ( n81990 , n81987 , n81989 );
nand ( n81991 , n80699 , n81245 );
not ( n81992 , n81991 );
and ( n81993 , n81990 , n81992 );
not ( n81994 , n81990 );
and ( n81995 , n81994 , n81991 );
nor ( n81996 , n81993 , n81995 );
nor ( n81997 , n81455 , n81709 );
not ( n81998 , n80547 );
not ( n81999 , n80563 );
nand ( n82000 , n81998 , n81999 );
and ( n82001 , n81997 , n82000 );
nand ( n82002 , n80628 , n82001 , n80578 );
not ( n82003 , n82002 );
not ( n82004 , n82003 );
not ( n82005 , n81776 );
or ( n82006 , n82004 , n82005 );
not ( n82007 , n82001 );
not ( n82008 , n80578 );
not ( n82009 , n81447 );
or ( n82010 , n82008 , n82009 );
nand ( n82011 , n82010 , n81453 );
not ( n82012 , n82011 );
or ( n82013 , n82007 , n82012 );
or ( n82014 , n81457 , n81709 );
nand ( n82015 , n82014 , n81711 );
and ( n82016 , n82015 , n82000 );
nor ( n82017 , n81998 , n81999 );
nor ( n82018 , n82016 , n82017 );
nand ( n82019 , n82013 , n82018 );
not ( n82020 , n82019 );
nand ( n82021 , n82006 , n82020 );
nor ( n82022 , n80567 , n80573 );
and ( n82023 , n80567 , n80573 );
nor ( n82024 , n82022 , n82023 );
and ( n82025 , n82021 , n82024 );
not ( n82026 , n82021 );
not ( n82027 , n82024 );
and ( n82028 , n82026 , n82027 );
nor ( n82029 , n82025 , n82028 );
not ( n82030 , n80628 );
nand ( n82031 , n80578 , n81997 );
nor ( n82032 , n82030 , n82031 );
not ( n82033 , n82032 );
not ( n82034 , n81776 );
or ( n82035 , n82033 , n82034 );
not ( n82036 , n82031 );
and ( n82037 , n81448 , n82036 );
not ( n82038 , n81710 );
or ( n82039 , n81453 , n81455 );
nand ( n82040 , n82039 , n81457 );
not ( n82041 , n82040 );
or ( n82042 , n82038 , n82041 );
nand ( n82043 , n82042 , n81711 );
nor ( n82044 , n82037 , n82043 );
nand ( n82045 , n82035 , n82044 );
not ( n82046 , n82017 );
nand ( n82047 , n82046 , n82000 );
not ( n82048 , n82047 );
and ( n82049 , n82045 , n82048 );
not ( n82050 , n82045 );
and ( n82051 , n82050 , n82047 );
nor ( n82052 , n82049 , n82051 );
not ( n82053 , n80624 );
nor ( n82054 , n82053 , n80622 );
and ( n82055 , n80618 , n82054 );
not ( n82056 , n82055 );
not ( n82057 , n81776 );
or ( n82058 , n82056 , n82057 );
not ( n82059 , n80622 );
not ( n82060 , n82059 );
not ( n82061 , n81427 );
or ( n82062 , n82060 , n82061 );
not ( n82063 , n81433 );
nand ( n82064 , n82062 , n82063 );
and ( n82065 , n82064 , n80624 );
not ( n82066 , n81438 );
nor ( n82067 , n82065 , n82066 );
nand ( n82068 , n82058 , n82067 );
nand ( n82069 , n80623 , n81440 );
not ( n82070 , n82069 );
and ( n82071 , n82068 , n82070 );
not ( n82072 , n82068 );
and ( n82073 , n82072 , n82069 );
nor ( n82074 , n82071 , n82073 );
not ( n82075 , n80717 );
buf ( n82076 , n80711 );
not ( n82077 , n82076 );
buf ( n82078 , n81196 );
not ( n82079 , n82078 );
or ( n82080 , n82077 , n82079 );
buf ( n82081 , n81211 );
not ( n82082 , n82081 );
nand ( n82083 , n82080 , n82082 );
not ( n82084 , n82083 );
or ( n82085 , n82075 , n82084 );
buf ( n82086 , n81215 );
nand ( n82087 , n82085 , n82086 );
nand ( n82088 , n81202 , n81219 );
not ( n82089 , n82088 );
and ( n82090 , n82087 , n82089 );
not ( n82091 , n82087 );
and ( n82092 , n82091 , n82088 );
nor ( n82093 , n82090 , n82092 );
nand ( n82094 , n81234 , n81989 );
not ( n82095 , n82094 );
and ( n82096 , n81985 , n82095 );
not ( n82097 , n81985 );
and ( n82098 , n82097 , n82094 );
nor ( n82099 , n82096 , n82098 );
and ( n82100 , n80706 , n81971 );
not ( n82101 , n82100 );
buf ( n82102 , n81978 );
not ( n82103 , n82102 );
or ( n82104 , n82101 , n82103 );
and ( n82105 , n81234 , n80699 );
not ( n82106 , n82105 );
not ( n82107 , n81983 );
or ( n82108 , n82106 , n82107 );
not ( n82109 , n81246 );
nand ( n82110 , n82108 , n82109 );
and ( n82111 , n82110 , n80702 );
nor ( n82112 , n82111 , n81239 );
nand ( n82113 , n82104 , n82112 );
nand ( n82114 , n80726 , n81248 );
not ( n82115 , n82114 );
and ( n82116 , n82113 , n82115 );
not ( n82117 , n82113 );
and ( n82118 , n82117 , n82114 );
nor ( n82119 , n82116 , n82118 );
not ( n82120 , n80630 );
buf ( n82121 , n81551 );
not ( n82122 , n82121 );
or ( n82123 , n82120 , n82122 );
buf ( n82124 , n81260 );
buf ( n82125 , n82124 );
nand ( n82126 , n82123 , n82125 );
nand ( n82127 , n80634 , n81262 );
not ( n82128 , n82127 );
and ( n82129 , n82126 , n82128 );
not ( n82130 , n82126 );
and ( n82131 , n82130 , n82127 );
nor ( n82132 , n82129 , n82131 );
nand ( n82133 , n80655 , n81276 );
not ( n82134 , n82133 );
and ( n82135 , n81662 , n82134 );
not ( n82136 , n81662 );
and ( n82137 , n82136 , n82133 );
nor ( n82138 , n82135 , n82137 );
nand ( n82139 , n80670 , n81917 );
not ( n82140 , n82139 );
and ( n82141 , n81745 , n82140 );
not ( n82142 , n81745 );
and ( n82143 , n82142 , n82139 );
nor ( n82144 , n82141 , n82143 );
not ( n82145 , n80735 );
not ( n82146 , n80731 );
buf ( n82147 , n81159 );
buf ( n82148 , n80771 );
nand ( n82149 , n82147 , n82148 , n81160 );
buf ( n82150 , n82149 );
not ( n82151 , n82150 );
or ( n82152 , n82146 , n82151 );
buf ( n82153 , n81186 );
not ( n82154 , n82153 );
nand ( n82155 , n82152 , n82154 );
not ( n82156 , n82155 );
or ( n82157 , n82145 , n82156 );
nand ( n82158 , n82157 , n81189 );
nand ( n82159 , n81193 , n80736 );
not ( n82160 , n82159 );
and ( n82161 , n82158 , n82160 );
not ( n82162 , n82158 );
and ( n82163 , n82162 , n82159 );
nor ( n82164 , n82161 , n82163 );
nand ( n82165 , n80630 , n82125 );
not ( n82166 , n82165 );
and ( n82167 , n82121 , n82166 );
not ( n82168 , n82121 );
and ( n82169 , n82168 , n82165 );
nor ( n82170 , n82167 , n82169 );
not ( n82171 , n80724 );
nand ( n82172 , n82171 , n81224 );
not ( n82173 , n82172 );
and ( n82174 , n82102 , n82173 );
not ( n82175 , n82102 );
and ( n82176 , n82175 , n82172 );
nor ( n82177 , n82174 , n82176 );
or ( n82178 , n81164 , n64914 );
not ( n82179 , n82178 );
buf ( n82180 , n80737 );
not ( n82181 , n82180 );
not ( n82182 , n82181 );
not ( n82183 , n82150 );
or ( n82184 , n82182 , n82183 );
and ( n82185 , n81191 , n81193 );
nand ( n82186 , n82184 , n82185 );
not ( n82187 , n82186 );
or ( n82188 , n82179 , n82187 );
nand ( n82189 , n82188 , n81192 );
or ( n82190 , n81172 , n81169 );
not ( n82191 , n82190 );
and ( n82192 , n82189 , n82191 );
not ( n82193 , n82189 );
and ( n82194 , n82193 , n82190 );
nor ( n82195 , n82192 , n82194 );
not ( n82196 , n80710 );
not ( n82197 , n82196 );
not ( n82198 , n82078 );
or ( n82199 , n82197 , n82198 );
buf ( n82200 , n81208 );
nand ( n82201 , n82199 , n82200 );
not ( n82202 , n80709 );
nand ( n82203 , n82202 , n81210 );
not ( n82204 , n82203 );
and ( n82205 , n82201 , n82204 );
not ( n82206 , n82201 );
and ( n82207 , n82206 , n82203 );
nor ( n82208 , n82205 , n82207 );
nand ( n82209 , n82196 , n82200 );
not ( n82210 , n82209 );
and ( n82211 , n82078 , n82210 );
not ( n82212 , n82078 );
and ( n82213 , n82212 , n82209 );
nor ( n82214 , n82211 , n82213 );
nand ( n82215 , n82178 , n81192 );
not ( n82216 , n82215 );
and ( n82217 , n82186 , n82216 );
not ( n82218 , n82186 );
and ( n82219 , n82218 , n82215 );
nor ( n82220 , n82217 , n82219 );
nand ( n82221 , n80735 , n81189 );
not ( n82222 , n82221 );
and ( n82223 , n82155 , n82222 );
not ( n82224 , n82155 );
and ( n82225 , n82224 , n82221 );
nor ( n82226 , n82223 , n82225 );
not ( n82227 , n80729 );
not ( n82228 , n82227 );
not ( n82229 , n82150 );
or ( n82230 , n82228 , n82229 );
buf ( n82231 , n81183 );
nand ( n82232 , n82230 , n82231 );
not ( n82233 , n80730 );
nand ( n82234 , n82233 , n81185 );
not ( n82235 , n82234 );
and ( n82236 , n82232 , n82235 );
not ( n82237 , n82232 );
and ( n82238 , n82237 , n82234 );
nor ( n82239 , n82236 , n82238 );
not ( n82240 , n80743 );
buf ( n82241 , n80764 );
buf ( n82242 , n82241 );
not ( n82243 , n82242 );
not ( n82244 , n81155 );
buf ( n82245 , n81145 );
nand ( n82246 , n82244 , n82245 );
nand ( n82247 , n82243 , n82246 );
not ( n82248 , n82247 );
or ( n82249 , n82240 , n82248 );
nand ( n82250 , n82249 , n80767 );
nand ( n82251 , n80770 , n81160 );
not ( n82252 , n82251 );
and ( n82253 , n82250 , n82252 );
not ( n82254 , n82250 );
and ( n82255 , n82254 , n82251 );
nor ( n82256 , n82253 , n82255 );
not ( n82257 , n81154 );
not ( n82258 , n81152 );
not ( n82259 , n82245 );
or ( n82260 , n82258 , n82259 );
buf ( n82261 , n80756 );
not ( n82262 , n82261 );
nand ( n82263 , n82260 , n82262 );
not ( n82264 , n82263 );
or ( n82265 , n82257 , n82264 );
nand ( n82266 , n82265 , n80759 );
not ( n82267 , n81146 );
nand ( n82268 , n82267 , n80763 );
not ( n82269 , n82268 );
and ( n82270 , n82266 , n82269 );
not ( n82271 , n82266 );
and ( n82272 , n82271 , n82268 );
nor ( n82273 , n82270 , n82272 );
nand ( n82274 , n80743 , n80767 );
not ( n82275 , n82274 );
and ( n82276 , n82247 , n82275 );
not ( n82277 , n82247 );
and ( n82278 , n82277 , n82274 );
nor ( n82279 , n82276 , n82278 );
not ( n82280 , n81150 );
not ( n82281 , n82280 );
not ( n82282 , n82245 );
or ( n82283 , n82281 , n82282 );
buf ( n82284 , n80753 );
nand ( n82285 , n82283 , n82284 );
not ( n82286 , n81151 );
buf ( n82287 , n80755 );
nand ( n82288 , n82286 , n82287 );
not ( n82289 , n82288 );
and ( n82290 , n82285 , n82289 );
not ( n82291 , n82285 );
and ( n82292 , n82291 , n82288 );
nor ( n82293 , n82290 , n82292 );
buf ( n82294 , n81117 );
not ( n82295 , n80776 );
and ( n82296 , n82294 , n82295 );
nor ( n82297 , n82296 , n81139 );
not ( n82298 , n80778 );
or ( n82299 , n82297 , n82298 );
nand ( n82300 , n82299 , n81142 );
not ( n82301 , n81124 );
buf ( n82302 , n81120 );
nand ( n82303 , n82301 , n82302 );
not ( n82304 , n82303 );
and ( n82305 , n82300 , n82304 );
not ( n82306 , n82300 );
and ( n82307 , n82306 , n82303 );
nor ( n82308 , n82305 , n82307 );
not ( n82309 , n80772 );
nand ( n82310 , n82309 , n82294 );
not ( n82311 , n80774 );
or ( n82312 , n82310 , n82311 );
not ( n82313 , n81135 );
nand ( n82314 , n82312 , n82313 );
nand ( n82315 , n80775 , n81138 );
not ( n82316 , n82315 );
and ( n82317 , n82314 , n82316 );
not ( n82318 , n82314 );
and ( n82319 , n82318 , n82315 );
nor ( n82320 , n82317 , n82319 );
not ( n82321 , n82297 );
nand ( n82322 , n81142 , n81140 );
not ( n82323 , n82322 );
and ( n82324 , n82321 , n82323 );
not ( n82325 , n82321 );
and ( n82326 , n82325 , n82322 );
nor ( n82327 , n82324 , n82326 );
buf ( n82328 , n81132 );
nand ( n82329 , n82328 , n82310 );
nand ( n82330 , n80774 , n81134 );
not ( n82331 , n82330 );
and ( n82332 , n82329 , n82331 );
not ( n82333 , n82329 );
and ( n82334 , n82333 , n82330 );
nor ( n82335 , n82332 , n82334 );
buf ( n82336 , n81099 );
not ( n82337 , n82336 );
not ( n82338 , n80784 );
or ( n82339 , n82337 , n82338 );
buf ( n82340 , n81110 );
not ( n82341 , n82340 );
nand ( n82342 , n82339 , n82341 );
buf ( n82343 , n81102 );
nand ( n82344 , n80788 , n82343 );
not ( n82345 , n82344 );
and ( n82346 , n82342 , n82345 );
not ( n82347 , n82342 );
and ( n82348 , n82347 , n82344 );
nor ( n82349 , n82346 , n82348 );
buf ( n82350 , n80783 );
not ( n82351 , n82350 );
not ( n82352 , n82351 );
not ( n82353 , n82336 );
or ( n82354 , n82352 , n82353 );
buf ( n82355 , n81107 );
nand ( n82356 , n82354 , n82355 );
not ( n82357 , n80782 );
nand ( n82358 , n82357 , n81109 );
not ( n82359 , n82358 );
and ( n82360 , n82356 , n82359 );
not ( n82361 , n82356 );
and ( n82362 , n82361 , n82358 );
nor ( n82363 , n82360 , n82362 );
buf ( n82364 , n81074 );
not ( n82365 , n80798 );
nand ( n82366 , n82364 , n82365 );
or ( n82367 , n82366 , n80797 );
not ( n82368 , n81081 );
nand ( n82369 , n82367 , n82368 );
not ( n82370 , n81084 );
nand ( n82371 , n82370 , n81082 );
not ( n82372 , n82371 );
and ( n82373 , n82369 , n82372 );
not ( n82374 , n82369 );
and ( n82375 , n82374 , n82371 );
nor ( n82376 , n82373 , n82375 );
not ( n82377 , n80793 );
not ( n82378 , n82377 );
buf ( n82379 , n81086 );
buf ( n82380 , n82379 );
not ( n82381 , n82380 );
or ( n82382 , n82378 , n82381 );
nand ( n82383 , n82382 , n81090 );
not ( n82384 , n81046 );
not ( n82385 , n82384 );
not ( n82386 , n80812 );
not ( n82387 , n81030 );
or ( n82388 , n82386 , n82387 );
nand ( n82389 , n82388 , n81042 );
buf ( n82390 , n82389 );
not ( n82391 , n82390 );
or ( n82392 , n82385 , n82391 );
nand ( n82393 , n82392 , n81055 );
buf ( n82394 , n81030 );
not ( n82395 , n80811 );
nand ( n82396 , n82394 , n82395 );
nand ( n82397 , n81033 , n82396 );
not ( n82398 , n80815 );
not ( n82399 , n82398 );
not ( n82400 , n81020 );
or ( n82401 , n82399 , n82400 );
nand ( n82402 , n82401 , n81024 );
buf ( n82403 , n80988 );
nand ( n82404 , n82403 , n80991 );
nand ( n82405 , n82284 , n82280 );
not ( n82406 , n82405 );
nand ( n82407 , n80717 , n82086 );
nand ( n82408 , n82309 , n82328 );
not ( n82409 , n80833 );
not ( n82410 , n82409 );
not ( n82411 , n80971 );
or ( n82412 , n82410 , n82411 );
not ( n82413 , n80975 );
nand ( n82414 , n82412 , n82413 );
not ( n82415 , n80677 );
not ( n82416 , n81334 );
not ( n82417 , n82416 );
or ( n82418 , n82415 , n82417 );
nand ( n82419 , n82418 , n81638 );
and ( n82420 , n82419 , n81338 );
not ( n82421 , n81347 );
nor ( n82422 , n82420 , n82421 );
nor ( n82423 , n80791 , n80793 );
not ( n82424 , n81223 );
buf ( n82425 , n81226 );
nand ( n82426 , n82424 , n82425 );
nand ( n82427 , n82351 , n82355 );
nand ( n82428 , n82377 , n81090 );
nand ( n82429 , n82365 , n81078 );
not ( n82430 , n81058 );
not ( n82431 , n80838 );
nand ( n82432 , n82431 , n80966 );
not ( n82433 , n82432 );
buf ( n82434 , n80963 );
not ( n82435 , n82434 );
or ( n82436 , n82433 , n82435 );
or ( n82437 , n82434 , n82432 );
nand ( n82438 , n82436 , n82437 );
nand ( n82439 , n82384 , n81055 );
not ( n82440 , n80810 );
nand ( n82441 , n82440 , n81038 );
nand ( n82442 , n80687 , n81327 );
not ( n82443 , n82442 );
nor ( n82444 , n82002 , n82022 );
nand ( n82445 , n81023 , n81027 );
nand ( n82446 , n81646 , n81341 );
buf ( n82447 , n80949 );
not ( n82448 , n80845 );
and ( n82449 , n82447 , n82448 );
not ( n82450 , n80952 );
nor ( n82451 , n82449 , n82450 );
not ( n82452 , n82451 );
and ( n82453 , n80957 , n80954 );
not ( n82454 , n82453 );
or ( n82455 , n82452 , n82454 );
or ( n82456 , n82453 , n82451 );
nand ( n82457 , n82455 , n82456 );
not ( n82458 , n81574 );
nand ( n82459 , n82398 , n81024 );
not ( n82460 , n81352 );
nand ( n82461 , n82460 , n81349 );
not ( n82462 , n82461 );
nand ( n82463 , n82448 , n80952 );
not ( n82464 , n82463 );
not ( n82465 , n82447 );
or ( n82466 , n82464 , n82465 );
or ( n82467 , n82447 , n82463 );
nand ( n82468 , n82466 , n82467 );
not ( n82469 , n80819 );
nand ( n82470 , n82469 , n81015 );
not ( n82471 , n80823 );
nand ( n82472 , n82471 , n81005 );
nand ( n82473 , n81004 , n81008 );
nand ( n82474 , n80993 , n81000 );
not ( n82475 , n80945 );
not ( n82476 , n82475 );
and ( n82477 , n80848 , n80948 );
not ( n82478 , n82477 );
or ( n82479 , n82476 , n82478 );
or ( n82480 , n82475 , n82477 );
nand ( n82481 , n82479 , n82480 );
not ( n82482 , n81364 );
nor ( n82483 , n82482 , n80580 );
not ( n82484 , n80990 );
nand ( n82485 , n82484 , n80996 );
not ( n82486 , n80983 );
nor ( n82487 , n82486 , n80986 );
nand ( n82488 , n80586 , n81370 );
nand ( n82489 , n82409 , n82413 );
nand ( n82490 , n80974 , n80977 );
nand ( n82491 , n80836 , n80970 );
and ( n82492 , n81433 , n80624 );
nor ( n82493 , n82492 , n82066 );
or ( n82494 , n82493 , n81437 );
nand ( n82495 , n82494 , n81440 );
not ( n82496 , n80937 );
not ( n82497 , n82496 );
and ( n82498 , n80852 , n80940 );
not ( n82499 , n82498 );
or ( n82500 , n82497 , n82499 );
or ( n82501 , n82496 , n82498 );
nand ( n82502 , n82500 , n82501 );
nand ( n82503 , n82054 , n80623 );
not ( n82504 , n82503 );
nand ( n82505 , n81727 , n81418 );
not ( n82506 , n82505 );
nand ( n82507 , n80854 , n80936 );
not ( n82508 , n82507 );
not ( n82509 , n80933 );
or ( n82510 , n82508 , n82509 );
or ( n82511 , n80933 , n82507 );
nand ( n82512 , n82510 , n82511 );
not ( n82513 , n80927 );
not ( n82514 , n82513 );
and ( n82515 , n80929 , n80932 );
not ( n82516 , n82515 );
or ( n82517 , n82514 , n82516 );
or ( n82518 , n82515 , n82513 );
nand ( n82519 , n82517 , n82518 );
nand ( n82520 , n80850 , n80944 );
not ( n82521 , n80856 );
nand ( n82522 , n82521 , n80926 );
not ( n82523 , n82522 );
not ( n82524 , n80924 );
not ( n82525 , n82524 );
or ( n82526 , n82523 , n82525 );
or ( n82527 , n82524 , n82522 );
nand ( n82528 , n82526 , n82527 );
nand ( n82529 , n80578 , n81453 );
not ( n82530 , n80921 );
not ( n82531 , n82530 );
not ( n82532 , n80857 );
nor ( n82533 , n82532 , n80923 );
not ( n82534 , n82533 );
or ( n82535 , n82531 , n82534 );
or ( n82536 , n82530 , n82533 );
nand ( n82537 , n82535 , n82536 );
nand ( n82538 , n80917 , n80920 );
not ( n82539 , n82538 );
not ( n82540 , n80915 );
or ( n82541 , n82539 , n82540 );
or ( n82542 , n80915 , n82538 );
nand ( n82543 , n82541 , n82542 );
xor ( n82544 , n45870 , n45929 );
xor ( n82545 , n82544 , n80912 );
xor ( n82546 , n45793 , n80908 );
xor ( n82547 , n82546 , n45866 );
not ( n82548 , n82022 );
not ( n82549 , n80895 );
nand ( n82550 , n80902 , n80907 );
not ( n82551 , n82550 );
or ( n82552 , n82549 , n82551 );
or ( n82553 , n80895 , n82550 );
nand ( n82554 , n82552 , n82553 );
xor ( n82555 , n80859 , n80872 );
xor ( n82556 , n82555 , n80892 );
xor ( n82557 , n80874 , n80886 );
xor ( n82558 , n82557 , n80890 );
and ( n82559 , n80882 , n80885 );
nor ( n82560 , n82559 , n80886 );
not ( n82561 , n80571 );
not ( n82562 , n80569 );
buf ( n82563 , n80788 );
not ( n82564 , n82563 );
not ( n82565 , n82342 );
or ( n82566 , n82564 , n82565 );
nand ( n82567 , n82566 , n82343 );
not ( n82568 , n81115 );
nor ( n82569 , n82568 , n81104 );
xor ( n82570 , n82567 , n82569 );
not ( n82571 , n80791 );
nand ( n82572 , n82571 , n81092 );
xnor ( n82573 , n82383 , n82572 );
xnor ( n82574 , n82380 , n82428 );
nand ( n82575 , n80641 , n81267 );
xnor ( n82576 , n81959 , n82575 );
xnor ( n82577 , n82364 , n82429 );
xnor ( n82578 , n80967 , n82491 );
not ( n82579 , n81045 );
nand ( n82580 , n82579 , n81057 );
xnor ( n82581 , n82393 , n82580 );
xnor ( n82582 , n82390 , n82439 );
xnor ( n82583 , n82397 , n82441 );
nand ( n82584 , n82395 , n81033 );
xnor ( n82585 , n82394 , n82584 );
xnor ( n82586 , n82402 , n82445 );
xnor ( n82587 , n81020 , n82459 );
not ( n82588 , n82469 );
not ( n82589 , n81011 );
or ( n82590 , n82588 , n82589 );
nand ( n82591 , n82590 , n81015 );
nor ( n82592 , n81018 , n80818 );
xor ( n82593 , n82591 , n82592 );
not ( n82594 , n82471 );
buf ( n82595 , n81001 );
not ( n82596 , n82595 );
or ( n82597 , n82594 , n82596 );
nand ( n82598 , n82597 , n81005 );
xnor ( n82599 , n82598 , n82473 );
not ( n82600 , n80998 );
nand ( n82601 , n82600 , n82404 );
xnor ( n82602 , n82601 , n82474 );
xnor ( n82603 , n82403 , n82485 );
not ( n82604 , n80829 );
not ( n82605 , n82604 );
not ( n82606 , n80980 );
or ( n82607 , n82605 , n82606 );
not ( n82608 , n80984 );
nand ( n82609 , n82607 , n82608 );
xor ( n82610 , n82609 , n82487 );
xnor ( n82611 , n81469 , n82488 );
nand ( n82612 , n82608 , n82604 );
xnor ( n82613 , n80980 , n82612 );
xnor ( n82614 , n80971 , n82489 );
xnor ( n82615 , n82414 , n82490 );
not ( n82616 , n80356 );
nor ( n82617 , n82616 , n42663 );
and ( n82618 , n71960 , n80356 );
nor ( n82619 , n82618 , n82562 );
xor ( n82620 , n82619 , n82617 );
xor ( n82621 , n82620 , n82561 );
xor ( n82622 , n42883 , n43049 );
and ( n82623 , n42914 , n42916 , n42911 );
nor ( n82624 , n82623 , n42131 );
not ( n82625 , n82624 );
xor ( n82626 , n82625 , n43064 );
xnor ( n82627 , n81635 , n82446 );
xor ( n82628 , n81776 , n82483 );
not ( n82629 , n82171 );
not ( n82630 , n81978 );
or ( n82631 , n82629 , n82630 );
nand ( n82632 , n82631 , n81224 );
xnor ( n82633 , n82632 , n82426 );
xnor ( n82634 , n82083 , n82407 );
xnor ( n82635 , n80941 , n82520 );
not ( n82636 , n81354 );
not ( n82637 , n82001 );
not ( n82638 , n82011 );
or ( n82639 , n82637 , n82638 );
nand ( n82640 , n82639 , n82018 );
and ( n82641 , n82640 , n82548 );
nor ( n82642 , n82641 , n82023 );
nor ( n82643 , n81067 , n81072 );
not ( n82644 , n80609 );
nor ( n82645 , n82644 , n81859 );
and ( n82646 , n82645 , n81510 );
not ( n82647 , n82646 );
not ( n82648 , n81745 );
or ( n82649 , n82647 , n82648 );
nor ( n82650 , n81547 , n81726 );
nand ( n82651 , n82458 , n82650 );
not ( n82652 , n81726 );
nand ( n82653 , n82652 , n82458 , n81562 , n81564 );
or ( n82654 , n81726 , n80609 );
nand ( n82655 , n82651 , n82653 , n82654 );
nand ( n82656 , n82649 , n82655 );
and ( n82657 , n82656 , n82506 );
not ( n82658 , n82656 );
and ( n82659 , n82658 , n82505 );
nor ( n82660 , n82657 , n82659 );
not ( n82661 , n82444 );
not ( n82662 , n81776 );
or ( n82663 , n82661 , n82662 );
nand ( n82664 , n82663 , n82642 );
not ( n82665 , n80577 );
not ( n82666 , n82621 );
or ( n82667 , n82665 , n82666 );
or ( n82668 , n82621 , n80577 );
nand ( n82669 , n82667 , n82668 );
not ( n82670 , n82669 );
and ( n82671 , n82664 , n82670 );
not ( n82672 , n82664 );
and ( n82673 , n82672 , n82669 );
nor ( n82674 , n82671 , n82673 );
not ( n82675 , n81449 );
nor ( n82676 , n82675 , n82529 );
not ( n82677 , n82676 );
not ( n82678 , n82636 );
nand ( n82679 , n81510 , n81527 );
not ( n82680 , n82679 );
or ( n82681 , n82678 , n82680 );
nand ( n82682 , n82681 , n80628 );
not ( n82683 , n82682 );
or ( n82684 , n82677 , n82683 );
and ( n82685 , n81449 , n82636 );
not ( n82686 , n82685 );
not ( n82687 , n82679 );
or ( n82688 , n82686 , n82687 );
not ( n82689 , n80628 );
and ( n82690 , n82689 , n81449 );
not ( n82691 , n82529 );
nor ( n82692 , n82690 , n82691 );
nand ( n82693 , n82688 , n82692 );
nand ( n82694 , n82684 , n82693 );
not ( n82695 , n81741 );
not ( n82696 , n81527 );
or ( n82697 , n82695 , n82696 );
buf ( n82698 , n81323 );
not ( n82699 , n82698 );
nand ( n82700 , n82697 , n82699 );
and ( n82701 , n82700 , n82443 );
not ( n82702 , n82700 );
and ( n82703 , n82702 , n82442 );
nor ( n82704 , n82701 , n82703 );
not ( n82705 , n82472 );
not ( n82706 , n82595 );
or ( n82707 , n82705 , n82706 );
or ( n82708 , n82472 , n82595 );
nand ( n82709 , n82707 , n82708 );
or ( n82710 , n80810 , n81033 );
nand ( n82711 , n82710 , n81038 );
and ( n82712 , n82380 , n82423 );
or ( n82713 , n81090 , n81089 );
nand ( n82714 , n82713 , n81092 );
nor ( n82715 , n82712 , n82714 );
and ( n82716 , n82245 , n82406 );
not ( n82717 , n82245 );
and ( n82718 , n82717 , n82405 );
nor ( n82719 , n82716 , n82718 );
not ( n82720 , n82408 );
not ( n82721 , n82294 );
or ( n82722 , n82720 , n82721 );
or ( n82723 , n82408 , n82294 );
nand ( n82724 , n82722 , n82723 );
not ( n82725 , n82427 );
not ( n82726 , n82336 );
or ( n82727 , n82725 , n82726 );
or ( n82728 , n82427 , n82336 );
nand ( n82729 , n82727 , n82728 );
not ( n82730 , n82059 );
not ( n82731 , n81536 );
or ( n82732 , n82730 , n82731 );
buf ( n82733 , n82063 );
nand ( n82734 , n82732 , n82733 );
nand ( n82735 , n80624 , n81438 );
not ( n82736 , n82735 );
and ( n82737 , n82734 , n82736 );
not ( n82738 , n82734 );
and ( n82739 , n82738 , n82735 );
nor ( n82740 , n82737 , n82739 );
nand ( n82741 , n51303 , n51630 );
nand ( n82742 , n80804 , n80805 );
buf ( n82743 , n81069 );
not ( n82744 , n81052 );
not ( n82745 , n81043 );
or ( n82746 , n82744 , n82745 );
buf ( n82747 , n81063 );
nand ( n82748 , n82746 , n82747 );
nand ( n82749 , n82742 , n82748 );
nand ( n82750 , n82743 , n82749 );
xor ( n82751 , n82750 , n82643 );
and ( n82752 , n81534 , n82504 );
nor ( n82753 , n82752 , n82495 );
not ( n82754 , n82503 );
nand ( n82755 , n82754 , n81527 , n81514 );
nand ( n82756 , n81154 , n80759 );
not ( n82757 , n82756 );
not ( n82758 , n82263 );
or ( n82759 , n82757 , n82758 );
or ( n82760 , n82756 , n82263 );
nand ( n82761 , n82759 , n82760 );
nand ( n82762 , n42281 , n42460 );
and ( n82763 , n82762 , n42402 );
not ( n82764 , n82762 );
and ( n82765 , n82764 , n42401 );
nor ( n82766 , n82763 , n82765 );
nand ( n82767 , n82755 , n82753 );
nand ( n82768 , n80625 , n81444 );
not ( n82769 , n82768 );
and ( n82770 , n82767 , n82769 );
not ( n82771 , n82767 );
and ( n82772 , n82771 , n82768 );
nor ( n82773 , n82770 , n82772 );
nand ( n82774 , n82227 , n82231 );
not ( n82775 , n82774 );
and ( n82776 , n82150 , n82775 );
not ( n82777 , n82150 );
and ( n82778 , n82777 , n82774 );
nor ( n82779 , n82776 , n82778 );
nand ( n82780 , n82394 , n82395 , n82440 );
not ( n82781 , n45152 );
not ( n82782 , n44149 );
or ( n82783 , n82781 , n82782 );
nand ( n82784 , n82783 , n44197 );
not ( n82785 , n82784 );
nand ( n82786 , n44118 , n44207 );
not ( n82787 , n82786 );
or ( n82788 , n82785 , n82787 );
or ( n82789 , n82786 , n82784 );
nand ( n82790 , n82788 , n82789 );
not ( n82791 , n80841 );
nand ( n82792 , n82791 , n80962 );
not ( n82793 , n82792 );
buf ( n82794 , n80959 );
not ( n82795 , n82794 );
or ( n82796 , n82793 , n82795 );
or ( n82797 , n82794 , n82792 );
nand ( n82798 , n82796 , n82797 );
not ( n82799 , n82715 );
and ( n82800 , n81094 , n81096 );
not ( n82801 , n82800 );
or ( n82802 , n82799 , n82801 );
or ( n82803 , n82800 , n82715 );
nand ( n82804 , n82802 , n82803 );
nand ( n82805 , n43689 , n43685 );
not ( n82806 , n82805 );
not ( n82807 , n44889 );
or ( n82808 , n82806 , n82807 );
or ( n82809 , n82805 , n44889 );
nand ( n82810 , n82808 , n82809 );
not ( n82811 , n81062 );
buf ( n82812 , n81060 );
nand ( n82813 , n82811 , n82812 );
not ( n82814 , n82813 );
not ( n82815 , n82390 );
not ( n82816 , n81047 );
or ( n82817 , n82815 , n82816 );
nand ( n82818 , n82817 , n82430 );
not ( n82819 , n82818 );
or ( n82820 , n82814 , n82819 );
or ( n82821 , n82813 , n82818 );
nand ( n82822 , n82820 , n82821 );
buf ( n82823 , n81041 );
nand ( n82824 , n82823 , n82741 );
not ( n82825 , n82824 );
not ( n82826 , n82711 );
nand ( n82827 , n82826 , n82780 );
not ( n82828 , n82827 );
or ( n82829 , n82825 , n82828 );
or ( n82830 , n82824 , n82827 );
nand ( n82831 , n82829 , n82830 );
nand ( n82832 , n40283 , n42208 );
not ( n82833 , n82832 );
nand ( n82834 , n42203 , n42752 );
not ( n82835 , n82834 );
or ( n82836 , n82833 , n82835 );
or ( n82837 , n82832 , n82834 );
nand ( n82838 , n82836 , n82837 );
nand ( n82839 , n82743 , n82742 );
not ( n82840 , n82839 );
and ( n82841 , n82748 , n82840 );
not ( n82842 , n82748 );
and ( n82843 , n82842 , n82839 );
nor ( n82844 , n82841 , n82843 );
not ( n82845 , n44738 );
nand ( n82846 , n82845 , n44760 );
not ( n82847 , n82846 );
nand ( n82848 , n44734 , n44755 );
not ( n82849 , n82848 );
or ( n82850 , n82847 , n82849 );
or ( n82851 , n82846 , n82848 );
nand ( n82852 , n82850 , n82851 );
nand ( n82853 , n44502 , n44580 );
not ( n82854 , n82853 );
not ( n82855 , n44510 );
not ( n82856 , n45071 );
or ( n82857 , n82855 , n82856 );
nand ( n82858 , n82857 , n45474 );
not ( n82859 , n82858 );
or ( n82860 , n82854 , n82859 );
or ( n82861 , n82853 , n82858 );
nand ( n82862 , n82860 , n82861 );
not ( n82863 , n80797 );
nand ( n82864 , n82863 , n81080 );
not ( n82865 , n82864 );
nand ( n82866 , n81078 , n82366 );
not ( n82867 , n82866 );
or ( n82868 , n82865 , n82867 );
or ( n82869 , n82864 , n82866 );
nand ( n82870 , n82868 , n82869 );
not ( n82871 , n41535 );
nand ( n82872 , n82871 , n42138 );
not ( n82873 , n82872 );
not ( n82874 , n42132 );
not ( n82875 , n82625 );
or ( n82876 , n82874 , n82875 );
nand ( n82877 , n82876 , n42134 );
not ( n82878 , n82877 );
or ( n82879 , n82873 , n82878 );
or ( n82880 , n82872 , n82877 );
nand ( n82881 , n82879 , n82880 );
not ( n82882 , n44379 );
nand ( n82883 , n82882 , n44410 );
not ( n82884 , n82883 );
nand ( n82885 , n45041 , n44404 );
not ( n82886 , n82885 );
or ( n82887 , n82884 , n82886 );
or ( n82888 , n82883 , n82885 );
nand ( n82889 , n82887 , n82888 );
nand ( n82890 , n42916 , n42128 );
not ( n82891 , n82890 );
not ( n82892 , n42914 );
or ( n82893 , n82891 , n82892 );
or ( n82894 , n82890 , n42914 );
nand ( n82895 , n82893 , n82894 );
or ( n82896 , n43567 , n44722 );
not ( n82897 , n82896 );
not ( n82898 , n44688 );
not ( n82899 , n44946 );
or ( n82900 , n82898 , n82899 );
nand ( n82901 , n82900 , n44711 );
not ( n82902 , n82901 );
or ( n82903 , n82897 , n82902 );
or ( n82904 , n82896 , n82901 );
nand ( n82905 , n82903 , n82904 );
not ( n82906 , n43470 );
not ( n82907 , n44778 );
or ( n82908 , n82906 , n82907 );
nand ( n82909 , n82908 , n44785 );
nor ( n82910 , n43476 , n44794 );
and ( n82911 , n82909 , n82910 );
not ( n82912 , n82909 );
not ( n82913 , n82910 );
and ( n82914 , n82912 , n82913 );
nor ( n82915 , n82911 , n82914 );
not ( n82916 , n80989 );
nand ( n82917 , n82916 , n80995 );
not ( n82918 , n82917 );
not ( n82919 , n82484 );
not ( n82920 , n82403 );
or ( n82921 , n82919 , n82920 );
nand ( n82922 , n82921 , n80996 );
not ( n82923 , n82922 );
or ( n82924 , n82918 , n82923 );
or ( n82925 , n82917 , n82922 );
nand ( n82926 , n82924 , n82925 );
not ( n82927 , n42073 );
nand ( n82928 , n42053 , n42076 );
not ( n82929 , n82928 );
or ( n82930 , n82927 , n82929 );
or ( n82931 , n42073 , n82928 );
nand ( n82932 , n82930 , n82931 );
not ( n82933 , n82424 );
not ( n82934 , n82632 );
or ( n82935 , n82933 , n82934 );
nand ( n82936 , n82935 , n82425 );
nand ( n82937 , n81228 , n81230 );
not ( n82938 , n82937 );
and ( n82939 , n82936 , n82938 );
not ( n82940 , n82936 );
and ( n82941 , n82940 , n82937 );
nor ( n82942 , n82939 , n82941 );
buf ( n82943 , n45587 );
buf ( n82944 , n44809 );
xor ( n82945 , n82943 , n82944 );
buf ( n82946 , n82945 );
not ( n82947 , n82105 );
not ( n82948 , n81985 );
or ( n82949 , n82947 , n82948 );
nand ( n82950 , n82949 , n82109 );
nand ( n82951 , n81238 , n80702 );
not ( n82952 , n82951 );
and ( n82953 , n82950 , n82952 );
not ( n82954 , n82950 );
and ( n82955 , n82954 , n82951 );
nor ( n82956 , n82953 , n82955 );
nand ( n82957 , n81585 , n81379 );
not ( n82958 , n82957 );
and ( n82959 , n81567 , n82958 );
not ( n82960 , n81567 );
and ( n82961 , n82960 , n82957 );
nor ( n82962 , n82959 , n82961 );
xor ( n82963 , n32034 , n46440 );
not ( n82964 , n42848 );
and ( n82965 , n42169 , n42172 );
not ( n82966 , n82965 );
or ( n82967 , n82964 , n82966 );
or ( n82968 , n82965 , n42848 );
nand ( n82969 , n82967 , n82968 );
xnor ( n82970 , n81011 , n82470 );
buf ( n82971 , n42038 );
buf ( n82972 , n44004 );
xor ( n82973 , n82971 , n82972 );
buf ( n82974 , n82973 );
xnor ( n82975 , n44855 , n45453 );
and ( n82976 , n81306 , n80677 , n81338 );
not ( n82977 , n82461 );
nand ( n82978 , n82977 , n82422 );
or ( n82979 , n82978 , n82700 );
not ( n82980 , n82976 );
nor ( n82981 , n82980 , n82462 );
nand ( n82982 , n82981 , n82700 );
not ( n82983 , n82422 );
not ( n82984 , n82462 );
and ( n82985 , n82983 , n82984 );
nor ( n82986 , n82976 , n82461 );
and ( n82987 , n82422 , n82986 );
nor ( n82988 , n82985 , n82987 );
nand ( n82989 , n82979 , n82982 , n82988 );
not ( C0n , n0 );
and ( C0 , C0n , n0 );
endmodule
