module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
 n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
 n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
 n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
 n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
 n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , 
 n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , 
 n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , 
 n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , 
 n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , 
 n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , 
 n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , 
 n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , 
 n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , 
 n361 , n362 , n363 , n364 , n365 , n366 , n367 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 ;
output n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
 n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
 n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
 n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
 n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
 n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , 
 n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , 
 n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , 
 n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , 
 n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , 
 n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , 
 n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , 
 n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , 
 n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , 
 n361 , n362 , n363 , n364 , n365 , n366 , n367 ;
wire n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , 
 n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , 
 n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , 
 n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , 
 n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , 
 n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , 
 n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , 
 n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , 
 n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , 
 n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , 
 n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , 
 n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , 
 n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , 
 n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , 
 n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , 
 n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , 
 n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , 
 n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , 
 n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , 
 n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , 
 n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , 
 n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , 
 n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , 
 n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , 
 n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , 
 n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , 
 n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , 
 n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , 
 n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , 
 n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , 
 n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , 
 n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , 
 n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , 
 n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , 
 n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , 
 n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , 
 n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , 
 n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , 
 n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , 
 n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , 
 n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , 
 n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , 
 n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , 
 n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , 
 n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , 
 n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , 
 n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , 
 n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , 
 n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , 
 n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , 
 n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , 
 n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , 
 n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , 
 n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , 
 n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , 
 n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , 
 n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , 
 n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , 
 n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , 
 n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , 
 n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , 
 n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , 
 n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , 
 n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , 
 n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , 
 n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , 
 n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , 
 n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , 
 n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , 
 n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , 
 n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , 
 n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , 
 n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , 
 n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , 
 n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , 
 n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , 
 n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , 
 n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , 
 n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , 
 n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , 
 n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , 
 n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , 
 n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , 
 n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , 
 n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , 
 n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , 
 n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , 
 n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , 
 n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , 
 n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , 
 n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , 
 n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , 
 n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , 
 n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , 
 n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , 
 n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , 
 n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , 
 n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , 
 n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , 
 n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , 
 n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , 
 n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , 
 n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , 
 n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , 
 n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , 
 n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , 
 n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , 
 n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , 
 n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , 
 n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , 
 n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , 
 n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , 
 n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , 
 n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , 
 n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , 
 n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , 
 n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , 
 n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , 
 n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , 
 n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , 
 n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , 
 n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , 
 n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , 
 n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , 
 n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , 
 n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , 
 n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , 
 n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , 
 n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , 
 n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , 
 n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , 
 n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , 
 n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , 
 n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , 
 n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , 
 n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , 
 n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , 
 n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , 
 n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , 
 n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , 
 n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , 
 n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , 
 n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , 
 n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , 
 n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , 
 n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , 
 n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , 
 n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , 
 n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , 
 n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , 
 n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , 
 n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , 
 n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , 
 n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , 
 n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , 
 n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , 
 n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , 
 n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , 
 n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , 
 n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , 
 n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , 
 n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , 
 n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , 
 n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , 
 n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , 
 n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , 
 n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , 
 n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , 
 n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , 
 n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , 
 n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , 
 n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , 
 n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , 
 n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , 
 n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , 
 n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , 
 n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , 
 n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , 
 n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , 
 n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , 
 n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , 
 n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , 
 n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , 
 n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , 
 n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , 
 n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , 
 n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , 
 n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , 
 n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , 
 n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , 
 n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , 
 n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , 
 n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , 
 n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , 
 n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , 
 n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , 
 n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , 
 n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , 
 n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , 
 n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , 
 n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , 
 n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , 
 n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , 
 n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , 
 n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , 
 n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , 
 n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , 
 n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , 
 n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , 
 n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , 
 n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , 
 n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , 
 n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , 
 n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , 
 n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , 
 n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , 
 n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , 
 n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , 
 n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , 
 n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , 
 n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , 
 n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , 
 n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , 
 n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , 
 n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , 
 n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , 
 n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , 
 n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , 
 n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , 
 n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , 
 n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , 
 n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , 
 n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , 
 n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , 
 n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , 
 n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , 
 n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , 
 n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , 
 n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , 
 n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , 
 n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , 
 n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , 
 n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , 
 n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , 
 n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , 
 n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , 
 n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , 
 n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , 
 n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , 
 n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , 
 n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , 
 n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , 
 n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , 
 n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , 
 n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , 
 n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , 
 n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , 
 n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , 
 n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , 
 n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , 
 n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , 
 n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , 
 n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , 
 n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , 
 n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , 
 n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , 
 n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , 
 n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , 
 n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , 
 n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , 
 n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , 
 n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , 
 n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , 
 n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , 
 n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , 
 n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , 
 n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , 
 n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , 
 n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , 
 n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , 
 n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , 
 n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , 
 n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , 
 n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , 
 n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , 
 n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , 
 n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , 
 n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , 
 n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , 
 n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , 
 n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , 
 n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , 
 n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , 
 n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , 
 n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , 
 n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , 
 n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , 
 n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , 
 n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , 
 n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , 
 n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , 
 n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , 
 n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , 
 n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , 
 n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , 
 n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , 
 n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , 
 n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , 
 n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , 
 n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , 
 n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , 
 n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , 
 n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , 
 n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , 
 n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , 
 n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , 
 n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , 
 n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , 
 n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , 
 n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , 
 n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , 
 n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , 
 n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , 
 n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , 
 n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , 
 n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , 
 n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , 
 n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , 
 n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , 
 n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , 
 n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , 
 n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , 
 n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , 
 n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , 
 n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , 
 n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , 
 n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , 
 n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , 
 n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , 
 n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , 
 n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , 
 n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , 
 n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , 
 n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , 
 n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , 
 n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , 
 n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , 
 n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , 
 n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , 
 n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , 
 n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , 
 n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , 
 n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , 
 n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , 
 n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , 
 n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , 
 n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , 
 n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , 
 n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , 
 n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , 
 n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , 
 n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , 
 n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , 
 n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , 
 n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , 
 n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , 
 n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , 
 n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , 
 n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , 
 n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , 
 n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , 
 n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , 
 n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , 
 n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , 
 n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , 
 n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , 
 n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , 
 n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , 
 n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , 
 n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , 
 n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , 
 n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , 
 n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , 
 n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , 
 n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , 
 n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , 
 n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , 
 n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , 
 n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , 
 n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , 
 n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , 
 n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , 
 n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , 
 n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , 
 n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , 
 n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , 
 n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , 
 n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , 
 n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , 
 n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , 
 n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , 
 n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , 
 n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , 
 n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , 
 n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , 
 n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , 
 n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , 
 n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , 
 n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , 
 n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , 
 n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , 
 n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , 
 n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , 
 n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , 
 n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , 
 n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , 
 n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , 
 n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , 
 n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , 
 n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , 
 n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , 
 n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , 
 n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , 
 n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , 
 n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , 
 n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , 
 n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , 
 n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , 
 n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , 
 n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , 
 n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , 
 n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , 
 n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , 
 n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , 
 n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , 
 n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , 
 n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , 
 n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , 
 n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , 
 n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , 
 n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , 
 n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , 
 n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , 
 n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , 
 n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , 
 n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , 
 n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , 
 n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , 
 n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , 
 n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , 
 n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , 
 n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , 
 n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , 
 n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , 
 n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , 
 n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , 
 n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , 
 n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , 
 n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , 
 n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , 
 n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , 
 n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , 
 n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , 
 n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , 
 n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , 
 n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , 
 n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , 
 n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , 
 n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , 
 n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , 
 n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , 
 n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , 
 n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , 
 n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , 
 n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , 
 n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , 
 n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , 
 n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , 
 n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , 
 n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , 
 n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , 
 n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , 
 n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , 
 n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , 
 n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , 
 n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , 
 n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , 
 n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , 
 n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , 
 n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , 
 n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , 
 n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , 
 n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , 
 n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , 
 n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , 
 n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , 
 n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , 
 n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , 
 n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , 
 n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , 
 n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , 
 n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , 
 n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , 
 n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , 
 n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , 
 n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , 
 n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , 
 n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , 
 n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , 
 n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , 
 n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , 
 n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , 
 n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , 
 n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , 
 n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , 
 n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , 
 n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , 
 n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , 
 n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , 
 n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , 
 n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , 
 n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , 
 n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , 
 n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , 
 n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , 
 n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , 
 n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , 
 n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , 
 n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , 
 n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , 
 n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , 
 n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , 
 n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , 
 n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , 
 n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , 
 n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , 
 n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , 
 n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , 
 n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , 
 n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , 
 n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , 
 n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , 
 n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , 
 n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , 
 n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , 
 n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , 
 n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , 
 n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , 
 n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , 
 n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , 
 n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , 
 n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , 
 n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , 
 n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , 
 n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , 
 n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , 
 n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , 
 n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , 
 n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , 
 n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , 
 n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , 
 n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , 
 n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , 
 n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , 
 n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , 
 n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , 
 n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , 
 n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , 
 n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , 
 n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , 
 n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , 
 n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , 
 n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , 
 n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , 
 n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , 
 n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , 
 n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , 
 n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , 
 n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , 
 n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , 
 n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , 
 n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , 
 n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , 
 n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , 
 n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , 
 n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , 
 n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , 
 n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , 
 n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , 
 n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , 
 n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , 
 n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , 
 n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , 
 n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , 
 n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , 
 n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , 
 n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , 
 n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , 
 n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , 
 n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , 
 n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , 
 n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , 
 n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , 
 n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , 
 n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , 
 n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , 
 n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , 
 n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , 
 n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , 
 n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , 
 n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , 
 n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , 
 n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , 
 n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , 
 n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , 
 n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , 
 n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , 
 n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , 
 n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , 
 n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , 
 n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , 
 n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , 
 n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , 
 n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , 
 n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , 
 n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , 
 n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , 
 n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , 
 n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , 
 n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , 
 n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , 
 n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , 
 n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , 
 n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , 
 n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , 
 n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , 
 n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , 
 n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , 
 n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , 
 n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , 
 n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , 
 n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , 
 n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , 
 n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , 
 n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , 
 n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , 
 n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , 
 n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , 
 n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , 
 n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , 
 n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , 
 n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , 
 n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , 
 n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , 
 n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , 
 n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , 
 n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , 
 n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , 
 n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , 
 n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , 
 n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , 
 n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , 
 n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , 
 n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , 
 n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , 
 n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , 
 n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , 
 n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , 
 n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , 
 n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , 
 n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , 
 n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , 
 n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , 
 n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , 
 n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , 
 n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , 
 n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , 
 n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , 
 n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , 
 n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , 
 n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , 
 n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , 
 n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , 
 n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , 
 n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , 
 n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , 
 n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , 
 n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , 
 n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , 
 n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , 
 n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , 
 n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , 
 n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , 
 n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , 
 n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , 
 n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , 
 n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , 
 n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , 
 n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , 
 n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , 
 n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , 
 n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , 
 n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , 
 n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , 
 n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , 
 n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , 
 n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , 
 n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , 
 n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , 
 n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , 
 n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , 
 n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , 
 n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , 
 n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , 
 n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , 
 n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , 
 n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , 
 n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , 
 n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , 
 n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , 
 n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , 
 n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , 
 n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , 
 n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , 
 n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , 
 n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , 
 n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , 
 n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , 
 n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , 
 n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , 
 n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , 
 n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , 
 n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , 
 n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , 
 n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , 
 n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , 
 n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , 
 n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , 
 n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , 
 n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , 
 n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , 
 n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , 
 n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , 
 n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , 
 n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , 
 n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , 
 n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , 
 n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , 
 n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , 
 n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , 
 n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , 
 n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , 
 n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , 
 n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , 
 n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , 
 n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , 
 n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , 
 n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , 
 n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , 
 n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , 
 n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , 
 n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , 
 n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , 
 n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , 
 n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , 
 n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , 
 n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , 
 n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , 
 n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , 
 n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , 
 n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , 
 n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , 
 n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , 
 n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , 
 n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , 
 n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , 
 n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , 
 n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , 
 n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , 
 n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , 
 n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , 
 n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , 
 n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , 
 n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , 
 n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , 
 n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , 
 n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , 
 n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , 
 n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , 
 n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , 
 n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , 
 n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , 
 n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , 
 n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , 
 n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , 
 n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , 
 n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , 
 n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , 
 n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , 
 n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , 
 n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , 
 n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , 
 n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , 
 n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , 
 n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , 
 n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , 
 n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , 
 n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , 
 n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , 
 n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , 
 n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , 
 n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , 
 n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , 
 n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , 
 n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , 
 n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , 
 n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , 
 n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , 
 n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , 
 n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , 
 n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , 
 n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , 
 n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , 
 n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , 
 n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , 
 n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , 
 n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , 
 n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , 
 n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , 
 n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , 
 n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , 
 n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , 
 n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , 
 n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , 
 n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , 
 n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , 
 n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , 
 n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , 
 n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , 
 n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , 
 n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , 
 n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , 
 n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , 
 n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , 
 n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , 
 n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , 
 n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , 
 n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , 
 n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , 
 n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , 
 n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , 
 n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , 
 n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , 
 n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , 
 n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , 
 n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , 
 n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , 
 n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , 
 n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , 
 n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , 
 n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , 
 n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , 
 n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , 
 n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , 
 n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , 
 n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , 
 n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , 
 n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , 
 n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , 
 n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , 
 n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , 
 n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , 
 n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , 
 n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , 
 n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , 
 n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , 
 n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , 
 n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , 
 n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , 
 n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , 
 n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , 
 n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , 
 n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , 
 n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , 
 n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , 
 n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , 
 n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , 
 n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , 
 n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , 
 n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , 
 n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , 
 n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , 
 n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , 
 n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , 
 n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , 
 n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , 
 n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , 
 n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , 
 n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , 
 n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , 
 n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , 
 n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , 
 n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , 
 n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , 
 n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , 
 n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , 
 n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , 
 n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , 
 n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , 
 n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , 
 n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , 
 n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , 
 n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , 
 n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , 
 n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , 
 n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , 
 n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , 
 n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , 
 n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , 
 n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , 
 n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , 
 n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , 
 n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , 
 n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , 
 n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , 
 n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , 
 n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , 
 n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , 
 n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , 
 n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , 
 n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , 
 n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , 
 n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , 
 n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , 
 n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , 
 n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , 
 n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , 
 n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , 
 n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , 
 n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , 
 n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , 
 n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , 
 n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , 
 n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , 
 n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , 
 n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , 
 n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , 
 n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , 
 n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , 
 n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , 
 n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , 
 n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , 
 n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , 
 n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , 
 n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , 
 n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , 
 n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , 
 n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , 
 n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , 
 n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , 
 n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , 
 n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , 
 n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , 
 n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , 
 n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , 
 n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , 
 n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , 
 n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , 
 n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , 
 n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , 
 n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , 
 n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , 
 n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , 
 n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , 
 n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , 
 n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , 
 n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , 
 n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , 
 n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , 
 n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , 
 n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , 
 n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , 
 n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , 
 n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , 
 n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , 
 n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , 
 n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , 
 n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , 
 n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , 
 n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , 
 n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , 
 n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , 
 n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , 
 n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , 
 n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , 
 n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , 
 n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , 
 n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , 
 n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , 
 n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , 
 n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , 
 n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , 
 n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , 
 n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , 
 n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , 
 n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , 
 n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , 
 n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , 
 n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , 
 n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , 
 n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , 
 n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , 
 n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , 
 n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , 
 n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , 
 n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , 
 n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , 
 n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , 
 n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , 
 n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , 
 n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , 
 n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , 
 n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , 
 n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , 
 n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , 
 n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , 
 n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , 
 n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , 
 n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , 
 n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , 
 n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , 
 n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , 
 n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , 
 n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , 
 n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , 
 n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , 
 n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , 
 n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , 
 n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , 
 n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , 
 n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , 
 n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , 
 n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , 
 n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , 
 n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , 
 n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , 
 n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , 
 n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , 
 n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , 
 n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , 
 n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , 
 n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , 
 n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , 
 n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , 
 n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , 
 n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , 
 n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , 
 n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , 
 n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , 
 n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , 
 n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , 
 n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , 
 n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , 
 n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , 
 n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , 
 n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , 
 n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , 
 n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , 
 n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , 
 n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , 
 n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , 
 n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , 
 n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , 
 n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , 
 n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , 
 n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , 
 n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , 
 n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , 
 n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , 
 n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , 
 n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , 
 n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , 
 n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , 
 n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , 
 n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , 
 n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , 
 n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , 
 n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , 
 n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , 
 n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , 
 n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , 
 n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , 
 n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , 
 n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , 
 n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , 
 n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , 
 n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , 
 n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , 
 n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , 
 n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , 
 n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , 
 n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , 
 n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , 
 n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , 
 n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , 
 n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , 
 n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , 
 n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , 
 n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , 
 n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , 
 n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , 
 n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , 
 n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , 
 n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , 
 n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , 
 n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , 
 n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , 
 n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , 
 n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , 
 n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , 
 n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , 
 n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , 
 n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , 
 n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , 
 n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , 
 n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , 
 n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , 
 n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , 
 n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , 
 n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , 
 n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , 
 n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , 
 n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , 
 n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , 
 n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , 
 n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , 
 n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , 
 n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , 
 n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , 
 n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , 
 n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , 
 n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , 
 n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , 
 n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , 
 n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , 
 n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , 
 n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , 
 n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , 
 n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , 
 n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , 
 n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , 
 n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , 
 n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , 
 n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , 
 n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , 
 n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , 
 n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , 
 n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , 
 n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , 
 n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , 
 n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , 
 n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , 
 n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , 
 n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , 
 n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , 
 n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , 
 n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , 
 n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , 
 n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , 
 n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , 
 n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , 
 n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , 
 n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , 
 n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , 
 n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , 
 n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , 
 n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , 
 n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , 
 n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , 
 n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , 
 n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , 
 n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , 
 n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , 
 n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , 
 n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , 
 n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , 
 n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , 
 n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , 
 n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , 
 n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , 
 n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , 
 n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , 
 n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , 
 n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , 
 n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , 
 n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , 
 n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , 
 n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , 
 n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , 
 n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , 
 n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , 
 n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , 
 n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , 
 n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , 
 n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , 
 n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , 
 n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , 
 n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , 
 n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , 
 n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , 
 n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , 
 n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , 
 n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , 
 n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , 
 n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , 
 n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , 
 n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , 
 n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , 
 n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , 
 n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , 
 n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , 
 n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , 
 n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , 
 n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , 
 n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , 
 n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , 
 n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , 
 n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , 
 n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , 
 n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , 
 n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , 
 n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , 
 n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , 
 n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , 
 n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , 
 n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , 
 n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , 
 n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , 
 n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , 
 n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , 
 n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , 
 n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , 
 n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , 
 n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , 
 n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , 
 n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , 
 n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , 
 n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , 
 n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , 
 n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , 
 n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , 
 n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , 
 n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , 
 n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , 
 n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , 
 n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , 
 n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , 
 n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , 
 n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , 
 n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , 
 n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , 
 n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , 
 n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , 
 n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , 
 n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , 
 n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , 
 n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , 
 n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , 
 n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , 
 n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , 
 n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , 
 n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , 
 n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , 
 n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , 
 n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , 
 n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , 
 n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , 
 n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , 
 n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , 
 n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , 
 n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , 
 n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , 
 n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , 
 n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , 
 n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , 
 n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , 
 n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , 
 n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , 
 n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , 
 n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , 
 n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , 
 n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , 
 n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , 
 n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , 
 n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , 
 n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , 
 n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , 
 n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , 
 n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , 
 n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , 
 n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , 
 n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , 
 n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , 
 n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , 
 n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , 
 n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , 
 n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , 
 n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , 
 n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , 
 n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , 
 n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , 
 n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , 
 n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , 
 n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , 
 n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , 
 n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , 
 n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , 
 n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , 
 n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , 
 n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , 
 n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , 
 n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , 
 n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , 
 n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , 
 n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , 
 n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , 
 n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , 
 n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , 
 n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , 
 n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , 
 n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , 
 n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , 
 n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , 
 n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , 
 n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , 
 n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , 
 n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , 
 n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , 
 n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , 
 n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , 
 n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , 
 n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , 
 n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , 
 n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , 
 n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , 
 n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , 
 n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , 
 n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , 
 n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , 
 n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , 
 n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , 
 n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , 
 n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , 
 n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , 
 n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , 
 n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , 
 n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , 
 n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , 
 n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , 
 n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , 
 n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , 
 n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , 
 n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , 
 n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , 
 n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , 
 n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , 
 n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , 
 n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , 
 n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , 
 n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , 
 n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , 
 n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , 
 n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , 
 n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , 
 n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , 
 n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , 
 n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , 
 n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , 
 n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , 
 n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , 
 n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , 
 n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , 
 n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , 
 n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , 
 n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , 
 n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , 
 n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , 
 n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , 
 n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , 
 n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , 
 n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , 
 n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , 
 n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , 
 n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , 
 n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , 
 n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , 
 n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , 
 n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , 
 n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , 
 n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , 
 n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , 
 n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , 
 n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , 
 n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , 
 n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , 
 n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , 
 n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , 
 n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , 
 n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , 
 n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , 
 n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , 
 n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , 
 n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , 
 n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , 
 n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , 
 n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , 
 n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , 
 n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , 
 n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , 
 n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , 
 n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , 
 n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , 
 n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , 
 n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , 
 n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , 
 n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , 
 n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , 
 n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , 
 n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , 
 n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , 
 n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , 
 n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , 
 n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , 
 n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , 
 n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , 
 n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , 
 n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , 
 n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , 
 n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , 
 n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , 
 n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , 
 n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , 
 n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , 
 n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , 
 n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , 
 n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , 
 n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , 
 n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , 
 n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , 
 n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , 
 n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , 
 n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , 
 n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , 
 n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , 
 n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , 
 n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , 
 n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , 
 n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , 
 n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , 
 n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , 
 n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , 
 n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , 
 n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , 
 n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , 
 n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , 
 n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , 
 n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , 
 n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , 
 n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , 
 n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , 
 n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , 
 n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , 
 n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , 
 n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , 
 n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , 
 n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , 
 n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , 
 n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , 
 n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , 
 n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , 
 n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , 
 n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , 
 n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , 
 n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , 
 n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , 
 n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , 
 n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , 
 n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , 
 n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , 
 n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , 
 n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , 
 n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , 
 n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , 
 n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , 
 n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , 
 n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , 
 n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , 
 n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , 
 n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , 
 n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , 
 n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , 
 n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , 
 n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , 
 n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , 
 n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , 
 n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , 
 n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , 
 n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , 
 n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , 
 n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , 
 n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , 
 n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , 
 n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , 
 n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , 
 n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , 
 n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , 
 n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , 
 n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , 
 n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , 
 n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , 
 n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , 
 n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , 
 n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , 
 n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , 
 n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , 
 n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , 
 n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , 
 n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , 
 n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , 
 n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , 
 n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , 
 n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , 
 n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , 
 n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , 
 n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , 
 n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , 
 n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , 
 n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , 
 n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , 
 n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , 
 n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , 
 n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , 
 n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , 
 n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , 
 n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , 
 n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , 
 n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , 
 n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , 
 n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , 
 n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , 
 n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , 
 n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , 
 n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , 
 n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , 
 n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , 
 n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , 
 n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , 
 n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , 
 n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , 
 n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , 
 n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , 
 n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , 
 n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , 
 n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , 
 n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , 
 n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , 
 n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , 
 n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , 
 n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , 
 n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , 
 n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , 
 n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , 
 n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , 
 n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , 
 n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , 
 n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , 
 n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , 
 n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , 
 n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , 
 n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , 
 n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , 
 n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , 
 n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , 
 n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , 
 n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , 
 n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , 
 n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , 
 n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , 
 n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , 
 n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , 
 n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , 
 n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , 
 n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , 
 n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , 
 n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , 
 n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , 
 n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , 
 n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , 
 n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , 
 n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , 
 n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , 
 n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , 
 n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , 
 n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , 
 n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , 
 n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , 
 n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , 
 n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , 
 n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , 
 n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , 
 n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , 
 n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , 
 n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , 
 n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , 
 n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , 
 n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , 
 n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , 
 n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , 
 n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , 
 n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , 
 n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , 
 n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , 
 n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , 
 n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , 
 n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , 
 n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , 
 n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , 
 n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , 
 n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , 
 n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , 
 n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , 
 n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , 
 n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , 
 n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , 
 n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , 
 n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , 
 n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , 
 n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , 
 n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , 
 n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , 
 n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , 
 n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , 
 n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , 
 n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , 
 n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , 
 n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , 
 n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , 
 n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , 
 n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , 
 n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , 
 n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , 
 n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , 
 n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , 
 n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , 
 n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , 
 n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , 
 n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , 
 n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , 
 n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , 
 n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , 
 n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , 
 n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , 
 n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , 
 n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , 
 n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , 
 n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , 
 n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , 
 n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , 
 n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , 
 n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , 
 n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , 
 n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , 
 n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , 
 n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , 
 n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , 
 n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , 
 n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , 
 n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , 
 n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , 
 n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , 
 n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , 
 n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , 
 n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , 
 n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , 
 n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , 
 n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , 
 n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , 
 n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , 
 n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , 
 n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , 
 n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , 
 n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , 
 n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , 
 n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , 
 n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , 
 n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , 
 n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , 
 n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , 
 n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , 
 n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , 
 n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , 
 n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , 
 n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , 
 n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , 
 n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , 
 n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , 
 n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , 
 n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , 
 n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , 
 n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , 
 n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , 
 n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , 
 n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , 
 n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , 
 n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , 
 n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , 
 n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , 
 n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , 
 n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , 
 n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , 
 n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , 
 n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , 
 n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , 
 n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , 
 n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , 
 n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , 
 n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , 
 n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , 
 n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , 
 n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , 
 n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , 
 n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , 
 n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , 
 n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , 
 n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , 
 n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , 
 n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , 
 n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , 
 n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , 
 n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , 
 n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , 
 n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , 
 n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , 
 n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , 
 n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , 
 n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , 
 n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , 
 n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , 
 n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , 
 n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , 
 n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , 
 n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , 
 n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , 
 n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , 
 n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , 
 n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , 
 n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , 
 n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , 
 n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , 
 n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , 
 n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , 
 n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , 
 n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , 
 n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , 
 n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , 
 n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , 
 n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , 
 n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , 
 n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , 
 n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , 
 n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , 
 n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , 
 n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , 
 n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , 
 n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , 
 n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , 
 n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , 
 n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , 
 n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , 
 n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , 
 n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , 
 n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , 
 n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , 
 n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , 
 n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , 
 n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , 
 n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , 
 n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , 
 n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , 
 n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , 
 n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , 
 n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , 
 n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , 
 n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , 
 n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , 
 n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , 
 n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , 
 n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , 
 n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , 
 n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , 
 n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , 
 n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , 
 n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , 
 n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , 
 n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , 
 n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , 
 n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , 
 n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , 
 n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , 
 n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , 
 n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , 
 n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , 
 n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , 
 n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , 
 n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , 
 n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , 
 n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , 
 n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , 
 n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , 
 n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , 
 n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , 
 n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , 
 n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , 
 n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , 
 n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , 
 n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , 
 n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , 
 n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , 
 n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , 
 n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , 
 n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , 
 n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , 
 n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , 
 n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , 
 n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , 
 n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , 
 n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , 
 n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , 
 n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , 
 n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , 
 n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , 
 n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , 
 n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , 
 n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , 
 n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , 
 n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , 
 n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , 
 n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , 
 n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , 
 n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , 
 n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , 
 n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , 
 n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , 
 n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , 
 n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , 
 n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , 
 n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , 
 n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , 
 n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , 
 n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , 
 n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , 
 n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , 
 n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , 
 n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , 
 n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , 
 n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , 
 n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , 
 n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , 
 n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , 
 n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , 
 n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , 
 n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , 
 n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , 
 n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , 
 n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , 
 n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , 
 n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , 
 n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , 
 n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , 
 n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , 
 n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , 
 n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , 
 n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , 
 n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , 
 n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , 
 n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , 
 n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , 
 n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , 
 n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , 
 n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , 
 n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , 
 n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , 
 n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , 
 n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , 
 n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , 
 n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , 
 n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , 
 n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , 
 n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , 
 n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , 
 n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , 
 n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , 
 n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , 
 n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , 
 n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , 
 n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , 
 n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , 
 n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , 
 n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , 
 n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , 
 n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , 
 n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , 
 n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , 
 n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , 
 n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , 
 n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , 
 n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , 
 n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , 
 n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , 
 n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , 
 n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , 
 n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , 
 n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , 
 n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , 
 n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , 
 n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , 
 n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , 
 n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , 
 n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , 
 n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , 
 n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , 
 n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , 
 n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , 
 n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , 
 n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , 
 n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , 
 n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , 
 n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , 
 n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , 
 n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , 
 n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , 
 n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , 
 n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , 
 n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , 
 n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , 
 n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , 
 n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , 
 n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , 
 n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , 
 n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , 
 n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , 
 n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , 
 n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , 
 n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , 
 n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , 
 n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , 
 n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , 
 n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , 
 n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , 
 n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , 
 n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , 
 n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , 
 n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , 
 n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , 
 n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , 
 n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , 
 n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , 
 n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , 
 n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , 
 n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , 
 n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , 
 n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , 
 n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , 
 n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , 
 n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , 
 n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , 
 n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , 
 n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , 
 n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , 
 n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , 
 n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , 
 n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , 
 n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , 
 n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , 
 n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , 
 n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , 
 n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , 
 n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , 
 n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , 
 n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , 
 n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , 
 n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , 
 n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , 
 n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , 
 n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , 
 n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , 
 n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , 
 n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , 
 n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , 
 n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , 
 n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , 
 n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , 
 n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , 
 n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , 
 n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , 
 n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , 
 n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , 
 n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , 
 n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , 
 n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , 
 n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , 
 n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , 
 n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , 
 n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , 
 n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , 
 n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , 
 n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , 
 n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , 
 n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , 
 n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , 
 n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , 
 n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , 
 n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , 
 n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , 
 n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , 
 n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , 
 n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , 
 n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , 
 n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , 
 n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , 
 n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , 
 n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , 
 n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , 
 n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , 
 n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , 
 n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , 
 n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , 
 n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , 
 n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , 
 n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , 
 n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , 
 n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , 
 n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , 
 n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , 
 n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , 
 n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , 
 n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , 
 n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , 
 n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , 
 n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , 
 n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , 
 n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , 
 n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , 
 n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , 
 n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , 
 n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , 
 n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , 
 n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , 
 n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , 
 n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , 
 n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , 
 n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , 
 n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , 
 n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , 
 n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , 
 n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , 
 n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , 
 n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , 
 n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , 
 n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , 
 n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , 
 n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , 
 n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , 
 n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , 
 n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , 
 n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , 
 n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , 
 n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , 
 n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , 
 n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , 
 n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , 
 n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , 
 n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , 
 n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , 
 n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , 
 n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , 
 n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , 
 n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , 
 n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , 
 n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , 
 n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , 
 n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , 
 n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , 
 n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , 
 n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , 
 n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , 
 n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , 
 n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , 
 n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , 
 n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , 
 n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , 
 n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , 
 n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , 
 n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , 
 n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , 
 n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , 
 n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , 
 n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , 
 n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , 
 n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , 
 n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , 
 n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , 
 n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , 
 n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , 
 n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , 
 n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , 
 n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , 
 n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , 
 n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , 
 n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , 
 n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , 
 n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , 
 n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , 
 n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , 
 n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , 
 n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , 
 n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , 
 n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , 
 n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , 
 n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , 
 n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , 
 n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , 
 n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , 
 n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , 
 n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , 
 n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , 
 n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , 
 n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , 
 n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , 
 n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , 
 n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , 
 n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , 
 n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , 
 n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , 
 n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , 
 n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , 
 n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , 
 n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , 
 n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , 
 n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , 
 n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , 
 n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , 
 n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , 
 n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , 
 n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , 
 n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , 
 n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , 
 n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , 
 n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , 
 n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , 
 n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , 
 n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , 
 n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , 
 n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , 
 n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , 
 n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , 
 n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , 
 n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , 
 n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , 
 n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , 
 n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , 
 n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , 
 n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , 
 n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , 
 n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , 
 n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , 
 n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , 
 n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , 
 n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , 
 n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , 
 n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , 
 n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , 
 n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , 
 n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , 
 n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , 
 n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , 
 n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , 
 n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , 
 n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , 
 n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , 
 n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , 
 n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , 
 n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , 
 n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , 
 n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , 
 n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , 
 n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , 
 n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , 
 n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , 
 n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , 
 n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , 
 n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , 
 n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , 
 n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , 
 n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , 
 n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , 
 n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , 
 n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , 
 n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , 
 n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , 
 n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , 
 n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , 
 n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , 
 n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , 
 n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , 
 n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , 
 n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , 
 n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , 
 n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , 
 n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , 
 n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , 
 n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , 
 n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , 
 n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , 
 n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , 
 n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , 
 n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , 
 n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , 
 n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , 
 n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , 
 n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , 
 n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , 
 n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , 
 n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , 
 n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , 
 n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , 
 n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , 
 n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , 
 n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , 
 n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , 
 n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , 
 n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , 
 n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , 
 n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , 
 n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , 
 n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , 
 n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , 
 n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , 
 n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , 
 n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , 
 n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , 
 n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , 
 n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , 
 n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , 
 n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , 
 n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , 
 n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , 
 n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , 
 n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , 
 n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , 
 n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , 
 n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , 
 n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , 
 n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , 
 n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , 
 n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , 
 n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , 
 n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , 
 n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , 
 n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , 
 n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , 
 n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , 
 n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , 
 n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , 
 n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , 
 n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , 
 n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , 
 n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , 
 n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , 
 n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , 
 n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , 
 n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , 
 n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , 
 n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , 
 n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , 
 n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , 
 n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , 
 n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , 
 n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , 
 n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , 
 n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , 
 n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , 
 n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , 
 n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , 
 n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , 
 n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , 
 n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , 
 n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , 
 n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , 
 n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , 
 n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , 
 n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , 
 n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , 
 n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , 
 n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , 
 n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , 
 n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , 
 n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , 
 n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , 
 n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , 
 n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , 
 n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , 
 n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , 
 n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , 
 n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , 
 n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , 
 n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , 
 n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , 
 n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , 
 n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , 
 n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , 
 n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , 
 n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , 
 n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , 
 n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , 
 n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , 
 n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , 
 n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , 
 n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , 
 n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , 
 n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , 
 n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , 
 n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , 
 n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , 
 n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , 
 n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , 
 n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , 
 n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , 
 n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , 
 n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , 
 n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , 
 n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , 
 n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , 
 n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , 
 n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , 
 n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , 
 n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , 
 n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , 
 n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , 
 n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , 
 n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , 
 n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , 
 n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , 
 n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , 
 n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , 
 n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , 
 n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , 
 n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , 
 n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , 
 n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , 
 n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , 
 n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , 
 n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , 
 n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , 
 n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , 
 n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , 
 n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , 
 n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , 
 n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , 
 n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , 
 n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , 
 n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , 
 n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , 
 n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , 
 n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , 
 n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , 
 n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , 
 n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , 
 n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , 
 n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , 
 n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , 
 n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , 
 n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , 
 n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , 
 n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , 
 n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , 
 n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , 
 n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , 
 n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , 
 n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , 
 n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , 
 n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , 
 n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , 
 n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , 
 n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , 
 n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , 
 n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , 
 n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , 
 n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , 
 n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , 
 n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , 
 n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , 
 n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , 
 n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , 
 n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , 
 n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , 
 n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , 
 n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , 
 n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , 
 n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , 
 n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , 
 n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , 
 n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , 
 n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , 
 n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , 
 n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , 
 n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , 
 n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , 
 n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , 
 n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , 
 n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , 
 n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , 
 n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , 
 n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , 
 n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , 
 n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , 
 n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , 
 n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , 
 n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , 
 n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , 
 n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , 
 n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , 
 n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , 
 n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , 
 n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , 
 n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , 
 n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , 
 n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , 
 n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , 
 n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , 
 n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , 
 n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , 
 n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , 
 n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , 
 n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , 
 n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , 
 n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , 
 n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , 
 n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , 
 n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , 
 n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , 
 n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , 
 n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , 
 n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , 
 n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , 
 n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , 
 n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , 
 n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , 
 n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , 
 n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , 
 n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , 
 n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , 
 n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , 
 n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , 
 n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , 
 n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , 
 n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , 
 n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , 
 n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , 
 n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , 
 n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , 
 n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , 
 n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , 
 n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , 
 n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , 
 n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , 
 n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , 
 n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , 
 n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , 
 n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , 
 n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , 
 n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , 
 n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , 
 n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , 
 n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , 
 n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , 
 n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , 
 n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , 
 n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , 
 n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , 
 n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , 
 n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , 
 n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , 
 n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , 
 n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , 
 n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , 
 n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , 
 n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , 
 n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , 
 n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , 
 n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , 
 n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , 
 n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , 
 n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , 
 n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , 
 n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , 
 n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , 
 n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , 
 n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , 
 n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , 
 n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , 
 n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , 
 n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , 
 n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , 
 n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , 
 n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , 
 n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , 
 n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , 
 n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , 
 n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , 
 n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , 
 n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , 
 n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , 
 n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , 
 n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , 
 n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , 
 n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , 
 n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , 
 n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , 
 n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , 
 n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , 
 n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , 
 n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , 
 n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , 
 n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , 
 n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , 
 n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , 
 n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , 
 n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , 
 n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , 
 n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , 
 n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , 
 n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , 
 n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , 
 n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , 
 n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , 
 n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , 
 n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , 
 n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , 
 n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , 
 n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , 
 n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , 
 n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , 
 n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , 
 n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , 
 n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , 
 n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , 
 n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , 
 n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , 
 n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , 
 n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , 
 n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , 
 n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , 
 n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , 
 n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , 
 n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , 
 n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , 
 n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , 
 n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , 
 n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , 
 n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , 
 n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , 
 n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , 
 n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , 
 n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , 
 n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , 
 n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , 
 n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , 
 n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , 
 n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , 
 n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , 
 n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , 
 n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , 
 n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , 
 n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , 
 n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , 
 n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , 
 n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , 
 n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , 
 n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , 
 n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , 
 n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , 
 n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , 
 n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , 
 n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , 
 n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , 
 n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , 
 n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , 
 n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , 
 n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , 
 n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , 
 n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , 
 n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , 
 n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , 
 n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , 
 n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , 
 n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , 
 n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , 
 n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , 
 n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , 
 n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , 
 n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , 
 n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , 
 n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , 
 n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , 
 n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , 
 n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , 
 n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , 
 n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , 
 n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , 
 n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , 
 n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , 
 n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , 
 n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , 
 n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , 
 n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , 
 n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , 
 n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , 
 n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , 
 n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , 
 n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , 
 n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , 
 n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , 
 n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , 
 n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , 
 n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , 
 n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , 
 n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , 
 n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , 
 n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , 
 n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , 
 n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , 
 n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , 
 n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , 
 n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , 
 n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , 
 n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , 
 n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , 
 n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , 
 n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , 
 n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , 
 n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , 
 n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , 
 n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , 
 n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , 
 n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , 
 n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , 
 n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , 
 n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , 
 n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , 
 n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , 
 n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , 
 n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , 
 n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , 
 n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , 
 n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , 
 n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , 
 n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , 
 n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , 
 n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , 
 n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , 
 n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , 
 n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , 
 n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , 
 n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , 
 n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , 
 n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , 
 n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , 
 n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , 
 n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , 
 n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , 
 n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , 
 n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , 
 n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , 
 n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , 
 n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , 
 n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , 
 n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , 
 n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , 
 n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , 
 n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , 
 n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , 
 n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , 
 n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , 
 n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , 
 n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , 
 n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , 
 n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , 
 n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , 
 n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , 
 n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , 
 n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , 
 n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , 
 n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , 
 n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , 
 n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , 
 n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , 
 n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , 
 n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , 
 n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , 
 n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , 
 n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , 
 n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , 
 n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , 
 n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , 
 n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , 
 n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , 
 n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , 
 n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , 
 n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , 
 n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , 
 n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , 
 n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , 
 n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , 
 n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , 
 n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , 
 n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , 
 n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , 
 n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , 
 n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , 
 n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , 
 n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , 
 n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , 
 n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , 
 n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , 
 n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , 
 n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , 
 n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , 
 n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , 
 n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , 
 n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , 
 n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , 
 n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , 
 n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , 
 n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , 
 n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , 
 n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , 
 n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , 
 n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , 
 n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , 
 n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , 
 n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , 
 n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , 
 n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , 
 n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , 
 n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , 
 n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , 
 n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , 
 n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , 
 n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , 
 n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , 
 n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , 
 n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , 
 n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , 
 n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , 
 n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , 
 n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , 
 n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , 
 n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , 
 n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , 
 n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , 
 n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , 
 n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , 
 n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , 
 n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , 
 n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , 
 n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , 
 n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , 
 n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , 
 n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , 
 n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , 
 n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , 
 n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , 
 n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , 
 n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , 
 n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , 
 n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , 
 n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , 
 n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , 
 n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , 
 n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , 
 n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , 
 n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , 
 n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , 
 n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , 
 n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , 
 n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , 
 n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , 
 n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , 
 n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , 
 n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , 
 n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , 
 n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , 
 n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , 
 n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , 
 n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , 
 n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , 
 n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , 
 n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , 
 n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , 
 n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , 
 n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , 
 n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , 
 n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , 
 n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , 
 n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , 
 n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , 
 n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , 
 n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , 
 n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , 
 n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , 
 n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , 
 n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , 
 n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , 
 n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , 
 n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , 
 n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , 
 n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , 
 n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , 
 n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , 
 n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , 
 n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , 
 n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , 
 n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , 
 n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , 
 n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , 
 n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , 
 n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , 
 n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , 
 n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , 
 n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , 
 n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , 
 n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , 
 n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , 
 n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , 
 n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , 
 n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , 
 n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , 
 n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , 
 n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , 
 n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , 
 n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , 
 n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , 
 n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , 
 n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , 
 n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , 
 n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , 
 n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , 
 n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , 
 n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , 
 n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , 
 n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , 
 n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , 
 n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , 
 n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , 
 n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , 
 n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , 
 n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , 
 n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , 
 n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , 
 n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , 
 n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , 
 n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , 
 n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , 
 n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , 
 n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , 
 n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , 
 n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , 
 n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , 
 n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , 
 n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , 
 n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , 
 n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , 
 n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , 
 n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , 
 n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , 
 n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , 
 n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , 
 n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , 
 n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , 
 n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , 
 n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , 
 n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , 
 n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , 
 n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , 
 n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , 
 n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , 
 n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , 
 n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , 
 n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , 
 n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , 
 n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , 
 n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , 
 n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , 
 n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , 
 n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , 
 n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , 
 n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , 
 n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , 
 n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , 
 n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , 
 n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , 
 n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , 
 n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , 
 n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , 
 n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , 
 n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , 
 n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , 
 n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , 
 n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , 
 n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , 
 n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , 
 n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , 
 n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , 
 n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , 
 n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , 
 n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , 
 n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , 
 n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , 
 n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , 
 n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , 
 n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , 
 n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , 
 n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , 
 n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , 
 n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , 
 n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , 
 n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , 
 n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , 
 n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , 
 n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , 
 n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , 
 n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , 
 n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , 
 n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , 
 n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , 
 n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , 
 n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , 
 n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , 
 n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , 
 n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , 
 n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , 
 n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , 
 n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , 
 n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , 
 n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , 
 n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , 
 n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , 
 n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , 
 n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , 
 n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , 
 n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , 
 n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , 
 n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , 
 n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , 
 n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , 
 n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , 
 n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , 
 n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , 
 n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , 
 n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , 
 n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , 
 n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , 
 n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , 
 n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , 
 n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , 
 n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , 
 n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , 
 n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , 
 n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , 
 n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , 
 n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , 
 n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , 
 n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , 
 n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , 
 n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , 
 n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , 
 n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , 
 n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , 
 n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , 
 n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , 
 n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , 
 n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , 
 n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , 
 n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , 
 n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , 
 n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , 
 n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , 
 n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , 
 n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , 
 n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , 
 n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , 
 n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , 
 n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , 
 n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , 
 n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , 
 n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , 
 n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , 
 n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , 
 n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , 
 n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , 
 n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , 
 n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , 
 n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , 
 n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , 
 n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , 
 n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , 
 n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , 
 n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , 
 n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , 
 n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , 
 n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , 
 n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , 
 n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , 
 n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , 
 n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , 
 n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , 
 n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , 
 n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , 
 n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , 
 n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , 
 n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , 
 n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , 
 n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , 
 n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , 
 n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , 
 n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , 
 n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , 
 n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , 
 n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , 
 n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , 
 n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , 
 n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , 
 n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , 
 n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , 
 n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , 
 n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , 
 n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , 
 n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , 
 n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , 
 n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , 
 n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , 
 n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , 
 n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , 
 n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , 
 n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , 
 n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , 
 n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , 
 n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , 
 n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , 
 n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , 
 n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , 
 n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , 
 n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , 
 n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , 
 n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , 
 n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , 
 n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , 
 n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , 
 n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , 
 n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , 
 n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , 
 n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , 
 n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , 
 n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , 
 n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , 
 n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , 
 n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , 
 n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , 
 n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , 
 n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , 
 n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , 
 n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , 
 n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , 
 n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , 
 n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , 
 n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , 
 n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , 
 n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , 
 n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , 
 n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , 
 n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , 
 n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , 
 n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , 
 n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , 
 n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , 
 n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , 
 n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , 
 n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , 
 n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , 
 n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , 
 n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , 
 n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , 
 n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , 
 n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , 
 n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , 
 n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , 
 n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , 
 n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , 
 n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , 
 n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , 
 n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , 
 n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , 
 n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , 
 n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , 
 n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , 
 n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , 
 n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , 
 n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , 
 n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , 
 n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , 
 n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , 
 n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , 
 n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , 
 n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , 
 n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , 
 n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , 
 n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , 
 n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , 
 n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , 
 n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , 
 n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , 
 n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , 
 n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , 
 n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , 
 n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , 
 n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , 
 n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , 
 n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , 
 n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , 
 n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , 
 n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , 
 n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , 
 n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , 
 n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , 
 n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , 
 n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , 
 n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , 
 n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , 
 n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , 
 n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , 
 n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , 
 n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , 
 n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , 
 n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , 
 n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , 
 n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , 
 n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , 
 n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , 
 n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , 
 n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , 
 n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , 
 n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , 
 n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , 
 n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , 
 n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , 
 n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , 
 n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , 
 n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , 
 n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , 
 n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , 
 n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , 
 n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , 
 n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , 
 n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , 
 n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , 
 n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , 
 n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , 
 n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , 
 n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , 
 n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , 
 n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , 
 n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , 
 n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , 
 n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , 
 n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , 
 n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , 
 n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , 
 n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , 
 n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , 
 n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , 
 n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , 
 n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , 
 n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , 
 n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , 
 n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , 
 n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , 
 n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , 
 n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , 
 n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , 
 n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , 
 n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , 
 n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , 
 n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , 
 n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , 
 n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , 
 n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , 
 n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , 
 n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , 
 n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , 
 n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , 
 n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , 
 n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , 
 n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , 
 n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , 
 n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , 
 n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , 
 n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , 
 n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , 
 n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , 
 n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , 
 n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , 
 n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , 
 n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , 
 n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , 
 n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , 
 n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , 
 n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , 
 n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , 
 n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , 
 n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , 
 n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , 
 n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , 
 n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , 
 n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , 
 n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , 
 n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , 
 n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , 
 n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , 
 n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , 
 n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , 
 n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , 
 n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , 
 n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , 
 n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , 
 n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , 
 n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , 
 n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , 
 n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , 
 n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , 
 n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , 
 n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , 
 n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , 
 n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , 
 n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , 
 n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , 
 n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , 
 n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , 
 n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , 
 n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , 
 n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , 
 n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , 
 n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , 
 n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , 
 n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , 
 n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , 
 n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , 
 n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , 
 n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , 
 n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , 
 n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , 
 n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , 
 n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , 
 n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , 
 n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , 
 n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , 
 n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , 
 n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , 
 n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , 
 n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , 
 n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , 
 n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , 
 n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , 
 n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , 
 n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , 
 n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , 
 n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , 
 n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , 
 n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , 
 n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , 
 n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , 
 n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , 
 n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , 
 n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , 
 n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , 
 n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , 
 n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , 
 n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , 
 n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , 
 n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , 
 n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , 
 n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , 
 n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , 
 n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , 
 n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , 
 n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , 
 n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , 
 n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , 
 n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , 
 n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , 
 n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , 
 n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , 
 n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , 
 n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , 
 n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , 
 n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , 
 n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , 
 n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , 
 n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , 
 n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , 
 n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , 
 n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , 
 n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , 
 n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , 
 n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , 
 n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , 
 n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , 
 n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , 
 n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , 
 n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , 
 n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , 
 n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , 
 n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , 
 n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , 
 n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , 
 n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , 
 n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , 
 n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , 
 n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , 
 n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , 
 n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , 
 n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , 
 n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , 
 n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , 
 n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , 
 n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , 
 n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , 
 n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , 
 n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , 
 n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , 
 n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , 
 n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , 
 n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , 
 n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , 
 n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , 
 n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , 
 n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , 
 n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , 
 n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , 
 n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , 
 n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , 
 n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , 
 n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , 
 n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , 
 n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , 
 n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , 
 n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , 
 n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , 
 n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , 
 n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , 
 n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , 
 n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , 
 n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , 
 n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , 
 n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , 
 n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , 
 n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , 
 n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , 
 n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , 
 n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , 
 n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , 
 n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , 
 n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , 
 n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , 
 n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , 
 n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , 
 n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , 
 n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , 
 n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , 
 n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , 
 n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , 
 n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , 
 n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , 
 n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , 
 n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , 
 n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , 
 n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , 
 n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , 
 n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , 
 n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , 
 n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , 
 n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , 
 n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , 
 n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , 
 n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , 
 n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , 
 n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , 
 n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , 
 n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , 
 n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , 
 n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , 
 n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , 
 n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , 
 n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , 
 n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , 
 n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , 
 n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , 
 n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , 
 n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , 
 n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , 
 n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , 
 n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , 
 n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , 
 n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , 
 n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , 
 n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , 
 n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , 
 n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , 
 n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , 
 n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , 
 n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , 
 n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , 
 n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , 
 n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , 
 n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , 
 n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , 
 n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , 
 n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , 
 n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , 
 n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , 
 n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , 
 n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , 
 n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , 
 n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , 
 n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , 
 n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , 
 n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , 
 n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , 
 n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , 
 n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , 
 n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , 
 n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , 
 n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , 
 n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , 
 n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , 
 n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , 
 n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , 
 n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , 
 n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , 
 n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , 
 n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , 
 n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , 
 n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , 
 n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , 
 n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , 
 n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , 
 n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , 
 n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , 
 n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , 
 n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , 
 n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , 
 n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , 
 n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , 
 n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , 
 n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , 
 n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , 
 n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , 
 n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , 
 n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , 
 n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , 
 n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , 
 n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , 
 n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , 
 n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , 
 n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , 
 n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , 
 n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , 
 n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , 
 n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , 
 n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , 
 n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , 
 n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , 
 n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , 
 n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , 
 n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , 
 n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , 
 n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , 
 n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , 
 n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , 
 n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , 
 n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , 
 n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , 
 n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , 
 n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , 
 n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , 
 n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , 
 n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , 
 n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , 
 n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , 
 n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , 
 n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , 
 n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , 
 n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , 
 n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , 
 n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , 
 n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , 
 n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , 
 n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , 
 n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , 
 n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , 
 n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , 
 n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , 
 n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , 
 n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , 
 n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , 
 n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , 
 n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , 
 n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , 
 n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , 
 n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , 
 n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , 
 n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , 
 n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , 
 n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , 
 n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , 
 n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , 
 n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , 
 n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , 
 n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , 
 n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , 
 n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , 
 n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , 
 n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , 
 n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , 
 n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , 
 n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , 
 n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , 
 n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , 
 n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , 
 n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , 
 n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , 
 n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , 
 n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , 
 n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , 
 n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , 
 n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , 
 n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , 
 n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , 
 n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , 
 n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , 
 n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , 
 n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , 
 n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , 
 n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , 
 n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , 
 n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , 
 n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , 
 n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , 
 n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , 
 n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , 
 n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , 
 n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , 
 n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , 
 n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , 
 n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , 
 n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , 
 n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , 
 n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , 
 n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , 
 n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , 
 n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , 
 n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , 
 n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , 
 n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , 
 n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , 
 n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , 
 n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , 
 n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , 
 n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , 
 n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , 
 n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , 
 n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , 
 n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , 
 n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , 
 n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , 
 n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , 
 n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , 
 n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , 
 n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , 
 n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , 
 n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , 
 n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , 
 n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , 
 n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , 
 n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , 
 n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , 
 n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , 
 n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , 
 n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , 
 n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , 
 n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , 
 n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , 
 n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , 
 n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , 
 n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , 
 n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , 
 n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , 
 n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , 
 n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , 
 n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , 
 n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , 
 n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , 
 n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , 
 n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , 
 n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , 
 n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , 
 n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , 
 n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , 
 n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , 
 n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , 
 n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , 
 n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , 
 n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , 
 n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , 
 n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , 
 n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , 
 n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , 
 n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , 
 n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , 
 n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , 
 n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , 
 n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , 
 n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , 
 n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , 
 n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , 
 n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , 
 n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , 
 n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , 
 n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , 
 n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , 
 n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , 
 n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , 
 n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , 
 n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , 
 n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , 
 n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , 
 n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , 
 n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , 
 n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , 
 n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , 
 n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , 
 n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , 
 n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , 
 n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , 
 n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , 
 n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , 
 n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , 
 n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , 
 n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , 
 n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , 
 n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , 
 n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , 
 n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , 
 n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , 
 n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , 
 n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , 
 n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , 
 n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , 
 n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , 
 n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , 
 n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , 
 n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , 
 n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , 
 n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , 
 n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , 
 n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , 
 n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , 
 n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , 
 n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , 
 n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , 
 n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , 
 n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , 
 n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , 
 n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , 
 n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , 
 n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , 
 n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , 
 n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , 
 n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , 
 n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , 
 n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , 
 n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , 
 n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , 
 n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , 
 n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , 
 n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , 
 n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , 
 n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , 
 n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , 
 n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , 
 n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , 
 n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , 
 n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , 
 n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , 
 n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , 
 n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , 
 n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , 
 n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , 
 n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , 
 n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , 
 n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , 
 n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , 
 n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , 
 n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , 
 n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , 
 n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , 
 n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , 
 n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , 
 n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , 
 n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , 
 n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , 
 n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , 
 n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , 
 n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , 
 n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , 
 n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , 
 n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , 
 n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , 
 n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , 
 n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , 
 n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , 
 n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , 
 n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , 
 n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , 
 n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , 
 n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , 
 n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , 
 n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , 
 n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , 
 n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , 
 n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , 
 n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , 
 n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , 
 n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , 
 n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , 
 n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , 
 n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , 
 n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , 
 n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , 
 n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , 
 n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , 
 n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , 
 n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , 
 n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , 
 n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , 
 n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , 
 n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , 
 n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , 
 n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , 
 n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , 
 n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , 
 n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , 
 n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , 
 n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , 
 n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , 
 n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , 
 n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , 
 n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , 
 n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , 
 n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , 
 n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , 
 n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , 
 n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , 
 n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , 
 n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , 
 n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , 
 n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , 
 n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , 
 n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , 
 n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , 
 n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , 
 n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , 
 n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , 
 n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , 
 n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , 
 n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , 
 n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , 
 n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , 
 n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , 
 n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , 
 n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , 
 n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , 
 n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , 
 n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , 
 n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , 
 n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , 
 n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , 
 n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , 
 n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , 
 n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , 
 n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , 
 n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , 
 n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , 
 n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , 
 n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , 
 n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , 
 n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , 
 n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , 
 n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , 
 n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , 
 n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , 
 n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , 
 n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , 
 n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , 
 n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , 
 n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , 
 n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , 
 n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , 
 n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , 
 n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , 
 n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , 
 n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , 
 n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , 
 n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , 
 n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , 
 n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , 
 n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , 
 n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , 
 n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , 
 n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , 
 n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , 
 n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , 
 n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , 
 n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , 
 n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , 
 n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , 
 n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , 
 n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , 
 n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , 
 n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , 
 n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , 
 n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , 
 n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , 
 n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , 
 n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , 
 n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , 
 n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , 
 n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , 
 n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , 
 n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , 
 n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , 
 n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , 
 n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , 
 n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , 
 n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , 
 n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , 
 n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , 
 n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , 
 n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , 
 n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , 
 n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , 
 n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , 
 n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , 
 n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , 
 n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , 
 n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , 
 n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , 
 n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , 
 n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , 
 n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , 
 n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , 
 n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , 
 n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , 
 n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , 
 n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , 
 n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , 
 n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , 
 n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , 
 n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , 
 n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , 
 n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , 
 n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , 
 n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , 
 n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , 
 n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , 
 n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , 
 n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , 
 n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , 
 n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , 
 n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , 
 n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , 
 n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , 
 n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , 
 n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , 
 n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , 
 n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , 
 n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , 
 n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , 
 n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , 
 n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , 
 n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , 
 n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , 
 n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , 
 n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , 
 n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , 
 n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , 
 n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , 
 n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , 
 n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , 
 n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , 
 n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , 
 n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , 
 n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , 
 n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , 
 n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , 
 n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , 
 n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , 
 n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , 
 n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , 
 n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , 
 n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , 
 n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , 
 n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , 
 n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , 
 n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , 
 n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , 
 n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , 
 n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , 
 n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , 
 n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , 
 n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , 
 n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , 
 n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , 
 n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , 
 n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , 
 n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , 
 n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , 
 n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , 
 n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , 
 n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , 
 n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , 
 n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , 
 n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , 
 n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , 
 n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , 
 n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , 
 n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , 
 n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , 
 n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , 
 n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , 
 n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , 
 n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , 
 n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , 
 n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , 
 n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , 
 n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , 
 n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , 
 n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , 
 n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , 
 n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , 
 n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , 
 n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , 
 n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , 
 n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , 
 n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , 
 n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , 
 n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , 
 n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , 
 n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , 
 n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , 
 n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , 
 n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , 
 n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , 
 n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , 
 n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , 
 n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , 
 n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , 
 n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , 
 n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , 
 n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , 
 n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , 
 n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , 
 n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , 
 n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , 
 n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , 
 n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , 
 n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , 
 n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , 
 n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , 
 n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , 
 n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , 
 n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , 
 n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , 
 n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , 
 n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , 
 n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , 
 n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , 
 n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , 
 n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , 
 n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , 
 n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , 
 n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , 
 n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , 
 n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , 
 n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , 
 n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , 
 n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , 
 n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , 
 n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , 
 n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , 
 n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , 
 n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , 
 n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , 
 n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , 
 n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , 
 n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , 
 n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , 
 n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , 
 n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , 
 n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , 
 n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , 
 n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , 
 n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , 
 n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , 
 n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , 
 n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , 
 n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , 
 n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , 
 n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , 
 n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , 
 n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , 
 n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , 
 n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , 
 n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , 
 n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , 
 n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , 
 n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , 
 n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , 
 n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , 
 n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , 
 n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , 
 n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , 
 n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , 
 n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , 
 n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , 
 n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , 
 n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , 
 n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , 
 n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , 
 n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , 
 n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , 
 n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , 
 n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , 
 n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , 
 n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , 
 n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , 
 n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , 
 n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , 
 n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , 
 n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , 
 n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , 
 n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , 
 n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , 
 n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , 
 n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , 
 n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , 
 n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , 
 n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , 
 n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , 
 n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , 
 n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , 
 n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , 
 n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , 
 n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , 
 n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , 
 n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , 
 n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , 
 n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , 
 n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , 
 n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , 
 n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , 
 n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , 
 n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , 
 n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , 
 n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , 
 n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , 
 n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , 
 n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , 
 n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , 
 n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , 
 n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , 
 n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , 
 n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , 
 n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , 
 n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , 
 n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , 
 n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , 
 n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , 
 n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , 
 n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , 
 n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , 
 n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , 
 n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , 
 n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , 
 n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , 
 n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , 
 n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , 
 n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , 
 n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , 
 n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , 
 n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , 
 n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , 
 n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , 
 n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , 
 n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , 
 n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , 
 n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , 
 n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , 
 n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , 
 n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , 
 n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , 
 n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , 
 n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , 
 n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , 
 n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , 
 n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , 
 n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , 
 n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , 
 n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , 
 n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , 
 n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , 
 n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , 
 n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , 
 n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , 
 n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , 
 n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , 
 n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , 
 n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , 
 n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , 
 n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , 
 n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , 
 n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , 
 n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , 
 n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , 
 n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , 
 n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , 
 n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , 
 n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , 
 n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , 
 n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , 
 n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , 
 n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , 
 n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , 
 n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , 
 n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , 
 n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , 
 n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , 
 n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , 
 n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , 
 n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , 
 n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , 
 n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , 
 n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , 
 n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , 
 n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , 
 n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , 
 n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , 
 n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , 
 n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , 
 n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , 
 n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , 
 n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , 
 n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , 
 n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , 
 n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , 
 n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , 
 n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , 
 n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , 
 n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , 
 n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , 
 n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , 
 n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , 
 n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , 
 n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , 
 n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , 
 n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , 
 n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , 
 n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , 
 n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , 
 n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , 
 n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , 
 n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , 
 n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , 
 n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , 
 n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , 
 n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , 
 n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , 
 n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , 
 n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , 
 n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , 
 n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , 
 n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , 
 n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , 
 n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , 
 n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , 
 n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , 
 n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , 
 n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , 
 n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , 
 n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , 
 n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , 
 n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , 
 n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , 
 n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , 
 n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , 
 n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , 
 n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , 
 n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , 
 n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , 
 n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , 
 n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , 
 n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , 
 n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , 
 n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , 
 n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , 
 n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , 
 n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , 
 n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , 
 n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , 
 n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , 
 n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , 
 n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , 
 n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , 
 n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , 
 n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , 
 n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , 
 n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , 
 n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , 
 n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , 
 n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , 
 n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , 
 n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , 
 n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , 
 n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , 
 n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , 
 n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , 
 n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , 
 n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , 
 n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , 
 n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , 
 n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , 
 n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , 
 n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , 
 n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , 
 n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , 
 n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , 
 n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , 
 n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , 
 n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , 
 n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , 
 n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , 
 n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , 
 n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , 
 n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , 
 n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , 
 n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , 
 n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , 
 n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , 
 n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , 
 n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , 
 n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , 
 n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , 
 n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , 
 n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , 
 n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , 
 n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , 
 n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , 
 n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , 
 n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , 
 n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , 
 n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , 
 n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , 
 n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , 
 n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , 
 n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , 
 n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , 
 n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , 
 n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , 
 n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , 
 n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , 
 n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , 
 n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , 
 n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , 
 n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , 
 n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , 
 n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , 
 n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , 
 n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , 
 n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , 
 n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , 
 n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , 
 n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , 
 n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , 
 n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , 
 n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , 
 n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , 
 n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , 
 n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , 
 n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , 
 n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , 
 n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , 
 n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , 
 n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , 
 n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , 
 n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , 
 n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , 
 n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , 
 n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , 
 n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , 
 n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , 
 n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , 
 n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , 
 n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , 
 n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , 
 n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , 
 n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , 
 n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , 
 n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , 
 n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , 
 n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , 
 n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , 
 n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , 
 n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , 
 n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , 
 n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , 
 n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , 
 n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , 
 n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , 
 n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , 
 n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , 
 n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , 
 n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , 
 n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , 
 n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , 
 n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , 
 n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , 
 n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , 
 n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , 
 n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , 
 n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , 
 n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , 
 n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , 
 n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , 
 n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , 
 n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , 
 n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , 
 n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , 
 n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , 
 n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , 
 n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , 
 n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , 
 n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , 
 n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , 
 n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , 
 n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , 
 n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , 
 n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , 
 n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , 
 n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , 
 n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , 
 n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , 
 n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , 
 n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , 
 n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , 
 n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , 
 n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , 
 n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , 
 n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , 
 n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , 
 n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , 
 n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , 
 n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , 
 n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , 
 n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , 
 n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , 
 n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , 
 n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , 
 n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , 
 n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , 
 n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , 
 n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , 
 n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , 
 n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , 
 n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , 
 n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , 
 n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , 
 n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , 
 n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , 
 n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , 
 n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , 
 n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , 
 n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , 
 n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , 
 n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , 
 n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , 
 n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , 
 n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , 
 n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , 
 n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , 
 n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , 
 n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , 
 n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , 
 n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , 
 n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , 
 n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , 
 n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , 
 n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , 
 n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , 
 n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , 
 n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , 
 n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , 
 n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , 
 n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , 
 n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , 
 n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , 
 n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , 
 n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , 
 n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , 
 n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , 
 n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , 
 n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , 
 n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , 
 n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , 
 n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , 
 n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , 
 n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , 
 n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , 
 n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , 
 n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , 
 n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , 
 n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , 
 n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , 
 n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , 
 n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , 
 n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , 
 n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , 
 n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , 
 n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , 
 n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , 
 n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , 
 n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , 
 n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , 
 n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , 
 n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , 
 n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , 
 n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , 
 n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , 
 n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , 
 n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , 
 n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , 
 n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , 
 n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , 
 n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , 
 n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , 
 n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , 
 n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , 
 n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , 
 n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , 
 n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , 
 n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , 
 n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , 
 n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , 
 n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , 
 n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , 
 n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , 
 n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , 
 n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , 
 n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , 
 n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , 
 n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , 
 n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , 
 n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , 
 n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , 
 n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , 
 n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , 
 n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , 
 n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , 
 n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , 
 n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , 
 n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , 
 n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , 
 n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , 
 n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , 
 n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , 
 n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , 
 n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , 
 n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , 
 n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , 
 n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , 
 n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , 
 n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , 
 n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , 
 n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , 
 n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , 
 n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , 
 n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , 
 n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , 
 n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , 
 n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , 
 n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , 
 n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , 
 n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , 
 n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , 
 n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , 
 n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , 
 n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , 
 n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , 
 n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , 
 n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , 
 n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , 
 n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , 
 n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , 
 n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , 
 n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , 
 n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , 
 n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , 
 n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , 
 n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , 
 n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , 
 n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , 
 n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , 
 n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , 
 n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , 
 n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , 
 n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , 
 n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , 
 n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , 
 n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , 
 n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , 
 n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , 
 n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , 
 n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , 
 n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , 
 n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , 
 n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , 
 n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , 
 n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , 
 n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , 
 n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , 
 n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , 
 n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , 
 n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , 
 n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , 
 n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , 
 n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , 
 n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , 
 n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , 
 n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , 
 n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , 
 n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , 
 n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , 
 n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , 
 n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , 
 n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , 
 n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , 
 n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , 
 n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , 
 n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , 
 n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , 
 n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , 
 n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , 
 n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , 
 n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , 
 n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , 
 n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , 
 n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , 
 n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , 
 n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , 
 n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , 
 n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , 
 n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , 
 n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , 
 n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , 
 n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , 
 n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , 
 n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , 
 n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , 
 n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , 
 n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , 
 n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , 
 n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , 
 n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , 
 n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , 
 n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , 
 n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , 
 n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , 
 n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , 
 n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , 
 n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , 
 n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , 
 n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , 
 n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , 
 n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , 
 n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , 
 n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , 
 n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , 
 n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , 
 n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , 
 n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , 
 n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , 
 n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , 
 n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , 
 n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , 
 n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , 
 n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , 
 n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , 
 n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , 
 n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , 
 n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , 
 n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , 
 n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , 
 n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , 
 n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , 
 n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , 
 n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , 
 n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , 
 n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , 
 n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , 
 n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , 
 n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , 
 n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , 
 n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , 
 n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , 
 n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , 
 n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , 
 n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , 
 n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , 
 n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , 
 n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , 
 n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , 
 n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , 
 n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , 
 n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , 
 n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , 
 n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , 
 n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , 
 n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , 
 n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , 
 n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , 
 n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , 
 n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , 
 n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , 
 n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , 
 n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , 
 n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , 
 n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , 
 n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , 
 n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , 
 n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , 
 n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , 
 n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , 
 n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , 
 n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , 
 n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , 
 n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , 
 n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , 
 n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , 
 n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , 
 n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , 
 n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , 
 n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , 
 n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , 
 n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , 
 n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , 
 n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , 
 n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , 
 n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , 
 n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , 
 n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , 
 n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , 
 n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , 
 n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , 
 n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , 
 n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , 
 n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , 
 n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , 
 n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , 
 n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , 
 n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , 
 n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , 
 n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , 
 n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , 
 n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , 
 n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , 
 n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , 
 n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , 
 n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , 
 n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , 
 n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , 
 n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , 
 n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , 
 n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , 
 n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , 
 n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , 
 n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , 
 n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , 
 n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , 
 n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , 
 n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , 
 n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , 
 n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , 
 n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , 
 n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , 
 n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , 
 n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , 
 n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , 
 n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , 
 n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , 
 n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , 
 n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , 
 n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , 
 n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , 
 n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , 
 n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , 
 n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , 
 n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , 
 n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , 
 n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , 
 n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , 
 n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , 
 n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , 
 n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , 
 n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , 
 n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , 
 n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , 
 n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , 
 n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , 
 n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , 
 n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , 
 n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , 
 n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , 
 n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , 
 n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , 
 n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , 
 n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , 
 n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , 
 n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , 
 n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , 
 n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , 
 n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , 
 n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , 
 n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , 
 n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , 
 n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , 
 n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , 
 n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , 
 n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , 
 n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , 
 n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , 
 n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , 
 n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , 
 n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , 
 n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , 
 n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , 
 n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , 
 n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , 
 n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , 
 n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , 
 n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , 
 n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , 
 n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , 
 n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , 
 n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , 
 n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , 
 n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , 
 n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , 
 n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , 
 n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , 
 n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , 
 n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , 
 n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , 
 n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , 
 n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , 
 n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , 
 n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , 
 n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , 
 n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , 
 n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , 
 n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , 
 n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , 
 n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , 
 n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , 
 n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , 
 n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , 
 n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , 
 n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , 
 n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , 
 n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , 
 n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , 
 n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , 
 n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , 
 n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , 
 n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , 
 n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , 
 n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , 
 n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , 
 n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , 
 n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , 
 n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , 
 n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , 
 n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , 
 n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , 
 n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , 
 n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , 
 n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , 
 n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , 
 n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , 
 n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , 
 n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , 
 n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , 
 n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , 
 n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , 
 n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , 
 n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , 
 n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , 
 n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , 
 n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , 
 n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , 
 n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , 
 n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , 
 n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , 
 n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , 
 n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , 
 n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , 
 n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , 
 n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , 
 n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , 
 n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , 
 n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , 
 n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , 
 n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , 
 n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , 
 n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , 
 n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , 
 n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , 
 n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , 
 n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , 
 n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , 
 n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , 
 n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , 
 n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , 
 n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , 
 n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , 
 n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , 
 n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , 
 n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , 
 n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , 
 n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , 
 n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , 
 n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , 
 n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , 
 n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , 
 n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , 
 n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , 
 n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , 
 n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , 
 n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , 
 n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , 
 n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , 
 n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , 
 n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , 
 n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , 
 n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , 
 n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , 
 n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , 
 n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , 
 n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , 
 n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , 
 n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , 
 n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , 
 n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , 
 n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , 
 n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , 
 n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , 
 n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , 
 n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , 
 n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , 
 n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , 
 n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , 
 n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , 
 n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , 
 n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , 
 n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , 
 n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , 
 n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , 
 n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , 
 n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , 
 n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , 
 n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , 
 n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , 
 n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , 
 n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , 
 n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , 
 n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , 
 n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , 
 n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , 
 n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , 
 n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , 
 n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , 
 n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , 
 n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , 
 n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , 
 n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , 
 n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , 
 n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , 
 n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , 
 n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , 
 n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , 
 n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , 
 n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , 
 n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , 
 n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , 
 n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , 
 n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , 
 n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , 
 n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , 
 n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , 
 n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , 
 n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , 
 n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , 
 n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , 
 n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , 
 n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , 
 n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , 
 n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , 
 n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , 
 n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , 
 n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , 
 n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , 
 n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , 
 n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , 
 n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , 
 n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , 
 n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , 
 n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , 
 n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , 
 n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , 
 n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , 
 n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , 
 n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , 
 n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , 
 n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , 
 n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , 
 n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , 
 n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , 
 n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , 
 n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , 
 n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , 
 n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , 
 n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , 
 n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , 
 n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , 
 n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , 
 n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , 
 n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , 
 n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , 
 n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , 
 n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , 
 n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , 
 n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , 
 n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , 
 n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , 
 n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , 
 n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , 
 n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , 
 n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , 
 n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , 
 n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , 
 n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , 
 n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , 
 n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , 
 n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , 
 n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , 
 n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , 
 n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , 
 n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , 
 n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , 
 n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , 
 n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , 
 n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , 
 n50737 , n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , 
 n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , 
 n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , 
 n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , 
 n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , 
 n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , 
 n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , 
 n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , 
 n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , 
 n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , 
 n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , 
 n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , 
 n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , 
 n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , 
 n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , 
 n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , 
 n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , 
 n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , 
 n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , 
 n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , 
 n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , 
 n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , 
 n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , 
 n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , 
 n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , 
 n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , 
 n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , 
 n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , 
 n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , 
 n51027 , n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , 
 n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , 
 n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , 
 n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , 
 n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , 
 n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , 
 n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , 
 n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , 
 n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , 
 n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , 
 n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , 
 n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , 
 n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , 
 n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , 
 n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , 
 n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , 
 n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , 
 n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , 
 n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , 
 n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , 
 n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , 
 n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , 
 n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , 
 n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , 
 n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , 
 n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , 
 n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , 
 n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , 
 n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , 
 n51317 , n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , 
 n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , 
 n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , 
 n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , 
 n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , 
 n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , 
 n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , 
 n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , 
 n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , 
 n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , 
 n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , 
 n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , 
 n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , 
 n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , 
 n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , 
 n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , 
 n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , 
 n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , 
 n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , 
 n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , 
 n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , 
 n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , 
 n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , 
 n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , 
 n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , 
 n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , 
 n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , 
 n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , 
 n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , 
 n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , 
 n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , 
 n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , 
 n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , 
 n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , 
 n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , 
 n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , 
 n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , 
 n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , 
 n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , 
 n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , 
 n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , 
 n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , 
 n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , 
 n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , 
 n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , 
 n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , 
 n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , 
 n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , 
 n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , 
 n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , 
 n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , 
 n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , 
 n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , 
 n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , 
 n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , 
 n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , 
 n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , 
 n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , 
 n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , 
 n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , 
 n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , 
 n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , 
 n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , 
 n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , 
 n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , 
 n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , 
 n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , 
 n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , 
 n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , 
 n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , 
 n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , 
 n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , 
 n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , 
 n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , 
 n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , 
 n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , 
 n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , 
 n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , 
 n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , 
 n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , 
 n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , 
 n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , 
 n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , 
 n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , 
 n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , 
 n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , 
 n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , 
 n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , 
 n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , 
 n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , 
 n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , 
 n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , 
 n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , 
 n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , 
 n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , 
 n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , 
 n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , 
 n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , 
 n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , 
 n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , 
 n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , 
 n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , 
 n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , 
 n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , 
 n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , 
 n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , 
 n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , 
 n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , 
 n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , 
 n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , 
 n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , 
 n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , 
 n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , 
 n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , 
 n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , 
 n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , 
 n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , 
 n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , 
 n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , 
 n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , 
 n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , 
 n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , 
 n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , 
 n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , 
 n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , 
 n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , 
 n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , 
 n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , 
 n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , 
 n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , 
 n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , 
 n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , 
 n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , 
 n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , 
 n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , 
 n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , 
 n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , 
 n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , 
 n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , 
 n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , 
 n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , 
 n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , 
 n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , 
 n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , 
 n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , 
 n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , 
 n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , 
 n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , 
 n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , 
 n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , 
 n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , 
 n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , 
 n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , 
 n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , 
 n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , 
 n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , 
 n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , 
 n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , 
 n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , 
 n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , 
 n52917 , n52918 , n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , 
 n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , 
 n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , 
 n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , 
 n52957 , n52958 , n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , 
 n52967 , n52968 , n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , 
 n52977 , n52978 , n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , 
 n52987 , n52988 , n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , 
 n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , 
 n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , 
 n53017 , n53018 , n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , 
 n53027 , n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , 
 n53037 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , 
 n53047 , n53048 , n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , 
 n53057 , n53058 , n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , 
 n53067 , n53068 , n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , 
 n53077 , n53078 , n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , 
 n53087 , n53088 , n53089 , n53090 , n53091 , n53092 , n53093 , n53094 , n53095 , n53096 , 
 n53097 , n53098 , n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , 
 n53107 , n53108 , n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , 
 n53117 , n53118 , n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , 
 n53127 , n53128 , n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , 
 n53137 , n53138 , n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , 
 n53147 , n53148 , n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , 
 n53157 , n53158 , n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , 
 n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , 
 n53177 , n53178 , n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , 
 n53187 , n53188 , n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , 
 n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , 
 n53207 , n53208 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , 
 n53217 , n53218 , n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , 
 n53227 , n53228 , n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , 
 n53237 , n53238 , n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , 
 n53247 , n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , 
 n53257 , n53258 , n53259 , n53260 , n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , 
 n53267 , n53268 , n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , 
 n53277 , n53278 , n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , 
 n53287 , n53288 , n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , 
 n53297 , n53298 , n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , 
 n53307 , n53308 , n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , 
 n53317 , n53318 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , 
 n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , 
 n53337 , n53338 , n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , 
 n53347 , n53348 , n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , 
 n53357 , n53358 , n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , 
 n53367 , n53368 , n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , 
 n53377 , n53378 , n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , 
 n53387 , n53388 , n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , 
 n53397 , n53398 , n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , 
 n53407 , n53408 , n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , 
 n53417 , n53418 , n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , 
 n53427 , n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , 
 n53437 , n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , 
 n53447 , n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , 
 n53457 , n53458 , n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , 
 n53467 , n53468 , n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , 
 n53477 , n53478 , n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , 
 n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , 
 n53497 , n53498 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , 
 n53507 , n53508 , n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , 
 n53517 , n53518 , n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , 
 n53527 , n53528 , n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , 
 n53537 , n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , 
 n53547 , n53548 , n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , 
 n53557 , n53558 , n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , 
 n53567 , n53568 , n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , 
 n53577 , n53578 , n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , 
 n53587 , n53588 , n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , 
 n53597 , n53598 , n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , 
 n53607 , n53608 , n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , 
 n53617 , n53618 , n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , 
 n53627 , n53628 , n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , 
 n53637 , n53638 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , 
 n53647 , n53648 , n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , 
 n53657 , n53658 , n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , 
 n53667 , n53668 , n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , 
 n53677 , n53678 , n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , 
 n53687 , n53688 , n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , 
 n53697 , n53698 , n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , 
 n53707 , n53708 , n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , 
 n53717 , n53718 , n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , 
 n53727 , n53728 , n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , 
 n53737 , n53738 , n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , 
 n53747 , n53748 , n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , 
 n53757 , n53758 , n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , 
 n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , 
 n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , 
 n53787 , n53788 , n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , 
 n53797 , n53798 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , 
 n53807 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , 
 n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , 
 n53827 , n53828 , n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , 
 n53837 , n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , 
 n53847 , n53848 , n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , 
 n53857 , n53858 , n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , 
 n53867 , n53868 , n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , 
 n53877 , n53878 , n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , 
 n53887 , n53888 , n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , 
 n53897 , n53898 , n53899 , n53900 , n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , 
 n53907 , n53908 , n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , 
 n53917 , n53918 , n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , 
 n53927 , n53928 , n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , 
 n53937 , n53938 , n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , 
 n53947 , n53948 , n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , 
 n53957 , n53958 , n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , 
 n53967 , n53968 , n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , 
 n53977 , n53978 , n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , 
 n53987 , n53988 , n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , 
 n53997 , n53998 , n53999 , n54000 , n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , 
 n54007 , n54008 , n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , 
 n54017 , n54018 , n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , 
 n54027 , n54028 , n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , 
 n54037 , n54038 , n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , 
 n54047 , n54048 , n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , 
 n54057 , n54058 , n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , 
 n54067 , n54068 , n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , 
 n54077 , n54078 , n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , 
 n54087 , n54088 , n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , 
 n54097 , n54098 , n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , 
 n54107 , n54108 , n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , 
 n54117 , n54118 , n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , 
 n54127 , n54128 , n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , 
 n54137 , n54138 , n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , 
 n54147 , n54148 , n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , 
 n54157 , n54158 , n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , 
 n54167 , n54168 , n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , 
 n54177 , n54178 , n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , 
 n54187 , n54188 , n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , 
 n54197 , n54198 , n54199 , n54200 , n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , 
 n54207 , n54208 , n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , 
 n54217 , n54218 , n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , 
 n54227 , n54228 , n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , 
 n54237 , n54238 , n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , 
 n54247 , n54248 , n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , 
 n54257 , n54258 , n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , 
 n54267 , n54268 , n54269 , n54270 , n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , 
 n54277 , n54278 , n54279 , n54280 , n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , 
 n54287 , n54288 , n54289 , n54290 , n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , 
 n54297 , n54298 , n54299 , n54300 , n54301 , n54302 , n54303 , n54304 , n54305 , n54306 , 
 n54307 , n54308 , n54309 , n54310 , n54311 , n54312 , n54313 , n54314 , n54315 , n54316 , 
 n54317 , n54318 , n54319 , n54320 , n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , 
 n54327 , n54328 , n54329 , n54330 , n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , 
 n54337 , n54338 , n54339 , n54340 , n54341 , n54342 , n54343 , n54344 , n54345 , n54346 , 
 n54347 , n54348 , n54349 , n54350 , n54351 , n54352 , n54353 , n54354 , n54355 , n54356 , 
 n54357 , n54358 , n54359 , n54360 , n54361 , n54362 , n54363 , n54364 , n54365 , n54366 , 
 n54367 , n54368 , n54369 , n54370 , n54371 , n54372 , n54373 , n54374 , n54375 , n54376 , 
 n54377 , n54378 , n54379 , n54380 , n54381 , n54382 , n54383 , n54384 , n54385 , n54386 , 
 n54387 , n54388 , n54389 , n54390 , n54391 , n54392 , n54393 , n54394 , n54395 , n54396 , 
 n54397 , n54398 , n54399 , n54400 , n54401 , n54402 , n54403 , n54404 , n54405 , n54406 , 
 n54407 , n54408 , n54409 , n54410 , n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , 
 n54417 , n54418 , n54419 , n54420 , n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , 
 n54427 , n54428 , n54429 , n54430 , n54431 , n54432 , n54433 , n54434 , n54435 , n54436 , 
 n54437 , n54438 , n54439 , n54440 , n54441 , n54442 , n54443 , n54444 , n54445 , n54446 , 
 n54447 , n54448 , n54449 , n54450 , n54451 , n54452 , n54453 , n54454 , n54455 , n54456 , 
 n54457 , n54458 , n54459 , n54460 , n54461 , n54462 , n54463 , n54464 , n54465 , n54466 , 
 n54467 , n54468 , n54469 , n54470 , n54471 , n54472 , n54473 , n54474 , n54475 , n54476 , 
 n54477 , n54478 , n54479 , n54480 , n54481 , n54482 , n54483 , n54484 , n54485 , n54486 , 
 n54487 , n54488 , n54489 , n54490 , n54491 , n54492 , n54493 , n54494 , n54495 , n54496 , 
 n54497 , n54498 , n54499 , n54500 , n54501 , n54502 , n54503 , n54504 , n54505 , n54506 , 
 n54507 , n54508 , n54509 , n54510 , n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , 
 n54517 , n54518 , n54519 , n54520 , n54521 , n54522 , n54523 , n54524 , n54525 , n54526 , 
 n54527 , n54528 , n54529 , n54530 , n54531 , n54532 , n54533 , n54534 , n54535 , n54536 , 
 n54537 , n54538 , n54539 , n54540 , n54541 , n54542 , n54543 , n54544 , n54545 , n54546 , 
 n54547 , n54548 , n54549 , n54550 , n54551 , n54552 , n54553 , n54554 , n54555 , n54556 , 
 n54557 , n54558 , n54559 , n54560 , n54561 , n54562 , n54563 , n54564 , n54565 , n54566 , 
 n54567 , n54568 , n54569 , n54570 , n54571 , n54572 , n54573 , n54574 , n54575 , n54576 , 
 n54577 , n54578 , n54579 , n54580 , n54581 , n54582 , n54583 , n54584 , n54585 , n54586 , 
 n54587 , n54588 , n54589 , n54590 , n54591 , n54592 , n54593 , n54594 , n54595 , n54596 , 
 n54597 , n54598 , n54599 , n54600 , n54601 , n54602 , n54603 , n54604 , n54605 , n54606 , 
 n54607 , n54608 , n54609 , n54610 , n54611 , n54612 , n54613 , n54614 , n54615 , n54616 , 
 n54617 , n54618 , n54619 , n54620 , n54621 , n54622 , n54623 , n54624 , n54625 , n54626 , 
 n54627 , n54628 , n54629 , n54630 , n54631 , n54632 , n54633 , n54634 , n54635 , n54636 , 
 n54637 , n54638 , n54639 , n54640 , n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , 
 n54647 , n54648 , n54649 , n54650 , n54651 , n54652 , n54653 , n54654 , n54655 , n54656 , 
 n54657 , n54658 , n54659 , n54660 , n54661 , n54662 , n54663 , n54664 , n54665 , n54666 , 
 n54667 , n54668 , n54669 , n54670 , n54671 , n54672 , n54673 , n54674 , n54675 , n54676 , 
 n54677 , n54678 , n54679 , n54680 , n54681 , n54682 , n54683 , n54684 , n54685 , n54686 , 
 n54687 , n54688 , n54689 , n54690 , n54691 , n54692 , n54693 , n54694 , n54695 , n54696 , 
 n54697 , n54698 , n54699 , n54700 , n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , 
 n54707 , n54708 , n54709 , n54710 , n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , 
 n54717 , n54718 , n54719 , n54720 , n54721 , n54722 , n54723 , n54724 , n54725 , n54726 , 
 n54727 , n54728 , n54729 , n54730 , n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , 
 n54737 , n54738 , n54739 , n54740 , n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , 
 n54747 , n54748 , n54749 , n54750 , n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , 
 n54757 , n54758 , n54759 , n54760 , n54761 , n54762 , n54763 , n54764 , n54765 , n54766 , 
 n54767 , n54768 , n54769 , n54770 , n54771 , n54772 , n54773 , n54774 , n54775 , n54776 , 
 n54777 , n54778 , n54779 , n54780 , n54781 , n54782 , n54783 , n54784 , n54785 , n54786 , 
 n54787 , n54788 , n54789 , n54790 , n54791 , n54792 , n54793 , n54794 , n54795 , n54796 , 
 n54797 , n54798 , n54799 , n54800 , n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , 
 n54807 , n54808 , n54809 , n54810 , n54811 , n54812 , n54813 , n54814 , n54815 , n54816 , 
 n54817 , n54818 , n54819 , n54820 , n54821 , n54822 , n54823 , n54824 , n54825 , n54826 , 
 n54827 , n54828 , n54829 , n54830 , n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , 
 n54837 , n54838 , n54839 , n54840 , n54841 , n54842 , n54843 , n54844 , n54845 , n54846 , 
 n54847 , n54848 , n54849 , n54850 , n54851 , n54852 , n54853 , n54854 , n54855 , n54856 , 
 n54857 , n54858 , n54859 , n54860 , n54861 , n54862 , n54863 , n54864 , n54865 , n54866 , 
 n54867 , n54868 , n54869 , n54870 , n54871 , n54872 , n54873 , n54874 , n54875 , n54876 , 
 n54877 , n54878 , n54879 , n54880 , n54881 , n54882 , n54883 , n54884 , n54885 , n54886 , 
 n54887 , n54888 , n54889 , n54890 , n54891 , n54892 , n54893 , n54894 , n54895 , n54896 , 
 n54897 , n54898 , n54899 , n54900 , n54901 , n54902 , n54903 , n54904 , n54905 , n54906 , 
 n54907 , n54908 , n54909 , n54910 , n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , 
 n54917 , n54918 , n54919 , n54920 , n54921 , n54922 , n54923 , n54924 , n54925 , n54926 , 
 n54927 , n54928 , n54929 , n54930 , n54931 , n54932 , n54933 , n54934 , n54935 , n54936 , 
 n54937 , n54938 , n54939 , n54940 , n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , 
 n54947 , n54948 , n54949 , n54950 , n54951 , n54952 , n54953 , n54954 , n54955 , n54956 , 
 n54957 , n54958 , n54959 , n54960 , n54961 , n54962 , n54963 , n54964 , n54965 , n54966 , 
 n54967 , n54968 , n54969 , n54970 , n54971 , n54972 , n54973 , n54974 , n54975 , n54976 , 
 n54977 , n54978 , n54979 , n54980 , n54981 , n54982 , n54983 , n54984 , n54985 , n54986 , 
 n54987 , n54988 , n54989 , n54990 , n54991 , n54992 , n54993 , n54994 , n54995 , n54996 , 
 n54997 , n54998 , n54999 , n55000 , n55001 , n55002 , n55003 , n55004 , n55005 , n55006 , 
 n55007 , n55008 , n55009 , n55010 , n55011 , n55012 , n55013 , n55014 , n55015 , n55016 , 
 n55017 , n55018 , n55019 , n55020 , n55021 , n55022 , n55023 , n55024 , n55025 , n55026 , 
 n55027 , n55028 , n55029 , n55030 , n55031 , n55032 , n55033 , n55034 , n55035 , n55036 , 
 n55037 , n55038 , n55039 , n55040 , n55041 , n55042 , n55043 , n55044 , n55045 , n55046 , 
 n55047 , n55048 , n55049 , n55050 , n55051 , n55052 , n55053 , n55054 , n55055 , n55056 , 
 n55057 , n55058 , n55059 , n55060 , n55061 , n55062 , n55063 , n55064 , n55065 , n55066 , 
 n55067 , n55068 , n55069 , n55070 , n55071 , n55072 , n55073 , n55074 , n55075 , n55076 , 
 n55077 , n55078 , n55079 , n55080 , n55081 , n55082 , n55083 , n55084 , n55085 , n55086 , 
 n55087 , n55088 , n55089 , n55090 , n55091 , n55092 , n55093 , n55094 , n55095 , n55096 , 
 n55097 , n55098 , n55099 , n55100 , n55101 , n55102 , n55103 , n55104 , n55105 , n55106 , 
 n55107 , n55108 , n55109 , n55110 , n55111 , n55112 , n55113 , n55114 , n55115 , n55116 , 
 n55117 , n55118 , n55119 , n55120 , n55121 , n55122 , n55123 , n55124 , n55125 , n55126 , 
 n55127 , n55128 , n55129 , n55130 , n55131 , n55132 , n55133 , n55134 , n55135 , n55136 , 
 n55137 , n55138 , n55139 , n55140 , n55141 , n55142 , n55143 , n55144 , n55145 , n55146 , 
 n55147 , n55148 , n55149 , n55150 , n55151 , n55152 , n55153 , n55154 , n55155 , n55156 , 
 n55157 , n55158 , n55159 , n55160 , n55161 , n55162 , n55163 , n55164 , n55165 , n55166 , 
 n55167 , n55168 , n55169 , n55170 , n55171 , n55172 , n55173 , n55174 , n55175 , n55176 , 
 n55177 , n55178 , n55179 , n55180 , n55181 , n55182 , n55183 , n55184 , n55185 , n55186 , 
 n55187 , n55188 , n55189 , n55190 , n55191 , n55192 , n55193 , n55194 , n55195 , n55196 , 
 n55197 , n55198 , n55199 , n55200 , n55201 , n55202 , n55203 , n55204 , n55205 , n55206 , 
 n55207 , n55208 , n55209 , n55210 , n55211 , n55212 , n55213 , n55214 , n55215 , n55216 , 
 n55217 , n55218 , n55219 , n55220 , n55221 , n55222 , n55223 , n55224 , n55225 , n55226 , 
 n55227 , n55228 , n55229 , n55230 , n55231 , n55232 , n55233 , n55234 , n55235 , n55236 , 
 n55237 , n55238 , n55239 , n55240 , n55241 , n55242 , n55243 , n55244 , n55245 , n55246 , 
 n55247 , n55248 , n55249 , n55250 , n55251 , n55252 , n55253 , n55254 , n55255 , n55256 , 
 n55257 , n55258 , n55259 , n55260 , n55261 , n55262 , n55263 , n55264 , n55265 , n55266 , 
 n55267 , n55268 , n55269 , n55270 , n55271 , n55272 , n55273 , n55274 , n55275 , n55276 , 
 n55277 , n55278 , n55279 , n55280 , n55281 , n55282 , n55283 , n55284 , n55285 , n55286 , 
 n55287 , n55288 , n55289 , n55290 , n55291 , n55292 , n55293 , n55294 , n55295 , n55296 , 
 n55297 , n55298 , n55299 , n55300 , n55301 , n55302 , n55303 , n55304 , n55305 , n55306 , 
 n55307 , n55308 , n55309 , n55310 , n55311 , n55312 , n55313 , n55314 , n55315 , n55316 , 
 n55317 , n55318 , n55319 , n55320 , n55321 , n55322 , n55323 , n55324 , n55325 , n55326 , 
 n55327 , n55328 , n55329 , n55330 , n55331 , n55332 , n55333 , n55334 , n55335 , n55336 , 
 n55337 , n55338 , n55339 , n55340 , n55341 , n55342 , n55343 , n55344 , n55345 , n55346 , 
 n55347 , n55348 , n55349 , n55350 , n55351 , n55352 , n55353 , n55354 , n55355 , n55356 , 
 n55357 , n55358 , n55359 , n55360 , n55361 , n55362 , n55363 , n55364 , n55365 , n55366 , 
 n55367 , n55368 , n55369 , n55370 , n55371 , n55372 , n55373 , n55374 , n55375 , n55376 , 
 n55377 , n55378 , n55379 , n55380 , n55381 , n55382 , n55383 , n55384 , n55385 , n55386 , 
 n55387 , n55388 , n55389 , n55390 , n55391 , n55392 , n55393 , n55394 , n55395 , n55396 , 
 n55397 , n55398 , n55399 , n55400 , n55401 , n55402 , n55403 , n55404 , n55405 , n55406 , 
 n55407 , n55408 , n55409 , n55410 , n55411 , n55412 , n55413 , n55414 , n55415 , n55416 , 
 n55417 , n55418 , n55419 , n55420 , n55421 , n55422 , n55423 , n55424 , n55425 , n55426 , 
 n55427 , n55428 , n55429 , n55430 , n55431 , n55432 , n55433 , n55434 , n55435 , n55436 , 
 n55437 , n55438 , n55439 , n55440 , n55441 , n55442 , n55443 , n55444 , n55445 , n55446 , 
 n55447 , n55448 , n55449 , n55450 , n55451 , n55452 , n55453 , n55454 , n55455 , n55456 , 
 n55457 , n55458 , n55459 , n55460 , n55461 , n55462 , n55463 , n55464 , n55465 , n55466 , 
 n55467 , n55468 , n55469 , n55470 , n55471 , n55472 , n55473 , n55474 , n55475 , n55476 , 
 n55477 , n55478 , n55479 , n55480 , n55481 , n55482 , n55483 , n55484 , n55485 , n55486 , 
 n55487 , n55488 , n55489 , n55490 , n55491 , n55492 , n55493 , n55494 , n55495 , n55496 , 
 n55497 , n55498 , n55499 , n55500 , n55501 , n55502 , n55503 , n55504 , n55505 , n55506 , 
 n55507 , n55508 , n55509 , n55510 , n55511 , n55512 , n55513 , n55514 , n55515 , n55516 , 
 n55517 , n55518 , n55519 , n55520 , n55521 , n55522 , n55523 , n55524 , n55525 , n55526 , 
 n55527 , n55528 , n55529 , n55530 , n55531 , n55532 , n55533 , n55534 , n55535 , n55536 , 
 n55537 , n55538 , n55539 , n55540 , n55541 , n55542 , n55543 , n55544 , n55545 , n55546 , 
 n55547 , n55548 , n55549 , n55550 , n55551 , n55552 , n55553 , n55554 , n55555 , n55556 , 
 n55557 , n55558 , n55559 , n55560 , n55561 , n55562 , n55563 , n55564 , n55565 , n55566 , 
 n55567 , n55568 , n55569 , n55570 , n55571 , n55572 , n55573 , n55574 , n55575 , n55576 , 
 n55577 , n55578 , n55579 , n55580 , n55581 , n55582 , n55583 , n55584 , n55585 , n55586 , 
 n55587 , n55588 , n55589 , n55590 , n55591 , n55592 , n55593 , n55594 , n55595 , n55596 , 
 n55597 , n55598 , n55599 , n55600 , n55601 , n55602 , n55603 , n55604 , n55605 , n55606 , 
 n55607 , n55608 , n55609 , n55610 , n55611 , n55612 , n55613 , n55614 , n55615 , n55616 , 
 n55617 , n55618 , n55619 , n55620 , n55621 , n55622 , n55623 , n55624 , n55625 , n55626 , 
 n55627 , n55628 , n55629 , n55630 , n55631 , n55632 , n55633 , n55634 , n55635 , n55636 , 
 n55637 , n55638 , n55639 , n55640 , n55641 , n55642 , n55643 , n55644 , n55645 , n55646 , 
 n55647 , n55648 , n55649 , n55650 , n55651 , n55652 , n55653 , n55654 , n55655 , n55656 , 
 n55657 , n55658 , n55659 , n55660 , n55661 , n55662 , n55663 , n55664 , n55665 , n55666 , 
 n55667 , n55668 , n55669 , n55670 , n55671 , n55672 , n55673 , n55674 , n55675 , n55676 , 
 n55677 , n55678 , n55679 , n55680 , n55681 , n55682 , n55683 , n55684 , n55685 , n55686 , 
 n55687 , n55688 , n55689 , n55690 , n55691 , n55692 , n55693 , n55694 , n55695 , n55696 , 
 n55697 , n55698 , n55699 , n55700 , n55701 , n55702 , n55703 , n55704 , n55705 , n55706 , 
 n55707 , n55708 , n55709 , n55710 , n55711 , n55712 , n55713 , n55714 , n55715 , n55716 , 
 n55717 , n55718 , n55719 , n55720 , n55721 , n55722 , n55723 , n55724 , n55725 , n55726 , 
 n55727 , n55728 , n55729 , n55730 , n55731 , n55732 , n55733 , n55734 , n55735 , n55736 , 
 n55737 , n55738 , n55739 , n55740 , n55741 , n55742 , n55743 , n55744 , n55745 , n55746 , 
 n55747 , n55748 , n55749 , n55750 , n55751 , n55752 , n55753 , n55754 , n55755 , n55756 , 
 n55757 , n55758 , n55759 , n55760 , n55761 , n55762 , n55763 , n55764 , n55765 , n55766 , 
 n55767 , n55768 , n55769 , n55770 , n55771 , n55772 , n55773 , n55774 , n55775 , n55776 , 
 n55777 , n55778 , n55779 , n55780 , n55781 , n55782 , n55783 , n55784 , n55785 , n55786 , 
 n55787 , n55788 , n55789 , n55790 , n55791 , n55792 , n55793 , n55794 , n55795 , n55796 , 
 n55797 , n55798 , n55799 , n55800 , n55801 , n55802 , n55803 , n55804 , n55805 , n55806 , 
 n55807 , n55808 , n55809 , n55810 , n55811 , n55812 , n55813 , n55814 , n55815 , n55816 , 
 n55817 , n55818 , n55819 , n55820 , n55821 , n55822 , n55823 , n55824 , n55825 , n55826 , 
 n55827 , n55828 , n55829 , n55830 , n55831 , n55832 , n55833 , n55834 , n55835 , n55836 , 
 n55837 , n55838 , n55839 , n55840 , n55841 , n55842 , n55843 , n55844 , n55845 , n55846 , 
 n55847 , n55848 , n55849 , n55850 , n55851 , n55852 , n55853 , n55854 , n55855 , n55856 , 
 n55857 , n55858 , n55859 , n55860 , n55861 , n55862 , n55863 , n55864 , n55865 , n55866 , 
 n55867 , n55868 , n55869 , n55870 , n55871 , n55872 , n55873 , n55874 , n55875 , n55876 , 
 n55877 , n55878 , n55879 , n55880 , n55881 , n55882 , n55883 , n55884 , n55885 , n55886 , 
 n55887 , n55888 , n55889 , n55890 , n55891 , n55892 , n55893 , n55894 , n55895 , n55896 , 
 n55897 , n55898 , n55899 , n55900 , n55901 , n55902 , n55903 , n55904 , n55905 , n55906 , 
 n55907 , n55908 , n55909 , n55910 , n55911 , n55912 , n55913 , n55914 , n55915 , n55916 , 
 n55917 , n55918 , n55919 , n55920 , n55921 , n55922 , n55923 , n55924 , n55925 , n55926 , 
 n55927 , n55928 , n55929 , n55930 , n55931 , n55932 , n55933 , n55934 , n55935 , n55936 , 
 n55937 , n55938 , n55939 , n55940 , n55941 , n55942 , n55943 , n55944 , n55945 , n55946 , 
 n55947 , n55948 , n55949 , n55950 , n55951 , n55952 , n55953 , n55954 , n55955 , n55956 , 
 n55957 , n55958 , n55959 , n55960 , n55961 , n55962 , n55963 , n55964 , n55965 , n55966 , 
 n55967 , n55968 , n55969 , n55970 , n55971 , n55972 , n55973 , n55974 , n55975 , n55976 , 
 n55977 , n55978 , n55979 , n55980 , n55981 , n55982 , n55983 , n55984 , n55985 , n55986 , 
 n55987 , n55988 , n55989 , n55990 , n55991 , n55992 , n55993 , n55994 , n55995 , n55996 , 
 n55997 , n55998 , n55999 , n56000 , n56001 , n56002 , n56003 , n56004 , n56005 , n56006 , 
 n56007 , n56008 , n56009 , n56010 , n56011 , n56012 , n56013 , n56014 , n56015 , n56016 , 
 n56017 , n56018 , n56019 , n56020 , n56021 , n56022 , n56023 , n56024 , n56025 , n56026 , 
 n56027 , n56028 , n56029 , n56030 , n56031 , n56032 , n56033 , n56034 , n56035 , n56036 , 
 n56037 , n56038 , n56039 , n56040 , n56041 , n56042 , n56043 , n56044 , n56045 , n56046 , 
 n56047 , n56048 , n56049 , n56050 , n56051 , n56052 , n56053 , n56054 , n56055 , n56056 , 
 n56057 , n56058 , n56059 , n56060 , n56061 , n56062 , n56063 , n56064 , n56065 , n56066 , 
 n56067 , n56068 , n56069 , n56070 , n56071 , n56072 , n56073 , n56074 , n56075 , n56076 , 
 n56077 , n56078 , n56079 , n56080 , n56081 , n56082 , n56083 , n56084 , n56085 , n56086 , 
 n56087 , n56088 , n56089 , n56090 , n56091 , n56092 , n56093 , n56094 , n56095 , n56096 , 
 n56097 , n56098 , n56099 , n56100 , n56101 , n56102 , n56103 , n56104 , n56105 , n56106 , 
 n56107 , n56108 , n56109 , n56110 , n56111 , n56112 , n56113 , n56114 , n56115 , n56116 , 
 n56117 , n56118 , n56119 , n56120 , n56121 , n56122 , n56123 , n56124 , n56125 , n56126 , 
 n56127 , n56128 , n56129 , n56130 , n56131 , n56132 , n56133 , n56134 , n56135 , n56136 , 
 n56137 , n56138 , n56139 , n56140 , n56141 , n56142 , n56143 , n56144 , n56145 , n56146 , 
 n56147 , n56148 , n56149 , n56150 , n56151 , n56152 , n56153 , n56154 , n56155 , n56156 , 
 n56157 , n56158 , n56159 , n56160 , n56161 , n56162 , n56163 , n56164 , n56165 , n56166 , 
 n56167 , n56168 , n56169 , n56170 , n56171 , n56172 , n56173 , n56174 , n56175 , n56176 , 
 n56177 , n56178 , n56179 , n56180 , n56181 , n56182 , n56183 , n56184 , n56185 , n56186 , 
 n56187 , n56188 , n56189 , n56190 , n56191 , n56192 , n56193 , n56194 , n56195 , n56196 , 
 n56197 , n56198 , n56199 , n56200 , n56201 , n56202 , n56203 , n56204 , n56205 , n56206 , 
 n56207 , n56208 , n56209 , n56210 , n56211 , n56212 , n56213 , n56214 , n56215 , n56216 , 
 n56217 , n56218 , n56219 , n56220 , n56221 , n56222 , n56223 , n56224 , n56225 , n56226 , 
 n56227 , n56228 , n56229 , n56230 , n56231 , n56232 , n56233 , n56234 , n56235 , n56236 , 
 n56237 , n56238 , n56239 , n56240 , n56241 , n56242 , n56243 , n56244 , n56245 , n56246 , 
 n56247 , n56248 , n56249 , n56250 , n56251 , n56252 , n56253 , n56254 , n56255 , n56256 , 
 n56257 , n56258 , n56259 , n56260 , n56261 , n56262 , n56263 , n56264 , n56265 , n56266 , 
 n56267 , n56268 , n56269 , n56270 , n56271 , n56272 , n56273 , n56274 , n56275 , n56276 , 
 n56277 , n56278 , n56279 , n56280 , n56281 , n56282 , n56283 , n56284 , n56285 , n56286 , 
 n56287 , n56288 , n56289 , n56290 , n56291 , n56292 , n56293 , n56294 , n56295 , n56296 , 
 n56297 , n56298 , n56299 , n56300 , n56301 , n56302 , n56303 , n56304 , n56305 , n56306 , 
 n56307 , n56308 , n56309 , n56310 , n56311 , n56312 , n56313 , n56314 , n56315 , n56316 , 
 n56317 , n56318 , n56319 , n56320 , n56321 , n56322 , n56323 , n56324 , n56325 , n56326 , 
 n56327 , n56328 , n56329 , n56330 , n56331 , n56332 , n56333 , n56334 , n56335 , n56336 , 
 n56337 , n56338 , n56339 , n56340 , n56341 , n56342 , n56343 , n56344 , n56345 , n56346 , 
 n56347 , n56348 , n56349 , n56350 , n56351 , n56352 , n56353 , n56354 , n56355 , n56356 , 
 n56357 , n56358 , n56359 , n56360 , n56361 , n56362 , n56363 , n56364 , n56365 , n56366 , 
 n56367 , n56368 , n56369 , n56370 , n56371 , n56372 , n56373 , n56374 , n56375 , n56376 , 
 n56377 , n56378 , n56379 , n56380 , n56381 , n56382 , n56383 , n56384 , n56385 , n56386 , 
 n56387 , n56388 , n56389 , n56390 , n56391 , n56392 , n56393 , n56394 , n56395 , n56396 , 
 n56397 , n56398 , n56399 , n56400 , n56401 , n56402 , n56403 , n56404 , n56405 , n56406 , 
 n56407 , n56408 , n56409 , n56410 , n56411 , n56412 , n56413 , n56414 , n56415 , n56416 , 
 n56417 , n56418 , n56419 , n56420 , n56421 , n56422 , n56423 , n56424 , n56425 , n56426 , 
 n56427 , n56428 , n56429 , n56430 , n56431 , n56432 , n56433 , n56434 , n56435 , n56436 , 
 n56437 , n56438 , n56439 , n56440 , n56441 , n56442 , n56443 , n56444 , n56445 , n56446 , 
 n56447 , n56448 , n56449 , n56450 , n56451 , n56452 , n56453 , n56454 , n56455 , n56456 , 
 n56457 , n56458 , n56459 , n56460 , n56461 , n56462 , n56463 , n56464 , n56465 , n56466 , 
 n56467 , n56468 , n56469 , n56470 , n56471 , n56472 , n56473 , n56474 , n56475 , n56476 , 
 n56477 , n56478 , n56479 , n56480 , n56481 , n56482 , n56483 , n56484 , n56485 , n56486 , 
 n56487 , n56488 , n56489 , n56490 , n56491 , n56492 , n56493 , n56494 , n56495 , n56496 , 
 n56497 , n56498 , n56499 , n56500 , n56501 , n56502 , n56503 , n56504 , n56505 , n56506 , 
 n56507 , n56508 , n56509 , n56510 , n56511 , n56512 , n56513 , n56514 , n56515 , n56516 , 
 n56517 , n56518 , n56519 , n56520 , n56521 , n56522 , n56523 , n56524 , n56525 , n56526 , 
 n56527 , n56528 , n56529 , n56530 , n56531 , n56532 , n56533 , n56534 , n56535 , n56536 , 
 n56537 , n56538 , n56539 , n56540 , n56541 , n56542 , n56543 , n56544 , n56545 , n56546 , 
 n56547 , n56548 , n56549 , n56550 , n56551 , n56552 , n56553 , n56554 , n56555 , n56556 , 
 n56557 , n56558 , n56559 , n56560 , n56561 , n56562 , n56563 , n56564 , n56565 , n56566 , 
 n56567 , n56568 , n56569 , n56570 , n56571 , n56572 , n56573 , n56574 , n56575 , n56576 , 
 n56577 , n56578 , n56579 , n56580 , n56581 , n56582 , n56583 , n56584 , n56585 , n56586 , 
 n56587 , n56588 , n56589 , n56590 , n56591 , n56592 , n56593 , n56594 , n56595 , n56596 , 
 n56597 , n56598 , n56599 , n56600 , n56601 , n56602 , n56603 , n56604 , n56605 , n56606 , 
 n56607 , n56608 , n56609 , n56610 , n56611 , n56612 , n56613 , n56614 , n56615 , n56616 , 
 n56617 , n56618 , n56619 , n56620 , n56621 , n56622 , n56623 , n56624 , n56625 , n56626 , 
 n56627 , n56628 , n56629 , n56630 , n56631 , n56632 , n56633 , n56634 , n56635 , n56636 , 
 n56637 , n56638 , n56639 , n56640 , n56641 , n56642 , n56643 , n56644 , n56645 , n56646 , 
 n56647 , n56648 , n56649 , n56650 , n56651 , n56652 , n56653 , n56654 , n56655 , n56656 , 
 n56657 , n56658 , n56659 , n56660 , n56661 , n56662 , n56663 , n56664 , n56665 , n56666 , 
 n56667 , n56668 , n56669 , n56670 , n56671 , n56672 , n56673 , n56674 , n56675 , n56676 , 
 n56677 , n56678 , n56679 , n56680 , n56681 , n56682 , n56683 , n56684 , n56685 , n56686 , 
 n56687 , n56688 , n56689 , n56690 , n56691 , n56692 , n56693 , n56694 , n56695 , n56696 , 
 n56697 , n56698 , n56699 , n56700 , n56701 , n56702 , n56703 , n56704 , n56705 , n56706 , 
 n56707 , n56708 , n56709 , n56710 , n56711 , n56712 , n56713 , n56714 , n56715 , n56716 , 
 n56717 , n56718 , n56719 , n56720 , n56721 , n56722 , n56723 , n56724 , n56725 , n56726 , 
 n56727 , n56728 , n56729 , n56730 , n56731 , n56732 , n56733 , n56734 , n56735 , n56736 , 
 n56737 , n56738 , n56739 , n56740 , n56741 , n56742 , n56743 , n56744 , n56745 , n56746 , 
 n56747 , n56748 , n56749 , n56750 , n56751 , n56752 , n56753 , n56754 , n56755 , n56756 , 
 n56757 , n56758 , n56759 , n56760 , n56761 , n56762 , n56763 , n56764 , n56765 , n56766 , 
 n56767 , n56768 , n56769 , n56770 , n56771 , n56772 , n56773 , n56774 , n56775 , n56776 , 
 n56777 , n56778 , n56779 , n56780 , n56781 , n56782 , n56783 , n56784 , n56785 , n56786 , 
 n56787 , n56788 , n56789 , n56790 , n56791 , n56792 , n56793 , n56794 , n56795 , n56796 , 
 n56797 , n56798 , n56799 , n56800 , n56801 , n56802 , n56803 , n56804 , n56805 , n56806 , 
 n56807 , n56808 , n56809 , n56810 , n56811 , n56812 , n56813 , n56814 , n56815 , n56816 , 
 n56817 , n56818 , n56819 , n56820 , n56821 , n56822 , n56823 , n56824 , n56825 , n56826 , 
 n56827 , n56828 , n56829 , n56830 , n56831 , n56832 , n56833 , n56834 , n56835 , n56836 , 
 n56837 , n56838 , n56839 , n56840 , n56841 , n56842 , n56843 , n56844 , n56845 , n56846 , 
 n56847 , n56848 , n56849 , n56850 , n56851 , n56852 , n56853 , n56854 , n56855 , n56856 , 
 n56857 , n56858 , n56859 , n56860 , n56861 , n56862 , n56863 , n56864 , n56865 , n56866 , 
 n56867 , n56868 , n56869 , n56870 , n56871 , n56872 , n56873 , n56874 , n56875 , n56876 , 
 n56877 , n56878 , n56879 , n56880 , n56881 , n56882 , n56883 , n56884 , n56885 , n56886 , 
 n56887 , n56888 , n56889 , n56890 , n56891 , n56892 , n56893 , n56894 , n56895 , n56896 , 
 n56897 , n56898 , n56899 , n56900 , n56901 , n56902 , n56903 , n56904 , n56905 , n56906 , 
 n56907 , n56908 , n56909 , n56910 , n56911 , n56912 , n56913 , n56914 , n56915 , n56916 , 
 n56917 , n56918 , n56919 , n56920 , n56921 , n56922 , n56923 , n56924 , n56925 , n56926 , 
 n56927 , n56928 , n56929 , n56930 , n56931 , n56932 , n56933 , n56934 , n56935 , n56936 , 
 n56937 , n56938 , n56939 , n56940 , n56941 , n56942 , n56943 , n56944 , n56945 , n56946 , 
 n56947 , n56948 , n56949 , n56950 , n56951 , n56952 , n56953 , n56954 , n56955 , n56956 , 
 n56957 , n56958 , n56959 , n56960 , n56961 , n56962 , n56963 , n56964 , n56965 , n56966 , 
 n56967 , n56968 , n56969 , n56970 , n56971 , n56972 , n56973 , n56974 , n56975 , n56976 , 
 n56977 , n56978 , n56979 , n56980 , n56981 , n56982 , n56983 , n56984 , n56985 , n56986 , 
 n56987 , n56988 , n56989 , n56990 , n56991 , n56992 , n56993 , n56994 , n56995 , n56996 , 
 n56997 , n56998 , n56999 , n57000 , n57001 , n57002 , n57003 , n57004 , n57005 , n57006 , 
 n57007 , n57008 , n57009 , n57010 , n57011 , n57012 , n57013 , n57014 , n57015 , n57016 , 
 n57017 , n57018 , n57019 , n57020 , n57021 , n57022 , n57023 , n57024 , n57025 , n57026 , 
 n57027 , n57028 , n57029 , n57030 , n57031 , n57032 , n57033 , n57034 , n57035 , n57036 , 
 n57037 , n57038 , n57039 , n57040 , n57041 , n57042 , n57043 , n57044 , n57045 , n57046 , 
 n57047 , n57048 , n57049 , n57050 , n57051 , n57052 , n57053 , n57054 , n57055 , n57056 , 
 n57057 , n57058 , n57059 , n57060 , n57061 , n57062 , n57063 , n57064 , n57065 , n57066 , 
 n57067 , n57068 , n57069 , n57070 , n57071 , n57072 , n57073 , n57074 , n57075 , n57076 , 
 n57077 , n57078 , n57079 , n57080 , n57081 , n57082 , n57083 , n57084 , n57085 , n57086 , 
 n57087 , n57088 , n57089 , n57090 , n57091 , n57092 , n57093 , n57094 , n57095 , n57096 , 
 n57097 , n57098 , n57099 , n57100 , n57101 , n57102 , n57103 , n57104 , n57105 , n57106 , 
 n57107 , n57108 , n57109 , n57110 , n57111 , n57112 , n57113 , n57114 , n57115 , n57116 , 
 n57117 , n57118 , n57119 , n57120 , n57121 , n57122 , n57123 , n57124 , n57125 , n57126 , 
 n57127 , n57128 , n57129 , n57130 , n57131 , n57132 , n57133 , n57134 , n57135 , n57136 , 
 n57137 , n57138 , n57139 , n57140 , n57141 , n57142 , n57143 , n57144 , n57145 , n57146 , 
 n57147 , n57148 , n57149 , n57150 , n57151 , n57152 , n57153 , n57154 , n57155 , n57156 , 
 n57157 , n57158 , n57159 , n57160 , n57161 , n57162 , n57163 , n57164 , n57165 , n57166 , 
 n57167 , n57168 , n57169 , n57170 , n57171 , n57172 , n57173 , n57174 , n57175 , n57176 , 
 n57177 , n57178 , n57179 , n57180 , n57181 , n57182 , n57183 , n57184 , n57185 , n57186 , 
 n57187 , n57188 , n57189 , n57190 , n57191 , n57192 , n57193 , n57194 , n57195 , n57196 , 
 n57197 , n57198 , n57199 , n57200 , n57201 , n57202 , n57203 , n57204 , n57205 , n57206 , 
 n57207 , n57208 , n57209 , n57210 , n57211 , n57212 , n57213 , n57214 , n57215 , n57216 , 
 n57217 , n57218 , n57219 , n57220 , n57221 , n57222 , n57223 , n57224 , n57225 , n57226 , 
 n57227 , n57228 , n57229 , n57230 , n57231 , n57232 , n57233 , n57234 , n57235 , n57236 , 
 n57237 , n57238 , n57239 , n57240 , n57241 , n57242 , n57243 , n57244 , n57245 , n57246 , 
 n57247 , n57248 , n57249 , n57250 , n57251 , n57252 , n57253 , n57254 , n57255 , n57256 , 
 n57257 , n57258 , n57259 , n57260 , n57261 , n57262 , n57263 , n57264 , n57265 , n57266 , 
 n57267 , n57268 , n57269 , n57270 , n57271 , n57272 , n57273 , n57274 , n57275 , n57276 , 
 n57277 , n57278 , n57279 , n57280 , n57281 , n57282 , n57283 , n57284 , n57285 , n57286 , 
 n57287 , n57288 , n57289 , n57290 , n57291 , n57292 , n57293 , n57294 , n57295 , n57296 , 
 n57297 , n57298 , n57299 , n57300 , n57301 , n57302 , n57303 , n57304 , n57305 , n57306 , 
 n57307 , n57308 , n57309 , n57310 , n57311 , n57312 , n57313 , n57314 , n57315 , n57316 , 
 n57317 , n57318 , n57319 , n57320 , n57321 , n57322 , n57323 , n57324 , n57325 , n57326 , 
 n57327 , n57328 , n57329 , n57330 , n57331 , n57332 , n57333 , n57334 , n57335 , n57336 , 
 n57337 , n57338 , n57339 , n57340 , n57341 , n57342 , n57343 , n57344 , n57345 , n57346 , 
 n57347 , n57348 , n57349 , n57350 , n57351 , n57352 , n57353 , n57354 , n57355 , n57356 , 
 n57357 , n57358 , n57359 , n57360 , n57361 , n57362 , n57363 , n57364 , n57365 , n57366 , 
 n57367 , n57368 , n57369 , n57370 , n57371 , n57372 , n57373 , n57374 , n57375 , n57376 , 
 n57377 , n57378 , n57379 , n57380 , n57381 , n57382 , n57383 , n57384 , n57385 , n57386 , 
 n57387 , n57388 , n57389 , n57390 , n57391 , n57392 , n57393 , n57394 , n57395 , n57396 , 
 n57397 , n57398 , n57399 , n57400 , n57401 , n57402 , n57403 , n57404 , n57405 , n57406 , 
 n57407 , n57408 , n57409 , n57410 , n57411 , n57412 , n57413 , n57414 , n57415 , n57416 , 
 n57417 , n57418 , n57419 , n57420 , n57421 , n57422 , n57423 , n57424 , n57425 , n57426 , 
 n57427 , n57428 , n57429 , n57430 , n57431 , n57432 , n57433 , n57434 , n57435 , n57436 , 
 n57437 , n57438 , n57439 , n57440 , n57441 , n57442 , n57443 , n57444 , n57445 , n57446 , 
 n57447 , n57448 , n57449 , n57450 , n57451 , n57452 , n57453 , n57454 , n57455 , n57456 , 
 n57457 , n57458 , n57459 , n57460 , n57461 , n57462 , n57463 , n57464 , n57465 , n57466 , 
 n57467 , n57468 , n57469 , n57470 , n57471 , n57472 , n57473 , n57474 , n57475 , n57476 , 
 n57477 , n57478 , n57479 , n57480 , n57481 , n57482 , n57483 , n57484 , n57485 , n57486 , 
 n57487 , n57488 , n57489 , n57490 , n57491 , n57492 , n57493 , n57494 , n57495 , n57496 , 
 n57497 , n57498 , n57499 , n57500 , n57501 , n57502 , n57503 , n57504 , n57505 , n57506 , 
 n57507 , n57508 , n57509 , n57510 , n57511 , n57512 , n57513 , n57514 , n57515 , n57516 , 
 n57517 , n57518 , n57519 , n57520 , n57521 , n57522 , n57523 , n57524 , n57525 , n57526 , 
 n57527 , n57528 , n57529 , n57530 , n57531 , n57532 , n57533 , n57534 , n57535 , n57536 , 
 n57537 , n57538 , n57539 , n57540 , n57541 , n57542 , n57543 , n57544 , n57545 , n57546 , 
 n57547 , n57548 , n57549 , n57550 , n57551 , n57552 , n57553 , n57554 , n57555 , n57556 , 
 n57557 , n57558 , n57559 , n57560 , n57561 , n57562 , n57563 , n57564 , n57565 , n57566 , 
 n57567 , n57568 , n57569 , n57570 , n57571 , n57572 , n57573 , n57574 , n57575 , n57576 , 
 n57577 , n57578 , n57579 , n57580 , n57581 , n57582 , n57583 , n57584 , n57585 , n57586 , 
 n57587 , n57588 , n57589 , n57590 , n57591 , n57592 , n57593 , n57594 , n57595 , n57596 , 
 n57597 , n57598 , n57599 , n57600 , n57601 , n57602 , n57603 , n57604 , n57605 , n57606 , 
 n57607 , n57608 , n57609 , n57610 , n57611 , n57612 , n57613 , n57614 , n57615 , n57616 , 
 n57617 , n57618 , n57619 , n57620 , n57621 , n57622 , n57623 , n57624 , n57625 , n57626 , 
 n57627 , n57628 , n57629 , n57630 , n57631 , n57632 , n57633 , n57634 , n57635 , n57636 , 
 n57637 , n57638 , n57639 , n57640 , n57641 , n57642 , n57643 , n57644 , n57645 , n57646 , 
 n57647 , n57648 , n57649 , n57650 , n57651 , n57652 , n57653 , n57654 , n57655 , n57656 , 
 n57657 , n57658 , n57659 , n57660 , n57661 , n57662 , n57663 , n57664 , n57665 , n57666 , 
 n57667 , n57668 , n57669 , n57670 , n57671 , n57672 , n57673 , n57674 , n57675 , n57676 , 
 n57677 , n57678 , n57679 , n57680 , n57681 , n57682 , n57683 , n57684 , n57685 , n57686 , 
 n57687 , n57688 , n57689 , n57690 , n57691 , n57692 , n57693 , n57694 , n57695 , n57696 , 
 n57697 , n57698 , n57699 , n57700 , n57701 , n57702 , n57703 , n57704 , n57705 , n57706 , 
 n57707 , n57708 , n57709 , n57710 , n57711 , n57712 , n57713 , n57714 , n57715 , n57716 , 
 n57717 , n57718 , n57719 , n57720 , n57721 , n57722 , n57723 , n57724 , n57725 , n57726 , 
 n57727 , n57728 , n57729 , n57730 , n57731 , n57732 , n57733 , n57734 , n57735 , n57736 , 
 n57737 , n57738 , n57739 , n57740 , n57741 , n57742 , n57743 , n57744 , n57745 , n57746 , 
 n57747 , n57748 , n57749 , n57750 , n57751 , n57752 , n57753 , n57754 , n57755 , n57756 , 
 n57757 , n57758 , n57759 , n57760 , n57761 , n57762 , n57763 , n57764 , n57765 , n57766 , 
 n57767 , n57768 , n57769 , n57770 , n57771 , n57772 , n57773 , n57774 , n57775 , n57776 , 
 n57777 , n57778 , n57779 , n57780 , n57781 , n57782 , n57783 , n57784 , n57785 , n57786 , 
 n57787 , n57788 , n57789 , n57790 , n57791 , n57792 , n57793 , n57794 , n57795 , n57796 , 
 n57797 , n57798 , n57799 , n57800 , n57801 , n57802 , n57803 , n57804 , n57805 , n57806 , 
 n57807 , n57808 , n57809 , n57810 , n57811 , n57812 , n57813 , n57814 , n57815 , n57816 , 
 n57817 , n57818 , n57819 , n57820 , n57821 , n57822 , n57823 , n57824 , n57825 , n57826 , 
 n57827 , n57828 , n57829 , n57830 , n57831 , n57832 , n57833 , n57834 , n57835 , n57836 , 
 n57837 , n57838 , n57839 , n57840 , n57841 , n57842 , n57843 , n57844 , n57845 , n57846 , 
 n57847 , n57848 , n57849 , n57850 , n57851 , n57852 , n57853 , n57854 , n57855 , n57856 , 
 n57857 , n57858 , n57859 , n57860 , n57861 , n57862 , n57863 , n57864 , n57865 , n57866 , 
 n57867 , n57868 , n57869 , n57870 , n57871 , n57872 , n57873 , n57874 , n57875 , n57876 , 
 n57877 , n57878 , n57879 , n57880 , n57881 , n57882 , n57883 , n57884 , n57885 , n57886 , 
 n57887 , n57888 , n57889 , n57890 , n57891 , n57892 , n57893 , n57894 , n57895 , n57896 , 
 n57897 , n57898 , n57899 , n57900 , n57901 , n57902 , n57903 , n57904 , n57905 , n57906 , 
 n57907 , n57908 , n57909 , n57910 , n57911 , n57912 , n57913 , n57914 , n57915 , n57916 , 
 n57917 , n57918 , n57919 , n57920 , n57921 , n57922 , n57923 , n57924 , n57925 , n57926 , 
 n57927 , n57928 , n57929 , n57930 , n57931 , n57932 , n57933 , n57934 , n57935 , n57936 , 
 n57937 , n57938 , n57939 , n57940 , n57941 , n57942 , n57943 , n57944 , n57945 , n57946 , 
 n57947 , n57948 , n57949 , n57950 , n57951 , n57952 , n57953 , n57954 , n57955 , n57956 , 
 n57957 , n57958 , n57959 , n57960 , n57961 , n57962 , n57963 , n57964 , n57965 , n57966 , 
 n57967 , n57968 , n57969 , n57970 , n57971 , n57972 , n57973 , n57974 , n57975 , n57976 , 
 n57977 , n57978 , n57979 , n57980 , n57981 , n57982 , n57983 , n57984 , n57985 , n57986 , 
 n57987 , n57988 , n57989 , n57990 , n57991 , n57992 , n57993 , n57994 , n57995 , n57996 , 
 n57997 , n57998 , n57999 , n58000 , n58001 , n58002 , n58003 , n58004 , n58005 , n58006 , 
 n58007 , n58008 , n58009 , n58010 , n58011 , n58012 , n58013 , n58014 , n58015 , n58016 , 
 n58017 , n58018 , n58019 , n58020 , n58021 , n58022 , n58023 , n58024 , n58025 , n58026 , 
 n58027 , n58028 , n58029 , n58030 , n58031 , n58032 , n58033 , n58034 , n58035 , n58036 , 
 n58037 , n58038 , n58039 , n58040 , n58041 , n58042 , n58043 , n58044 , n58045 , n58046 , 
 n58047 , n58048 , n58049 , n58050 , n58051 , n58052 , n58053 , n58054 , n58055 , n58056 , 
 n58057 , n58058 , n58059 , n58060 , n58061 , n58062 , n58063 , n58064 , n58065 , n58066 , 
 n58067 , n58068 , n58069 , n58070 , n58071 , n58072 , n58073 , n58074 , n58075 , n58076 , 
 n58077 , n58078 , n58079 , n58080 , n58081 , n58082 , n58083 , n58084 , n58085 , n58086 , 
 n58087 , n58088 , n58089 , n58090 , n58091 , n58092 , n58093 , n58094 , n58095 , n58096 , 
 n58097 , n58098 , n58099 , n58100 , n58101 , n58102 , n58103 , n58104 , n58105 , n58106 , 
 n58107 , n58108 , n58109 , n58110 , n58111 , n58112 , n58113 , n58114 , n58115 , n58116 , 
 n58117 , n58118 , n58119 , n58120 , n58121 , n58122 , n58123 , n58124 , n58125 , n58126 , 
 n58127 , n58128 , n58129 , n58130 , n58131 , n58132 , n58133 , n58134 , n58135 , n58136 , 
 n58137 , n58138 , n58139 , n58140 , n58141 , n58142 , n58143 , n58144 , n58145 , n58146 , 
 n58147 , n58148 , n58149 , n58150 , n58151 , n58152 , n58153 , n58154 , n58155 , n58156 , 
 n58157 , n58158 , n58159 , n58160 , n58161 , n58162 , n58163 , n58164 , n58165 , n58166 , 
 n58167 , n58168 , n58169 , n58170 , n58171 , n58172 , n58173 , n58174 , n58175 , n58176 , 
 n58177 , n58178 , n58179 , n58180 , n58181 , n58182 , n58183 , n58184 , n58185 , n58186 , 
 n58187 , n58188 , n58189 , n58190 , n58191 , n58192 , n58193 , n58194 , n58195 , n58196 , 
 n58197 , n58198 , n58199 , n58200 , n58201 , n58202 , n58203 , n58204 , n58205 , n58206 , 
 n58207 , n58208 , n58209 , n58210 , n58211 , n58212 , n58213 , n58214 , n58215 , n58216 , 
 n58217 , n58218 , n58219 , n58220 , n58221 , n58222 , n58223 , n58224 , n58225 , n58226 , 
 n58227 , n58228 , n58229 , n58230 , n58231 , n58232 , n58233 , n58234 , n58235 , n58236 , 
 n58237 , n58238 , n58239 , n58240 , n58241 , n58242 , n58243 , n58244 , n58245 , n58246 , 
 n58247 , n58248 , n58249 , n58250 , n58251 , n58252 , n58253 , n58254 , n58255 , n58256 , 
 n58257 , n58258 , n58259 , n58260 , n58261 , n58262 , n58263 , n58264 , n58265 , n58266 , 
 n58267 , n58268 , n58269 , n58270 , n58271 , n58272 , n58273 , n58274 , n58275 , n58276 , 
 n58277 , n58278 , n58279 , n58280 , n58281 , n58282 , n58283 , n58284 , n58285 , n58286 , 
 n58287 , n58288 , n58289 , n58290 , n58291 , n58292 , n58293 , n58294 , n58295 , n58296 , 
 n58297 , n58298 , n58299 , n58300 , n58301 , n58302 , n58303 , n58304 , n58305 , n58306 , 
 n58307 , n58308 , n58309 , n58310 , n58311 , n58312 , n58313 , n58314 , n58315 , n58316 , 
 n58317 , n58318 , n58319 , n58320 , n58321 , n58322 , n58323 , n58324 , n58325 , n58326 , 
 n58327 , n58328 , n58329 , n58330 , n58331 , n58332 , n58333 , n58334 , n58335 , n58336 , 
 n58337 , n58338 , n58339 , n58340 , n58341 , n58342 , n58343 , n58344 , n58345 , n58346 , 
 n58347 , n58348 , n58349 , n58350 , n58351 , n58352 , n58353 , n58354 , n58355 , n58356 , 
 n58357 , n58358 , n58359 , n58360 , n58361 , n58362 , n58363 , n58364 , n58365 , n58366 , 
 n58367 , n58368 , n58369 , n58370 , n58371 , n58372 , n58373 , n58374 , n58375 , n58376 , 
 n58377 , n58378 , n58379 , n58380 , n58381 , n58382 , n58383 , n58384 , n58385 , n58386 , 
 n58387 , n58388 , n58389 , n58390 , n58391 , n58392 , n58393 , n58394 , n58395 , n58396 , 
 n58397 , n58398 , n58399 , n58400 , n58401 , n58402 , n58403 , n58404 , n58405 , n58406 , 
 n58407 , n58408 , n58409 , n58410 , n58411 , n58412 , n58413 , n58414 , n58415 , n58416 , 
 n58417 , n58418 , n58419 , n58420 , n58421 , n58422 , n58423 , n58424 , n58425 , n58426 , 
 n58427 , n58428 , n58429 , n58430 , n58431 , n58432 , n58433 , n58434 , n58435 , n58436 , 
 n58437 , n58438 , n58439 , n58440 , n58441 , n58442 , n58443 , n58444 , n58445 , n58446 , 
 n58447 , n58448 , n58449 , n58450 , n58451 , n58452 , n58453 , n58454 , n58455 , n58456 , 
 n58457 , n58458 , n58459 , n58460 , n58461 , n58462 , n58463 , n58464 , n58465 , n58466 , 
 n58467 , n58468 , n58469 , n58470 , n58471 , n58472 , n58473 , n58474 , n58475 , n58476 , 
 n58477 , n58478 , n58479 , n58480 , n58481 , n58482 , n58483 , n58484 , n58485 , n58486 , 
 n58487 , n58488 , n58489 , n58490 , n58491 , n58492 , n58493 , n58494 , n58495 , n58496 , 
 n58497 , n58498 , n58499 , n58500 , n58501 , n58502 , n58503 , n58504 , n58505 , n58506 , 
 n58507 , n58508 , n58509 , n58510 , n58511 , n58512 , n58513 , n58514 , n58515 , n58516 , 
 n58517 , n58518 , n58519 , n58520 , n58521 , n58522 , n58523 , n58524 , n58525 , n58526 , 
 n58527 , n58528 , n58529 , n58530 , n58531 , n58532 , n58533 , n58534 , n58535 , n58536 , 
 n58537 , n58538 , n58539 , n58540 , n58541 , n58542 , n58543 , n58544 , n58545 , n58546 , 
 n58547 , n58548 , n58549 , n58550 , n58551 , n58552 , n58553 , n58554 , n58555 , n58556 , 
 n58557 , n58558 , n58559 , n58560 , n58561 , n58562 , n58563 , n58564 , n58565 , n58566 , 
 n58567 , n58568 , n58569 , n58570 , n58571 , n58572 , n58573 , n58574 , n58575 , n58576 , 
 n58577 , n58578 , n58579 , n58580 , n58581 , n58582 , n58583 , n58584 , n58585 , n58586 , 
 n58587 , n58588 , n58589 , n58590 , n58591 , n58592 , n58593 , n58594 , n58595 , n58596 , 
 n58597 , n58598 , n58599 , n58600 , n58601 , n58602 , n58603 , n58604 , n58605 , n58606 , 
 n58607 , n58608 , n58609 , n58610 , n58611 , n58612 , n58613 , n58614 , n58615 , n58616 , 
 n58617 , n58618 , n58619 , n58620 , n58621 , n58622 , n58623 , n58624 , n58625 , n58626 , 
 n58627 , n58628 , n58629 , n58630 , n58631 , n58632 , n58633 , n58634 , n58635 , n58636 , 
 n58637 , n58638 , n58639 , n58640 , n58641 , n58642 , n58643 , n58644 , n58645 , n58646 , 
 n58647 , n58648 , n58649 , n58650 , n58651 , n58652 , n58653 , n58654 , n58655 , n58656 , 
 n58657 , n58658 , n58659 , n58660 , n58661 , n58662 , n58663 , n58664 , n58665 , n58666 , 
 n58667 , n58668 , n58669 , n58670 , n58671 , n58672 , n58673 , n58674 , n58675 , n58676 , 
 n58677 , n58678 , n58679 , n58680 , n58681 , n58682 , n58683 , n58684 , n58685 , n58686 , 
 n58687 , n58688 , n58689 , n58690 , n58691 , n58692 , n58693 , n58694 , n58695 , n58696 , 
 n58697 , n58698 , n58699 , n58700 , n58701 , n58702 , n58703 , n58704 , n58705 , n58706 , 
 n58707 , n58708 , n58709 , n58710 , n58711 , n58712 , n58713 , n58714 , n58715 , n58716 , 
 n58717 , n58718 , n58719 , n58720 , n58721 , n58722 , n58723 , n58724 , n58725 , n58726 , 
 n58727 , n58728 , n58729 , n58730 , n58731 , n58732 , n58733 , n58734 , n58735 , n58736 , 
 n58737 , n58738 , n58739 , n58740 , n58741 , n58742 , n58743 , n58744 , n58745 , n58746 , 
 n58747 , n58748 , n58749 , n58750 , n58751 , n58752 , n58753 , n58754 , n58755 , n58756 , 
 n58757 , n58758 , n58759 , n58760 , n58761 , n58762 , n58763 , n58764 , n58765 , n58766 , 
 n58767 , n58768 , n58769 , n58770 , n58771 , n58772 , n58773 , n58774 , n58775 , n58776 , 
 n58777 , n58778 , n58779 , n58780 , n58781 , n58782 , n58783 , n58784 , n58785 , n58786 , 
 n58787 , n58788 , n58789 , n58790 , n58791 , n58792 , n58793 , n58794 , n58795 , n58796 , 
 n58797 , n58798 , n58799 , n58800 , n58801 , n58802 , n58803 , n58804 , n58805 , n58806 , 
 n58807 , n58808 , n58809 , n58810 , n58811 , n58812 , n58813 , n58814 , n58815 , n58816 , 
 n58817 , n58818 , n58819 , n58820 , n58821 , n58822 , n58823 , n58824 , n58825 , n58826 , 
 n58827 , n58828 , n58829 , n58830 , n58831 , n58832 , n58833 , n58834 , n58835 , n58836 , 
 n58837 , n58838 , n58839 , n58840 , n58841 , n58842 , n58843 , n58844 , n58845 , n58846 , 
 n58847 , n58848 , n58849 , n58850 , n58851 , n58852 , n58853 , n58854 , n58855 , n58856 , 
 n58857 , n58858 , n58859 , n58860 , n58861 , n58862 , n58863 , n58864 , n58865 , n58866 , 
 n58867 , n58868 , n58869 , n58870 , n58871 , n58872 , n58873 , n58874 , n58875 , n58876 , 
 n58877 , n58878 , n58879 , n58880 , n58881 , n58882 , n58883 , n58884 , n58885 , n58886 , 
 n58887 , n58888 , n58889 , n58890 , n58891 , n58892 , n58893 , n58894 , n58895 , n58896 , 
 n58897 , n58898 , n58899 , n58900 , n58901 , n58902 , n58903 , n58904 , n58905 , n58906 , 
 n58907 , n58908 , n58909 , n58910 , n58911 , n58912 , n58913 , n58914 , n58915 , n58916 , 
 n58917 , n58918 , n58919 , n58920 , n58921 , n58922 , n58923 , n58924 , n58925 , n58926 , 
 n58927 , n58928 , n58929 , n58930 , n58931 , n58932 , n58933 , n58934 , n58935 , n58936 , 
 n58937 , n58938 , n58939 , n58940 , n58941 , n58942 , n58943 , n58944 , n58945 , n58946 , 
 n58947 , n58948 , n58949 , n58950 , n58951 , n58952 , n58953 , n58954 , n58955 , n58956 , 
 n58957 , n58958 , n58959 , n58960 , n58961 , n58962 , n58963 , n58964 , n58965 , n58966 , 
 n58967 , n58968 , n58969 , n58970 , n58971 , n58972 , n58973 , n58974 , n58975 , n58976 , 
 n58977 , n58978 , n58979 , n58980 , n58981 , n58982 , n58983 , n58984 , n58985 , n58986 , 
 n58987 , n58988 , n58989 , n58990 , n58991 , n58992 , n58993 , n58994 , n58995 , n58996 , 
 n58997 , n58998 , n58999 , n59000 , n59001 , n59002 , n59003 , n59004 , n59005 , n59006 , 
 n59007 , n59008 , n59009 , n59010 , n59011 , n59012 , n59013 , n59014 , n59015 , n59016 , 
 n59017 , n59018 , n59019 , n59020 , n59021 , n59022 , n59023 , n59024 , n59025 , n59026 , 
 n59027 , n59028 , n59029 , n59030 , n59031 , n59032 , n59033 , n59034 , n59035 , n59036 , 
 n59037 , n59038 , n59039 , n59040 , n59041 , n59042 , n59043 , n59044 , n59045 , n59046 , 
 n59047 , n59048 , n59049 , n59050 , n59051 , n59052 , n59053 , n59054 , n59055 , n59056 , 
 n59057 , n59058 , n59059 , n59060 , n59061 , n59062 , n59063 , n59064 , n59065 , n59066 , 
 n59067 , n59068 , n59069 , n59070 , n59071 , n59072 , n59073 , n59074 , n59075 , n59076 , 
 n59077 , n59078 , n59079 , n59080 , n59081 , n59082 , n59083 , n59084 , n59085 , n59086 , 
 n59087 , n59088 , n59089 , n59090 , n59091 , n59092 , n59093 , n59094 , n59095 , n59096 , 
 n59097 , n59098 , n59099 , n59100 , n59101 , n59102 , n59103 , n59104 , n59105 , n59106 , 
 n59107 , n59108 , n59109 , n59110 , n59111 , n59112 , n59113 , n59114 , n59115 , n59116 , 
 n59117 , n59118 , n59119 , n59120 , n59121 , n59122 , n59123 , n59124 , n59125 , n59126 , 
 n59127 , n59128 , n59129 , n59130 , n59131 , n59132 , n59133 , n59134 , n59135 , n59136 , 
 n59137 , n59138 , n59139 , n59140 , n59141 , n59142 , n59143 , n59144 , n59145 , n59146 , 
 n59147 , n59148 , n59149 , n59150 , n59151 , n59152 , n59153 , n59154 , n59155 , n59156 , 
 n59157 , n59158 , n59159 , n59160 , n59161 , n59162 , n59163 , n59164 , n59165 , n59166 , 
 n59167 , n59168 , n59169 , n59170 , n59171 , n59172 , n59173 , n59174 , n59175 , n59176 , 
 n59177 , n59178 , n59179 , n59180 , n59181 , n59182 , n59183 , n59184 , n59185 , n59186 , 
 n59187 , n59188 , n59189 , n59190 , n59191 , n59192 , n59193 , n59194 , n59195 , n59196 , 
 n59197 , n59198 , n59199 , n59200 , n59201 , n59202 , n59203 , n59204 , n59205 , n59206 , 
 n59207 , n59208 , n59209 , n59210 , n59211 , n59212 , n59213 , n59214 , n59215 , n59216 , 
 n59217 , n59218 , n59219 , n59220 , n59221 , n59222 , n59223 , n59224 , n59225 , n59226 , 
 n59227 , n59228 , n59229 , n59230 , n59231 , n59232 , n59233 , n59234 , n59235 , n59236 , 
 n59237 , n59238 , n59239 , n59240 , n59241 , n59242 , n59243 , n59244 , n59245 , n59246 , 
 n59247 , n59248 , n59249 , n59250 , n59251 , n59252 , n59253 , n59254 , n59255 , n59256 , 
 n59257 , n59258 , n59259 , n59260 , n59261 , n59262 , n59263 , n59264 , n59265 , n59266 , 
 n59267 , n59268 , n59269 , n59270 , n59271 , n59272 , n59273 , n59274 , n59275 , n59276 , 
 n59277 , n59278 , n59279 , n59280 , n59281 , n59282 , n59283 , n59284 , n59285 , n59286 , 
 n59287 , n59288 , n59289 , n59290 , n59291 , n59292 , n59293 , n59294 , n59295 , n59296 , 
 n59297 , n59298 , n59299 , n59300 , n59301 , n59302 , n59303 , n59304 , n59305 , n59306 , 
 n59307 , n59308 , n59309 , n59310 , n59311 , n59312 , n59313 , n59314 , n59315 , n59316 , 
 n59317 , n59318 , n59319 , n59320 , n59321 , n59322 , n59323 , n59324 , n59325 , n59326 , 
 n59327 , n59328 , n59329 , n59330 , n59331 , n59332 , n59333 , n59334 , n59335 , n59336 , 
 n59337 , n59338 , n59339 , n59340 , n59341 , n59342 , n59343 , n59344 , n59345 , n59346 , 
 n59347 , n59348 , n59349 , n59350 , n59351 , n59352 , n59353 , n59354 , n59355 , n59356 , 
 n59357 , n59358 , n59359 , n59360 , n59361 , n59362 , n59363 , n59364 , n59365 , n59366 , 
 n59367 , n59368 , n59369 , n59370 , n59371 , n59372 , n59373 , n59374 , n59375 , n59376 , 
 n59377 , n59378 , n59379 , n59380 , n59381 , n59382 , n59383 , n59384 , n59385 , n59386 , 
 n59387 , n59388 , n59389 , n59390 , n59391 , n59392 , n59393 , n59394 , n59395 , n59396 , 
 n59397 , n59398 , n59399 , n59400 , n59401 , n59402 , n59403 , n59404 , n59405 , n59406 , 
 n59407 , n59408 , n59409 , n59410 , n59411 , n59412 , n59413 , n59414 , n59415 , n59416 , 
 n59417 , n59418 , n59419 , n59420 , n59421 , n59422 , n59423 , n59424 , n59425 , n59426 , 
 n59427 , n59428 , n59429 , n59430 , n59431 , n59432 , n59433 , n59434 , n59435 , n59436 , 
 n59437 , n59438 , n59439 , n59440 , n59441 , n59442 , n59443 , n59444 , n59445 , n59446 , 
 n59447 , n59448 , n59449 , n59450 , n59451 , n59452 , n59453 , n59454 , n59455 , n59456 , 
 n59457 , n59458 , n59459 , n59460 , n59461 , n59462 , n59463 , n59464 , n59465 , n59466 , 
 n59467 , n59468 , n59469 , n59470 , n59471 , n59472 , n59473 , n59474 , n59475 , n59476 , 
 n59477 , n59478 , n59479 , n59480 , n59481 , n59482 , n59483 , n59484 , n59485 , n59486 , 
 n59487 , n59488 , n59489 , n59490 , n59491 , n59492 , n59493 , n59494 , n59495 , n59496 , 
 n59497 , n59498 , n59499 , n59500 , n59501 , n59502 , n59503 , n59504 , n59505 , n59506 , 
 n59507 , n59508 , n59509 , n59510 , n59511 , n59512 , n59513 , n59514 , n59515 , n59516 , 
 n59517 , n59518 , n59519 , n59520 , n59521 , n59522 , n59523 , n59524 , n59525 , n59526 , 
 n59527 , n59528 , n59529 , n59530 , n59531 , n59532 , n59533 , n59534 , n59535 , n59536 , 
 n59537 , n59538 , n59539 , n59540 , n59541 , n59542 , n59543 , n59544 , n59545 , n59546 , 
 n59547 , n59548 , n59549 , n59550 , n59551 , n59552 , n59553 , n59554 , n59555 , n59556 , 
 n59557 , n59558 , n59559 , n59560 , n59561 , n59562 , n59563 , n59564 , n59565 , n59566 , 
 n59567 , n59568 , n59569 , n59570 , n59571 , n59572 , n59573 , n59574 , n59575 , n59576 , 
 n59577 , n59578 , n59579 , n59580 , n59581 , n59582 , n59583 , n59584 , n59585 , n59586 , 
 n59587 , n59588 , n59589 , n59590 , n59591 , n59592 , n59593 , n59594 , n59595 , n59596 , 
 n59597 , n59598 , n59599 , n59600 , n59601 , n59602 , n59603 , n59604 , n59605 , n59606 , 
 n59607 , n59608 , n59609 , n59610 , n59611 , n59612 , n59613 , n59614 , n59615 , n59616 , 
 n59617 , n59618 , n59619 , n59620 , n59621 , n59622 , n59623 , n59624 , n59625 , n59626 , 
 n59627 , n59628 , n59629 , n59630 , n59631 , n59632 , n59633 , n59634 , n59635 , n59636 , 
 n59637 , n59638 , n59639 , n59640 , n59641 , n59642 , n59643 , n59644 , n59645 , n59646 , 
 n59647 , n59648 , n59649 , n59650 , n59651 , n59652 , n59653 , n59654 , n59655 , n59656 , 
 n59657 , n59658 , n59659 , n59660 , n59661 , n59662 , n59663 , n59664 , n59665 , n59666 , 
 n59667 , n59668 , n59669 , n59670 , n59671 , n59672 , n59673 , n59674 , n59675 , n59676 , 
 n59677 , n59678 , n59679 , n59680 , n59681 , n59682 , n59683 , n59684 , n59685 , n59686 , 
 n59687 , n59688 , n59689 , n59690 , n59691 , n59692 , n59693 , n59694 , n59695 , n59696 , 
 n59697 , n59698 , n59699 , n59700 , n59701 , n59702 , n59703 , n59704 , n59705 , n59706 , 
 n59707 , n59708 , n59709 , n59710 , n59711 , n59712 , n59713 , n59714 , n59715 , n59716 , 
 n59717 , n59718 , n59719 , n59720 , n59721 , n59722 , n59723 , n59724 , n59725 , n59726 , 
 n59727 , n59728 , n59729 , n59730 , n59731 , n59732 , n59733 , n59734 , n59735 , n59736 , 
 n59737 , n59738 , n59739 , n59740 , n59741 , n59742 , n59743 , n59744 , n59745 , n59746 , 
 n59747 , n59748 , n59749 , n59750 , n59751 , n59752 , n59753 , n59754 , n59755 , n59756 , 
 n59757 , n59758 , n59759 , n59760 , n59761 , n59762 , n59763 , n59764 , n59765 , n59766 , 
 n59767 , n59768 , n59769 , n59770 , n59771 , n59772 , n59773 , n59774 , n59775 , n59776 , 
 n59777 , n59778 , n59779 , n59780 , n59781 , n59782 , n59783 , n59784 , n59785 , n59786 , 
 n59787 , n59788 , n59789 , n59790 , n59791 , n59792 , n59793 , n59794 , n59795 , n59796 , 
 n59797 , n59798 , n59799 , n59800 , n59801 , n59802 , n59803 , n59804 , n59805 , n59806 , 
 n59807 , n59808 , n59809 , n59810 , n59811 , n59812 , n59813 , n59814 , n59815 , n59816 , 
 n59817 , n59818 , n59819 , n59820 , n59821 , n59822 , n59823 , n59824 , n59825 , n59826 , 
 n59827 , n59828 , n59829 , n59830 , n59831 , n59832 , n59833 , n59834 , n59835 , n59836 , 
 n59837 , n59838 , n59839 , n59840 , n59841 , n59842 , n59843 , n59844 , n59845 , n59846 , 
 n59847 , n59848 , n59849 , n59850 , n59851 , n59852 , n59853 , n59854 , n59855 , n59856 , 
 n59857 , n59858 , n59859 , n59860 , n59861 , n59862 , n59863 , n59864 , n59865 , n59866 , 
 n59867 , n59868 , n59869 , n59870 , n59871 , n59872 , n59873 , n59874 , n59875 , n59876 , 
 n59877 , n59878 , n59879 , n59880 , n59881 , n59882 , n59883 , n59884 , n59885 , n59886 , 
 n59887 , n59888 , n59889 , n59890 , n59891 , n59892 , n59893 , n59894 , n59895 , n59896 , 
 n59897 , n59898 , n59899 , n59900 , n59901 , n59902 , n59903 , n59904 , n59905 , n59906 , 
 n59907 , n59908 , n59909 , n59910 , n59911 , n59912 , n59913 , n59914 , n59915 , n59916 , 
 n59917 , n59918 , n59919 , n59920 , n59921 , n59922 , n59923 , n59924 , n59925 , n59926 , 
 n59927 , n59928 , n59929 , n59930 , n59931 , n59932 , n59933 , n59934 , n59935 , n59936 , 
 n59937 , n59938 , n59939 , n59940 , n59941 , n59942 , n59943 , n59944 , n59945 , n59946 , 
 n59947 , n59948 , n59949 , n59950 , n59951 , n59952 , n59953 , n59954 , n59955 , n59956 , 
 n59957 , n59958 , n59959 , n59960 , n59961 , n59962 , n59963 , n59964 , n59965 , n59966 , 
 n59967 , n59968 , n59969 , n59970 , n59971 , n59972 , n59973 , n59974 , n59975 , n59976 , 
 n59977 , n59978 , n59979 , n59980 , n59981 , n59982 , n59983 , n59984 , n59985 , n59986 , 
 n59987 , n59988 , n59989 , n59990 , n59991 , n59992 , n59993 , n59994 , n59995 , n59996 , 
 n59997 , n59998 , n59999 , n60000 , n60001 , n60002 , n60003 , n60004 , n60005 , n60006 , 
 n60007 , n60008 , n60009 , n60010 , n60011 , n60012 , n60013 , n60014 , n60015 , n60016 , 
 n60017 , n60018 , n60019 , n60020 , n60021 , n60022 , n60023 , n60024 , n60025 , n60026 , 
 n60027 , n60028 , n60029 , n60030 , n60031 , n60032 , n60033 , n60034 , n60035 , n60036 , 
 n60037 , n60038 , n60039 , n60040 , n60041 , n60042 , n60043 , n60044 , n60045 , n60046 , 
 n60047 , n60048 , n60049 , n60050 , n60051 , n60052 , n60053 , n60054 , n60055 , n60056 , 
 n60057 , n60058 , n60059 , n60060 , n60061 , n60062 , n60063 , n60064 , n60065 , n60066 , 
 n60067 , n60068 , n60069 , n60070 , n60071 , n60072 , n60073 , n60074 , n60075 , n60076 , 
 n60077 , n60078 , n60079 , n60080 , n60081 , n60082 , n60083 , n60084 , n60085 , n60086 , 
 n60087 , n60088 , n60089 , n60090 , n60091 , n60092 , n60093 , n60094 , n60095 , n60096 , 
 n60097 , n60098 , n60099 , n60100 , n60101 , n60102 , n60103 , n60104 , n60105 , n60106 , 
 n60107 , n60108 , n60109 , n60110 , n60111 , n60112 , n60113 , n60114 , n60115 , n60116 , 
 n60117 , n60118 , n60119 , n60120 , n60121 , n60122 , n60123 , n60124 , n60125 , n60126 , 
 n60127 , n60128 , n60129 , n60130 , n60131 , n60132 , n60133 , n60134 , n60135 , n60136 , 
 n60137 , n60138 , n60139 , n60140 , n60141 , n60142 , n60143 , n60144 , n60145 , n60146 , 
 n60147 , n60148 , n60149 , n60150 , n60151 , n60152 , n60153 , n60154 , n60155 , n60156 , 
 n60157 , n60158 , n60159 , n60160 , n60161 , n60162 , n60163 , n60164 , n60165 , n60166 , 
 n60167 , n60168 , n60169 , n60170 , n60171 , n60172 , n60173 , n60174 , n60175 , n60176 , 
 n60177 , n60178 , n60179 , n60180 , n60181 , n60182 , n60183 , n60184 , n60185 , n60186 , 
 n60187 , n60188 , n60189 , n60190 , n60191 , n60192 , n60193 , n60194 , n60195 , n60196 , 
 n60197 , n60198 , n60199 , n60200 , n60201 , n60202 , n60203 , n60204 , n60205 , n60206 , 
 n60207 , n60208 , n60209 , n60210 , n60211 , n60212 , n60213 , n60214 , n60215 , n60216 , 
 n60217 , n60218 , n60219 , n60220 , n60221 , n60222 , n60223 , n60224 , n60225 , n60226 , 
 n60227 , n60228 , n60229 , n60230 , n60231 , n60232 , n60233 , n60234 , n60235 , n60236 , 
 n60237 , n60238 , n60239 , n60240 , n60241 , n60242 , n60243 , n60244 , n60245 , n60246 , 
 n60247 , n60248 , n60249 , n60250 , n60251 , n60252 , n60253 , n60254 , n60255 , n60256 , 
 n60257 , n60258 , n60259 , n60260 , n60261 , n60262 , n60263 , n60264 , n60265 , n60266 , 
 n60267 , n60268 , n60269 , n60270 , n60271 , n60272 , n60273 , n60274 , n60275 , n60276 , 
 n60277 , n60278 , n60279 , n60280 , n60281 , n60282 , n60283 , n60284 , n60285 , n60286 , 
 n60287 , n60288 , n60289 , n60290 , n60291 , n60292 , n60293 , n60294 , n60295 , n60296 , 
 n60297 , n60298 , n60299 , n60300 , n60301 , n60302 , n60303 , n60304 , n60305 , n60306 , 
 n60307 , n60308 , n60309 , n60310 , n60311 , n60312 , n60313 , n60314 , n60315 , n60316 , 
 n60317 , n60318 , n60319 , n60320 , n60321 , n60322 , n60323 , n60324 , n60325 , n60326 , 
 n60327 , n60328 , n60329 , n60330 , n60331 , n60332 , n60333 , n60334 , n60335 , n60336 , 
 n60337 , n60338 , n60339 , n60340 , n60341 , n60342 , n60343 , n60344 , n60345 , n60346 , 
 n60347 , n60348 , n60349 , n60350 , n60351 , n60352 , n60353 , n60354 , n60355 , n60356 , 
 n60357 , n60358 , n60359 , n60360 , n60361 , n60362 , n60363 , n60364 , n60365 , n60366 , 
 n60367 , n60368 , n60369 , n60370 , n60371 , n60372 , n60373 , n60374 , n60375 , n60376 , 
 n60377 , n60378 , n60379 , n60380 , n60381 , n60382 , n60383 , n60384 , n60385 , n60386 , 
 n60387 , n60388 , n60389 , n60390 , n60391 , n60392 , n60393 , n60394 , n60395 , n60396 , 
 n60397 , n60398 , n60399 , n60400 , n60401 , n60402 , n60403 , n60404 , n60405 , n60406 , 
 n60407 , n60408 , n60409 , n60410 , n60411 , n60412 , n60413 , n60414 , n60415 , n60416 , 
 n60417 , n60418 , n60419 , n60420 , n60421 , n60422 , n60423 , n60424 , n60425 , n60426 , 
 n60427 , n60428 , n60429 , n60430 , n60431 , n60432 , n60433 , n60434 , n60435 , n60436 , 
 n60437 , n60438 , n60439 , n60440 , n60441 , n60442 , n60443 , n60444 , n60445 , n60446 , 
 n60447 , n60448 , n60449 , n60450 , n60451 , n60452 , n60453 , n60454 , n60455 , n60456 , 
 n60457 , n60458 , n60459 , n60460 , n60461 , n60462 , n60463 , n60464 , n60465 , n60466 , 
 n60467 , n60468 , n60469 , n60470 , n60471 , n60472 , n60473 , n60474 , n60475 , n60476 , 
 n60477 , n60478 , n60479 , n60480 , n60481 , n60482 , n60483 , n60484 , n60485 , n60486 , 
 n60487 , n60488 , n60489 , n60490 , n60491 , n60492 , n60493 , n60494 , n60495 , n60496 , 
 n60497 , n60498 , n60499 , n60500 , n60501 , n60502 , n60503 , n60504 , n60505 , n60506 , 
 n60507 , n60508 , n60509 , n60510 , n60511 , n60512 , n60513 , n60514 , n60515 , n60516 , 
 n60517 , n60518 , n60519 , n60520 , n60521 , n60522 , n60523 , n60524 , n60525 , n60526 , 
 n60527 , n60528 , n60529 , n60530 , n60531 , n60532 , n60533 , n60534 , n60535 , n60536 , 
 n60537 , n60538 , n60539 , n60540 , n60541 , n60542 , n60543 , n60544 , n60545 , n60546 , 
 n60547 , n60548 , n60549 , n60550 , n60551 , n60552 , n60553 , n60554 , n60555 , n60556 , 
 n60557 , n60558 , n60559 , n60560 , n60561 , n60562 , n60563 , n60564 , n60565 , n60566 , 
 n60567 , n60568 , n60569 , n60570 , n60571 , n60572 , n60573 , n60574 , n60575 , n60576 , 
 n60577 , n60578 , n60579 , n60580 , n60581 , n60582 , n60583 , n60584 , n60585 , n60586 , 
 n60587 , n60588 , n60589 , n60590 , n60591 , n60592 , n60593 , n60594 , n60595 , n60596 , 
 n60597 , n60598 , n60599 , n60600 , n60601 , n60602 , n60603 , n60604 , n60605 , n60606 , 
 n60607 , n60608 , n60609 , n60610 , n60611 , n60612 , n60613 , n60614 , n60615 , n60616 , 
 n60617 , n60618 , n60619 , n60620 , n60621 , n60622 , n60623 , n60624 , n60625 , n60626 , 
 n60627 , n60628 , n60629 , n60630 , n60631 , n60632 , n60633 , n60634 , n60635 , n60636 , 
 n60637 , n60638 , n60639 , n60640 , n60641 , n60642 , n60643 , n60644 , n60645 , n60646 , 
 n60647 , n60648 , n60649 , n60650 , n60651 , n60652 , n60653 , n60654 , n60655 , n60656 , 
 n60657 , n60658 , n60659 , n60660 , n60661 , n60662 , n60663 , n60664 , n60665 , n60666 , 
 n60667 , n60668 , n60669 , n60670 , n60671 , n60672 , n60673 , n60674 , n60675 , n60676 , 
 n60677 , n60678 , n60679 , n60680 , n60681 , n60682 , n60683 , n60684 , n60685 , n60686 , 
 n60687 , n60688 , n60689 , n60690 , n60691 , n60692 , n60693 , n60694 , n60695 , n60696 , 
 n60697 , n60698 , n60699 , n60700 , n60701 , n60702 , n60703 , n60704 , n60705 , n60706 , 
 n60707 , n60708 , n60709 , n60710 , n60711 , n60712 , n60713 , n60714 , n60715 , n60716 , 
 n60717 , n60718 , n60719 , n60720 , n60721 , n60722 , n60723 , n60724 , n60725 , n60726 , 
 n60727 , n60728 , n60729 , n60730 , n60731 , n60732 , n60733 , n60734 , n60735 , n60736 , 
 n60737 , n60738 , n60739 , n60740 , n60741 , n60742 , n60743 , n60744 , n60745 , n60746 , 
 n60747 , n60748 , n60749 , n60750 , n60751 , n60752 , n60753 , n60754 , n60755 , n60756 , 
 n60757 , n60758 , n60759 , n60760 , n60761 , n60762 , n60763 , n60764 , n60765 , n60766 , 
 n60767 , n60768 , n60769 , n60770 , n60771 , n60772 , n60773 , n60774 , n60775 , n60776 , 
 n60777 , n60778 , n60779 , n60780 , n60781 , n60782 , n60783 , n60784 , n60785 , n60786 , 
 n60787 , n60788 , n60789 , n60790 , n60791 , n60792 , n60793 , n60794 , n60795 , n60796 , 
 n60797 , n60798 , n60799 , n60800 , n60801 , n60802 , n60803 , n60804 , n60805 , n60806 , 
 n60807 , n60808 , n60809 , n60810 , n60811 , n60812 , n60813 , n60814 , n60815 , n60816 , 
 n60817 , n60818 , n60819 , n60820 , n60821 , n60822 , n60823 , n60824 , n60825 , n60826 , 
 n60827 , n60828 , n60829 , n60830 , n60831 , n60832 , n60833 , n60834 , n60835 , n60836 , 
 n60837 , n60838 , n60839 , n60840 , n60841 , n60842 , n60843 , n60844 , n60845 , n60846 , 
 n60847 , n60848 , n60849 , n60850 , n60851 , n60852 , n60853 , n60854 , n60855 , n60856 , 
 n60857 , n60858 , n60859 , n60860 , n60861 , n60862 , n60863 , n60864 , n60865 , n60866 , 
 n60867 , n60868 , n60869 , n60870 , n60871 , n60872 , n60873 , n60874 , n60875 , n60876 , 
 n60877 , n60878 , n60879 , n60880 , n60881 , n60882 , n60883 , n60884 , n60885 , n60886 , 
 n60887 , n60888 , n60889 , n60890 , n60891 , n60892 , n60893 , n60894 , n60895 , n60896 , 
 n60897 , n60898 , n60899 , n60900 , n60901 , n60902 , n60903 , n60904 , n60905 , n60906 , 
 n60907 , n60908 , n60909 , n60910 , n60911 , n60912 , n60913 , n60914 , n60915 , n60916 , 
 n60917 , n60918 , n60919 , n60920 , n60921 , n60922 , n60923 , n60924 , n60925 , n60926 , 
 n60927 , n60928 , n60929 , n60930 , n60931 , n60932 , n60933 , n60934 , n60935 , n60936 , 
 n60937 , n60938 , n60939 , n60940 , n60941 , n60942 , n60943 , n60944 , n60945 , n60946 , 
 n60947 , n60948 , n60949 , n60950 , n60951 , n60952 , n60953 , n60954 , n60955 , n60956 , 
 n60957 , n60958 , n60959 , n60960 , n60961 , n60962 , n60963 , n60964 , n60965 , n60966 , 
 n60967 , n60968 , n60969 , n60970 , n60971 , n60972 , n60973 , n60974 , n60975 , n60976 , 
 n60977 , n60978 , n60979 , n60980 , n60981 , n60982 , n60983 , n60984 , n60985 , n60986 , 
 n60987 , n60988 , n60989 , n60990 , n60991 , n60992 , n60993 , n60994 , n60995 , n60996 , 
 n60997 , n60998 , n60999 , n61000 , n61001 , n61002 , n61003 , n61004 , n61005 , n61006 , 
 n61007 , n61008 , n61009 , n61010 , n61011 , n61012 , n61013 , n61014 , n61015 , n61016 , 
 n61017 , n61018 , n61019 , n61020 , n61021 , n61022 , n61023 , n61024 , n61025 , n61026 , 
 n61027 , n61028 , n61029 , n61030 , n61031 , n61032 , n61033 , n61034 , n61035 , n61036 , 
 n61037 , n61038 , n61039 , n61040 , n61041 , n61042 , n61043 , n61044 , n61045 , n61046 , 
 n61047 , n61048 , n61049 , n61050 , n61051 , n61052 , n61053 , n61054 , n61055 , n61056 , 
 n61057 , n61058 , n61059 , n61060 , n61061 , n61062 , n61063 , n61064 , n61065 , n61066 , 
 n61067 , n61068 , n61069 , n61070 , n61071 , n61072 , n61073 , n61074 , n61075 , n61076 , 
 n61077 , n61078 , n61079 , n61080 , n61081 , n61082 , n61083 , n61084 , n61085 , n61086 , 
 n61087 , n61088 , n61089 , n61090 , n61091 , n61092 , n61093 , n61094 , n61095 , n61096 , 
 n61097 , n61098 , n61099 , n61100 , n61101 , n61102 , n61103 , n61104 , n61105 , n61106 , 
 n61107 , n61108 , n61109 , n61110 , n61111 , n61112 , n61113 , n61114 , n61115 , n61116 , 
 n61117 , n61118 , n61119 , n61120 , n61121 , n61122 , n61123 , n61124 , n61125 , n61126 , 
 n61127 , n61128 , n61129 , n61130 , n61131 , n61132 , n61133 , n61134 , n61135 , n61136 , 
 n61137 , n61138 , n61139 , n61140 , n61141 , n61142 , n61143 , n61144 , n61145 , n61146 , 
 n61147 , n61148 , n61149 , n61150 , n61151 , n61152 , n61153 , n61154 , n61155 , n61156 , 
 n61157 , n61158 , n61159 , n61160 , n61161 , n61162 , n61163 , n61164 , n61165 , n61166 , 
 n61167 , n61168 , n61169 , n61170 , n61171 , n61172 , n61173 , n61174 , n61175 , n61176 , 
 n61177 , n61178 , n61179 , n61180 , n61181 , n61182 , n61183 , n61184 , n61185 , n61186 , 
 n61187 , n61188 , n61189 , n61190 , n61191 , n61192 , n61193 , n61194 , n61195 , n61196 , 
 n61197 , n61198 , n61199 , n61200 , n61201 , n61202 , n61203 , n61204 , n61205 , n61206 , 
 n61207 , n61208 , n61209 , n61210 , n61211 , n61212 , n61213 , n61214 , n61215 , n61216 , 
 n61217 , n61218 , n61219 , n61220 , n61221 , n61222 , n61223 , n61224 , n61225 , n61226 , 
 n61227 , n61228 , n61229 , n61230 , n61231 , n61232 , n61233 , n61234 , n61235 , n61236 , 
 n61237 , n61238 , n61239 , n61240 , n61241 , n61242 , n61243 , n61244 , n61245 , n61246 , 
 n61247 , n61248 , n61249 , n61250 , n61251 , n61252 , n61253 , n61254 , n61255 , n61256 , 
 n61257 , n61258 , n61259 , n61260 , n61261 , n61262 , n61263 , n61264 , n61265 , n61266 , 
 n61267 , n61268 , n61269 , n61270 , n61271 , n61272 , n61273 , n61274 , n61275 , n61276 , 
 n61277 , n61278 , n61279 , n61280 , n61281 , n61282 , n61283 , n61284 , n61285 , n61286 , 
 n61287 , n61288 , n61289 , n61290 , n61291 , n61292 , n61293 , n61294 , n61295 , n61296 , 
 n61297 , n61298 , n61299 , n61300 , n61301 , n61302 , n61303 , n61304 , n61305 , n61306 , 
 n61307 , n61308 , n61309 , n61310 , n61311 , n61312 , n61313 , n61314 , n61315 , n61316 , 
 n61317 , n61318 , n61319 , n61320 , n61321 , n61322 , n61323 , n61324 , n61325 , n61326 , 
 n61327 , n61328 , n61329 , n61330 , n61331 , n61332 , n61333 , n61334 , n61335 , n61336 , 
 n61337 , n61338 , n61339 , n61340 , n61341 , n61342 , n61343 , n61344 , n61345 , n61346 , 
 n61347 , n61348 , n61349 , n61350 , n61351 , n61352 , n61353 , n61354 , n61355 , n61356 , 
 n61357 , n61358 , n61359 , n61360 , n61361 , n61362 , n61363 , n61364 , n61365 , n61366 , 
 n61367 , n61368 , n61369 , n61370 , n61371 , n61372 , n61373 , n61374 , n61375 , n61376 , 
 n61377 , n61378 , n61379 , n61380 , n61381 , n61382 , n61383 , n61384 , n61385 , n61386 , 
 n61387 , n61388 , n61389 , n61390 , n61391 , n61392 , n61393 , n61394 , n61395 , n61396 , 
 n61397 , n61398 , n61399 , n61400 , n61401 , n61402 , n61403 , n61404 , n61405 , n61406 , 
 n61407 , n61408 , n61409 , n61410 , n61411 , n61412 , n61413 , n61414 , n61415 , n61416 , 
 n61417 , n61418 , n61419 , n61420 , n61421 , n61422 , n61423 , n61424 , n61425 , n61426 , 
 n61427 , n61428 , n61429 , n61430 , n61431 , n61432 , n61433 , n61434 , n61435 , n61436 , 
 n61437 , n61438 , n61439 , n61440 , n61441 , n61442 , n61443 , n61444 , n61445 , n61446 , 
 n61447 , n61448 , n61449 , n61450 , n61451 , n61452 , n61453 , n61454 , n61455 , n61456 , 
 n61457 , n61458 , n61459 , n61460 , n61461 , n61462 , n61463 , n61464 , n61465 , n61466 , 
 n61467 , n61468 , n61469 , n61470 , n61471 , n61472 , n61473 , n61474 , n61475 , n61476 , 
 n61477 , n61478 , n61479 , n61480 , n61481 , n61482 , n61483 , n61484 , n61485 , n61486 , 
 n61487 , n61488 , n61489 , n61490 , n61491 , n61492 , n61493 , n61494 , n61495 , n61496 , 
 n61497 , n61498 , n61499 , n61500 , n61501 , n61502 , n61503 , n61504 , n61505 , n61506 , 
 n61507 , n61508 , n61509 , n61510 , n61511 , n61512 , n61513 , n61514 , n61515 , n61516 , 
 n61517 , n61518 , n61519 , n61520 , n61521 , n61522 , n61523 , n61524 , n61525 , n61526 , 
 n61527 , n61528 , n61529 , n61530 , n61531 , n61532 , n61533 , n61534 , n61535 , n61536 , 
 n61537 , n61538 , n61539 , n61540 , n61541 , n61542 , n61543 , n61544 , n61545 , n61546 , 
 n61547 , n61548 , n61549 , n61550 , n61551 , n61552 , n61553 , n61554 , n61555 , n61556 , 
 n61557 , n61558 , n61559 , n61560 , n61561 , n61562 , n61563 , n61564 , n61565 , n61566 , 
 n61567 , n61568 , n61569 , n61570 , n61571 , n61572 , n61573 , n61574 , n61575 , n61576 , 
 n61577 , n61578 , n61579 , n61580 , n61581 , n61582 , n61583 , n61584 , n61585 , n61586 , 
 n61587 , n61588 , n61589 , n61590 , n61591 , n61592 , n61593 , n61594 , n61595 , n61596 , 
 n61597 , n61598 , n61599 , n61600 , n61601 , n61602 , n61603 , n61604 , n61605 , n61606 , 
 n61607 , n61608 , n61609 , n61610 , n61611 , n61612 , n61613 , n61614 , n61615 , n61616 , 
 n61617 , n61618 , n61619 , n61620 , n61621 , n61622 , n61623 , n61624 , n61625 , n61626 , 
 n61627 , n61628 , n61629 , n61630 , n61631 , n61632 , n61633 , n61634 , n61635 , n61636 , 
 n61637 , n61638 , n61639 , n61640 , n61641 , n61642 , n61643 , n61644 , n61645 , n61646 , 
 n61647 , n61648 , n61649 , n61650 , n61651 , n61652 , n61653 , n61654 , n61655 , n61656 , 
 n61657 , n61658 , n61659 , n61660 , n61661 , n61662 , n61663 , n61664 , n61665 , n61666 , 
 n61667 , n61668 , n61669 , n61670 , n61671 , n61672 , n61673 , n61674 , n61675 , n61676 , 
 n61677 , n61678 , n61679 , n61680 , n61681 , n61682 , n61683 , n61684 , n61685 , n61686 , 
 n61687 , n61688 , n61689 , n61690 , n61691 , n61692 , n61693 , n61694 , n61695 , n61696 , 
 n61697 , n61698 , n61699 , n61700 , n61701 , n61702 , n61703 , n61704 , n61705 , n61706 , 
 n61707 , n61708 , n61709 , n61710 , n61711 , n61712 , n61713 , n61714 , n61715 , n61716 , 
 n61717 , n61718 , n61719 , n61720 , n61721 , n61722 , n61723 , n61724 , n61725 , n61726 , 
 n61727 , n61728 , n61729 , n61730 , n61731 , n61732 , n61733 , n61734 , n61735 , n61736 , 
 n61737 , n61738 , n61739 , n61740 , n61741 , n61742 , n61743 , n61744 , n61745 , n61746 , 
 n61747 , n61748 , n61749 , n61750 , n61751 , n61752 , n61753 , n61754 , n61755 , n61756 , 
 n61757 , n61758 , n61759 , n61760 , n61761 , n61762 , n61763 , n61764 , n61765 , n61766 , 
 n61767 , n61768 , n61769 , n61770 , n61771 , n61772 , n61773 , n61774 , n61775 , n61776 , 
 n61777 , n61778 , n61779 , n61780 , n61781 , n61782 , n61783 , n61784 , n61785 , n61786 , 
 n61787 , n61788 , n61789 , n61790 , n61791 , n61792 , n61793 , n61794 , n61795 , n61796 , 
 n61797 , n61798 , n61799 , n61800 , n61801 , n61802 , n61803 , n61804 , n61805 , n61806 , 
 n61807 , n61808 , n61809 , n61810 , n61811 , n61812 , n61813 , n61814 , n61815 , n61816 , 
 n61817 , n61818 , n61819 , n61820 , n61821 , n61822 , n61823 , n61824 , n61825 , n61826 , 
 n61827 , n61828 , n61829 , n61830 , n61831 , n61832 , n61833 , n61834 , n61835 , n61836 , 
 n61837 , n61838 , n61839 , n61840 , n61841 , n61842 , n61843 , n61844 , n61845 , n61846 , 
 n61847 , n61848 , n61849 , n61850 , n61851 , n61852 , n61853 , n61854 , n61855 , n61856 , 
 n61857 , n61858 , n61859 , n61860 , n61861 , n61862 , n61863 , n61864 , n61865 , n61866 , 
 n61867 , n61868 , n61869 , n61870 , n61871 , n61872 , n61873 , n61874 , n61875 , n61876 , 
 n61877 , n61878 , n61879 , n61880 , n61881 , n61882 , n61883 , n61884 , n61885 , n61886 , 
 n61887 , n61888 , n61889 , n61890 , n61891 , n61892 , n61893 , n61894 , n61895 , n61896 , 
 n61897 , n61898 , n61899 , n61900 , n61901 , n61902 , n61903 , n61904 , n61905 , n61906 , 
 n61907 , n61908 , n61909 , n61910 , n61911 , n61912 , n61913 , n61914 , n61915 , n61916 , 
 n61917 , n61918 , n61919 , n61920 , n61921 , n61922 , n61923 , n61924 , n61925 , n61926 , 
 n61927 , n61928 , n61929 , n61930 , n61931 , n61932 , n61933 , n61934 , n61935 , n61936 , 
 n61937 , n61938 , n61939 , n61940 , n61941 , n61942 , n61943 , n61944 , n61945 , n61946 , 
 n61947 , n61948 , n61949 , n61950 , n61951 , n61952 , n61953 , n61954 , n61955 , n61956 , 
 n61957 , n61958 , n61959 , n61960 , n61961 , n61962 , n61963 , n61964 , n61965 , n61966 , 
 n61967 , n61968 , n61969 , n61970 , n61971 , n61972 , n61973 , n61974 , n61975 , n61976 , 
 n61977 , n61978 , n61979 , n61980 , n61981 , n61982 , n61983 , n61984 , n61985 , n61986 , 
 n61987 , n61988 , n61989 , n61990 , n61991 , n61992 , n61993 , n61994 , n61995 , n61996 , 
 n61997 , n61998 , n61999 , n62000 , n62001 , n62002 , n62003 , n62004 , n62005 , n62006 , 
 n62007 , n62008 , n62009 , n62010 , n62011 , n62012 , n62013 , n62014 , n62015 , n62016 , 
 n62017 , n62018 , n62019 , n62020 , n62021 , n62022 , n62023 , n62024 , n62025 , n62026 , 
 n62027 , n62028 , n62029 , n62030 , n62031 , n62032 , n62033 , n62034 , n62035 , n62036 , 
 n62037 , n62038 , n62039 , n62040 , n62041 , n62042 , n62043 , n62044 , n62045 , n62046 , 
 n62047 , n62048 , n62049 , n62050 , n62051 , n62052 , n62053 , n62054 , n62055 , n62056 , 
 n62057 , n62058 , n62059 , n62060 , n62061 , n62062 , n62063 , n62064 , n62065 , n62066 , 
 n62067 , n62068 , n62069 , n62070 , n62071 , n62072 , n62073 , n62074 , n62075 , n62076 , 
 n62077 , n62078 , n62079 , n62080 , n62081 , n62082 , n62083 , n62084 , n62085 , n62086 , 
 n62087 , n62088 , n62089 , n62090 , n62091 , n62092 , n62093 , n62094 , n62095 , n62096 , 
 n62097 , n62098 , n62099 , n62100 , n62101 , n62102 , n62103 , n62104 , n62105 , n62106 , 
 n62107 , n62108 , n62109 , n62110 , n62111 , n62112 , n62113 , n62114 , n62115 , n62116 , 
 n62117 , n62118 , n62119 , n62120 , n62121 , n62122 , n62123 , n62124 , n62125 , n62126 , 
 n62127 , n62128 , n62129 , n62130 , n62131 , n62132 , n62133 , n62134 , n62135 , n62136 , 
 n62137 , n62138 , n62139 , n62140 , n62141 , n62142 , n62143 , n62144 , n62145 , n62146 , 
 n62147 , n62148 , n62149 , n62150 , n62151 , n62152 , n62153 , n62154 , n62155 , n62156 , 
 n62157 , n62158 , n62159 , n62160 , n62161 , n62162 , n62163 , n62164 , n62165 , n62166 , 
 n62167 , n62168 , n62169 , n62170 , n62171 , n62172 , n62173 , n62174 , n62175 , n62176 , 
 n62177 , n62178 , n62179 , n62180 , n62181 , n62182 , n62183 , n62184 , n62185 , n62186 , 
 n62187 , n62188 , n62189 , n62190 , n62191 , n62192 , n62193 , n62194 , n62195 , n62196 , 
 n62197 , n62198 , n62199 , n62200 , n62201 , n62202 , n62203 , n62204 , n62205 , n62206 , 
 n62207 , n62208 , n62209 , n62210 , n62211 , n62212 , n62213 , n62214 , n62215 , n62216 , 
 n62217 , n62218 , n62219 , n62220 , n62221 , n62222 , n62223 , n62224 , n62225 , n62226 , 
 n62227 , n62228 , n62229 , n62230 , n62231 , n62232 , n62233 , n62234 , n62235 , n62236 , 
 n62237 , n62238 , n62239 , n62240 , n62241 , n62242 , n62243 , n62244 , n62245 , n62246 , 
 n62247 , n62248 , n62249 , n62250 , n62251 , n62252 , n62253 , n62254 , n62255 , n62256 , 
 n62257 , n62258 , n62259 , n62260 , n62261 , n62262 , n62263 , n62264 , n62265 , n62266 , 
 n62267 , n62268 , n62269 , n62270 , n62271 , n62272 , n62273 , n62274 , n62275 , n62276 , 
 n62277 , n62278 , n62279 , n62280 , n62281 , n62282 , n62283 , n62284 , n62285 , n62286 , 
 n62287 , n62288 , n62289 , n62290 , n62291 , n62292 , n62293 , n62294 , n62295 , n62296 , 
 n62297 , n62298 , n62299 , n62300 , n62301 , n62302 , n62303 , n62304 , n62305 , n62306 , 
 n62307 , n62308 , n62309 , n62310 , n62311 , n62312 , n62313 , n62314 , n62315 , n62316 , 
 n62317 , n62318 , n62319 , n62320 , n62321 , n62322 , n62323 , n62324 , n62325 , n62326 , 
 n62327 , n62328 , n62329 , n62330 , n62331 , n62332 , n62333 , n62334 , n62335 , n62336 , 
 n62337 , n62338 , n62339 , n62340 , n62341 , n62342 , n62343 , n62344 , n62345 , n62346 , 
 n62347 , n62348 , n62349 , n62350 , n62351 , n62352 , n62353 , n62354 , n62355 , n62356 , 
 n62357 , n62358 , n62359 , n62360 , n62361 , n62362 , n62363 , n62364 , n62365 , n62366 , 
 n62367 , n62368 , n62369 , n62370 , n62371 , n62372 , n62373 , n62374 , n62375 , n62376 , 
 n62377 , n62378 , n62379 , n62380 , n62381 , n62382 , n62383 , n62384 , n62385 , n62386 , 
 n62387 , n62388 , n62389 , n62390 , n62391 , n62392 , n62393 , n62394 , n62395 , n62396 , 
 n62397 , n62398 , n62399 , n62400 , n62401 , n62402 , n62403 , n62404 , n62405 , n62406 , 
 n62407 , n62408 , n62409 , n62410 , n62411 , n62412 , n62413 , n62414 , n62415 , n62416 , 
 n62417 , n62418 , n62419 , n62420 , n62421 , n62422 , n62423 , n62424 , n62425 , n62426 , 
 n62427 , n62428 , n62429 , n62430 , n62431 , n62432 , n62433 , n62434 , n62435 , n62436 , 
 n62437 , n62438 , n62439 , n62440 , n62441 , n62442 , n62443 , n62444 , n62445 , n62446 , 
 n62447 , n62448 , n62449 , n62450 , n62451 , n62452 , n62453 , n62454 , n62455 , n62456 , 
 n62457 , n62458 , n62459 , n62460 , n62461 , n62462 , n62463 , n62464 , n62465 , n62466 , 
 n62467 , n62468 , n62469 , n62470 , n62471 , n62472 , n62473 , n62474 , n62475 , n62476 , 
 n62477 , n62478 , n62479 , n62480 , n62481 , n62482 , n62483 , n62484 , n62485 , n62486 , 
 n62487 , n62488 , n62489 , n62490 , n62491 , n62492 , n62493 , n62494 , n62495 , n62496 , 
 n62497 , n62498 , n62499 , n62500 , n62501 , n62502 , n62503 , n62504 , n62505 , n62506 , 
 n62507 , n62508 , n62509 , n62510 , n62511 , n62512 , n62513 , n62514 , n62515 , n62516 , 
 n62517 , n62518 , n62519 , n62520 , n62521 , n62522 , n62523 , n62524 , n62525 , n62526 , 
 n62527 , n62528 , n62529 , n62530 , n62531 , n62532 , n62533 , n62534 , n62535 , n62536 , 
 n62537 , n62538 , n62539 , n62540 , n62541 , n62542 , n62543 , n62544 , n62545 , n62546 , 
 n62547 , n62548 , n62549 , n62550 , n62551 , n62552 , n62553 , n62554 , n62555 , n62556 , 
 n62557 , n62558 , n62559 , n62560 , n62561 , n62562 , n62563 , n62564 , n62565 , n62566 , 
 n62567 , n62568 , n62569 , n62570 , n62571 , n62572 , n62573 , n62574 , n62575 , n62576 , 
 n62577 , n62578 , n62579 , n62580 , n62581 , n62582 , n62583 , n62584 , n62585 , n62586 , 
 n62587 , n62588 , n62589 , n62590 , n62591 , n62592 , n62593 , n62594 , n62595 , n62596 , 
 n62597 , n62598 , n62599 , n62600 , n62601 , n62602 , n62603 , n62604 , n62605 , n62606 , 
 n62607 , n62608 , n62609 , n62610 , n62611 , n62612 , n62613 , n62614 , n62615 , n62616 , 
 n62617 , n62618 , n62619 , n62620 , n62621 , n62622 , n62623 , n62624 , n62625 , n62626 , 
 n62627 , n62628 , n62629 , n62630 , n62631 , n62632 , n62633 , n62634 , n62635 , n62636 , 
 n62637 , n62638 , n62639 , n62640 , n62641 , n62642 , n62643 , n62644 , n62645 , n62646 , 
 n62647 , n62648 , n62649 , n62650 , n62651 , n62652 , n62653 , n62654 , n62655 , n62656 , 
 n62657 , n62658 , n62659 , n62660 , n62661 , n62662 , n62663 , n62664 , n62665 , n62666 , 
 n62667 , n62668 , n62669 , n62670 , n62671 , n62672 , n62673 , n62674 , n62675 , n62676 , 
 n62677 , n62678 , n62679 , n62680 , n62681 , n62682 , n62683 , n62684 , n62685 , n62686 , 
 n62687 , n62688 , n62689 , n62690 , n62691 , n62692 , n62693 , n62694 , n62695 , n62696 , 
 n62697 , n62698 , n62699 , n62700 , n62701 , n62702 , n62703 , n62704 , n62705 , n62706 , 
 n62707 , n62708 , n62709 , n62710 , n62711 , n62712 , n62713 , n62714 , n62715 , n62716 , 
 n62717 , n62718 , n62719 , n62720 , n62721 , n62722 , n62723 , n62724 , n62725 , n62726 , 
 n62727 , n62728 , n62729 , n62730 , n62731 , n62732 , n62733 , n62734 , n62735 , n62736 , 
 n62737 , n62738 , n62739 , n62740 , n62741 , n62742 , n62743 , n62744 , n62745 , n62746 , 
 n62747 , n62748 , n62749 , n62750 , n62751 , n62752 , n62753 , n62754 , n62755 , n62756 , 
 n62757 , n62758 , n62759 , n62760 , n62761 , n62762 , n62763 , n62764 , n62765 , n62766 , 
 n62767 , n62768 , n62769 , n62770 , n62771 , n62772 , n62773 , n62774 , n62775 , n62776 , 
 n62777 , n62778 , n62779 , n62780 , n62781 , n62782 , n62783 , n62784 , n62785 , n62786 , 
 n62787 , n62788 , n62789 , n62790 , n62791 , n62792 , n62793 , n62794 , n62795 , n62796 , 
 n62797 , n62798 , n62799 , n62800 , n62801 , n62802 , n62803 , n62804 , n62805 , n62806 , 
 n62807 , n62808 , n62809 , n62810 , n62811 , n62812 , n62813 , n62814 , n62815 , n62816 , 
 n62817 , n62818 , n62819 , n62820 , n62821 , n62822 , n62823 , n62824 , n62825 , n62826 , 
 n62827 , n62828 , n62829 , n62830 , n62831 , n62832 , n62833 , n62834 , n62835 , n62836 , 
 n62837 , n62838 , n62839 , n62840 , n62841 , n62842 , n62843 , n62844 , n62845 , n62846 , 
 n62847 , n62848 , n62849 , n62850 , n62851 , n62852 , n62853 , n62854 , n62855 , n62856 , 
 n62857 , n62858 , n62859 , n62860 , n62861 , n62862 , n62863 , n62864 , n62865 , n62866 , 
 n62867 , n62868 , n62869 , n62870 , n62871 , n62872 , n62873 , n62874 , n62875 , n62876 , 
 n62877 , n62878 , n62879 , n62880 , n62881 , n62882 , n62883 , n62884 , n62885 , n62886 , 
 n62887 , n62888 , n62889 , n62890 , n62891 , n62892 , n62893 , n62894 , n62895 , n62896 , 
 n62897 , n62898 , n62899 , n62900 , n62901 , n62902 , n62903 , n62904 , n62905 , n62906 , 
 n62907 , n62908 , n62909 , n62910 , n62911 , n62912 , n62913 , n62914 , n62915 , n62916 , 
 n62917 , n62918 , n62919 , n62920 , n62921 , n62922 , n62923 , n62924 , n62925 , n62926 , 
 n62927 , n62928 , n62929 , n62930 , n62931 , n62932 , n62933 , n62934 , n62935 , n62936 , 
 n62937 , n62938 , n62939 , n62940 , n62941 , n62942 , n62943 , n62944 , n62945 , n62946 , 
 n62947 , n62948 , n62949 , n62950 , n62951 , n62952 , n62953 , n62954 , n62955 , n62956 , 
 n62957 , n62958 , n62959 , n62960 , n62961 , n62962 , n62963 , n62964 , n62965 , n62966 , 
 n62967 , n62968 , n62969 , n62970 , n62971 , n62972 , n62973 , n62974 , n62975 , n62976 , 
 n62977 , n62978 , n62979 , n62980 , n62981 , n62982 , n62983 , n62984 , n62985 , n62986 , 
 n62987 , n62988 , n62989 , n62990 , n62991 , n62992 , n62993 , n62994 , n62995 , n62996 , 
 n62997 , n62998 , n62999 , n63000 , n63001 , n63002 , n63003 , n63004 , n63005 , n63006 , 
 n63007 , n63008 , n63009 , n63010 , n63011 , n63012 , n63013 , n63014 , n63015 , n63016 , 
 n63017 , n63018 , n63019 , n63020 , n63021 , n63022 , n63023 , n63024 , n63025 , n63026 , 
 n63027 , n63028 , n63029 , n63030 , n63031 , n63032 , n63033 , n63034 , n63035 , n63036 , 
 n63037 , n63038 , n63039 , n63040 , n63041 , n63042 , n63043 , n63044 , n63045 , n63046 , 
 n63047 , n63048 , n63049 , n63050 , n63051 , n63052 , n63053 , n63054 , n63055 , n63056 , 
 n63057 , n63058 , n63059 , n63060 , n63061 , n63062 , n63063 , n63064 , n63065 , n63066 , 
 n63067 , n63068 , n63069 , n63070 , n63071 , n63072 , n63073 , n63074 , n63075 , n63076 , 
 n63077 , n63078 , n63079 , n63080 , n63081 , n63082 , n63083 , n63084 , n63085 , n63086 , 
 n63087 , n63088 , n63089 , n63090 , n63091 , n63092 , n63093 , n63094 , n63095 , n63096 , 
 n63097 , n63098 , n63099 , n63100 , n63101 , n63102 , n63103 , n63104 , n63105 , n63106 , 
 n63107 , n63108 , n63109 , n63110 , n63111 , n63112 , n63113 , n63114 , n63115 , n63116 , 
 n63117 , n63118 , n63119 , n63120 , n63121 , n63122 , n63123 , n63124 , n63125 , n63126 , 
 n63127 , n63128 , n63129 , n63130 , n63131 , n63132 , n63133 , n63134 , n63135 , n63136 , 
 n63137 , n63138 , n63139 , n63140 , n63141 , n63142 , n63143 , n63144 , n63145 , n63146 , 
 n63147 , n63148 , n63149 , n63150 , n63151 , n63152 , n63153 , n63154 , n63155 , n63156 , 
 n63157 , n63158 , n63159 , n63160 , n63161 , n63162 , n63163 , n63164 , n63165 , n63166 , 
 n63167 , n63168 , n63169 , n63170 , n63171 , n63172 , n63173 , n63174 , n63175 , n63176 , 
 n63177 , n63178 , n63179 , n63180 , n63181 , n63182 , n63183 , n63184 , n63185 , n63186 , 
 n63187 , n63188 , n63189 , n63190 , n63191 , n63192 , n63193 , n63194 , n63195 , n63196 , 
 n63197 , n63198 , n63199 , n63200 , n63201 , n63202 , n63203 , n63204 , n63205 , n63206 , 
 n63207 , n63208 , n63209 , n63210 , n63211 , n63212 , n63213 , n63214 , n63215 , n63216 , 
 n63217 , n63218 , n63219 , n63220 , n63221 , n63222 , n63223 , n63224 , n63225 , n63226 , 
 n63227 , n63228 , n63229 , n63230 , n63231 , n63232 , n63233 , n63234 , n63235 , n63236 , 
 n63237 , n63238 , n63239 , n63240 , n63241 , n63242 , n63243 , n63244 , n63245 , n63246 , 
 n63247 , n63248 , n63249 , n63250 , n63251 , n63252 , n63253 , n63254 , n63255 , n63256 , 
 n63257 , n63258 , n63259 , n63260 , n63261 , n63262 , n63263 , n63264 , n63265 , n63266 , 
 n63267 , n63268 , n63269 , n63270 , n63271 , n63272 , n63273 , n63274 , n63275 , n63276 , 
 n63277 , n63278 , n63279 , n63280 , n63281 , n63282 , n63283 , n63284 , n63285 , n63286 , 
 n63287 , n63288 , n63289 , n63290 , n63291 , n63292 , n63293 , n63294 , n63295 , n63296 , 
 n63297 , n63298 , n63299 , n63300 , n63301 , n63302 , n63303 , n63304 , n63305 , n63306 , 
 n63307 , n63308 , n63309 , n63310 , n63311 , n63312 , n63313 , n63314 , n63315 , n63316 , 
 n63317 , n63318 , n63319 , n63320 , n63321 , n63322 , n63323 , n63324 , n63325 , n63326 , 
 n63327 , n63328 , n63329 , n63330 , n63331 , n63332 , n63333 , n63334 , n63335 , n63336 , 
 n63337 , n63338 , n63339 , n63340 , n63341 , n63342 , n63343 , n63344 , n63345 , n63346 , 
 n63347 , n63348 , n63349 , n63350 , n63351 , n63352 , n63353 , n63354 , n63355 , n63356 , 
 n63357 , n63358 , n63359 , n63360 , n63361 , n63362 , n63363 , n63364 , n63365 , n63366 , 
 n63367 , n63368 , n63369 , n63370 , n63371 , n63372 , n63373 , n63374 , n63375 , n63376 , 
 n63377 , n63378 , n63379 , n63380 , n63381 , n63382 , n63383 , n63384 , n63385 , n63386 , 
 n63387 , n63388 , n63389 , n63390 , n63391 , n63392 , n63393 , n63394 , n63395 , n63396 , 
 n63397 , n63398 , n63399 , n63400 , n63401 , n63402 , n63403 , n63404 , n63405 , n63406 , 
 n63407 , n63408 , n63409 , n63410 , n63411 , n63412 , n63413 , n63414 , n63415 , n63416 , 
 n63417 , n63418 , n63419 , n63420 , n63421 , n63422 , n63423 , n63424 , n63425 , n63426 , 
 n63427 , n63428 , n63429 , n63430 , n63431 , n63432 , n63433 , n63434 , n63435 , n63436 , 
 n63437 , n63438 , n63439 , n63440 , n63441 , n63442 , n63443 , n63444 , n63445 , n63446 , 
 n63447 , n63448 , n63449 , n63450 , n63451 , n63452 , n63453 , n63454 , n63455 , n63456 , 
 n63457 , n63458 , n63459 , n63460 , n63461 , n63462 , n63463 , n63464 , n63465 , n63466 , 
 n63467 , n63468 , n63469 , n63470 , n63471 , n63472 , n63473 , n63474 , n63475 , n63476 , 
 n63477 , n63478 , n63479 , n63480 , n63481 , n63482 , n63483 , n63484 , n63485 , n63486 , 
 n63487 , n63488 , n63489 , n63490 , n63491 , n63492 , n63493 , n63494 , n63495 , n63496 , 
 n63497 , n63498 , n63499 , n63500 , n63501 , n63502 , n63503 , n63504 , n63505 , n63506 , 
 n63507 , n63508 , n63509 , n63510 , n63511 , n63512 , n63513 , n63514 , n63515 , n63516 , 
 n63517 , n63518 , n63519 , n63520 , n63521 , n63522 , n63523 , n63524 , n63525 , n63526 , 
 n63527 , n63528 , n63529 , n63530 , n63531 , n63532 , n63533 , n63534 , n63535 , n63536 , 
 n63537 , n63538 , n63539 , n63540 , n63541 , n63542 , n63543 , n63544 , n63545 , n63546 , 
 n63547 , n63548 , n63549 , n63550 , n63551 , n63552 , n63553 , n63554 , n63555 , n63556 , 
 n63557 , n63558 , n63559 , n63560 , n63561 , n63562 , n63563 , n63564 , n63565 , n63566 , 
 n63567 , n63568 , n63569 , n63570 , n63571 , n63572 , n63573 , n63574 , n63575 , n63576 , 
 n63577 , n63578 , n63579 , n63580 , n63581 , n63582 , n63583 , n63584 , n63585 , n63586 , 
 n63587 , n63588 , n63589 , n63590 , n63591 , n63592 , n63593 , n63594 , n63595 , n63596 , 
 n63597 , n63598 , n63599 , n63600 , n63601 , n63602 , n63603 , n63604 , n63605 , n63606 , 
 n63607 , n63608 , n63609 , n63610 , n63611 , n63612 , n63613 , n63614 , n63615 , n63616 , 
 n63617 , n63618 , n63619 , n63620 , n63621 , n63622 , n63623 , n63624 , n63625 , n63626 , 
 n63627 , n63628 , n63629 , n63630 , n63631 , n63632 , n63633 , n63634 , n63635 , n63636 , 
 n63637 , n63638 , n63639 , n63640 , n63641 , n63642 , n63643 , n63644 , n63645 , n63646 , 
 n63647 , n63648 , n63649 , n63650 , n63651 , n63652 , n63653 , n63654 , n63655 , n63656 , 
 n63657 , n63658 , n63659 , n63660 , n63661 , n63662 , n63663 , n63664 , n63665 , n63666 , 
 n63667 , n63668 , n63669 , n63670 , n63671 , n63672 , n63673 , n63674 , n63675 , n63676 , 
 n63677 , n63678 , n63679 , n63680 , n63681 , n63682 , n63683 , n63684 , n63685 , n63686 , 
 n63687 , n63688 , n63689 , n63690 , n63691 , n63692 , n63693 , n63694 , n63695 , n63696 , 
 n63697 , n63698 , n63699 , n63700 , n63701 , n63702 , n63703 , n63704 , n63705 , n63706 , 
 n63707 , n63708 , n63709 , n63710 , n63711 , n63712 , n63713 , n63714 , n63715 , n63716 , 
 n63717 , n63718 , n63719 , n63720 , n63721 , n63722 , n63723 , n63724 , n63725 , n63726 , 
 n63727 , n63728 , n63729 , n63730 , n63731 , n63732 , n63733 , n63734 , n63735 , n63736 , 
 n63737 , n63738 , n63739 , n63740 , n63741 , n63742 , n63743 , n63744 , n63745 , n63746 , 
 n63747 , n63748 , n63749 , n63750 , n63751 , n63752 , n63753 , n63754 , n63755 , n63756 , 
 n63757 , n63758 , n63759 , n63760 , n63761 , n63762 , n63763 , n63764 , n63765 , n63766 , 
 n63767 , n63768 , n63769 , n63770 , n63771 , n63772 , n63773 , n63774 , n63775 , n63776 , 
 n63777 , n63778 , n63779 , n63780 , n63781 , n63782 , n63783 , n63784 , n63785 , n63786 , 
 n63787 , n63788 , n63789 , n63790 , n63791 , n63792 , n63793 , n63794 , n63795 , n63796 , 
 n63797 , n63798 , n63799 , n63800 , n63801 , n63802 , n63803 , n63804 , n63805 , n63806 , 
 n63807 , n63808 , n63809 , n63810 , n63811 , n63812 , n63813 , n63814 , n63815 , n63816 , 
 n63817 , n63818 , n63819 , n63820 , n63821 , n63822 , n63823 , n63824 , n63825 , n63826 , 
 n63827 , n63828 , n63829 , n63830 , n63831 , n63832 , n63833 , n63834 , n63835 , n63836 , 
 n63837 , n63838 , n63839 , n63840 , n63841 , n63842 , n63843 , n63844 , n63845 , n63846 , 
 n63847 , n63848 , n63849 , n63850 , n63851 , n63852 , n63853 , n63854 , n63855 , n63856 , 
 n63857 , n63858 , n63859 , n63860 , n63861 , n63862 , n63863 , n63864 , n63865 , n63866 , 
 n63867 , n63868 , n63869 , n63870 , n63871 , n63872 , n63873 , n63874 , n63875 , n63876 , 
 n63877 , n63878 , n63879 , n63880 , n63881 , n63882 , n63883 , n63884 , n63885 , n63886 , 
 n63887 , n63888 , n63889 , n63890 , n63891 , n63892 , n63893 , n63894 , n63895 , n63896 , 
 n63897 , n63898 , n63899 , n63900 , n63901 , n63902 , n63903 , n63904 , n63905 , n63906 , 
 n63907 , n63908 , n63909 , n63910 , n63911 , n63912 , n63913 , n63914 , n63915 , n63916 , 
 n63917 , n63918 , n63919 , n63920 , n63921 , n63922 , n63923 , n63924 , n63925 , n63926 , 
 n63927 , n63928 , n63929 , n63930 , n63931 , n63932 , n63933 , n63934 , n63935 , n63936 , 
 n63937 , n63938 , n63939 , n63940 , n63941 , n63942 , n63943 , n63944 , n63945 , n63946 , 
 n63947 , n63948 , n63949 , n63950 , n63951 , n63952 , n63953 , n63954 , n63955 , n63956 , 
 n63957 , n63958 , n63959 , n63960 , n63961 , n63962 , n63963 , n63964 , n63965 , n63966 , 
 n63967 , n63968 , n63969 , n63970 , n63971 , n63972 , n63973 , n63974 , n63975 , n63976 , 
 n63977 , n63978 , n63979 , n63980 , n63981 , n63982 , n63983 , n63984 , n63985 , n63986 , 
 n63987 , n63988 , n63989 , n63990 , n63991 , n63992 , n63993 , n63994 , n63995 , n63996 , 
 n63997 , n63998 , n63999 , n64000 , n64001 , n64002 , n64003 , n64004 , n64005 , n64006 , 
 n64007 , n64008 , n64009 , n64010 , n64011 , n64012 , n64013 , n64014 , n64015 , n64016 , 
 n64017 , n64018 , n64019 , n64020 , n64021 , n64022 , n64023 , n64024 , n64025 , n64026 , 
 n64027 , n64028 , n64029 , n64030 , n64031 , n64032 , n64033 , n64034 , n64035 , n64036 , 
 n64037 , n64038 , n64039 , n64040 , n64041 , n64042 , n64043 , n64044 , n64045 , n64046 , 
 n64047 , n64048 , n64049 , n64050 , n64051 , n64052 , n64053 , n64054 , n64055 , n64056 , 
 n64057 , n64058 , n64059 , n64060 , n64061 , n64062 , n64063 , n64064 , n64065 , n64066 , 
 n64067 , n64068 , n64069 , n64070 , n64071 , n64072 , n64073 , n64074 , n64075 , n64076 , 
 n64077 , n64078 , n64079 , n64080 , n64081 , n64082 , n64083 , n64084 , n64085 , n64086 , 
 n64087 , n64088 , n64089 , n64090 , n64091 , n64092 , n64093 , n64094 , n64095 , n64096 , 
 n64097 , n64098 , n64099 , n64100 , n64101 , n64102 , n64103 , n64104 , n64105 , n64106 , 
 n64107 , n64108 , n64109 , n64110 , n64111 , n64112 , n64113 , n64114 , n64115 , n64116 , 
 n64117 , n64118 , n64119 , n64120 , n64121 , n64122 , n64123 , n64124 , n64125 , n64126 , 
 n64127 , n64128 , n64129 , n64130 , n64131 , n64132 , n64133 , n64134 , n64135 , n64136 , 
 n64137 , n64138 , n64139 , n64140 , n64141 , n64142 , n64143 , n64144 , n64145 , n64146 , 
 n64147 , n64148 , n64149 , n64150 , n64151 , n64152 , n64153 , n64154 , n64155 , n64156 , 
 n64157 , n64158 , n64159 , n64160 , n64161 , n64162 , n64163 , n64164 , n64165 , n64166 , 
 n64167 , n64168 , n64169 , n64170 , n64171 , n64172 , n64173 , n64174 , n64175 , n64176 , 
 n64177 , n64178 , n64179 , n64180 , n64181 , n64182 , n64183 , n64184 , n64185 , n64186 , 
 n64187 , n64188 , n64189 , n64190 , n64191 , n64192 , n64193 , n64194 , n64195 , n64196 , 
 n64197 , n64198 , n64199 , n64200 , n64201 , n64202 , n64203 , n64204 , n64205 , n64206 , 
 n64207 , n64208 , n64209 , n64210 , n64211 , n64212 , n64213 , n64214 , n64215 , n64216 , 
 n64217 , n64218 , n64219 , n64220 , n64221 , n64222 , n64223 , n64224 , n64225 , n64226 , 
 n64227 , n64228 , n64229 , n64230 , n64231 , n64232 , n64233 , n64234 , n64235 , n64236 , 
 n64237 , n64238 , n64239 , n64240 , n64241 , n64242 , n64243 , n64244 , n64245 , n64246 , 
 n64247 , n64248 , n64249 , n64250 , n64251 , n64252 , n64253 , n64254 , n64255 , n64256 , 
 n64257 , n64258 , n64259 , n64260 , n64261 , n64262 , n64263 , n64264 , n64265 , n64266 , 
 n64267 , n64268 , n64269 , n64270 , n64271 , n64272 , n64273 , n64274 , n64275 , n64276 , 
 n64277 , n64278 , n64279 , n64280 , n64281 , n64282 , n64283 , n64284 , n64285 , n64286 , 
 n64287 , n64288 , n64289 , n64290 , n64291 , n64292 , n64293 , n64294 , n64295 , n64296 , 
 n64297 , n64298 , n64299 , n64300 , n64301 , n64302 , n64303 , n64304 , n64305 , n64306 , 
 n64307 , n64308 , n64309 , n64310 , n64311 , n64312 , n64313 , n64314 , n64315 , n64316 , 
 n64317 , n64318 , n64319 , n64320 , n64321 , n64322 , n64323 , n64324 , n64325 , n64326 , 
 n64327 , n64328 , n64329 , n64330 , n64331 , n64332 , n64333 , n64334 , n64335 , n64336 , 
 n64337 , n64338 , n64339 , n64340 , n64341 , n64342 , n64343 , n64344 , n64345 , n64346 , 
 n64347 , n64348 , n64349 , n64350 , n64351 , n64352 , n64353 , n64354 , n64355 , n64356 , 
 n64357 , n64358 , n64359 , n64360 , n64361 , n64362 , n64363 , n64364 , n64365 , n64366 , 
 n64367 , n64368 , n64369 , n64370 , n64371 , n64372 , n64373 , n64374 , n64375 , n64376 , 
 n64377 , n64378 , n64379 , n64380 , n64381 , n64382 , n64383 , n64384 , n64385 , n64386 , 
 n64387 , n64388 , n64389 , n64390 , n64391 , n64392 , n64393 , n64394 , n64395 , n64396 , 
 n64397 , n64398 , n64399 , n64400 , n64401 , n64402 , n64403 , n64404 , n64405 , n64406 , 
 n64407 , n64408 , n64409 , n64410 , n64411 , n64412 , n64413 , n64414 , n64415 , n64416 , 
 n64417 , n64418 , n64419 , n64420 , n64421 , n64422 , n64423 , n64424 , n64425 , n64426 , 
 n64427 , n64428 , n64429 , n64430 , n64431 , n64432 , n64433 , n64434 , n64435 , n64436 , 
 n64437 , n64438 , n64439 , n64440 , n64441 , n64442 , n64443 , n64444 , n64445 , n64446 , 
 n64447 , n64448 , n64449 , n64450 , n64451 , n64452 , n64453 , n64454 , n64455 , n64456 , 
 n64457 , n64458 , n64459 , n64460 , n64461 , n64462 , n64463 , n64464 , n64465 , n64466 , 
 n64467 , n64468 , n64469 , n64470 , n64471 , n64472 , n64473 , n64474 , n64475 , n64476 , 
 n64477 , n64478 , n64479 , n64480 , n64481 , n64482 , n64483 , n64484 , n64485 , n64486 , 
 n64487 , n64488 , n64489 , n64490 , n64491 , n64492 , n64493 , n64494 , n64495 , n64496 , 
 n64497 , n64498 , n64499 , n64500 , n64501 , n64502 , n64503 , n64504 , n64505 , n64506 , 
 n64507 , n64508 , n64509 , n64510 , n64511 , n64512 , n64513 , n64514 , n64515 , n64516 , 
 n64517 , n64518 , n64519 , n64520 , n64521 , n64522 , n64523 , n64524 , n64525 , n64526 , 
 n64527 , n64528 , n64529 , n64530 , n64531 , n64532 , n64533 , n64534 , n64535 , n64536 , 
 n64537 , n64538 , n64539 , n64540 , n64541 , n64542 , n64543 , n64544 , n64545 , n64546 , 
 n64547 , n64548 , n64549 , n64550 , n64551 , n64552 , n64553 , n64554 , n64555 , n64556 , 
 n64557 , n64558 , n64559 , n64560 , n64561 , n64562 , n64563 , n64564 , n64565 , n64566 , 
 n64567 , n64568 , n64569 , n64570 , n64571 , n64572 , n64573 , n64574 , n64575 , n64576 , 
 n64577 , n64578 , n64579 , n64580 , n64581 , n64582 , n64583 , n64584 , n64585 , n64586 , 
 n64587 , n64588 , n64589 , n64590 , n64591 , n64592 , n64593 , n64594 , n64595 , n64596 , 
 n64597 , n64598 , n64599 , n64600 , n64601 , n64602 , n64603 , n64604 , n64605 , n64606 , 
 n64607 , n64608 , n64609 , n64610 , n64611 , n64612 , n64613 , n64614 , n64615 , n64616 , 
 n64617 , n64618 , n64619 , n64620 , n64621 , n64622 , n64623 , n64624 , n64625 , n64626 , 
 n64627 , n64628 , n64629 , n64630 , n64631 , n64632 , n64633 , n64634 , n64635 , n64636 , 
 n64637 , n64638 , n64639 , n64640 , n64641 , n64642 , n64643 , n64644 , n64645 , n64646 , 
 n64647 , n64648 , n64649 , n64650 , n64651 , n64652 , n64653 , n64654 , n64655 , n64656 , 
 n64657 , n64658 , n64659 , n64660 , n64661 , n64662 , n64663 , n64664 , n64665 , n64666 , 
 n64667 , n64668 , n64669 , n64670 , n64671 , n64672 , n64673 , n64674 , n64675 , n64676 , 
 n64677 , n64678 , n64679 , n64680 , n64681 , n64682 , n64683 , n64684 , n64685 , n64686 , 
 n64687 , n64688 , n64689 , n64690 , n64691 , n64692 , n64693 , n64694 , n64695 , n64696 , 
 n64697 , n64698 , n64699 , n64700 , n64701 , n64702 , n64703 , n64704 , n64705 , n64706 , 
 n64707 , n64708 , n64709 , n64710 , n64711 , n64712 , n64713 , n64714 , n64715 , n64716 , 
 n64717 , n64718 , n64719 , n64720 , n64721 , n64722 , n64723 , n64724 , n64725 , n64726 , 
 n64727 , n64728 , n64729 , n64730 , n64731 , n64732 , n64733 , n64734 , n64735 , n64736 , 
 n64737 , n64738 , n64739 , n64740 , n64741 , n64742 , n64743 , n64744 , n64745 , n64746 , 
 n64747 , n64748 , n64749 , n64750 , n64751 , n64752 , n64753 , n64754 , n64755 , n64756 , 
 n64757 , n64758 , n64759 , n64760 , n64761 , n64762 , n64763 , n64764 , n64765 , n64766 , 
 n64767 , n64768 , n64769 , n64770 , n64771 , n64772 , n64773 , n64774 , n64775 , n64776 , 
 n64777 , n64778 , n64779 , n64780 , n64781 , n64782 , n64783 , n64784 , n64785 , n64786 , 
 n64787 , n64788 , n64789 , n64790 , n64791 , n64792 , n64793 , n64794 , n64795 , n64796 , 
 n64797 , n64798 , n64799 , n64800 , n64801 , n64802 , n64803 , n64804 , n64805 , n64806 , 
 n64807 , n64808 , n64809 , n64810 , n64811 , n64812 , n64813 , n64814 , n64815 , n64816 , 
 n64817 , n64818 , n64819 , n64820 , n64821 , n64822 , n64823 , n64824 , n64825 , n64826 , 
 n64827 , n64828 , n64829 , n64830 , n64831 , n64832 , n64833 , n64834 , n64835 , n64836 , 
 n64837 , n64838 , n64839 , n64840 , n64841 , n64842 , n64843 , n64844 , n64845 , n64846 , 
 n64847 , n64848 , n64849 , n64850 , n64851 , n64852 , n64853 , n64854 , n64855 , n64856 , 
 n64857 , n64858 , n64859 , n64860 , n64861 , n64862 , n64863 , n64864 , n64865 , n64866 , 
 n64867 , n64868 , n64869 , n64870 , n64871 , n64872 , n64873 , n64874 , n64875 , n64876 , 
 n64877 , n64878 , n64879 , n64880 , n64881 , n64882 , n64883 , n64884 , n64885 , n64886 , 
 n64887 , n64888 , n64889 , n64890 , n64891 , n64892 , n64893 , n64894 , n64895 , n64896 , 
 n64897 , n64898 , n64899 , n64900 , n64901 , n64902 , n64903 , n64904 , n64905 , n64906 , 
 n64907 , n64908 , n64909 , n64910 , n64911 , n64912 , n64913 , n64914 , n64915 , n64916 , 
 n64917 , n64918 , n64919 , n64920 , n64921 , n64922 , n64923 , n64924 , n64925 , n64926 , 
 n64927 , n64928 , n64929 , n64930 , n64931 , n64932 , n64933 , n64934 , n64935 , n64936 , 
 n64937 , n64938 , n64939 , n64940 , n64941 , n64942 , n64943 , n64944 , n64945 , n64946 , 
 n64947 , n64948 , n64949 , n64950 , n64951 , n64952 , n64953 , n64954 , n64955 , n64956 , 
 n64957 , n64958 , n64959 , n64960 , n64961 , n64962 , n64963 , n64964 , n64965 , n64966 , 
 n64967 , n64968 , n64969 , n64970 , n64971 , n64972 , n64973 , n64974 , n64975 , n64976 , 
 n64977 , n64978 , n64979 , n64980 , n64981 , n64982 , n64983 , n64984 , n64985 , n64986 , 
 n64987 , n64988 , n64989 , n64990 , n64991 , n64992 , n64993 , n64994 , n64995 , n64996 , 
 n64997 , n64998 , n64999 , n65000 , n65001 , n65002 , n65003 , n65004 , n65005 , n65006 , 
 n65007 , n65008 , n65009 , n65010 , n65011 , n65012 , n65013 , n65014 , n65015 , n65016 , 
 n65017 , n65018 , n65019 , n65020 , n65021 , n65022 , n65023 , n65024 , n65025 , n65026 , 
 n65027 , n65028 , n65029 , n65030 , n65031 , n65032 , n65033 , n65034 , n65035 , n65036 , 
 n65037 , n65038 , n65039 , n65040 , n65041 , n65042 , n65043 , n65044 , n65045 , n65046 , 
 n65047 , n65048 , n65049 , n65050 , n65051 , n65052 , n65053 , n65054 , n65055 , n65056 , 
 n65057 , n65058 , n65059 , n65060 , n65061 , n65062 , n65063 , n65064 , n65065 , n65066 , 
 n65067 , n65068 , n65069 , n65070 , n65071 , n65072 , n65073 , n65074 , n65075 , n65076 , 
 n65077 , n65078 , n65079 , n65080 , n65081 , n65082 , n65083 , n65084 , n65085 , n65086 , 
 n65087 , n65088 , n65089 , n65090 , n65091 , n65092 , n65093 , n65094 , n65095 , n65096 , 
 n65097 , n65098 , n65099 , n65100 , n65101 , n65102 , n65103 , n65104 , n65105 , n65106 , 
 n65107 , n65108 , n65109 , n65110 , n65111 , n65112 , n65113 , n65114 , n65115 , n65116 , 
 n65117 , n65118 , n65119 , n65120 , n65121 , n65122 , n65123 , n65124 , n65125 , n65126 , 
 n65127 , n65128 , n65129 , n65130 , n65131 , n65132 , n65133 , n65134 , n65135 , n65136 , 
 n65137 , n65138 , n65139 , n65140 , n65141 , n65142 , n65143 , n65144 , n65145 , n65146 , 
 n65147 , n65148 , n65149 , n65150 , n65151 , n65152 , n65153 , n65154 , n65155 , n65156 , 
 n65157 , n65158 , n65159 , n65160 , n65161 , n65162 , n65163 , n65164 , n65165 , n65166 , 
 n65167 , n65168 , n65169 , n65170 , n65171 , n65172 , n65173 , n65174 , n65175 , n65176 , 
 n65177 , n65178 , n65179 , n65180 , n65181 , n65182 , n65183 , n65184 , n65185 , n65186 , 
 n65187 , n65188 , n65189 , n65190 , n65191 , n65192 , n65193 , n65194 , n65195 , n65196 , 
 n65197 , n65198 , n65199 , n65200 , n65201 , n65202 , n65203 , n65204 , n65205 , n65206 , 
 n65207 , n65208 , n65209 , n65210 , n65211 , n65212 , n65213 , n65214 , n65215 , n65216 , 
 n65217 , n65218 , n65219 , n65220 , n65221 , n65222 , n65223 , n65224 , n65225 , n65226 , 
 n65227 , n65228 , n65229 , n65230 , n65231 , n65232 , n65233 , n65234 , n65235 , n65236 , 
 n65237 , n65238 , n65239 , n65240 , n65241 , n65242 , n65243 , n65244 , n65245 , n65246 , 
 n65247 , n65248 , n65249 , n65250 , n65251 , n65252 , n65253 , n65254 , n65255 , n65256 , 
 n65257 , n65258 , n65259 , n65260 , n65261 , n65262 , n65263 , n65264 , n65265 , n65266 , 
 n65267 , n65268 , n65269 , n65270 , n65271 , n65272 , n65273 , n65274 , n65275 , n65276 , 
 n65277 , n65278 , n65279 , n65280 , n65281 , n65282 , n65283 , n65284 , n65285 , n65286 , 
 n65287 , n65288 , n65289 , n65290 , n65291 , n65292 , n65293 , n65294 , n65295 , n65296 , 
 n65297 , n65298 , n65299 , n65300 , n65301 , n65302 , n65303 , n65304 , n65305 , n65306 , 
 n65307 , n65308 , n65309 , n65310 , n65311 , n65312 , n65313 , n65314 , n65315 , n65316 , 
 n65317 , n65318 , n65319 , n65320 , n65321 , n65322 , n65323 , n65324 , n65325 , n65326 , 
 n65327 , n65328 , n65329 , n65330 , n65331 , n65332 , n65333 , n65334 , n65335 , n65336 , 
 n65337 , n65338 , n65339 , n65340 , n65341 , n65342 , n65343 , n65344 , n65345 , n65346 , 
 n65347 , n65348 , n65349 , n65350 , n65351 , n65352 , n65353 , n65354 , n65355 , n65356 , 
 n65357 , n65358 , n65359 , n65360 , n65361 , n65362 , n65363 , n65364 , n65365 , n65366 , 
 n65367 , n65368 , n65369 , n65370 , n65371 , n65372 , n65373 , n65374 , n65375 , n65376 , 
 n65377 , n65378 , n65379 , n65380 , n65381 , n65382 , n65383 , n65384 , n65385 , n65386 , 
 n65387 , n65388 , n65389 , n65390 , n65391 , n65392 , n65393 , n65394 , n65395 , n65396 , 
 n65397 , n65398 , n65399 , n65400 , n65401 , n65402 , n65403 , n65404 , n65405 , n65406 , 
 n65407 , n65408 , n65409 , n65410 , n65411 , n65412 , n65413 , n65414 , n65415 , n65416 , 
 n65417 , n65418 , n65419 , n65420 , n65421 , n65422 , n65423 , n65424 , n65425 , n65426 , 
 n65427 , n65428 , n65429 , n65430 , n65431 , n65432 , n65433 , n65434 , n65435 , n65436 , 
 n65437 , n65438 , n65439 , n65440 , n65441 , n65442 , n65443 , n65444 , n65445 , n65446 , 
 n65447 , n65448 , n65449 , n65450 , n65451 , n65452 , n65453 , n65454 , n65455 , n65456 , 
 n65457 , n65458 , n65459 , n65460 , n65461 , n65462 , n65463 , n65464 , n65465 , n65466 , 
 n65467 , n65468 , n65469 , n65470 , n65471 , n65472 , n65473 , n65474 , n65475 , n65476 , 
 n65477 , n65478 , n65479 , n65480 , n65481 , n65482 , n65483 , n65484 , n65485 , n65486 , 
 n65487 , n65488 , n65489 , n65490 , n65491 , n65492 , n65493 , n65494 , n65495 , n65496 , 
 n65497 , n65498 , n65499 , n65500 , n65501 , n65502 , n65503 , n65504 , n65505 , n65506 , 
 n65507 , n65508 , n65509 , n65510 , n65511 , n65512 , n65513 , n65514 , n65515 , n65516 , 
 n65517 , n65518 , n65519 , n65520 , n65521 , n65522 , n65523 , n65524 , n65525 , n65526 , 
 n65527 , n65528 , n65529 , n65530 , n65531 , n65532 , n65533 , n65534 , n65535 , n65536 , 
 n65537 , n65538 , n65539 , n65540 , n65541 , n65542 , n65543 , n65544 , n65545 , n65546 , 
 n65547 , n65548 , n65549 , n65550 , n65551 , n65552 , n65553 , n65554 , n65555 , n65556 , 
 n65557 , n65558 , n65559 , n65560 , n65561 , n65562 , n65563 , n65564 , n65565 , n65566 , 
 n65567 , n65568 , n65569 , n65570 , n65571 , n65572 , n65573 , n65574 , n65575 , n65576 , 
 n65577 , n65578 , n65579 , n65580 , n65581 , n65582 , n65583 , n65584 , n65585 , n65586 , 
 n65587 , n65588 , n65589 , n65590 , n65591 , n65592 , n65593 , n65594 , n65595 , n65596 , 
 n65597 , n65598 , n65599 , n65600 , n65601 , n65602 , n65603 , n65604 , n65605 , n65606 , 
 n65607 , n65608 , n65609 , n65610 , n65611 , n65612 , n65613 , n65614 , n65615 , n65616 , 
 n65617 , n65618 , n65619 , n65620 , n65621 , n65622 , n65623 , n65624 , n65625 , n65626 , 
 n65627 , n65628 , n65629 , n65630 , n65631 , n65632 , n65633 , n65634 , n65635 , n65636 , 
 n65637 , n65638 , n65639 , n65640 , n65641 , n65642 , n65643 , n65644 , n65645 , n65646 , 
 n65647 , n65648 , n65649 , n65650 , n65651 , n65652 , n65653 , n65654 , n65655 , n65656 , 
 n65657 , n65658 , n65659 , n65660 , n65661 , n65662 , n65663 , n65664 , n65665 , n65666 , 
 n65667 , n65668 , n65669 , n65670 , n65671 , n65672 , n65673 , n65674 , n65675 , n65676 , 
 n65677 , n65678 , n65679 , n65680 , n65681 , n65682 , n65683 , n65684 , n65685 , n65686 , 
 n65687 , n65688 , n65689 , n65690 , n65691 , n65692 , n65693 , n65694 , n65695 , n65696 , 
 n65697 , n65698 , n65699 , n65700 , n65701 , n65702 , n65703 , n65704 , n65705 , n65706 , 
 n65707 , n65708 , n65709 , n65710 , n65711 , n65712 , n65713 , n65714 , n65715 , n65716 , 
 n65717 , n65718 , n65719 , n65720 , n65721 , n65722 , n65723 , n65724 , n65725 , n65726 , 
 n65727 , n65728 , n65729 , n65730 , n65731 , n65732 , n65733 , n65734 , n65735 , n65736 , 
 n65737 , n65738 , n65739 , n65740 , n65741 , n65742 , n65743 , n65744 , n65745 , n65746 , 
 n65747 , n65748 , n65749 , n65750 , n65751 , n65752 , n65753 , n65754 , n65755 , n65756 , 
 n65757 , n65758 , n65759 , n65760 , n65761 , n65762 , n65763 , n65764 , n65765 , n65766 , 
 n65767 , n65768 , n65769 , n65770 , n65771 , n65772 , n65773 , n65774 , n65775 , n65776 , 
 n65777 , n65778 , n65779 , n65780 , n65781 , n65782 , n65783 , n65784 , n65785 , n65786 , 
 n65787 , n65788 , n65789 , n65790 , n65791 , n65792 , n65793 , n65794 , n65795 , n65796 , 
 n65797 , n65798 , n65799 , n65800 , n65801 , n65802 , n65803 , n65804 , n65805 , n65806 , 
 n65807 , n65808 , n65809 , n65810 , n65811 , n65812 , n65813 , n65814 , n65815 , n65816 , 
 n65817 , n65818 , n65819 , n65820 , n65821 , n65822 , n65823 , n65824 , n65825 , n65826 , 
 n65827 , n65828 , n65829 , n65830 , n65831 , n65832 , n65833 , n65834 , n65835 , n65836 , 
 n65837 , n65838 , n65839 , n65840 , n65841 , n65842 , n65843 , n65844 , n65845 , n65846 , 
 n65847 , n65848 , n65849 , n65850 , n65851 , n65852 , n65853 , n65854 , n65855 , n65856 , 
 n65857 , n65858 , n65859 , n65860 , n65861 , n65862 , n65863 , n65864 , n65865 , n65866 , 
 n65867 , n65868 , n65869 , n65870 , n65871 , n65872 , n65873 , n65874 , n65875 , n65876 , 
 n65877 , n65878 , n65879 , n65880 , n65881 , n65882 , n65883 , n65884 , n65885 , n65886 , 
 n65887 , n65888 , n65889 , n65890 , n65891 , n65892 , n65893 , n65894 , n65895 , n65896 , 
 n65897 , n65898 , n65899 , n65900 , n65901 , n65902 , n65903 , n65904 , n65905 , n65906 , 
 n65907 , n65908 , n65909 , n65910 , n65911 , n65912 , n65913 , n65914 , n65915 , n65916 , 
 n65917 , n65918 , n65919 , n65920 , n65921 , n65922 , n65923 , n65924 , n65925 , n65926 , 
 n65927 , n65928 , n65929 , n65930 , n65931 , n65932 , n65933 , n65934 , n65935 , n65936 , 
 n65937 , n65938 , n65939 , n65940 , n65941 , n65942 , n65943 , n65944 , n65945 , n65946 , 
 n65947 , n65948 , n65949 , n65950 , n65951 , n65952 , n65953 , n65954 , n65955 , n65956 , 
 n65957 , n65958 , n65959 , n65960 , n65961 , n65962 , n65963 , n65964 , n65965 , n65966 , 
 n65967 , n65968 , n65969 , n65970 , n65971 , n65972 , n65973 , n65974 , n65975 , n65976 , 
 n65977 , n65978 , n65979 , n65980 , n65981 , n65982 , n65983 , n65984 , n65985 , n65986 , 
 n65987 , n65988 , n65989 , n65990 , n65991 , n65992 , n65993 , n65994 , n65995 , n65996 , 
 n65997 , n65998 , n65999 , n66000 , n66001 , n66002 , n66003 , n66004 , n66005 , n66006 , 
 n66007 , n66008 , n66009 , n66010 , n66011 , n66012 , n66013 , n66014 , n66015 , n66016 , 
 n66017 , n66018 , n66019 , n66020 , n66021 , n66022 , n66023 , n66024 , n66025 , n66026 , 
 n66027 , n66028 , n66029 , n66030 , n66031 , n66032 , n66033 , n66034 , n66035 , n66036 , 
 n66037 , n66038 , n66039 , n66040 , n66041 , n66042 , n66043 , n66044 , n66045 , n66046 , 
 n66047 , n66048 , n66049 , n66050 , n66051 , n66052 , n66053 , n66054 , n66055 , n66056 , 
 n66057 , n66058 , n66059 , n66060 , n66061 , n66062 , n66063 , n66064 , n66065 , n66066 , 
 n66067 , n66068 , n66069 , n66070 , n66071 , n66072 , n66073 , n66074 , n66075 , n66076 , 
 n66077 , n66078 , n66079 , n66080 , n66081 , n66082 , n66083 , n66084 , n66085 , n66086 , 
 n66087 , n66088 , n66089 , n66090 , n66091 , n66092 , n66093 , n66094 , n66095 , n66096 , 
 n66097 , n66098 , n66099 , n66100 , n66101 , n66102 , n66103 , n66104 , n66105 , n66106 , 
 n66107 , n66108 , n66109 , n66110 , n66111 , n66112 , n66113 , n66114 , n66115 , n66116 , 
 n66117 , n66118 , n66119 , n66120 , n66121 , n66122 , n66123 , n66124 , n66125 , n66126 , 
 n66127 , n66128 , n66129 , n66130 , n66131 , n66132 , n66133 , n66134 , n66135 , n66136 , 
 n66137 , n66138 , n66139 , n66140 , n66141 , n66142 , n66143 , n66144 , n66145 , n66146 , 
 n66147 , n66148 , n66149 , n66150 , n66151 , n66152 , n66153 , n66154 , n66155 , n66156 , 
 n66157 , n66158 , n66159 , n66160 , n66161 , n66162 , n66163 , n66164 , n66165 , n66166 , 
 n66167 , n66168 , n66169 , n66170 , n66171 , n66172 , n66173 , n66174 , n66175 , n66176 , 
 n66177 , n66178 , n66179 , n66180 , n66181 , n66182 , n66183 , n66184 , n66185 , n66186 , 
 n66187 , n66188 , n66189 , n66190 , n66191 , n66192 , n66193 , n66194 , n66195 , n66196 , 
 n66197 , n66198 , n66199 , n66200 , n66201 , n66202 , n66203 , n66204 , n66205 , n66206 , 
 n66207 , n66208 , n66209 , n66210 , n66211 , n66212 , n66213 , n66214 , n66215 , n66216 , 
 n66217 , n66218 , n66219 , n66220 , n66221 , n66222 , n66223 , n66224 , n66225 , n66226 , 
 n66227 , n66228 , n66229 , n66230 , n66231 , n66232 , n66233 , n66234 , n66235 , n66236 , 
 n66237 , n66238 , n66239 , n66240 , n66241 , n66242 , n66243 , n66244 , n66245 , n66246 , 
 n66247 , n66248 , n66249 , n66250 , n66251 , n66252 , n66253 , n66254 , n66255 , n66256 , 
 n66257 , n66258 , n66259 , n66260 , n66261 , n66262 , n66263 , n66264 , n66265 , n66266 , 
 n66267 , n66268 , n66269 , n66270 , n66271 , n66272 , n66273 , n66274 , n66275 , n66276 , 
 n66277 , n66278 , n66279 , n66280 , n66281 , n66282 , n66283 , n66284 , n66285 , n66286 , 
 n66287 , n66288 , n66289 , n66290 , n66291 , n66292 , n66293 , n66294 , n66295 , n66296 , 
 n66297 , n66298 , n66299 , n66300 , n66301 , n66302 , n66303 , n66304 , n66305 , n66306 , 
 n66307 , n66308 , n66309 , n66310 , n66311 , n66312 , n66313 , n66314 , n66315 , n66316 , 
 n66317 , n66318 , n66319 , n66320 , n66321 , n66322 , n66323 , n66324 , n66325 , n66326 , 
 n66327 , n66328 , n66329 , n66330 , n66331 , n66332 , n66333 , n66334 , n66335 , n66336 , 
 n66337 , n66338 , n66339 , n66340 , n66341 , n66342 , n66343 , n66344 , n66345 , n66346 , 
 n66347 , n66348 , n66349 , n66350 , n66351 , n66352 , n66353 , n66354 , n66355 , n66356 , 
 n66357 , n66358 , n66359 , n66360 , n66361 , n66362 , n66363 , n66364 , n66365 , n66366 , 
 n66367 , n66368 , n66369 , n66370 , n66371 , n66372 , n66373 , n66374 , n66375 , n66376 , 
 n66377 , n66378 , n66379 , n66380 , n66381 , n66382 , n66383 , n66384 , n66385 , n66386 , 
 n66387 , n66388 , n66389 , n66390 , n66391 , n66392 , n66393 , n66394 , n66395 , n66396 , 
 n66397 , n66398 , n66399 , n66400 , n66401 , n66402 , n66403 , n66404 , n66405 , n66406 , 
 n66407 , n66408 , n66409 , n66410 , n66411 , n66412 , n66413 , n66414 , n66415 , n66416 , 
 n66417 , n66418 , n66419 , n66420 , n66421 , n66422 , n66423 , n66424 , n66425 , n66426 , 
 n66427 , n66428 , n66429 , n66430 , n66431 , n66432 , n66433 , n66434 , n66435 , n66436 , 
 n66437 , n66438 , n66439 , n66440 , n66441 , n66442 , n66443 , n66444 , n66445 , n66446 , 
 n66447 , n66448 , n66449 , n66450 , n66451 , n66452 , n66453 , n66454 , n66455 , n66456 , 
 n66457 , n66458 , n66459 , n66460 , n66461 , n66462 , n66463 , n66464 , n66465 , n66466 , 
 n66467 , n66468 , n66469 , n66470 , n66471 , n66472 , n66473 , n66474 , n66475 , n66476 , 
 n66477 , n66478 , n66479 , n66480 , n66481 , n66482 , n66483 , n66484 , n66485 , n66486 , 
 n66487 , n66488 , n66489 , n66490 , n66491 , n66492 , n66493 , n66494 , n66495 , n66496 , 
 n66497 , n66498 , n66499 , n66500 , n66501 , n66502 , n66503 , n66504 , n66505 , n66506 , 
 n66507 , n66508 , n66509 , n66510 , n66511 , n66512 , n66513 , n66514 , n66515 , n66516 , 
 n66517 , n66518 , n66519 , n66520 , n66521 , n66522 , n66523 , n66524 , n66525 , n66526 , 
 n66527 , n66528 , n66529 , n66530 , n66531 , n66532 , n66533 , n66534 , n66535 , n66536 , 
 n66537 , n66538 , n66539 , n66540 , n66541 , n66542 , n66543 , n66544 , n66545 , n66546 , 
 n66547 , n66548 , n66549 , n66550 , n66551 , n66552 , n66553 , n66554 , n66555 , n66556 , 
 n66557 , n66558 , n66559 , n66560 , n66561 , n66562 , n66563 , n66564 , n66565 , n66566 , 
 n66567 , n66568 , n66569 , n66570 , n66571 , n66572 , n66573 , n66574 , n66575 , n66576 , 
 n66577 , n66578 , n66579 , n66580 , n66581 , n66582 , n66583 , n66584 , n66585 , n66586 , 
 n66587 , n66588 , n66589 , n66590 , n66591 , n66592 , n66593 , n66594 , n66595 , n66596 , 
 n66597 , n66598 , n66599 , n66600 , n66601 , n66602 , n66603 , n66604 , n66605 , n66606 , 
 n66607 , n66608 , n66609 , n66610 , n66611 , n66612 , n66613 , n66614 , n66615 , n66616 , 
 n66617 , n66618 , n66619 , n66620 , n66621 , n66622 , n66623 , n66624 , n66625 , n66626 , 
 n66627 , n66628 , n66629 , n66630 , n66631 , n66632 , n66633 , n66634 , n66635 , n66636 , 
 n66637 , n66638 , n66639 , n66640 , n66641 , n66642 , n66643 , n66644 , n66645 , n66646 , 
 n66647 , n66648 , n66649 , n66650 , n66651 , n66652 , n66653 , n66654 , n66655 , n66656 , 
 n66657 , n66658 , n66659 , n66660 , n66661 , n66662 , n66663 , n66664 , n66665 , n66666 , 
 n66667 , n66668 , n66669 , n66670 , n66671 , n66672 , n66673 , n66674 , n66675 , n66676 , 
 n66677 , n66678 , n66679 , n66680 , n66681 , n66682 , n66683 , n66684 , n66685 , n66686 , 
 n66687 , n66688 , n66689 , n66690 , n66691 , n66692 , n66693 , n66694 , n66695 , n66696 , 
 n66697 , n66698 , n66699 , n66700 , n66701 , n66702 , n66703 , n66704 , n66705 , n66706 , 
 n66707 , n66708 , n66709 , n66710 , n66711 , n66712 , n66713 , n66714 , n66715 , n66716 , 
 n66717 , n66718 , n66719 , n66720 , n66721 , n66722 , n66723 , n66724 , n66725 , n66726 , 
 n66727 , n66728 , n66729 , n66730 , n66731 , n66732 , n66733 , n66734 , n66735 , n66736 , 
 n66737 , n66738 , n66739 , n66740 , n66741 , n66742 , n66743 , n66744 , n66745 , n66746 , 
 n66747 , n66748 , n66749 , n66750 , n66751 , n66752 , n66753 , n66754 , n66755 , n66756 , 
 n66757 , n66758 , n66759 , n66760 , n66761 , n66762 , n66763 , n66764 , n66765 , n66766 , 
 n66767 , n66768 , n66769 , n66770 , n66771 , n66772 , n66773 , n66774 , n66775 , n66776 , 
 n66777 , n66778 , n66779 , n66780 , n66781 , n66782 , n66783 , n66784 , n66785 , n66786 , 
 n66787 , n66788 , n66789 , n66790 , n66791 , n66792 , n66793 , n66794 , n66795 , n66796 , 
 n66797 , n66798 , n66799 , n66800 , n66801 , n66802 , n66803 , n66804 , n66805 , n66806 , 
 n66807 , n66808 , n66809 , n66810 , n66811 , n66812 , n66813 , n66814 , n66815 , n66816 , 
 n66817 , n66818 , n66819 , n66820 , n66821 , n66822 , n66823 , n66824 , n66825 , n66826 , 
 n66827 , n66828 , n66829 , n66830 , n66831 , n66832 , n66833 , n66834 , n66835 , n66836 , 
 n66837 , n66838 , n66839 , n66840 , n66841 , n66842 , n66843 , n66844 , n66845 , n66846 , 
 n66847 , n66848 , n66849 , n66850 , n66851 , n66852 , n66853 , n66854 , n66855 , n66856 , 
 n66857 , n66858 , n66859 , n66860 , n66861 , n66862 , n66863 , n66864 , n66865 , n66866 , 
 n66867 , n66868 , n66869 , n66870 , n66871 , n66872 , n66873 , n66874 , n66875 , n66876 , 
 n66877 , n66878 , n66879 , n66880 , n66881 , n66882 , n66883 , n66884 , n66885 , n66886 , 
 n66887 , n66888 , n66889 , n66890 , n66891 , n66892 , n66893 , n66894 , n66895 , n66896 , 
 n66897 , n66898 , n66899 , n66900 , n66901 , n66902 , n66903 , n66904 , n66905 , n66906 , 
 n66907 , n66908 , n66909 , n66910 , n66911 , n66912 , n66913 , n66914 , n66915 , n66916 , 
 n66917 , n66918 , n66919 , n66920 , n66921 , n66922 , n66923 , n66924 , n66925 , n66926 , 
 n66927 , n66928 , n66929 , n66930 , n66931 , n66932 , n66933 , n66934 , n66935 , n66936 , 
 n66937 , n66938 , n66939 , n66940 , n66941 , n66942 , n66943 , n66944 , n66945 , n66946 , 
 n66947 , n66948 , n66949 , n66950 , n66951 , n66952 , n66953 , n66954 , n66955 , n66956 , 
 n66957 , n66958 , n66959 , n66960 , n66961 , n66962 , n66963 , n66964 , n66965 , n66966 , 
 n66967 , n66968 , n66969 , n66970 , n66971 , n66972 , n66973 , n66974 , n66975 , n66976 , 
 n66977 , n66978 , n66979 , n66980 , n66981 , n66982 , n66983 , n66984 , n66985 , n66986 , 
 n66987 , n66988 , n66989 , n66990 , n66991 , n66992 , n66993 , n66994 , n66995 , n66996 , 
 n66997 , n66998 , n66999 , n67000 , n67001 , n67002 , n67003 , n67004 , n67005 , n67006 , 
 n67007 , n67008 , n67009 , n67010 , n67011 , n67012 , n67013 , n67014 , n67015 , n67016 , 
 n67017 , n67018 , n67019 , n67020 , n67021 , n67022 , n67023 , n67024 , n67025 , n67026 , 
 n67027 , n67028 , n67029 , n67030 , n67031 , n67032 , n67033 , n67034 , n67035 , n67036 , 
 n67037 , n67038 , n67039 , n67040 , n67041 , n67042 , n67043 , n67044 , n67045 , n67046 , 
 n67047 , n67048 , n67049 , n67050 , n67051 , n67052 , n67053 , n67054 , n67055 , n67056 , 
 n67057 , n67058 , n67059 , n67060 , n67061 , n67062 , n67063 , n67064 , n67065 , n67066 , 
 n67067 , n67068 , n67069 , n67070 , n67071 , n67072 , n67073 , n67074 , n67075 , n67076 , 
 n67077 , n67078 , n67079 , n67080 , n67081 , n67082 , n67083 , n67084 , n67085 , n67086 , 
 n67087 , n67088 , n67089 , n67090 , n67091 , n67092 , n67093 , n67094 , n67095 , n67096 , 
 n67097 , n67098 , n67099 , n67100 , n67101 , n67102 , n67103 , n67104 , n67105 , n67106 , 
 n67107 , n67108 , n67109 , n67110 , n67111 , n67112 , n67113 , n67114 , n67115 , n67116 , 
 n67117 , n67118 , n67119 , n67120 , n67121 , n67122 , n67123 , n67124 , n67125 , n67126 , 
 n67127 , n67128 , n67129 , n67130 , n67131 , n67132 , n67133 , n67134 , n67135 , n67136 , 
 n67137 , n67138 , n67139 , n67140 , n67141 , n67142 , n67143 , n67144 , n67145 , n67146 , 
 n67147 , n67148 , n67149 , n67150 , n67151 , n67152 , n67153 , n67154 , n67155 , n67156 , 
 n67157 , n67158 , n67159 , n67160 , n67161 , n67162 , n67163 , n67164 , n67165 , n67166 , 
 n67167 , n67168 , n67169 , n67170 , n67171 , n67172 , n67173 , n67174 , n67175 , n67176 , 
 n67177 , n67178 , n67179 , n67180 , n67181 , n67182 , n67183 , n67184 , n67185 , n67186 , 
 n67187 , n67188 , n67189 , n67190 , n67191 , n67192 , n67193 , n67194 , n67195 , n67196 , 
 n67197 , n67198 , n67199 , n67200 , n67201 , n67202 , n67203 , n67204 , n67205 , n67206 , 
 n67207 , n67208 , n67209 , n67210 , n67211 , n67212 , n67213 , n67214 , n67215 , n67216 , 
 n67217 , n67218 , n67219 , n67220 , n67221 , n67222 , n67223 , n67224 , n67225 , n67226 , 
 n67227 , n67228 , n67229 , n67230 , n67231 , n67232 , n67233 , n67234 , n67235 , n67236 , 
 n67237 , n67238 , n67239 , n67240 , n67241 , n67242 , n67243 , n67244 , n67245 , n67246 , 
 n67247 , n67248 , n67249 , n67250 , n67251 , n67252 , n67253 , n67254 , n67255 , n67256 , 
 n67257 , n67258 , n67259 , n67260 , n67261 , n67262 , n67263 , n67264 , n67265 , n67266 , 
 n67267 , n67268 , n67269 , n67270 , n67271 , n67272 , n67273 , n67274 , n67275 , n67276 , 
 n67277 , n67278 , n67279 , n67280 , n67281 , n67282 , n67283 , n67284 , n67285 , n67286 , 
 n67287 , n67288 , n67289 , n67290 , n67291 , n67292 , n67293 , n67294 , n67295 , n67296 , 
 n67297 , n67298 , n67299 , n67300 , n67301 , n67302 , n67303 , n67304 , n67305 , n67306 , 
 n67307 , n67308 , n67309 , n67310 , n67311 , n67312 , n67313 , n67314 , n67315 , n67316 , 
 n67317 , n67318 , n67319 , n67320 , n67321 , n67322 , n67323 , n67324 , n67325 , n67326 , 
 n67327 , n67328 , n67329 , n67330 , n67331 , n67332 , n67333 , n67334 , n67335 , n67336 , 
 n67337 , n67338 , n67339 , n67340 , n67341 , n67342 , n67343 , n67344 , n67345 , n67346 , 
 n67347 , n67348 , n67349 , n67350 , n67351 , n67352 , n67353 , n67354 , n67355 , n67356 , 
 n67357 , n67358 , n67359 , n67360 , n67361 , n67362 , n67363 , n67364 , n67365 , n67366 , 
 n67367 , n67368 , n67369 , n67370 , n67371 , n67372 , n67373 , n67374 , n67375 , n67376 , 
 n67377 , n67378 , n67379 , n67380 , n67381 , n67382 , n67383 , n67384 , n67385 , n67386 , 
 n67387 , n67388 , n67389 , n67390 , n67391 , n67392 , n67393 , n67394 , n67395 , n67396 , 
 n67397 , n67398 , n67399 , n67400 , n67401 , n67402 , n67403 , n67404 , n67405 , n67406 , 
 n67407 , n67408 , n67409 , n67410 , n67411 , n67412 , n67413 , n67414 , n67415 , n67416 , 
 n67417 , n67418 , n67419 , n67420 , n67421 , n67422 , n67423 , n67424 , n67425 , n67426 , 
 n67427 , n67428 , n67429 , n67430 , n67431 , n67432 , n67433 , n67434 , n67435 , n67436 , 
 n67437 , n67438 , n67439 , n67440 , n67441 , n67442 , n67443 , n67444 , n67445 , n67446 , 
 n67447 , n67448 , n67449 , n67450 , n67451 , n67452 , n67453 , n67454 , n67455 , n67456 , 
 n67457 , n67458 , n67459 , n67460 , n67461 , n67462 , n67463 , n67464 , n67465 , n67466 , 
 n67467 , n67468 , n67469 , n67470 , n67471 , n67472 , n67473 , n67474 , n67475 , n67476 , 
 n67477 , n67478 , n67479 , n67480 , n67481 , n67482 , n67483 , n67484 , n67485 , n67486 , 
 n67487 , n67488 , n67489 , n67490 , n67491 , n67492 , n67493 , n67494 , n67495 , n67496 , 
 n67497 , n67498 , n67499 , n67500 , n67501 , n67502 , n67503 , n67504 , n67505 , n67506 , 
 n67507 , n67508 , n67509 , n67510 , n67511 , n67512 , n67513 , n67514 , n67515 , n67516 , 
 n67517 , n67518 , n67519 , n67520 , n67521 , n67522 , n67523 , n67524 , n67525 , n67526 , 
 n67527 , n67528 , n67529 , n67530 , n67531 , n67532 , n67533 , n67534 , n67535 , n67536 , 
 n67537 , n67538 , n67539 , n67540 , n67541 , n67542 , n67543 , n67544 , n67545 , n67546 , 
 n67547 , n67548 , n67549 , n67550 , n67551 , n67552 , n67553 , n67554 , n67555 , n67556 , 
 n67557 , n67558 , n67559 , n67560 , n67561 , n67562 , n67563 , n67564 , n67565 , n67566 , 
 n67567 , n67568 , n67569 , n67570 , n67571 , n67572 , n67573 , n67574 , n67575 , n67576 , 
 n67577 , n67578 , n67579 , n67580 , n67581 , n67582 , n67583 , n67584 , n67585 , n67586 , 
 n67587 , n67588 , n67589 , n67590 , n67591 , n67592 , n67593 , n67594 , n67595 , n67596 , 
 n67597 , n67598 , n67599 , n67600 , n67601 , n67602 , n67603 , n67604 , n67605 , n67606 , 
 n67607 , n67608 , n67609 , n67610 , n67611 , n67612 , n67613 , n67614 , n67615 , n67616 , 
 n67617 , n67618 , n67619 , n67620 , n67621 , n67622 , n67623 , n67624 , n67625 , n67626 , 
 n67627 , n67628 , n67629 , n67630 , n67631 , n67632 , n67633 , n67634 , n67635 , n67636 , 
 n67637 , n67638 , n67639 , n67640 , n67641 , n67642 , n67643 , n67644 , n67645 , n67646 , 
 n67647 , n67648 , n67649 , n67650 , n67651 , n67652 , n67653 , n67654 , n67655 , n67656 , 
 n67657 , n67658 , n67659 , n67660 , n67661 , n67662 , n67663 , n67664 , n67665 , n67666 , 
 n67667 , n67668 , n67669 , n67670 , n67671 , n67672 , n67673 , n67674 , n67675 , n67676 , 
 n67677 , n67678 , n67679 , n67680 , n67681 , n67682 , n67683 , n67684 , n67685 , n67686 , 
 n67687 , n67688 , n67689 , n67690 , n67691 , n67692 , n67693 , n67694 , n67695 , n67696 , 
 n67697 , n67698 , n67699 , n67700 , n67701 , n67702 , n67703 , n67704 , n67705 , n67706 , 
 n67707 , n67708 , n67709 , n67710 , n67711 , n67712 , n67713 , n67714 , n67715 , n67716 , 
 n67717 , n67718 , n67719 , n67720 , n67721 , n67722 , n67723 , n67724 , n67725 , n67726 , 
 n67727 , n67728 , n67729 , n67730 , n67731 , n67732 , n67733 , n67734 , n67735 , n67736 , 
 n67737 , n67738 , n67739 , n67740 , n67741 , n67742 , n67743 , n67744 , n67745 , n67746 , 
 n67747 , n67748 , n67749 , n67750 , n67751 , n67752 , n67753 , n67754 , n67755 , n67756 , 
 n67757 , n67758 , n67759 , n67760 , n67761 , n67762 , n67763 , n67764 , n67765 , n67766 , 
 n67767 , n67768 , n67769 , n67770 , n67771 , n67772 , n67773 , n67774 , n67775 , n67776 , 
 n67777 , n67778 , n67779 , n67780 , n67781 , n67782 , n67783 , n67784 , n67785 , n67786 , 
 n67787 , n67788 , n67789 , n67790 , n67791 , n67792 , n67793 , n67794 , n67795 , n67796 , 
 n67797 , n67798 , n67799 , n67800 , n67801 , n67802 , n67803 , n67804 , n67805 , n67806 , 
 n67807 , n67808 , n67809 , n67810 , n67811 , n67812 , n67813 , n67814 , n67815 , n67816 , 
 n67817 , n67818 , n67819 , n67820 , n67821 , n67822 , n67823 , n67824 , n67825 , n67826 , 
 n67827 , n67828 , n67829 , n67830 , n67831 , n67832 , n67833 , n67834 , n67835 , n67836 , 
 n67837 , n67838 , n67839 , n67840 , n67841 , n67842 , n67843 , n67844 , n67845 , n67846 , 
 n67847 , n67848 , n67849 , n67850 , n67851 , n67852 , n67853 , n67854 , n67855 , n67856 , 
 n67857 , n67858 , n67859 , n67860 , n67861 , n67862 , n67863 , n67864 , n67865 , n67866 , 
 n67867 , n67868 , n67869 , n67870 , n67871 , n67872 , n67873 , n67874 , n67875 , n67876 , 
 n67877 , n67878 , n67879 , n67880 , n67881 , n67882 , n67883 , n67884 , n67885 , n67886 , 
 n67887 , n67888 , n67889 , n67890 , n67891 , n67892 , n67893 , n67894 , n67895 , n67896 , 
 n67897 , n67898 , n67899 , n67900 , n67901 , n67902 , n67903 , n67904 , n67905 , n67906 , 
 n67907 , n67908 , n67909 , n67910 , n67911 , n67912 , n67913 , n67914 , n67915 , n67916 , 
 n67917 , n67918 , n67919 , n67920 , n67921 , n67922 , n67923 , n67924 , n67925 , n67926 , 
 n67927 , n67928 , n67929 , n67930 , n67931 , n67932 , n67933 , n67934 , n67935 , n67936 , 
 n67937 , n67938 , n67939 , n67940 , n67941 , n67942 , n67943 , n67944 , n67945 , n67946 , 
 n67947 , n67948 , n67949 , n67950 , n67951 , n67952 , n67953 , n67954 , n67955 , n67956 , 
 n67957 , n67958 , n67959 , n67960 , n67961 , n67962 , n67963 , n67964 , n67965 , n67966 , 
 n67967 , n67968 , n67969 , n67970 , n67971 , n67972 , n67973 , n67974 , n67975 , n67976 , 
 n67977 , n67978 , n67979 , n67980 , n67981 , n67982 , n67983 , n67984 , n67985 , n67986 , 
 n67987 , n67988 , n67989 , n67990 , n67991 , n67992 , n67993 , n67994 , n67995 , n67996 , 
 n67997 , n67998 , n67999 , n68000 , n68001 , n68002 , n68003 , n68004 , n68005 , n68006 , 
 n68007 , n68008 , n68009 , n68010 , n68011 , n68012 , n68013 , n68014 , n68015 , n68016 , 
 n68017 , n68018 , n68019 , n68020 , n68021 , n68022 , n68023 , n68024 , n68025 , n68026 , 
 n68027 , n68028 , n68029 , n68030 , n68031 , n68032 , n68033 , n68034 , n68035 , n68036 , 
 n68037 , n68038 , n68039 , n68040 , n68041 , n68042 , n68043 , n68044 , n68045 , n68046 , 
 n68047 , n68048 , n68049 , n68050 , n68051 , n68052 , n68053 , n68054 , n68055 , n68056 , 
 n68057 , n68058 , n68059 , n68060 , n68061 , n68062 , n68063 , n68064 , n68065 , n68066 , 
 n68067 , n68068 , n68069 , n68070 , n68071 , n68072 , n68073 , n68074 , n68075 , n68076 , 
 n68077 , n68078 , n68079 , n68080 , n68081 , n68082 , n68083 , n68084 , n68085 , n68086 , 
 n68087 , n68088 , n68089 , n68090 , n68091 , n68092 , n68093 , n68094 , n68095 , n68096 , 
 n68097 , n68098 , n68099 , n68100 , n68101 , n68102 , n68103 , n68104 , n68105 , n68106 , 
 n68107 , n68108 , n68109 , n68110 , n68111 , n68112 , n68113 , n68114 , n68115 , n68116 , 
 n68117 , n68118 , n68119 , n68120 , n68121 , n68122 , n68123 , n68124 , n68125 , n68126 , 
 n68127 , n68128 , n68129 , n68130 , n68131 , n68132 , n68133 , n68134 , n68135 , n68136 , 
 n68137 , n68138 , n68139 , n68140 , n68141 , n68142 , n68143 , n68144 , n68145 , n68146 , 
 n68147 , n68148 , n68149 , n68150 , n68151 , n68152 , n68153 , n68154 , n68155 , n68156 , 
 n68157 , n68158 , n68159 , n68160 , n68161 , n68162 , n68163 , n68164 , n68165 , n68166 , 
 n68167 , n68168 , n68169 , n68170 , n68171 , n68172 , n68173 , n68174 , n68175 , n68176 , 
 n68177 , n68178 , n68179 , n68180 , n68181 , n68182 , n68183 , n68184 , n68185 , n68186 , 
 n68187 , n68188 , n68189 , n68190 , n68191 , n68192 , n68193 , n68194 , n68195 , n68196 , 
 n68197 , n68198 , n68199 , n68200 , n68201 , n68202 , n68203 , n68204 , n68205 , n68206 , 
 n68207 , n68208 , n68209 , n68210 , n68211 , n68212 , n68213 , n68214 , n68215 , n68216 , 
 n68217 , n68218 , n68219 , n68220 , n68221 , n68222 , n68223 , n68224 , n68225 , n68226 , 
 n68227 , n68228 , n68229 , n68230 , n68231 , n68232 , n68233 , n68234 , n68235 , n68236 , 
 n68237 , n68238 , n68239 , n68240 , n68241 , n68242 , n68243 , n68244 , n68245 , n68246 , 
 n68247 , n68248 , n68249 , n68250 , n68251 , n68252 , n68253 , n68254 , n68255 , n68256 , 
 n68257 , n68258 , n68259 , n68260 , n68261 , n68262 , n68263 , n68264 , n68265 , n68266 , 
 n68267 , n68268 , n68269 , n68270 , n68271 , n68272 , n68273 , n68274 , n68275 , n68276 , 
 n68277 , n68278 , n68279 , n68280 , n68281 , n68282 , n68283 , n68284 , n68285 , n68286 , 
 n68287 , n68288 , n68289 , n68290 , n68291 , n68292 , n68293 , n68294 , n68295 , n68296 , 
 n68297 , n68298 , n68299 , n68300 , n68301 , n68302 , n68303 , n68304 , n68305 , n68306 , 
 n68307 , n68308 , n68309 , n68310 , n68311 , n68312 , n68313 , n68314 , n68315 , n68316 , 
 n68317 , n68318 , n68319 , n68320 , n68321 , n68322 , n68323 , n68324 , n68325 , n68326 , 
 n68327 , n68328 , n68329 , n68330 , n68331 , n68332 , n68333 , n68334 , n68335 , n68336 , 
 n68337 , n68338 , n68339 , n68340 , n68341 , n68342 , n68343 , n68344 , n68345 , n68346 , 
 n68347 , n68348 , n68349 , n68350 , n68351 , n68352 , n68353 , n68354 , n68355 , n68356 , 
 n68357 , n68358 , n68359 , n68360 , n68361 , n68362 , n68363 , n68364 , n68365 , n68366 , 
 n68367 , n68368 , n68369 , n68370 , n68371 , n68372 , n68373 , n68374 , n68375 , n68376 , 
 n68377 , n68378 , n68379 , n68380 , n68381 , n68382 , n68383 , n68384 , n68385 , n68386 , 
 n68387 , n68388 , n68389 , n68390 , n68391 , n68392 , n68393 , n68394 , n68395 , n68396 , 
 n68397 , n68398 , n68399 , n68400 , n68401 , n68402 , n68403 , n68404 , n68405 , n68406 , 
 n68407 , n68408 , n68409 , n68410 , n68411 , n68412 , n68413 , n68414 , n68415 , n68416 , 
 n68417 , n68418 , n68419 , n68420 , n68421 , n68422 , n68423 , n68424 , n68425 , n68426 , 
 n68427 , n68428 , n68429 , n68430 , n68431 , n68432 , n68433 , n68434 , n68435 , n68436 , 
 n68437 , n68438 , n68439 , n68440 , n68441 , n68442 , n68443 , n68444 , n68445 , n68446 , 
 n68447 , n68448 , n68449 , n68450 , n68451 , n68452 , n68453 , n68454 , n68455 , n68456 , 
 n68457 , n68458 , n68459 , n68460 , n68461 , n68462 , n68463 , n68464 , n68465 , n68466 , 
 n68467 , n68468 , n68469 , n68470 , n68471 , n68472 , n68473 , n68474 , n68475 , n68476 , 
 n68477 , n68478 , n68479 , n68480 , n68481 , n68482 , n68483 , n68484 , n68485 , n68486 , 
 n68487 , n68488 , n68489 , n68490 , n68491 , n68492 , n68493 , n68494 , n68495 , n68496 , 
 n68497 , n68498 , n68499 , n68500 , n68501 , n68502 , n68503 , n68504 , n68505 , n68506 , 
 n68507 , n68508 , n68509 , n68510 , n68511 , n68512 , n68513 , n68514 , n68515 , n68516 , 
 n68517 , n68518 , n68519 , n68520 , n68521 , n68522 , n68523 , n68524 , n68525 , n68526 , 
 n68527 , n68528 , n68529 , n68530 , n68531 , n68532 , n68533 , n68534 , n68535 , n68536 , 
 n68537 , n68538 , n68539 , n68540 , n68541 , n68542 , n68543 , n68544 , n68545 , n68546 , 
 n68547 , n68548 , n68549 , n68550 , n68551 , n68552 , n68553 , n68554 , n68555 , n68556 , 
 n68557 , n68558 , n68559 , n68560 , n68561 , n68562 , n68563 , n68564 , n68565 , n68566 , 
 n68567 , n68568 , n68569 , n68570 , n68571 , n68572 , n68573 , n68574 , n68575 , n68576 , 
 n68577 , n68578 , n68579 , n68580 , n68581 , n68582 , n68583 , n68584 , n68585 , n68586 , 
 n68587 , n68588 , n68589 , n68590 , n68591 , n68592 , n68593 , n68594 , n68595 , n68596 , 
 n68597 , n68598 , n68599 , n68600 , n68601 , n68602 , n68603 , n68604 , n68605 , n68606 , 
 n68607 , n68608 , n68609 , n68610 , n68611 , n68612 , n68613 , n68614 , n68615 , n68616 , 
 n68617 , n68618 , n68619 , n68620 , n68621 , n68622 , n68623 , n68624 , n68625 , n68626 , 
 n68627 , n68628 , n68629 , n68630 , n68631 , n68632 , n68633 , n68634 , n68635 , n68636 , 
 n68637 , n68638 , n68639 , n68640 , n68641 , n68642 , n68643 , n68644 , n68645 , n68646 , 
 n68647 , n68648 , n68649 , n68650 , n68651 , n68652 , n68653 , n68654 , n68655 , n68656 , 
 n68657 , n68658 , n68659 , n68660 , n68661 , n68662 , n68663 , n68664 , n68665 , n68666 , 
 n68667 , n68668 , n68669 , n68670 , n68671 , n68672 , n68673 , n68674 , n68675 , n68676 , 
 n68677 , n68678 , n68679 , n68680 , n68681 , n68682 , n68683 , n68684 , n68685 , n68686 , 
 n68687 , n68688 , n68689 , n68690 , n68691 , n68692 , n68693 , n68694 , n68695 , n68696 , 
 n68697 , n68698 , n68699 , n68700 , n68701 , n68702 , n68703 , n68704 , n68705 , n68706 , 
 n68707 , n68708 , n68709 , n68710 , n68711 , n68712 , n68713 , n68714 , n68715 , n68716 , 
 n68717 , n68718 , n68719 , n68720 , n68721 , n68722 , n68723 , n68724 , n68725 , n68726 , 
 n68727 , n68728 , n68729 , n68730 , n68731 , n68732 , n68733 , n68734 , n68735 , n68736 , 
 n68737 , n68738 , n68739 , n68740 , n68741 , n68742 , n68743 , n68744 , n68745 , n68746 , 
 n68747 , n68748 , n68749 , n68750 , n68751 , n68752 , n68753 , n68754 , n68755 , n68756 , 
 n68757 , n68758 , n68759 , n68760 , n68761 , n68762 , n68763 , n68764 , n68765 , n68766 , 
 n68767 , n68768 , n68769 , n68770 , n68771 , n68772 , n68773 , n68774 , n68775 , n68776 , 
 n68777 , n68778 , n68779 , n68780 , n68781 , n68782 , n68783 , n68784 , n68785 , n68786 , 
 n68787 , n68788 , n68789 , n68790 , n68791 , n68792 , n68793 , n68794 , n68795 , n68796 , 
 n68797 , n68798 , n68799 , n68800 , n68801 , n68802 , n68803 , n68804 , n68805 , n68806 , 
 n68807 , n68808 , n68809 , n68810 , n68811 , n68812 , n68813 , n68814 , n68815 , n68816 , 
 n68817 , n68818 , n68819 , n68820 , n68821 , n68822 , n68823 , n68824 , n68825 , n68826 , 
 n68827 , n68828 , n68829 , n68830 , n68831 , n68832 , n68833 , n68834 , n68835 , n68836 , 
 n68837 , n68838 , n68839 , n68840 , n68841 , n68842 , n68843 , n68844 , n68845 , n68846 , 
 n68847 , n68848 , n68849 , n68850 , n68851 , n68852 , n68853 , n68854 , n68855 , n68856 , 
 n68857 , n68858 , n68859 , n68860 , n68861 , n68862 , n68863 , n68864 , n68865 , n68866 , 
 n68867 , n68868 , n68869 , n68870 , n68871 , n68872 , n68873 , n68874 , n68875 , n68876 , 
 n68877 , n68878 , n68879 , n68880 , n68881 , n68882 , n68883 , n68884 , n68885 , n68886 , 
 n68887 , n68888 , n68889 , n68890 , n68891 , n68892 , n68893 , n68894 , n68895 , n68896 , 
 n68897 , n68898 , n68899 , n68900 , n68901 , n68902 , n68903 , n68904 , n68905 , n68906 , 
 n68907 , n68908 , n68909 , n68910 , n68911 , n68912 , n68913 , n68914 , n68915 , n68916 , 
 n68917 , n68918 , n68919 , n68920 , n68921 , n68922 , n68923 , n68924 , n68925 , n68926 , 
 n68927 , n68928 , n68929 , n68930 , n68931 , n68932 , n68933 , n68934 , n68935 , n68936 , 
 n68937 , n68938 , n68939 , n68940 , n68941 , n68942 , n68943 , n68944 , n68945 , n68946 , 
 n68947 , n68948 , n68949 , n68950 , n68951 , n68952 , n68953 , n68954 , n68955 , n68956 , 
 n68957 , n68958 , n68959 , n68960 , n68961 , n68962 , n68963 , n68964 , n68965 , n68966 , 
 n68967 , n68968 , n68969 , n68970 , n68971 , n68972 , n68973 , n68974 , n68975 , n68976 , 
 n68977 , n68978 , n68979 , n68980 , n68981 , n68982 , n68983 , n68984 , n68985 , n68986 , 
 n68987 , n68988 , n68989 , n68990 , n68991 , n68992 , n68993 , n68994 , n68995 , n68996 , 
 n68997 , n68998 , n68999 , n69000 , n69001 , n69002 , n69003 , n69004 , n69005 , n69006 , 
 n69007 , n69008 , n69009 , n69010 , n69011 , n69012 , n69013 , n69014 , n69015 , n69016 , 
 n69017 , n69018 , n69019 , n69020 , n69021 , n69022 , n69023 , n69024 , n69025 , n69026 , 
 n69027 , n69028 , n69029 , n69030 , n69031 , n69032 , n69033 , n69034 , n69035 , n69036 , 
 n69037 , n69038 , n69039 , n69040 , n69041 , n69042 , n69043 , n69044 , n69045 , n69046 , 
 n69047 , n69048 , n69049 , n69050 , n69051 , n69052 , n69053 , n69054 , n69055 , n69056 , 
 n69057 , n69058 , n69059 , n69060 , n69061 , n69062 , n69063 , n69064 , n69065 , n69066 , 
 n69067 , n69068 , n69069 , n69070 , n69071 , n69072 , n69073 , n69074 , n69075 , n69076 , 
 n69077 , n69078 , n69079 , n69080 , n69081 , n69082 , n69083 , n69084 , n69085 , n69086 , 
 n69087 , n69088 , n69089 , n69090 , n69091 , n69092 , n69093 , n69094 , n69095 , n69096 , 
 n69097 , n69098 , n69099 , n69100 , n69101 , n69102 , n69103 , n69104 , n69105 , n69106 , 
 n69107 , n69108 , n69109 , n69110 , n69111 , n69112 , n69113 , n69114 , n69115 , n69116 , 
 n69117 , n69118 , n69119 , n69120 , n69121 , n69122 , n69123 , n69124 , n69125 , n69126 , 
 n69127 , n69128 , n69129 , n69130 , n69131 , n69132 , n69133 , n69134 , n69135 , n69136 , 
 n69137 , n69138 , n69139 , n69140 , n69141 , n69142 , n69143 , n69144 , n69145 , n69146 , 
 n69147 , n69148 , n69149 , n69150 , n69151 , n69152 , n69153 , n69154 , n69155 , n69156 , 
 n69157 , n69158 , n69159 , n69160 , n69161 , n69162 , n69163 , n69164 , n69165 , n69166 , 
 n69167 , n69168 , n69169 , n69170 , n69171 , n69172 , n69173 , n69174 , n69175 , n69176 , 
 n69177 , n69178 , n69179 , n69180 , n69181 , n69182 , n69183 , n69184 , n69185 , n69186 , 
 n69187 , n69188 , n69189 , n69190 , n69191 , n69192 , n69193 , n69194 , n69195 , n69196 , 
 n69197 , n69198 , n69199 , n69200 , n69201 , n69202 , n69203 , n69204 , n69205 , n69206 , 
 n69207 , n69208 , n69209 , n69210 , n69211 , n69212 , n69213 , n69214 , n69215 , n69216 , 
 n69217 , n69218 , n69219 , n69220 , n69221 , n69222 , n69223 , n69224 , n69225 , n69226 , 
 n69227 , n69228 , n69229 , n69230 , n69231 , n69232 , n69233 , n69234 , n69235 , n69236 , 
 n69237 , n69238 , n69239 , n69240 , n69241 , n69242 , n69243 , n69244 , n69245 , n69246 , 
 n69247 , n69248 , n69249 , n69250 , n69251 , n69252 , n69253 , n69254 , n69255 , n69256 , 
 n69257 , n69258 , n69259 , n69260 , n69261 , n69262 , n69263 , n69264 , n69265 , n69266 , 
 n69267 , n69268 , n69269 , n69270 , n69271 , n69272 , n69273 , n69274 , n69275 , n69276 , 
 n69277 , n69278 , n69279 , n69280 , n69281 , n69282 , n69283 , n69284 , n69285 , n69286 , 
 n69287 , n69288 , n69289 , n69290 , n69291 , n69292 , n69293 , n69294 , n69295 , n69296 , 
 n69297 , n69298 , n69299 , n69300 , n69301 , n69302 , n69303 , n69304 , n69305 , n69306 , 
 n69307 , n69308 , n69309 , n69310 , n69311 , n69312 , n69313 , n69314 , n69315 , n69316 , 
 n69317 , n69318 , n69319 , n69320 , n69321 , n69322 , n69323 , n69324 , n69325 , n69326 , 
 n69327 , n69328 , n69329 , n69330 , n69331 , n69332 , n69333 , n69334 , n69335 , n69336 , 
 n69337 , n69338 , n69339 , n69340 , n69341 , n69342 , n69343 , n69344 , n69345 , n69346 , 
 n69347 , n69348 , n69349 , n69350 , n69351 , n69352 , n69353 , n69354 , n69355 , n69356 , 
 n69357 , n69358 , n69359 , n69360 , n69361 , n69362 , n69363 , n69364 , n69365 , n69366 , 
 n69367 , n69368 , n69369 , n69370 , n69371 , n69372 , n69373 , n69374 , n69375 , n69376 , 
 n69377 , n69378 , n69379 , n69380 , n69381 , n69382 , n69383 , n69384 , n69385 , n69386 , 
 n69387 , n69388 , n69389 , n69390 , n69391 , n69392 , n69393 , n69394 , n69395 , n69396 , 
 n69397 , n69398 , n69399 , n69400 , n69401 , n69402 , n69403 , n69404 , n69405 , n69406 , 
 n69407 , n69408 , n69409 , n69410 , n69411 , n69412 , n69413 , n69414 , n69415 , n69416 , 
 n69417 , n69418 , n69419 , n69420 , n69421 , n69422 , n69423 , n69424 , n69425 , n69426 , 
 n69427 , n69428 , n69429 , n69430 , n69431 , n69432 , n69433 , n69434 , n69435 , n69436 , 
 n69437 , n69438 , n69439 , n69440 , n69441 , n69442 , n69443 , n69444 , n69445 , n69446 , 
 n69447 , n69448 , n69449 , n69450 , n69451 , n69452 , n69453 , n69454 , n69455 , n69456 , 
 n69457 , n69458 , n69459 , n69460 , n69461 , n69462 , n69463 , n69464 , n69465 , n69466 , 
 n69467 , n69468 , n69469 , n69470 , n69471 , n69472 , n69473 , n69474 , n69475 , n69476 , 
 n69477 , n69478 , n69479 , n69480 , n69481 , n69482 , n69483 , n69484 , n69485 , n69486 , 
 n69487 , n69488 , n69489 , n69490 , n69491 , n69492 , n69493 , n69494 , n69495 , n69496 , 
 n69497 , n69498 , n69499 , n69500 , n69501 , n69502 , n69503 , n69504 , n69505 , n69506 , 
 n69507 , n69508 , n69509 , n69510 , n69511 , n69512 , n69513 , n69514 , n69515 , n69516 , 
 n69517 , n69518 , n69519 , n69520 , n69521 , n69522 , n69523 , n69524 , n69525 , n69526 , 
 n69527 , n69528 , n69529 , n69530 , n69531 , n69532 , n69533 , n69534 , n69535 , n69536 , 
 n69537 , n69538 , n69539 , n69540 , n69541 , n69542 , n69543 , n69544 , n69545 , n69546 , 
 n69547 , n69548 , n69549 , n69550 , n69551 , n69552 , n69553 , n69554 , n69555 , n69556 , 
 n69557 , n69558 , n69559 , n69560 , n69561 , n69562 , n69563 , n69564 , n69565 , n69566 , 
 n69567 , n69568 , n69569 , n69570 , n69571 , n69572 , n69573 , n69574 , n69575 , n69576 , 
 n69577 , n69578 , n69579 , n69580 , n69581 , n69582 , n69583 , n69584 , n69585 , n69586 , 
 n69587 , n69588 , n69589 , n69590 , n69591 , n69592 , n69593 , n69594 , n69595 , n69596 , 
 n69597 , n69598 , n69599 , n69600 , n69601 , n69602 , n69603 , n69604 , n69605 , n69606 , 
 n69607 , n69608 , n69609 , n69610 , n69611 , n69612 , n69613 , n69614 , n69615 , n69616 , 
 n69617 , n69618 , n69619 , n69620 , n69621 , n69622 , n69623 , n69624 , n69625 , n69626 , 
 n69627 , n69628 , n69629 , n69630 , n69631 , n69632 , n69633 , n69634 , n69635 , n69636 , 
 n69637 , n69638 , n69639 , n69640 , n69641 , n69642 , n69643 , n69644 , n69645 , n69646 , 
 n69647 , n69648 , n69649 , n69650 , n69651 , n69652 , n69653 , n69654 , n69655 , n69656 , 
 n69657 , n69658 , n69659 , n69660 , n69661 , n69662 , n69663 , n69664 , n69665 , n69666 , 
 n69667 , n69668 , n69669 , n69670 , n69671 , n69672 , n69673 , n69674 , n69675 , n69676 , 
 n69677 , n69678 , n69679 , n69680 , n69681 , n69682 , n69683 , n69684 , n69685 , n69686 , 
 n69687 , n69688 , n69689 , n69690 , n69691 , n69692 , n69693 , n69694 , n69695 , n69696 , 
 n69697 , n69698 , n69699 , n69700 , n69701 , n69702 , n69703 , n69704 , n69705 , n69706 , 
 n69707 , n69708 , n69709 , n69710 , n69711 , n69712 , n69713 , n69714 , n69715 , n69716 , 
 n69717 , n69718 , n69719 , n69720 , n69721 , n69722 , n69723 , n69724 , n69725 , n69726 , 
 n69727 , n69728 , n69729 , n69730 , n69731 , n69732 , n69733 , n69734 , n69735 , n69736 , 
 n69737 , n69738 , n69739 , n69740 , n69741 , n69742 , n69743 , n69744 , n69745 , n69746 , 
 n69747 , n69748 , n69749 , n69750 , n69751 , n69752 , n69753 , n69754 , n69755 , n69756 , 
 n69757 , n69758 , n69759 , n69760 , n69761 , n69762 , n69763 , n69764 , n69765 , n69766 , 
 n69767 , n69768 , n69769 , n69770 , n69771 , n69772 , n69773 , n69774 , n69775 , n69776 , 
 n69777 , n69778 , n69779 , n69780 , n69781 , n69782 , n69783 , n69784 , n69785 , n69786 , 
 n69787 , n69788 , n69789 , n69790 , n69791 , n69792 , n69793 , n69794 , n69795 , n69796 , 
 n69797 , n69798 , n69799 , n69800 , n69801 , n69802 , n69803 , n69804 , n69805 , n69806 , 
 n69807 , n69808 , n69809 , n69810 , n69811 , n69812 , n69813 , n69814 , n69815 , n69816 , 
 n69817 , n69818 , n69819 , n69820 , n69821 , n69822 , n69823 , n69824 , n69825 , n69826 , 
 n69827 , n69828 , n69829 , n69830 , n69831 , n69832 , n69833 , n69834 , n69835 , n69836 , 
 n69837 , n69838 , n69839 , n69840 , n69841 , n69842 , n69843 , n69844 , n69845 , n69846 , 
 n69847 , n69848 , n69849 , n69850 , n69851 , n69852 , n69853 , n69854 , n69855 , n69856 , 
 n69857 , n69858 , n69859 , n69860 , n69861 , n69862 , n69863 , n69864 , n69865 , n69866 , 
 n69867 , n69868 , n69869 , n69870 , n69871 , n69872 , n69873 , n69874 , n69875 , n69876 , 
 n69877 , n69878 , n69879 , n69880 , n69881 , n69882 , n69883 , n69884 , n69885 , n69886 , 
 n69887 , n69888 , n69889 , n69890 , n69891 , n69892 , n69893 , n69894 , n69895 , n69896 , 
 n69897 , n69898 , n69899 , n69900 , n69901 , n69902 , n69903 , n69904 , n69905 , n69906 , 
 n69907 , n69908 , n69909 , n69910 , n69911 , n69912 , n69913 , n69914 , n69915 , n69916 , 
 n69917 , n69918 , n69919 , n69920 , n69921 , n69922 , n69923 , n69924 , n69925 , n69926 , 
 n69927 , n69928 , n69929 , n69930 , n69931 , n69932 , n69933 , n69934 , n69935 , n69936 , 
 n69937 , n69938 , n69939 , n69940 , n69941 , n69942 , n69943 , n69944 , n69945 , n69946 , 
 n69947 , n69948 , n69949 , n69950 , n69951 , n69952 , n69953 , n69954 , n69955 , n69956 , 
 n69957 , n69958 , n69959 , n69960 , n69961 , n69962 , n69963 , n69964 , n69965 , n69966 , 
 n69967 , n69968 , n69969 , n69970 , n69971 , n69972 , n69973 , n69974 , n69975 , n69976 , 
 n69977 , n69978 , n69979 , n69980 , n69981 , n69982 , n69983 , n69984 , n69985 , n69986 , 
 n69987 , n69988 , n69989 , n69990 , n69991 , n69992 , n69993 , n69994 , n69995 , n69996 , 
 n69997 , n69998 , n69999 , n70000 , n70001 , n70002 , n70003 , n70004 , n70005 , n70006 , 
 n70007 , n70008 , n70009 , n70010 , n70011 , n70012 , n70013 , n70014 , n70015 , n70016 , 
 n70017 , n70018 , n70019 , n70020 , n70021 , n70022 , n70023 , n70024 , n70025 , n70026 , 
 n70027 , n70028 , n70029 , n70030 , n70031 , n70032 , n70033 , n70034 , n70035 , n70036 , 
 n70037 , n70038 , n70039 , n70040 , n70041 , n70042 , n70043 , n70044 , n70045 , n70046 , 
 n70047 , n70048 , n70049 , n70050 , n70051 , n70052 , n70053 , n70054 , n70055 , n70056 , 
 n70057 , n70058 , n70059 , n70060 , n70061 , n70062 , n70063 , n70064 , n70065 , n70066 , 
 n70067 , n70068 , n70069 , n70070 , n70071 , n70072 , n70073 , n70074 , n70075 , n70076 , 
 n70077 , n70078 , n70079 , n70080 , n70081 , n70082 , n70083 , n70084 , n70085 , n70086 , 
 n70087 , n70088 , n70089 , n70090 , n70091 , n70092 , n70093 , n70094 , n70095 , n70096 , 
 n70097 , n70098 , n70099 , n70100 , n70101 , n70102 , n70103 , n70104 , n70105 , n70106 , 
 n70107 , n70108 , n70109 , n70110 , n70111 , n70112 , n70113 , n70114 , n70115 , n70116 , 
 n70117 , n70118 , n70119 , n70120 , n70121 , n70122 , n70123 , n70124 , n70125 , n70126 , 
 n70127 , n70128 , n70129 , n70130 , n70131 , n70132 , n70133 , n70134 , n70135 , n70136 , 
 n70137 , n70138 , n70139 , n70140 , n70141 , n70142 , n70143 , n70144 , n70145 , n70146 , 
 n70147 , n70148 , n70149 , n70150 , n70151 , n70152 , n70153 , n70154 , n70155 , n70156 , 
 n70157 , n70158 , n70159 , n70160 , n70161 , n70162 , n70163 , n70164 , n70165 , n70166 , 
 n70167 , n70168 , n70169 , n70170 , n70171 , n70172 , n70173 , n70174 , n70175 , n70176 , 
 n70177 , n70178 , n70179 , n70180 , n70181 , n70182 , n70183 , n70184 , n70185 , n70186 , 
 n70187 , n70188 , n70189 , n70190 , n70191 , n70192 , n70193 , n70194 , n70195 , n70196 , 
 n70197 , n70198 , n70199 , n70200 , n70201 , n70202 , n70203 , n70204 , n70205 , n70206 , 
 n70207 , n70208 , n70209 , n70210 , n70211 , n70212 , n70213 , n70214 , n70215 , n70216 , 
 n70217 , n70218 , n70219 , n70220 , n70221 , n70222 , n70223 , n70224 , n70225 , n70226 , 
 n70227 , n70228 , n70229 , n70230 , n70231 , n70232 , n70233 , n70234 , n70235 , n70236 , 
 n70237 , n70238 , n70239 , n70240 , n70241 , n70242 , n70243 , n70244 , n70245 , n70246 , 
 n70247 , n70248 , n70249 , n70250 , n70251 , n70252 , n70253 , n70254 , n70255 , n70256 , 
 n70257 , n70258 , n70259 , n70260 , n70261 , n70262 , n70263 , n70264 , n70265 , n70266 , 
 n70267 , n70268 , n70269 , n70270 , n70271 , n70272 , n70273 , n70274 , n70275 , n70276 , 
 n70277 , n70278 , n70279 , n70280 , n70281 , n70282 , n70283 , n70284 , n70285 , n70286 , 
 n70287 , n70288 , n70289 , n70290 , n70291 , n70292 , n70293 , n70294 , n70295 , n70296 , 
 n70297 , n70298 , n70299 , n70300 , n70301 , n70302 , n70303 , n70304 , n70305 , n70306 , 
 n70307 , n70308 , n70309 , n70310 , n70311 , n70312 , n70313 , n70314 , n70315 , n70316 , 
 n70317 , n70318 , n70319 , n70320 , n70321 , n70322 , n70323 , n70324 , n70325 , n70326 , 
 n70327 , n70328 , n70329 , n70330 , n70331 , n70332 , n70333 , n70334 , n70335 , n70336 , 
 n70337 , n70338 , n70339 , n70340 , n70341 , n70342 , n70343 , n70344 , n70345 , n70346 , 
 n70347 , n70348 , n70349 , n70350 , n70351 , n70352 , n70353 , n70354 , n70355 , n70356 , 
 n70357 , n70358 , n70359 , n70360 , n70361 , n70362 , n70363 , n70364 , n70365 , n70366 , 
 n70367 , n70368 , n70369 , n70370 , n70371 , n70372 , n70373 , n70374 , n70375 , n70376 , 
 n70377 , n70378 , n70379 , n70380 , n70381 , n70382 , n70383 , n70384 , n70385 , n70386 , 
 n70387 , n70388 , n70389 , n70390 , n70391 , n70392 , n70393 , n70394 , n70395 , n70396 , 
 n70397 , n70398 , n70399 , n70400 , n70401 , n70402 , n70403 , n70404 , n70405 , n70406 , 
 n70407 , n70408 , n70409 , n70410 , n70411 , n70412 , n70413 , n70414 , n70415 , n70416 , 
 n70417 , n70418 , n70419 , n70420 , n70421 , n70422 , n70423 , n70424 , n70425 , n70426 , 
 n70427 , n70428 , n70429 , n70430 , n70431 , n70432 , n70433 , n70434 , n70435 , n70436 , 
 n70437 , n70438 , n70439 , n70440 , n70441 , n70442 , n70443 , n70444 , n70445 , n70446 , 
 n70447 , n70448 , n70449 , n70450 , n70451 , n70452 , n70453 , n70454 , n70455 , n70456 , 
 n70457 , n70458 , n70459 , n70460 , n70461 , n70462 , n70463 , n70464 , n70465 , n70466 , 
 n70467 , n70468 , n70469 , n70470 , n70471 , n70472 , n70473 , n70474 , n70475 , n70476 , 
 n70477 , n70478 , n70479 , n70480 , n70481 , n70482 , n70483 , n70484 , n70485 , n70486 , 
 n70487 , n70488 , n70489 , n70490 , n70491 , n70492 , n70493 , n70494 , n70495 , n70496 , 
 n70497 , n70498 , n70499 , n70500 , n70501 , n70502 , n70503 , n70504 , n70505 , n70506 , 
 n70507 , n70508 , n70509 , n70510 , n70511 , n70512 , n70513 , n70514 , n70515 , n70516 , 
 n70517 , n70518 , n70519 , n70520 , n70521 , n70522 , n70523 , n70524 , n70525 , n70526 , 
 n70527 , n70528 , n70529 , n70530 , n70531 , n70532 , n70533 , n70534 , n70535 , n70536 , 
 n70537 , n70538 , n70539 , n70540 , n70541 , n70542 , n70543 , n70544 , n70545 , n70546 , 
 n70547 , n70548 , n70549 , n70550 , n70551 , n70552 , n70553 , n70554 , n70555 , n70556 , 
 n70557 , n70558 , n70559 , n70560 , n70561 , n70562 , n70563 , n70564 , n70565 , n70566 , 
 n70567 , n70568 , n70569 , n70570 , n70571 , n70572 , n70573 , n70574 , n70575 , n70576 , 
 n70577 , n70578 , n70579 , n70580 , n70581 , n70582 , n70583 , n70584 , n70585 , n70586 , 
 n70587 , n70588 , n70589 , n70590 , n70591 , n70592 , n70593 , n70594 , n70595 , n70596 , 
 n70597 , n70598 , n70599 , n70600 , n70601 , n70602 , n70603 , n70604 , n70605 , n70606 , 
 n70607 , n70608 , n70609 , n70610 , n70611 , n70612 , n70613 , n70614 , n70615 , n70616 , 
 n70617 , n70618 , n70619 , n70620 , n70621 , n70622 , n70623 , n70624 , n70625 , n70626 , 
 n70627 , n70628 , n70629 , n70630 , n70631 , n70632 , n70633 , n70634 , n70635 , n70636 , 
 n70637 , n70638 , n70639 , n70640 , n70641 , n70642 , n70643 , n70644 , n70645 , n70646 , 
 n70647 , n70648 , n70649 , n70650 , n70651 , n70652 , n70653 , n70654 , n70655 , n70656 , 
 n70657 , n70658 , n70659 , n70660 , n70661 , n70662 , n70663 , n70664 , n70665 , n70666 , 
 n70667 , n70668 , n70669 , n70670 , n70671 , n70672 , n70673 , n70674 , n70675 , n70676 , 
 n70677 , n70678 , n70679 , n70680 , n70681 , n70682 , n70683 , n70684 , n70685 , n70686 , 
 n70687 , n70688 , n70689 , n70690 , n70691 , n70692 , n70693 , n70694 , n70695 , n70696 , 
 n70697 , n70698 , n70699 , n70700 , n70701 , n70702 , n70703 , n70704 , n70705 , n70706 , 
 n70707 , n70708 , n70709 , n70710 , n70711 , n70712 , n70713 , n70714 , n70715 , n70716 , 
 n70717 , n70718 , n70719 , n70720 , n70721 , n70722 , n70723 , n70724 , n70725 , n70726 , 
 n70727 , n70728 , n70729 , n70730 , n70731 , n70732 , n70733 , n70734 , n70735 , n70736 , 
 n70737 , n70738 , n70739 , n70740 , n70741 , n70742 , n70743 , n70744 , n70745 , n70746 , 
 n70747 , n70748 , n70749 , n70750 , n70751 , n70752 , n70753 , n70754 , n70755 , n70756 , 
 n70757 , n70758 , n70759 , n70760 , n70761 , n70762 , n70763 , n70764 , n70765 , n70766 , 
 n70767 , n70768 , n70769 , n70770 , n70771 , n70772 , n70773 , n70774 , n70775 , n70776 , 
 n70777 , n70778 , n70779 , n70780 , n70781 , n70782 , n70783 , n70784 , n70785 , n70786 , 
 n70787 , n70788 , n70789 , n70790 , n70791 , n70792 , n70793 , n70794 , n70795 , n70796 , 
 n70797 , n70798 , n70799 , n70800 , n70801 , n70802 , n70803 , n70804 , n70805 , n70806 , 
 n70807 , n70808 , n70809 , n70810 , n70811 , n70812 , n70813 , n70814 , n70815 , n70816 , 
 n70817 , n70818 , n70819 , n70820 , n70821 , n70822 , n70823 , n70824 , n70825 , n70826 , 
 n70827 , n70828 , n70829 , n70830 , n70831 , n70832 , n70833 , n70834 , n70835 , n70836 , 
 n70837 , n70838 , n70839 , n70840 , n70841 , n70842 , n70843 , n70844 , n70845 , n70846 , 
 n70847 , n70848 , n70849 , n70850 , n70851 , n70852 , n70853 , n70854 , n70855 , n70856 , 
 n70857 , n70858 , n70859 , n70860 , n70861 , n70862 , n70863 , n70864 , n70865 , n70866 , 
 n70867 , n70868 , n70869 , n70870 , n70871 , n70872 , n70873 , n70874 , n70875 , n70876 , 
 n70877 , n70878 , n70879 , n70880 , n70881 , n70882 , n70883 , n70884 , n70885 , n70886 , 
 n70887 , n70888 , n70889 , n70890 , n70891 , n70892 , n70893 , n70894 , n70895 , n70896 , 
 n70897 , n70898 , n70899 , n70900 , n70901 , n70902 , n70903 , n70904 , n70905 , n70906 , 
 n70907 , n70908 , n70909 , n70910 , n70911 , n70912 , n70913 , n70914 , n70915 , n70916 , 
 n70917 , n70918 , n70919 , n70920 , n70921 , n70922 , n70923 , n70924 , n70925 , n70926 , 
 n70927 , n70928 , n70929 , n70930 , n70931 , n70932 , n70933 , n70934 , n70935 , n70936 , 
 n70937 , n70938 , n70939 , n70940 , n70941 , n70942 , n70943 , n70944 , n70945 , n70946 , 
 n70947 , n70948 , n70949 , n70950 , n70951 , n70952 , n70953 , n70954 , n70955 , n70956 , 
 n70957 , n70958 , n70959 , n70960 , n70961 , n70962 , n70963 , n70964 , n70965 , n70966 , 
 n70967 , n70968 , n70969 , n70970 , n70971 , n70972 , n70973 , n70974 , n70975 , n70976 , 
 n70977 , n70978 , n70979 , n70980 , n70981 , n70982 , n70983 , n70984 , n70985 , n70986 , 
 n70987 , n70988 , n70989 , n70990 , n70991 , n70992 , n70993 , n70994 , n70995 , n70996 , 
 n70997 , n70998 , n70999 , n71000 , n71001 , n71002 , n71003 , n71004 , n71005 , n71006 , 
 n71007 , n71008 , n71009 , n71010 , n71011 , n71012 , n71013 , n71014 , n71015 , n71016 , 
 n71017 , n71018 , n71019 , n71020 , n71021 , n71022 , n71023 , n71024 , n71025 , n71026 , 
 n71027 , n71028 , n71029 , n71030 , n71031 , n71032 , n71033 , n71034 , n71035 , n71036 , 
 n71037 , n71038 , n71039 , n71040 , n71041 , n71042 , n71043 , n71044 , n71045 , n71046 , 
 n71047 , n71048 , n71049 , n71050 , n71051 , n71052 , n71053 , n71054 , n71055 , n71056 , 
 n71057 , n71058 , n71059 , n71060 , n71061 , n71062 , n71063 , n71064 , n71065 , n71066 , 
 n71067 , n71068 , n71069 , n71070 , n71071 , n71072 , n71073 , n71074 , n71075 , n71076 , 
 n71077 , n71078 , n71079 , n71080 , n71081 , n71082 , n71083 , n71084 , n71085 , n71086 , 
 n71087 , n71088 , n71089 , n71090 , n71091 , n71092 , n71093 , n71094 , n71095 , n71096 , 
 n71097 , n71098 , n71099 , n71100 , n71101 , n71102 , n71103 , n71104 , n71105 , n71106 , 
 n71107 , n71108 , n71109 , n71110 , n71111 , n71112 , n71113 , n71114 , n71115 , n71116 , 
 n71117 , n71118 , n71119 , n71120 , n71121 , n71122 , n71123 , n71124 , n71125 , n71126 , 
 n71127 , n71128 , n71129 , n71130 , n71131 , n71132 , n71133 , n71134 , n71135 , n71136 , 
 n71137 , n71138 , n71139 , n71140 , n71141 , n71142 , n71143 , n71144 , n71145 , n71146 , 
 n71147 , n71148 , n71149 , n71150 , n71151 , n71152 , n71153 , n71154 , n71155 , n71156 , 
 n71157 , n71158 , n71159 , n71160 , n71161 , n71162 , n71163 , n71164 , n71165 , n71166 , 
 n71167 , n71168 , n71169 , n71170 , n71171 , n71172 , n71173 , n71174 , n71175 , n71176 , 
 n71177 , n71178 , n71179 , n71180 , n71181 , n71182 , n71183 , n71184 , n71185 , n71186 , 
 n71187 , n71188 , n71189 , n71190 , n71191 , n71192 , n71193 , n71194 , n71195 , n71196 , 
 n71197 , n71198 , n71199 , n71200 , n71201 , n71202 , n71203 , n71204 , n71205 , n71206 , 
 n71207 , n71208 , n71209 , n71210 , n71211 , n71212 , n71213 , n71214 , n71215 , n71216 , 
 n71217 , n71218 , n71219 , n71220 , n71221 , n71222 , n71223 , n71224 , n71225 , n71226 , 
 n71227 , n71228 , n71229 , n71230 , n71231 , n71232 , n71233 , n71234 , n71235 , n71236 , 
 n71237 , n71238 , n71239 , n71240 , n71241 , n71242 , n71243 , n71244 , n71245 , n71246 , 
 n71247 , n71248 , n71249 , n71250 , n71251 , n71252 , n71253 , n71254 , n71255 , n71256 , 
 n71257 , n71258 , n71259 , n71260 , n71261 , n71262 , n71263 , n71264 , n71265 , n71266 , 
 n71267 , n71268 , n71269 , n71270 , n71271 , n71272 , n71273 , n71274 , n71275 , n71276 , 
 n71277 , n71278 , n71279 , n71280 , n71281 , n71282 , n71283 , n71284 , n71285 , n71286 , 
 n71287 , n71288 , n71289 , n71290 , n71291 , n71292 , n71293 , n71294 , n71295 , n71296 , 
 n71297 , n71298 , n71299 , n71300 , n71301 , n71302 , n71303 , n71304 , n71305 , n71306 , 
 n71307 , n71308 , n71309 , n71310 , n71311 , n71312 , n71313 , n71314 , n71315 , n71316 , 
 n71317 , n71318 , n71319 , n71320 , n71321 , n71322 , n71323 , n71324 , n71325 , n71326 , 
 n71327 , n71328 , n71329 , n71330 , n71331 , n71332 , n71333 , n71334 , n71335 , n71336 , 
 n71337 , n71338 , n71339 , n71340 , n71341 , n71342 , n71343 , n71344 , n71345 , n71346 , 
 n71347 , n71348 , n71349 , n71350 , n71351 , n71352 , n71353 , n71354 , n71355 , n71356 , 
 n71357 , n71358 , n71359 , n71360 , n71361 , n71362 , n71363 , n71364 , n71365 , n71366 , 
 n71367 , n71368 , n71369 , n71370 , n71371 , n71372 , n71373 , n71374 , n71375 , n71376 , 
 n71377 , n71378 , n71379 , n71380 , n71381 , n71382 , n71383 , n71384 , n71385 , n71386 , 
 n71387 , n71388 , n71389 , n71390 , n71391 , n71392 , n71393 , n71394 , n71395 , n71396 , 
 n71397 , n71398 , n71399 , n71400 , n71401 , n71402 , n71403 , n71404 , n71405 , n71406 , 
 n71407 , n71408 , n71409 , n71410 , n71411 , n71412 , n71413 , n71414 , n71415 , n71416 , 
 n71417 , n71418 , n71419 , n71420 , n71421 , n71422 , n71423 , n71424 , n71425 , n71426 , 
 n71427 , n71428 , n71429 , n71430 , n71431 , n71432 , n71433 , n71434 , n71435 , n71436 , 
 n71437 , n71438 , n71439 , n71440 , n71441 , n71442 , n71443 , n71444 , n71445 , n71446 , 
 n71447 , n71448 , n71449 , n71450 , n71451 , n71452 , n71453 , n71454 , n71455 , n71456 , 
 n71457 , n71458 , n71459 , n71460 , n71461 , n71462 , n71463 , n71464 , n71465 , n71466 , 
 n71467 , n71468 , n71469 , n71470 , n71471 , n71472 , n71473 , n71474 , n71475 , n71476 , 
 n71477 , n71478 , n71479 , n71480 , n71481 , n71482 , n71483 , n71484 , n71485 , n71486 , 
 n71487 , n71488 , n71489 , n71490 , n71491 , n71492 , n71493 , n71494 , n71495 , n71496 , 
 n71497 , n71498 , n71499 , n71500 , n71501 , n71502 , n71503 , n71504 , n71505 , n71506 , 
 n71507 , n71508 , n71509 , n71510 , n71511 , n71512 , n71513 , n71514 , n71515 , n71516 , 
 n71517 , n71518 , n71519 , n71520 , n71521 , n71522 , n71523 , n71524 , n71525 , n71526 , 
 n71527 , n71528 , n71529 , n71530 , n71531 , n71532 , n71533 , n71534 , n71535 , n71536 , 
 n71537 , n71538 , n71539 , n71540 , n71541 , n71542 , n71543 , n71544 , n71545 , n71546 , 
 n71547 , n71548 , n71549 , n71550 , n71551 , n71552 , n71553 , n71554 , n71555 , n71556 , 
 n71557 , n71558 , n71559 , n71560 , n71561 , n71562 , n71563 , n71564 , n71565 , n71566 , 
 n71567 , n71568 , n71569 , n71570 , n71571 , n71572 , n71573 , n71574 , n71575 , n71576 , 
 n71577 , n71578 , n71579 , n71580 , n71581 , n71582 , n71583 , n71584 , n71585 , n71586 , 
 n71587 , n71588 , n71589 , n71590 , n71591 , n71592 , n71593 , n71594 , n71595 , n71596 , 
 n71597 , n71598 , n71599 , n71600 , n71601 , n71602 , n71603 , n71604 , n71605 , n71606 , 
 n71607 , n71608 , n71609 , n71610 , n71611 , n71612 , n71613 , n71614 , n71615 , n71616 , 
 n71617 , n71618 , n71619 , n71620 , n71621 , n71622 , n71623 , n71624 , n71625 , n71626 , 
 n71627 , n71628 , n71629 , n71630 , n71631 , n71632 , n71633 , n71634 , n71635 , n71636 , 
 n71637 , n71638 , n71639 , n71640 , n71641 , n71642 , n71643 , n71644 , n71645 , n71646 , 
 n71647 , n71648 , n71649 , n71650 , n71651 , n71652 , n71653 , n71654 , n71655 , n71656 , 
 n71657 , n71658 , n71659 , n71660 , n71661 , n71662 , n71663 , n71664 , n71665 , n71666 , 
 n71667 , n71668 , n71669 , n71670 , n71671 , n71672 , n71673 , n71674 , n71675 , n71676 , 
 n71677 , n71678 , n71679 , n71680 , n71681 , n71682 , n71683 , n71684 , n71685 , n71686 , 
 n71687 , n71688 , n71689 , n71690 , n71691 , n71692 , n71693 , n71694 , n71695 , n71696 , 
 n71697 , n71698 , n71699 , n71700 , n71701 , n71702 , n71703 , n71704 , n71705 , n71706 , 
 n71707 , n71708 , n71709 , n71710 , n71711 , n71712 , n71713 , n71714 , n71715 , n71716 , 
 n71717 , n71718 , n71719 , n71720 , n71721 , n71722 , n71723 , n71724 , n71725 , n71726 , 
 n71727 , n71728 , n71729 , n71730 , n71731 , n71732 , n71733 , n71734 , n71735 , n71736 , 
 n71737 , n71738 , n71739 , n71740 , n71741 , n71742 , n71743 , n71744 , n71745 , n71746 , 
 n71747 , n71748 , n71749 , n71750 , n71751 , n71752 , n71753 , n71754 , n71755 , n71756 , 
 n71757 , n71758 , n71759 , n71760 , n71761 , n71762 , n71763 , n71764 , n71765 , n71766 , 
 n71767 , n71768 , n71769 , n71770 , n71771 , n71772 , n71773 , n71774 , n71775 , n71776 , 
 n71777 , n71778 , n71779 , n71780 , n71781 , n71782 , n71783 , n71784 , n71785 , n71786 , 
 n71787 , n71788 , n71789 , n71790 , n71791 , n71792 , n71793 , n71794 , n71795 , n71796 , 
 n71797 , n71798 , n71799 , n71800 , n71801 , n71802 , n71803 , n71804 , n71805 , n71806 , 
 n71807 , n71808 , n71809 , n71810 , n71811 , n71812 , n71813 , n71814 , n71815 , n71816 , 
 n71817 , n71818 , n71819 , n71820 , n71821 , n71822 , n71823 , n71824 , n71825 , n71826 , 
 n71827 , n71828 , n71829 , n71830 , n71831 , n71832 , n71833 , n71834 , n71835 , n71836 , 
 n71837 , n71838 , n71839 , n71840 , n71841 , n71842 , n71843 , n71844 , n71845 , n71846 , 
 n71847 , n71848 , n71849 , n71850 , n71851 , n71852 , n71853 , n71854 , n71855 , n71856 , 
 n71857 , n71858 , n71859 , n71860 , n71861 , n71862 , n71863 , n71864 , n71865 , n71866 , 
 n71867 , n71868 , n71869 , n71870 , n71871 , n71872 , n71873 , n71874 , n71875 , n71876 , 
 n71877 , n71878 , n71879 , n71880 , n71881 , n71882 , n71883 , n71884 , n71885 , n71886 , 
 n71887 , n71888 , n71889 , n71890 , n71891 , n71892 , n71893 , n71894 , n71895 , n71896 , 
 n71897 , n71898 , n71899 , n71900 , n71901 , n71902 , n71903 , n71904 , n71905 , n71906 , 
 n71907 , n71908 , n71909 , n71910 , n71911 , n71912 , n71913 , n71914 , n71915 , n71916 , 
 n71917 , n71918 , n71919 , n71920 , n71921 , n71922 , n71923 , n71924 , n71925 , n71926 , 
 n71927 , n71928 , n71929 , n71930 , n71931 , n71932 , n71933 , n71934 , n71935 , n71936 , 
 n71937 , n71938 , n71939 , n71940 , n71941 , n71942 , n71943 , n71944 , n71945 , n71946 , 
 n71947 , n71948 , n71949 , n71950 , n71951 , n71952 , n71953 , n71954 , n71955 , n71956 , 
 n71957 , n71958 , n71959 , n71960 , n71961 , n71962 , n71963 , n71964 , n71965 , n71966 , 
 n71967 , n71968 , n71969 , n71970 , n71971 , n71972 , n71973 , n71974 , n71975 , n71976 , 
 n71977 , n71978 , n71979 , n71980 , n71981 , n71982 , n71983 , n71984 , n71985 , n71986 , 
 n71987 , n71988 , n71989 , n71990 , n71991 , n71992 , n71993 , n71994 , n71995 , n71996 , 
 n71997 , n71998 , n71999 , n72000 , n72001 , n72002 , n72003 , n72004 , n72005 , n72006 , 
 n72007 , n72008 , n72009 , n72010 , n72011 , n72012 , n72013 , n72014 , n72015 , n72016 , 
 n72017 , n72018 , n72019 , n72020 , n72021 , n72022 , n72023 , n72024 , n72025 , n72026 , 
 n72027 , n72028 , n72029 , n72030 , n72031 , n72032 , n72033 , n72034 , n72035 , n72036 , 
 n72037 , n72038 , n72039 , n72040 , n72041 , n72042 , n72043 , n72044 , n72045 , n72046 , 
 n72047 , n72048 , n72049 , n72050 , n72051 , n72052 , n72053 , n72054 , n72055 , n72056 , 
 n72057 , n72058 , n72059 , n72060 , n72061 , n72062 , n72063 , n72064 , n72065 , n72066 , 
 n72067 , n72068 , n72069 , n72070 , n72071 , n72072 , n72073 , n72074 , n72075 , n72076 , 
 n72077 , n72078 , n72079 , n72080 , n72081 , n72082 , n72083 , n72084 , n72085 , n72086 , 
 n72087 , n72088 , n72089 , n72090 , n72091 , n72092 , n72093 , n72094 , n72095 , n72096 , 
 n72097 , n72098 , n72099 , n72100 , n72101 , n72102 , n72103 , n72104 , n72105 , n72106 , 
 n72107 , n72108 , n72109 , n72110 , n72111 , n72112 , n72113 , n72114 , n72115 , n72116 , 
 n72117 , n72118 , n72119 , n72120 , n72121 , n72122 , n72123 , n72124 , n72125 , n72126 , 
 n72127 , n72128 , n72129 , n72130 , n72131 , n72132 , n72133 , n72134 , n72135 , n72136 , 
 n72137 , n72138 , n72139 , n72140 , n72141 , n72142 , n72143 , n72144 , n72145 , n72146 , 
 n72147 , n72148 , n72149 , n72150 , n72151 , n72152 , n72153 , n72154 , n72155 , n72156 , 
 n72157 , n72158 , n72159 , n72160 , n72161 , n72162 , n72163 , n72164 , n72165 , n72166 , 
 n72167 , n72168 , n72169 , n72170 , n72171 , n72172 , n72173 , n72174 , n72175 , n72176 , 
 n72177 , n72178 , n72179 , n72180 , n72181 , n72182 , n72183 , n72184 , n72185 , n72186 , 
 n72187 , n72188 , n72189 , n72190 , n72191 , n72192 , n72193 , n72194 , n72195 , n72196 , 
 n72197 , n72198 , n72199 , n72200 , n72201 , n72202 , n72203 , n72204 , n72205 , n72206 , 
 n72207 , n72208 , n72209 , n72210 , n72211 , n72212 , n72213 , n72214 , n72215 , n72216 , 
 n72217 , n72218 , n72219 , n72220 , n72221 , n72222 , n72223 , n72224 , n72225 , n72226 , 
 n72227 , n72228 , n72229 , n72230 , n72231 , n72232 , n72233 , n72234 , n72235 , n72236 , 
 n72237 , n72238 , n72239 , n72240 , n72241 , n72242 , n72243 , n72244 , n72245 , n72246 , 
 n72247 , n72248 , n72249 , n72250 , n72251 , n72252 , n72253 , n72254 , n72255 , n72256 , 
 n72257 , n72258 , n72259 , n72260 , n72261 , n72262 , n72263 , n72264 , n72265 , n72266 , 
 n72267 , n72268 , n72269 , n72270 , n72271 , n72272 , n72273 , n72274 , n72275 , n72276 , 
 n72277 , n72278 , n72279 , n72280 , n72281 , n72282 , n72283 , n72284 , n72285 , n72286 , 
 n72287 , n72288 , n72289 , n72290 , n72291 , n72292 , n72293 , n72294 , n72295 , n72296 , 
 n72297 , n72298 , n72299 , n72300 , n72301 , n72302 , n72303 , n72304 , n72305 , n72306 , 
 n72307 , n72308 , n72309 , n72310 , n72311 , n72312 , n72313 , n72314 , n72315 , n72316 , 
 n72317 , n72318 , n72319 , n72320 , n72321 , n72322 , n72323 , n72324 , n72325 , n72326 , 
 n72327 , n72328 , n72329 , n72330 , n72331 , n72332 , n72333 , n72334 , n72335 , n72336 , 
 n72337 , n72338 , n72339 , n72340 , n72341 , n72342 , n72343 , n72344 , n72345 , n72346 , 
 n72347 , n72348 , n72349 , n72350 , n72351 , n72352 , n72353 , n72354 , n72355 , n72356 , 
 n72357 , n72358 , n72359 , n72360 , n72361 , n72362 , n72363 , n72364 , n72365 , n72366 , 
 n72367 , n72368 , n72369 , n72370 , n72371 , n72372 , n72373 , n72374 , n72375 , n72376 , 
 n72377 , n72378 , n72379 , n72380 , n72381 , n72382 , n72383 , n72384 , n72385 , n72386 , 
 n72387 , n72388 , n72389 , n72390 , n72391 , n72392 , n72393 , n72394 , n72395 , n72396 , 
 n72397 , n72398 , n72399 , n72400 , n72401 , n72402 , n72403 , n72404 , n72405 , n72406 , 
 n72407 , n72408 , n72409 , n72410 , n72411 , n72412 , n72413 , n72414 , n72415 , n72416 , 
 n72417 , n72418 , n72419 , n72420 , n72421 , n72422 , n72423 , n72424 , n72425 , n72426 , 
 n72427 , n72428 , n72429 , n72430 , n72431 , n72432 , n72433 , n72434 , n72435 , n72436 , 
 n72437 , n72438 , n72439 , n72440 , n72441 , n72442 , n72443 , n72444 , n72445 , n72446 , 
 n72447 , n72448 , n72449 , n72450 , n72451 , n72452 , n72453 , n72454 , n72455 , n72456 , 
 n72457 , n72458 , n72459 , n72460 , n72461 , n72462 , n72463 , n72464 , n72465 , n72466 , 
 n72467 , n72468 , n72469 , n72470 , n72471 , n72472 , n72473 , n72474 , n72475 , n72476 , 
 n72477 , n72478 , n72479 , n72480 , n72481 , n72482 , n72483 , n72484 , n72485 , n72486 , 
 n72487 , n72488 , n72489 , n72490 , n72491 , n72492 , n72493 , n72494 , n72495 , n72496 , 
 n72497 , n72498 , n72499 , n72500 , n72501 , n72502 , n72503 , n72504 , n72505 , n72506 , 
 n72507 , n72508 , n72509 , n72510 , n72511 , n72512 , n72513 , n72514 , n72515 , n72516 , 
 n72517 , n72518 , n72519 , n72520 , n72521 , n72522 , n72523 , n72524 , n72525 , n72526 , 
 n72527 , n72528 , n72529 , n72530 , n72531 , n72532 , n72533 , n72534 , n72535 , n72536 , 
 n72537 , n72538 , n72539 , n72540 , n72541 , n72542 , n72543 , n72544 , n72545 , n72546 , 
 n72547 , n72548 , n72549 , n72550 , n72551 , n72552 , n72553 , n72554 , n72555 , n72556 , 
 n72557 , n72558 , n72559 , n72560 , n72561 , n72562 , n72563 , n72564 , n72565 , n72566 , 
 n72567 , n72568 , n72569 , n72570 , n72571 , n72572 , n72573 , n72574 , n72575 , n72576 , 
 n72577 , n72578 , n72579 , n72580 , n72581 , n72582 , n72583 , n72584 , n72585 , n72586 , 
 n72587 , n72588 , n72589 , n72590 , n72591 , n72592 , n72593 , n72594 , n72595 , n72596 , 
 n72597 , n72598 , n72599 , n72600 , n72601 , n72602 , n72603 , n72604 , n72605 , n72606 , 
 n72607 , n72608 , n72609 , n72610 , n72611 , n72612 , n72613 , n72614 , n72615 , n72616 , 
 n72617 , n72618 , n72619 , n72620 , n72621 , n72622 , n72623 , n72624 , n72625 , n72626 , 
 n72627 , n72628 , n72629 , n72630 , n72631 , n72632 , n72633 , n72634 , n72635 , n72636 , 
 n72637 , n72638 , n72639 , n72640 , n72641 , n72642 , n72643 , n72644 , n72645 , n72646 , 
 n72647 , n72648 , n72649 , n72650 , n72651 , n72652 , n72653 , n72654 , n72655 , n72656 , 
 n72657 , n72658 , n72659 , n72660 , n72661 , n72662 , n72663 , n72664 , n72665 , n72666 , 
 n72667 , n72668 , n72669 , n72670 , n72671 , n72672 , n72673 , n72674 , n72675 , n72676 , 
 n72677 , n72678 , n72679 , n72680 , n72681 , n72682 , n72683 , n72684 , n72685 , n72686 , 
 n72687 , n72688 , n72689 , n72690 , n72691 , n72692 , n72693 , n72694 , n72695 , n72696 , 
 n72697 , n72698 , n72699 , n72700 , n72701 , n72702 , n72703 , n72704 , n72705 , n72706 , 
 n72707 , n72708 , n72709 , n72710 , n72711 , n72712 , n72713 , n72714 , n72715 , n72716 , 
 n72717 , n72718 , n72719 , n72720 , n72721 , n72722 , n72723 , n72724 , n72725 , n72726 , 
 n72727 , n72728 , n72729 , n72730 , n72731 , n72732 , n72733 , n72734 , n72735 , n72736 , 
 n72737 , n72738 , n72739 , n72740 , n72741 , n72742 , n72743 , n72744 , n72745 , n72746 , 
 n72747 , n72748 , n72749 , n72750 , n72751 , n72752 , n72753 , n72754 , n72755 , n72756 , 
 n72757 , n72758 , n72759 , n72760 , n72761 , n72762 , n72763 , n72764 , n72765 , n72766 , 
 n72767 , n72768 , n72769 , n72770 , n72771 , n72772 , n72773 , n72774 , n72775 , n72776 , 
 n72777 , n72778 , n72779 , n72780 , n72781 , n72782 , n72783 , n72784 , n72785 , n72786 , 
 n72787 , n72788 , n72789 , n72790 , n72791 , n72792 , n72793 , n72794 , n72795 , n72796 , 
 n72797 , n72798 , n72799 , n72800 , n72801 , n72802 , n72803 , n72804 , n72805 , n72806 , 
 n72807 , n72808 , n72809 , n72810 , n72811 , n72812 , n72813 , n72814 , n72815 , n72816 , 
 n72817 , n72818 , n72819 , n72820 , n72821 , n72822 , n72823 , n72824 , n72825 , n72826 , 
 n72827 , n72828 , n72829 , n72830 , n72831 , n72832 , n72833 , n72834 , n72835 , n72836 , 
 n72837 , n72838 , n72839 , n72840 , n72841 , n72842 , n72843 , n72844 , n72845 , n72846 , 
 n72847 , n72848 , n72849 , n72850 , n72851 , n72852 , n72853 , n72854 , n72855 , n72856 , 
 n72857 , n72858 , n72859 , n72860 , n72861 , n72862 , n72863 , n72864 , n72865 , n72866 , 
 n72867 , n72868 , n72869 , n72870 , n72871 , n72872 , n72873 , n72874 , n72875 , n72876 , 
 n72877 , n72878 , n72879 , n72880 , n72881 , n72882 , n72883 , n72884 , n72885 , n72886 , 
 n72887 , n72888 , n72889 , n72890 , n72891 , n72892 , n72893 , n72894 , n72895 , n72896 , 
 n72897 , n72898 , n72899 , n72900 , n72901 , n72902 , n72903 , n72904 , n72905 , n72906 , 
 n72907 , n72908 , n72909 , n72910 , n72911 , n72912 , n72913 , n72914 , n72915 , n72916 , 
 n72917 , n72918 , n72919 , n72920 , n72921 , n72922 , n72923 , n72924 , n72925 , n72926 , 
 n72927 , n72928 , n72929 , n72930 , n72931 , n72932 , n72933 , n72934 , n72935 , n72936 , 
 n72937 , n72938 , n72939 , n72940 , n72941 , n72942 , n72943 , n72944 , n72945 , n72946 , 
 n72947 , n72948 , n72949 , n72950 , n72951 , n72952 , n72953 , n72954 , n72955 , n72956 , 
 n72957 , n72958 , n72959 , n72960 , n72961 , n72962 , n72963 , n72964 , n72965 , n72966 , 
 n72967 , n72968 , n72969 , n72970 , n72971 , n72972 , n72973 , n72974 , n72975 , n72976 , 
 n72977 , n72978 , n72979 , n72980 , n72981 , n72982 , n72983 , n72984 , n72985 , n72986 , 
 n72987 , n72988 , n72989 , n72990 , n72991 , n72992 , n72993 , n72994 , n72995 , n72996 , 
 n72997 , n72998 , n72999 , n73000 , n73001 , n73002 , n73003 , n73004 , n73005 , n73006 , 
 n73007 , n73008 , n73009 , n73010 , n73011 , n73012 , n73013 , n73014 , n73015 , n73016 , 
 n73017 , n73018 , n73019 , n73020 , n73021 , n73022 , n73023 , n73024 , n73025 , n73026 , 
 n73027 , n73028 , n73029 , n73030 , n73031 , n73032 , n73033 , n73034 , n73035 , n73036 , 
 n73037 , n73038 , n73039 , n73040 , n73041 , n73042 , n73043 , n73044 , n73045 , n73046 , 
 n73047 , n73048 , n73049 , n73050 , n73051 , n73052 , n73053 , n73054 , n73055 , n73056 , 
 n73057 , n73058 , n73059 , n73060 , n73061 , n73062 , n73063 , n73064 , n73065 , n73066 , 
 n73067 , n73068 , n73069 , n73070 , n73071 , n73072 , n73073 , n73074 , n73075 , n73076 , 
 n73077 , n73078 , n73079 , n73080 , n73081 , n73082 , n73083 , n73084 , n73085 , n73086 , 
 n73087 , n73088 , n73089 , n73090 , n73091 , n73092 , n73093 , n73094 , n73095 , n73096 , 
 n73097 , n73098 , n73099 , n73100 , n73101 , n73102 , n73103 , n73104 , n73105 , n73106 , 
 n73107 , n73108 , n73109 , n73110 , n73111 , n73112 , n73113 , n73114 , n73115 , n73116 , 
 n73117 , n73118 , n73119 , n73120 , n73121 , n73122 , n73123 , n73124 , n73125 , n73126 , 
 n73127 , n73128 , n73129 , n73130 , n73131 , n73132 , n73133 , n73134 , n73135 , n73136 , 
 n73137 , n73138 , n73139 , n73140 , n73141 , n73142 , n73143 , n73144 , n73145 , n73146 , 
 n73147 , n73148 , n73149 , n73150 , n73151 , n73152 , n73153 , n73154 , n73155 , n73156 , 
 n73157 , n73158 , n73159 , n73160 , n73161 , n73162 , n73163 , n73164 , n73165 , n73166 , 
 n73167 , n73168 , n73169 , n73170 , n73171 , n73172 , n73173 , n73174 , n73175 , n73176 , 
 n73177 , n73178 , n73179 , n73180 , n73181 , n73182 , n73183 , n73184 , n73185 , n73186 , 
 n73187 , n73188 , n73189 , n73190 , n73191 , n73192 , n73193 , n73194 , n73195 , n73196 , 
 n73197 , n73198 , n73199 , n73200 , n73201 , n73202 , n73203 , n73204 , n73205 , n73206 , 
 n73207 , n73208 , n73209 , n73210 , n73211 , n73212 , n73213 , n73214 , n73215 , n73216 , 
 n73217 , n73218 , n73219 , n73220 , n73221 , n73222 , n73223 , n73224 , n73225 , n73226 , 
 n73227 , n73228 , n73229 , n73230 , n73231 , n73232 , n73233 , n73234 , n73235 , n73236 , 
 n73237 , n73238 , n73239 , n73240 , n73241 , n73242 , n73243 , n73244 , n73245 , n73246 , 
 n73247 , n73248 , n73249 , n73250 , n73251 , n73252 , n73253 , n73254 , n73255 , n73256 , 
 n73257 , n73258 , n73259 , n73260 , n73261 , n73262 , n73263 , n73264 , n73265 , n73266 , 
 n73267 , n73268 , n73269 , n73270 , n73271 , n73272 , n73273 , n73274 , n73275 , n73276 , 
 n73277 , n73278 , n73279 , n73280 , n73281 , n73282 , n73283 , n73284 , n73285 , n73286 , 
 n73287 , n73288 , n73289 , n73290 , n73291 , n73292 , n73293 , n73294 , n73295 , n73296 , 
 n73297 , n73298 , n73299 , n73300 , n73301 , n73302 , n73303 , n73304 , n73305 , n73306 , 
 n73307 , n73308 , n73309 , n73310 , n73311 , n73312 , n73313 , n73314 , n73315 , n73316 , 
 n73317 , n73318 , n73319 , n73320 , n73321 , n73322 , n73323 , n73324 , n73325 , n73326 , 
 n73327 , n73328 , n73329 , n73330 , n73331 , n73332 , n73333 , n73334 , n73335 , n73336 , 
 n73337 , n73338 , n73339 , n73340 , n73341 , n73342 , n73343 , n73344 , n73345 , n73346 , 
 n73347 , n73348 , n73349 , n73350 , n73351 , n73352 , n73353 , n73354 , n73355 , n73356 , 
 n73357 , n73358 , n73359 , n73360 , n73361 , n73362 , n73363 , n73364 , n73365 , n73366 , 
 n73367 , n73368 , n73369 , n73370 , n73371 , n73372 , n73373 , n73374 , n73375 , n73376 , 
 n73377 , n73378 , n73379 , n73380 , n73381 , n73382 , n73383 , n73384 , n73385 , n73386 , 
 n73387 , n73388 , n73389 , n73390 , n73391 , n73392 , n73393 , n73394 , n73395 , n73396 , 
 n73397 , n73398 , n73399 , n73400 , n73401 , n73402 , n73403 , n73404 , n73405 , n73406 , 
 n73407 , n73408 , n73409 , n73410 , n73411 , n73412 , n73413 , n73414 , n73415 , n73416 , 
 n73417 , n73418 , n73419 , n73420 , n73421 , n73422 , n73423 , n73424 , n73425 , n73426 , 
 n73427 , n73428 , n73429 , n73430 , n73431 , n73432 , n73433 , n73434 , n73435 , n73436 , 
 n73437 , n73438 , n73439 , n73440 , n73441 , n73442 , n73443 , n73444 , n73445 , n73446 , 
 n73447 , n73448 , n73449 , n73450 , n73451 , n73452 , n73453 , n73454 , n73455 , n73456 , 
 n73457 , n73458 , n73459 , n73460 , n73461 , n73462 , n73463 , n73464 , n73465 , n73466 , 
 n73467 , n73468 , n73469 , n73470 , n73471 , n73472 , n73473 , n73474 , n73475 , n73476 , 
 n73477 , n73478 , n73479 , n73480 , n73481 , n73482 , n73483 , n73484 , n73485 , n73486 , 
 n73487 , n73488 , n73489 , n73490 , n73491 , n73492 , n73493 , n73494 , n73495 , n73496 , 
 n73497 , n73498 , n73499 , n73500 , n73501 , n73502 , n73503 , n73504 , n73505 , n73506 , 
 n73507 , n73508 , n73509 , n73510 , n73511 , n73512 , n73513 , n73514 , n73515 , n73516 , 
 n73517 , n73518 , n73519 , n73520 , n73521 , n73522 , n73523 , n73524 , n73525 , n73526 , 
 n73527 , n73528 , n73529 , n73530 , n73531 , n73532 , n73533 , n73534 , n73535 , n73536 , 
 n73537 , n73538 , n73539 , n73540 , n73541 , n73542 , n73543 , n73544 , n73545 , n73546 , 
 n73547 , n73548 , n73549 , n73550 , n73551 , n73552 , n73553 , n73554 , n73555 , n73556 , 
 n73557 , n73558 , n73559 , n73560 , n73561 , n73562 , n73563 , n73564 , n73565 , n73566 , 
 n73567 , n73568 , n73569 , n73570 , n73571 , n73572 , n73573 , n73574 , n73575 , n73576 , 
 n73577 , n73578 , n73579 , n73580 , n73581 , n73582 , n73583 , n73584 , n73585 , n73586 , 
 n73587 , n73588 , n73589 , n73590 , n73591 , n73592 , n73593 , n73594 , n73595 , n73596 , 
 n73597 , n73598 , n73599 , n73600 , n73601 , n73602 , n73603 , n73604 , n73605 , n73606 , 
 n73607 , n73608 , n73609 , n73610 , n73611 , n73612 , n73613 , n73614 , n73615 , n73616 , 
 n73617 , n73618 , n73619 , n73620 , n73621 , n73622 , n73623 , n73624 , n73625 , n73626 , 
 n73627 , n73628 , n73629 , n73630 , n73631 , n73632 , n73633 , n73634 , n73635 , n73636 , 
 n73637 , n73638 , n73639 , n73640 , n73641 , n73642 , n73643 , n73644 , n73645 , n73646 , 
 n73647 , n73648 , n73649 , n73650 , n73651 , n73652 , n73653 , n73654 , n73655 , n73656 , 
 n73657 , n73658 , n73659 , n73660 , n73661 , n73662 , n73663 , n73664 , n73665 , n73666 , 
 n73667 , n73668 , n73669 , n73670 , n73671 , n73672 , n73673 , n73674 , n73675 , n73676 , 
 n73677 , n73678 , n73679 , n73680 , n73681 , n73682 , n73683 , n73684 , n73685 , n73686 , 
 n73687 , n73688 , n73689 , n73690 , n73691 , n73692 , n73693 , n73694 , n73695 , n73696 , 
 n73697 , n73698 , n73699 , n73700 , n73701 , n73702 , n73703 , n73704 , n73705 , n73706 , 
 n73707 , n73708 , n73709 , n73710 , n73711 , n73712 , n73713 , n73714 , n73715 , n73716 , 
 n73717 , n73718 , n73719 , n73720 , n73721 , n73722 , n73723 , n73724 , n73725 , n73726 , 
 n73727 , n73728 , n73729 , n73730 , n73731 , n73732 , n73733 , n73734 , n73735 , n73736 , 
 n73737 , n73738 , n73739 , n73740 , n73741 , n73742 , n73743 , n73744 , n73745 , n73746 , 
 n73747 , n73748 , n73749 , n73750 , n73751 , n73752 , n73753 , n73754 , n73755 , n73756 , 
 n73757 , n73758 , n73759 , n73760 , n73761 , n73762 , n73763 , n73764 , n73765 , n73766 , 
 n73767 , n73768 , n73769 , n73770 , n73771 , n73772 , n73773 , n73774 , n73775 , n73776 , 
 n73777 , n73778 , n73779 , n73780 , n73781 , n73782 , n73783 , n73784 , n73785 , n73786 , 
 n73787 , n73788 , n73789 , n73790 , n73791 , n73792 , n73793 , n73794 , n73795 , n73796 , 
 n73797 , n73798 , n73799 , n73800 , n73801 , n73802 , n73803 , n73804 , n73805 , n73806 , 
 n73807 , n73808 , n73809 , n73810 , n73811 , n73812 , n73813 , n73814 , n73815 , n73816 , 
 n73817 , n73818 , n73819 , n73820 , n73821 , n73822 , n73823 , n73824 , n73825 , n73826 , 
 n73827 , n73828 , n73829 , n73830 , n73831 , n73832 , n73833 , n73834 , n73835 , n73836 , 
 n73837 , n73838 , n73839 , n73840 , n73841 , n73842 , n73843 , n73844 , n73845 , n73846 , 
 n73847 , n73848 , n73849 , n73850 , n73851 , n73852 , n73853 , n73854 , n73855 , n73856 , 
 n73857 , n73858 , n73859 , n73860 , n73861 , n73862 , n73863 , n73864 , n73865 , n73866 , 
 n73867 , n73868 , n73869 , n73870 , n73871 , n73872 , n73873 , n73874 , n73875 , n73876 , 
 n73877 , n73878 , n73879 , n73880 , n73881 , n73882 , n73883 , n73884 , n73885 , n73886 , 
 n73887 , n73888 , n73889 , n73890 , n73891 , n73892 , n73893 , n73894 , n73895 , n73896 , 
 n73897 , n73898 , n73899 , n73900 , n73901 , n73902 , n73903 , n73904 , n73905 , n73906 , 
 n73907 , n73908 , n73909 , n73910 , n73911 , n73912 , n73913 , n73914 , n73915 , n73916 , 
 n73917 , n73918 , n73919 , n73920 , n73921 , n73922 , n73923 , n73924 , n73925 , n73926 , 
 n73927 , n73928 , n73929 , n73930 , n73931 , n73932 , n73933 , n73934 , n73935 , n73936 , 
 n73937 , n73938 , n73939 , n73940 , n73941 , n73942 , n73943 , n73944 , n73945 , n73946 , 
 n73947 , n73948 , n73949 , n73950 , n73951 , n73952 , n73953 , n73954 , n73955 , n73956 , 
 n73957 , n73958 , n73959 , n73960 , n73961 , n73962 , n73963 , n73964 , n73965 , n73966 , 
 n73967 , n73968 , n73969 , n73970 , n73971 , n73972 , n73973 , n73974 , n73975 , n73976 , 
 n73977 , n73978 , n73979 , n73980 , n73981 , n73982 , n73983 , n73984 , n73985 , n73986 , 
 n73987 , n73988 , n73989 , n73990 , n73991 , n73992 , n73993 , n73994 , n73995 , n73996 , 
 n73997 , n73998 , n73999 , n74000 , n74001 , n74002 , n74003 , n74004 , n74005 , n74006 , 
 n74007 , n74008 , n74009 , n74010 , n74011 , n74012 , n74013 , n74014 , n74015 , n74016 , 
 n74017 , n74018 , n74019 , n74020 , n74021 , n74022 , n74023 , n74024 , n74025 , n74026 , 
 n74027 , n74028 , n74029 , n74030 , n74031 , n74032 , n74033 , n74034 , n74035 , n74036 , 
 n74037 , n74038 , n74039 , n74040 , n74041 , n74042 , n74043 , n74044 , n74045 , n74046 , 
 n74047 , n74048 , n74049 , n74050 , n74051 , n74052 , n74053 , n74054 , n74055 , n74056 , 
 n74057 , n74058 , n74059 , n74060 , n74061 , n74062 , n74063 , n74064 , n74065 , n74066 , 
 n74067 , n74068 , n74069 , n74070 , n74071 , n74072 , n74073 , n74074 , n74075 , n74076 , 
 n74077 , n74078 , n74079 , n74080 , n74081 , n74082 , n74083 , n74084 , n74085 , n74086 , 
 n74087 , n74088 , n74089 , n74090 , n74091 , n74092 , n74093 , n74094 , n74095 , n74096 , 
 n74097 , n74098 , n74099 , n74100 , n74101 , n74102 , n74103 , n74104 , n74105 , n74106 , 
 n74107 , n74108 , n74109 , n74110 , n74111 , n74112 , n74113 , n74114 , n74115 , n74116 , 
 n74117 , n74118 , n74119 , n74120 , n74121 , n74122 , n74123 , n74124 , n74125 , n74126 , 
 n74127 , n74128 , n74129 , n74130 , n74131 , n74132 , n74133 , n74134 , n74135 , n74136 , 
 n74137 , n74138 , n74139 , n74140 , n74141 , n74142 , n74143 , n74144 , n74145 , n74146 , 
 n74147 , n74148 , n74149 , n74150 , n74151 , n74152 , n74153 , n74154 , n74155 , n74156 , 
 n74157 , n74158 , n74159 , n74160 , n74161 , n74162 , n74163 , n74164 , n74165 , n74166 , 
 n74167 , n74168 , n74169 , n74170 , n74171 , n74172 , n74173 , n74174 , n74175 , n74176 , 
 n74177 , n74178 , n74179 , n74180 , n74181 , n74182 , n74183 , n74184 , n74185 , n74186 , 
 n74187 , n74188 , n74189 , n74190 , n74191 , n74192 , n74193 , n74194 , n74195 , n74196 , 
 n74197 , n74198 , n74199 , n74200 , n74201 , n74202 , n74203 , n74204 , n74205 , n74206 , 
 n74207 , n74208 , n74209 , n74210 , n74211 , n74212 , n74213 , n74214 , n74215 , n74216 , 
 n74217 , n74218 , n74219 , n74220 , n74221 , n74222 , n74223 , n74224 , n74225 , n74226 , 
 n74227 , n74228 , n74229 , n74230 , n74231 , n74232 , n74233 , n74234 , n74235 , n74236 , 
 n74237 , n74238 , n74239 , n74240 , n74241 , n74242 , n74243 , n74244 , n74245 , n74246 , 
 n74247 , n74248 , n74249 , n74250 , n74251 , n74252 , n74253 , n74254 , n74255 , n74256 , 
 n74257 , n74258 , n74259 , n74260 , n74261 , n74262 , n74263 , n74264 , n74265 , n74266 , 
 n74267 , n74268 , n74269 , n74270 , n74271 , n74272 , n74273 , n74274 , n74275 , n74276 , 
 n74277 , n74278 , n74279 , n74280 , n74281 , n74282 , n74283 , n74284 , n74285 , n74286 , 
 n74287 , n74288 , n74289 , n74290 , n74291 , n74292 , n74293 , n74294 , n74295 , n74296 , 
 n74297 , n74298 , n74299 , n74300 , n74301 , n74302 , n74303 , n74304 , n74305 , n74306 , 
 n74307 , n74308 , n74309 , n74310 , n74311 , n74312 , n74313 , n74314 , n74315 , n74316 , 
 n74317 , n74318 , n74319 , n74320 , n74321 , n74322 , n74323 , n74324 , n74325 , n74326 , 
 n74327 , n74328 , n74329 , n74330 , n74331 , n74332 , n74333 , n74334 , n74335 , n74336 , 
 n74337 , n74338 , n74339 , n74340 , n74341 , n74342 , n74343 , n74344 , n74345 , n74346 , 
 n74347 , n74348 , n74349 , n74350 , n74351 , n74352 , n74353 , n74354 , n74355 , n74356 , 
 n74357 , n74358 , n74359 , n74360 , n74361 , n74362 , n74363 , n74364 , n74365 , n74366 , 
 n74367 , n74368 , n74369 , n74370 , n74371 , n74372 , n74373 , n74374 , n74375 , n74376 , 
 n74377 , n74378 , n74379 , n74380 , n74381 , n74382 , n74383 , n74384 , n74385 , n74386 , 
 n74387 , n74388 , n74389 , n74390 , n74391 , n74392 , n74393 , n74394 , n74395 , n74396 , 
 n74397 , n74398 , n74399 , n74400 , n74401 , n74402 , n74403 , n74404 , n74405 , n74406 , 
 n74407 , n74408 , n74409 , n74410 , n74411 , n74412 , n74413 , n74414 , n74415 , n74416 , 
 n74417 , n74418 , n74419 , n74420 , n74421 , n74422 , n74423 , n74424 , n74425 , n74426 , 
 n74427 , n74428 , n74429 , n74430 , n74431 , n74432 , n74433 , n74434 , n74435 , n74436 , 
 n74437 , n74438 , n74439 , n74440 , n74441 , n74442 , n74443 , n74444 , n74445 , n74446 , 
 n74447 , n74448 , n74449 , n74450 , n74451 , n74452 , n74453 , n74454 , n74455 , n74456 , 
 n74457 , n74458 , n74459 , n74460 , n74461 , n74462 , n74463 , n74464 , n74465 , n74466 , 
 n74467 , n74468 , n74469 , n74470 , n74471 , n74472 , n74473 , n74474 , n74475 , n74476 , 
 n74477 , n74478 , n74479 , n74480 , n74481 , n74482 , n74483 , n74484 , n74485 , n74486 , 
 n74487 , n74488 , n74489 , n74490 , n74491 , n74492 , n74493 , n74494 , n74495 , n74496 , 
 n74497 , n74498 , n74499 , n74500 , n74501 , n74502 , n74503 , n74504 , n74505 , n74506 , 
 n74507 , n74508 , n74509 , n74510 , n74511 , n74512 , n74513 , n74514 , n74515 , n74516 , 
 n74517 , n74518 , n74519 , n74520 , n74521 , n74522 , n74523 , n74524 , n74525 , n74526 , 
 n74527 , n74528 , n74529 , n74530 , n74531 , n74532 , n74533 , n74534 , n74535 , n74536 , 
 n74537 , n74538 , n74539 , n74540 , n74541 , n74542 , n74543 , n74544 , n74545 , n74546 , 
 n74547 , n74548 , n74549 , n74550 , n74551 , n74552 , n74553 , n74554 , n74555 , n74556 , 
 n74557 , n74558 , n74559 , n74560 , n74561 , n74562 , n74563 , n74564 , n74565 , n74566 , 
 n74567 , n74568 , n74569 , n74570 , n74571 , n74572 , n74573 , n74574 , n74575 , n74576 , 
 n74577 , n74578 , n74579 , n74580 , n74581 , n74582 , n74583 , n74584 , n74585 , n74586 , 
 n74587 , n74588 , n74589 , n74590 , n74591 , n74592 , n74593 , n74594 , n74595 , n74596 , 
 n74597 , n74598 , n74599 , n74600 , n74601 , n74602 , n74603 , n74604 , n74605 , n74606 , 
 n74607 , n74608 , n74609 , n74610 , n74611 , n74612 , n74613 , n74614 , n74615 , n74616 , 
 n74617 , n74618 , n74619 , n74620 , n74621 , n74622 , n74623 , n74624 , n74625 , n74626 , 
 n74627 , n74628 , n74629 , n74630 , n74631 , n74632 , n74633 , n74634 , n74635 , n74636 , 
 n74637 , n74638 , n74639 , n74640 , n74641 , n74642 , n74643 , n74644 , n74645 , n74646 , 
 n74647 , n74648 , n74649 , n74650 , n74651 , n74652 , n74653 , n74654 , n74655 , n74656 , 
 n74657 , n74658 , n74659 , n74660 , n74661 , n74662 , n74663 , n74664 , n74665 , n74666 , 
 n74667 , n74668 , n74669 , n74670 , n74671 , n74672 , n74673 , n74674 , n74675 , n74676 , 
 n74677 , n74678 , n74679 , n74680 , n74681 , n74682 , n74683 , n74684 , n74685 , n74686 , 
 n74687 , n74688 , n74689 , n74690 , n74691 , n74692 , n74693 , n74694 , n74695 , n74696 , 
 n74697 , n74698 , n74699 , n74700 , n74701 , n74702 , n74703 , n74704 , n74705 , n74706 , 
 n74707 , n74708 , n74709 , n74710 , n74711 , n74712 , n74713 , n74714 , n74715 , n74716 , 
 n74717 , n74718 , n74719 , n74720 , n74721 , n74722 , n74723 , n74724 , n74725 , n74726 , 
 n74727 , n74728 , n74729 , n74730 , n74731 , n74732 , n74733 , n74734 , n74735 , n74736 , 
 n74737 , n74738 , n74739 , n74740 , n74741 , n74742 , n74743 , n74744 , n74745 , n74746 , 
 n74747 , n74748 , n74749 , n74750 , n74751 , n74752 , n74753 , n74754 , n74755 , n74756 , 
 n74757 , n74758 , n74759 , n74760 , n74761 , n74762 , n74763 , n74764 , n74765 , n74766 , 
 n74767 , n74768 , n74769 , n74770 , n74771 , n74772 , n74773 , n74774 , n74775 , n74776 , 
 n74777 , n74778 , n74779 , n74780 , n74781 , n74782 , n74783 , n74784 , n74785 , n74786 , 
 n74787 , n74788 , n74789 , n74790 , n74791 , n74792 , n74793 , n74794 , n74795 , n74796 , 
 n74797 , n74798 , n74799 , n74800 , n74801 , n74802 , n74803 , n74804 , n74805 , n74806 , 
 n74807 , n74808 , n74809 , n74810 , n74811 , n74812 , n74813 , n74814 , n74815 , n74816 , 
 n74817 , n74818 , n74819 , n74820 , n74821 , n74822 , n74823 , n74824 , n74825 , n74826 , 
 n74827 , n74828 , n74829 , n74830 , n74831 , n74832 , n74833 , n74834 , n74835 , n74836 , 
 n74837 , n74838 , n74839 , n74840 , n74841 , n74842 , n74843 , n74844 , n74845 , n74846 , 
 n74847 , n74848 , n74849 , n74850 , n74851 , n74852 , n74853 , n74854 , n74855 , n74856 , 
 n74857 , n74858 , n74859 , n74860 , n74861 , n74862 , n74863 , n74864 , n74865 , n74866 , 
 n74867 , n74868 , n74869 , n74870 , n74871 , n74872 , n74873 , n74874 , n74875 , n74876 , 
 n74877 , n74878 , n74879 , n74880 , n74881 , n74882 , n74883 , n74884 , n74885 , n74886 , 
 n74887 , n74888 , n74889 , n74890 , n74891 , n74892 , n74893 , n74894 , n74895 , n74896 , 
 n74897 , n74898 , n74899 , n74900 , n74901 , n74902 , n74903 , n74904 , n74905 , n74906 , 
 n74907 , n74908 , n74909 , n74910 , n74911 , n74912 , n74913 , n74914 , n74915 , n74916 , 
 n74917 , n74918 , n74919 , n74920 , n74921 , n74922 , n74923 , n74924 , n74925 , n74926 , 
 n74927 , n74928 , n74929 , n74930 , n74931 , n74932 , n74933 , n74934 , n74935 , n74936 , 
 n74937 , n74938 , n74939 , n74940 , n74941 , n74942 , n74943 , n74944 , n74945 , n74946 , 
 n74947 , n74948 , n74949 , n74950 , n74951 , n74952 , n74953 , n74954 , n74955 , n74956 , 
 n74957 , n74958 , n74959 , n74960 , n74961 , n74962 , n74963 , n74964 , n74965 , n74966 , 
 n74967 , n74968 , n74969 , n74970 , n74971 , n74972 , n74973 , n74974 , n74975 , n74976 , 
 n74977 , n74978 , n74979 , n74980 , n74981 , n74982 , n74983 , n74984 , n74985 , n74986 , 
 n74987 , n74988 , n74989 , n74990 , n74991 , n74992 , n74993 , n74994 , n74995 , n74996 , 
 n74997 , n74998 , n74999 , n75000 , n75001 , n75002 , n75003 , n75004 , n75005 , n75006 , 
 n75007 , n75008 , n75009 , n75010 , n75011 , n75012 , n75013 , n75014 , n75015 , n75016 , 
 n75017 , n75018 , n75019 , n75020 , n75021 , n75022 , n75023 , n75024 , n75025 , n75026 , 
 n75027 , n75028 , n75029 , n75030 , n75031 , n75032 , n75033 , n75034 , n75035 , n75036 , 
 n75037 , n75038 , n75039 , n75040 , n75041 , n75042 , n75043 , n75044 , n75045 , n75046 , 
 n75047 , n75048 , n75049 , n75050 , n75051 , n75052 , n75053 , n75054 , n75055 , n75056 , 
 n75057 , n75058 , n75059 , n75060 , n75061 , n75062 , n75063 , n75064 , n75065 , n75066 , 
 n75067 , n75068 , n75069 , n75070 , n75071 , n75072 , n75073 , n75074 , n75075 , n75076 , 
 n75077 , n75078 , n75079 , n75080 , n75081 , n75082 , n75083 , n75084 , n75085 , n75086 , 
 n75087 , n75088 , n75089 , n75090 , n75091 , n75092 , n75093 , n75094 , n75095 , n75096 , 
 n75097 , n75098 , n75099 , n75100 , n75101 , n75102 , n75103 , n75104 , n75105 , n75106 , 
 n75107 , n75108 , n75109 , n75110 , n75111 , n75112 , n75113 , n75114 , n75115 , n75116 , 
 n75117 , n75118 , n75119 , n75120 , n75121 , n75122 , n75123 , n75124 , n75125 , n75126 , 
 n75127 , n75128 , n75129 , n75130 , n75131 , n75132 , n75133 , n75134 , n75135 , n75136 , 
 n75137 , n75138 , n75139 , n75140 , n75141 , n75142 , n75143 , n75144 , n75145 , n75146 , 
 n75147 , n75148 , n75149 , n75150 , n75151 , n75152 , n75153 , n75154 , n75155 , n75156 , 
 n75157 , n75158 , n75159 , n75160 , n75161 , n75162 , n75163 , n75164 , n75165 , n75166 , 
 n75167 , n75168 , n75169 , n75170 , n75171 , n75172 , n75173 , n75174 , n75175 , n75176 , 
 n75177 , n75178 , n75179 , n75180 , n75181 , n75182 , n75183 , n75184 , n75185 , n75186 , 
 n75187 , n75188 , n75189 , n75190 , n75191 , n75192 , n75193 , n75194 , n75195 , n75196 , 
 n75197 , n75198 , n75199 , n75200 , n75201 , n75202 , n75203 , n75204 , n75205 , n75206 , 
 n75207 , n75208 , n75209 , n75210 , n75211 , n75212 , n75213 , n75214 , n75215 , n75216 , 
 n75217 , n75218 , n75219 , n75220 , n75221 , n75222 , n75223 , n75224 , n75225 , n75226 , 
 n75227 , n75228 , n75229 , n75230 , n75231 , n75232 , n75233 , n75234 , n75235 , n75236 , 
 n75237 , n75238 , n75239 , n75240 , n75241 , n75242 , n75243 , n75244 , n75245 , n75246 , 
 n75247 , n75248 , n75249 , n75250 , n75251 , n75252 , n75253 , n75254 , n75255 , n75256 , 
 n75257 , n75258 , n75259 , n75260 , n75261 , n75262 , n75263 , n75264 , n75265 , n75266 , 
 n75267 , n75268 , n75269 , n75270 , n75271 , n75272 , n75273 , n75274 , n75275 , n75276 , 
 n75277 , n75278 , n75279 , n75280 , n75281 , n75282 , n75283 , n75284 , n75285 , n75286 , 
 n75287 , n75288 , n75289 , n75290 , n75291 , n75292 , n75293 , n75294 , n75295 , n75296 , 
 n75297 , n75298 , n75299 , n75300 , n75301 , n75302 , n75303 , n75304 , n75305 , n75306 , 
 n75307 , n75308 , n75309 , n75310 , n75311 , n75312 , n75313 , n75314 , n75315 , n75316 , 
 n75317 , n75318 , n75319 , n75320 , n75321 , n75322 , n75323 , n75324 , n75325 , n75326 , 
 n75327 , n75328 , n75329 , n75330 , n75331 , n75332 , n75333 , n75334 , n75335 , n75336 , 
 n75337 , n75338 , n75339 , n75340 , n75341 , n75342 , n75343 , n75344 , n75345 , n75346 , 
 n75347 , n75348 , n75349 , n75350 , n75351 , n75352 , n75353 , n75354 , n75355 , n75356 , 
 n75357 , n75358 , n75359 , n75360 , n75361 , n75362 , n75363 , n75364 , n75365 , n75366 , 
 n75367 , n75368 , n75369 , n75370 , n75371 , n75372 , n75373 , n75374 , n75375 , n75376 , 
 n75377 , n75378 , n75379 , n75380 , n75381 , n75382 , n75383 , n75384 , n75385 , n75386 , 
 n75387 , n75388 , n75389 , n75390 , n75391 , n75392 , n75393 , n75394 , n75395 , n75396 , 
 n75397 , n75398 , n75399 , n75400 , n75401 , n75402 , n75403 , n75404 , n75405 , n75406 , 
 n75407 , n75408 , n75409 , n75410 , n75411 , n75412 , n75413 , n75414 , n75415 , n75416 , 
 n75417 , n75418 , n75419 , n75420 , n75421 , n75422 , n75423 , n75424 , n75425 , n75426 , 
 n75427 , n75428 , n75429 , n75430 , n75431 , n75432 , n75433 , n75434 , n75435 , n75436 , 
 n75437 , n75438 , n75439 , n75440 , n75441 , n75442 , n75443 , n75444 , n75445 , n75446 , 
 n75447 , n75448 , n75449 , n75450 , n75451 , n75452 , n75453 , n75454 , n75455 , n75456 , 
 n75457 , n75458 , n75459 , n75460 , n75461 , n75462 , n75463 , n75464 , n75465 , n75466 , 
 n75467 , n75468 , n75469 , n75470 , n75471 , n75472 , n75473 , n75474 , n75475 , n75476 , 
 n75477 , n75478 , n75479 , n75480 , n75481 , n75482 , n75483 , n75484 , n75485 , n75486 , 
 n75487 , n75488 , n75489 , n75490 , n75491 , n75492 , n75493 , n75494 , n75495 , n75496 , 
 n75497 , n75498 , n75499 , n75500 , n75501 , n75502 , n75503 , n75504 , n75505 , n75506 , 
 n75507 , n75508 , n75509 , n75510 , n75511 , n75512 , n75513 , n75514 , n75515 , n75516 , 
 n75517 , n75518 , n75519 , n75520 , n75521 , n75522 , n75523 , n75524 , n75525 , n75526 , 
 n75527 , n75528 , n75529 , n75530 , n75531 , n75532 , n75533 , n75534 , n75535 , n75536 , 
 n75537 , n75538 , n75539 , n75540 , n75541 , n75542 , n75543 , n75544 , n75545 , n75546 , 
 n75547 , n75548 , n75549 , n75550 , n75551 , n75552 , n75553 , n75554 , n75555 , n75556 , 
 n75557 , n75558 , n75559 , n75560 , n75561 , n75562 , n75563 , n75564 , n75565 , n75566 , 
 n75567 , n75568 , n75569 , n75570 , n75571 , n75572 , n75573 , n75574 , n75575 , n75576 , 
 n75577 , n75578 , n75579 , n75580 , n75581 , n75582 , n75583 , n75584 , n75585 , n75586 , 
 n75587 , n75588 , n75589 , n75590 , n75591 , n75592 , n75593 , n75594 , n75595 , n75596 , 
 n75597 , n75598 , n75599 , n75600 , n75601 , n75602 , n75603 , n75604 , n75605 , n75606 , 
 n75607 , n75608 , n75609 , n75610 , n75611 , n75612 , n75613 , n75614 , n75615 , n75616 , 
 n75617 , n75618 , n75619 , n75620 , n75621 , n75622 , n75623 , n75624 , n75625 , n75626 , 
 n75627 , n75628 , n75629 , n75630 , n75631 , n75632 , n75633 , n75634 , n75635 , n75636 , 
 n75637 , n75638 , n75639 , n75640 , n75641 , n75642 , n75643 , n75644 , n75645 , n75646 , 
 n75647 , n75648 , n75649 , n75650 , n75651 , n75652 , n75653 , n75654 , n75655 , n75656 , 
 n75657 , n75658 , n75659 , n75660 , n75661 , n75662 , n75663 , n75664 , n75665 , n75666 , 
 n75667 , n75668 , n75669 , n75670 , n75671 , n75672 , n75673 , n75674 , n75675 , n75676 , 
 n75677 , n75678 , n75679 , n75680 , n75681 , n75682 , n75683 , n75684 , n75685 , n75686 , 
 n75687 , n75688 , n75689 , n75690 , n75691 , n75692 , n75693 , n75694 , n75695 , n75696 , 
 n75697 , n75698 , n75699 , n75700 , n75701 , n75702 , n75703 , n75704 , n75705 , n75706 , 
 n75707 , n75708 , n75709 , n75710 , n75711 , n75712 , n75713 , n75714 , n75715 , n75716 , 
 n75717 , n75718 , n75719 , n75720 , n75721 , n75722 , n75723 , n75724 , n75725 , n75726 , 
 n75727 , n75728 , n75729 , n75730 , n75731 , n75732 , n75733 , n75734 , n75735 , n75736 , 
 n75737 , n75738 , n75739 , n75740 , n75741 , n75742 , n75743 , n75744 , n75745 , n75746 , 
 n75747 , n75748 , n75749 , n75750 , n75751 , n75752 , n75753 , n75754 , n75755 , n75756 , 
 n75757 , n75758 , n75759 , n75760 , n75761 , n75762 , n75763 , n75764 , n75765 , n75766 , 
 n75767 , n75768 , n75769 , n75770 , n75771 , n75772 , n75773 , n75774 , n75775 , n75776 , 
 n75777 , n75778 , n75779 , n75780 , n75781 , n75782 , n75783 , n75784 , n75785 , n75786 , 
 n75787 , n75788 , n75789 , n75790 , n75791 , n75792 , n75793 , n75794 , n75795 , n75796 , 
 n75797 , n75798 , n75799 , n75800 , n75801 , n75802 , n75803 , n75804 , n75805 , n75806 , 
 n75807 , n75808 , n75809 , n75810 , n75811 , n75812 , n75813 , n75814 , n75815 , n75816 , 
 n75817 , n75818 , n75819 , n75820 , n75821 , n75822 , n75823 , n75824 , n75825 , n75826 , 
 n75827 , n75828 , n75829 , n75830 , n75831 , n75832 , n75833 , n75834 , n75835 , n75836 , 
 n75837 , n75838 , n75839 , n75840 , n75841 , n75842 , n75843 , n75844 , n75845 , n75846 , 
 n75847 , n75848 , n75849 , n75850 , n75851 , n75852 , n75853 , n75854 , n75855 , n75856 , 
 n75857 , n75858 , n75859 , n75860 , n75861 , n75862 , n75863 , n75864 , n75865 , n75866 , 
 n75867 , n75868 , n75869 , n75870 , n75871 , n75872 , n75873 , n75874 , n75875 , n75876 , 
 n75877 , n75878 , n75879 , n75880 , n75881 , n75882 , n75883 , n75884 , n75885 , n75886 , 
 n75887 , n75888 , n75889 , n75890 , n75891 , n75892 , n75893 , n75894 , n75895 , n75896 , 
 n75897 , n75898 , n75899 , n75900 , n75901 , n75902 , n75903 , n75904 , n75905 , n75906 , 
 n75907 , n75908 , n75909 , n75910 , n75911 , n75912 , n75913 , n75914 , n75915 , n75916 , 
 n75917 , n75918 , n75919 , n75920 , n75921 , n75922 , n75923 , n75924 , n75925 , n75926 , 
 n75927 , n75928 , n75929 , n75930 , n75931 , n75932 , n75933 , n75934 , n75935 , n75936 , 
 n75937 , n75938 , n75939 , n75940 , n75941 , n75942 , n75943 , n75944 , n75945 , n75946 , 
 n75947 , n75948 , n75949 , n75950 , n75951 , n75952 , n75953 , n75954 , n75955 , n75956 , 
 n75957 , n75958 , n75959 , n75960 , n75961 , n75962 , n75963 , n75964 , n75965 , n75966 , 
 n75967 , n75968 , n75969 , n75970 , n75971 , n75972 , n75973 , n75974 , n75975 , n75976 , 
 n75977 , n75978 , n75979 , n75980 , n75981 , n75982 , n75983 , n75984 , n75985 , n75986 , 
 n75987 , n75988 , n75989 , n75990 , n75991 , n75992 , n75993 , n75994 , n75995 , n75996 , 
 n75997 , n75998 , n75999 , n76000 , n76001 , n76002 , n76003 , n76004 , n76005 , n76006 , 
 n76007 , n76008 , n76009 , n76010 , n76011 , n76012 , n76013 , n76014 , n76015 , n76016 , 
 n76017 , n76018 , n76019 , n76020 , n76021 , n76022 , n76023 , n76024 , n76025 , n76026 , 
 n76027 , n76028 , n76029 , n76030 , n76031 , n76032 , n76033 , n76034 , n76035 , n76036 , 
 n76037 , n76038 , n76039 , n76040 , n76041 , n76042 , n76043 , n76044 , n76045 , n76046 , 
 n76047 , n76048 , n76049 , n76050 , n76051 , n76052 , n76053 , n76054 , n76055 , n76056 , 
 n76057 , n76058 , n76059 , n76060 , n76061 , n76062 , n76063 , n76064 , n76065 , n76066 , 
 n76067 , n76068 , n76069 , n76070 , n76071 , n76072 , n76073 , n76074 , n76075 , n76076 , 
 n76077 , n76078 , n76079 , n76080 , n76081 , n76082 , n76083 , n76084 , n76085 , n76086 , 
 n76087 , n76088 , n76089 , n76090 , n76091 , n76092 , n76093 , n76094 , n76095 , n76096 , 
 n76097 , n76098 , n76099 , n76100 , n76101 , n76102 , n76103 , n76104 , n76105 , n76106 , 
 n76107 , n76108 , n76109 , n76110 , n76111 , n76112 , n76113 , n76114 , n76115 , n76116 , 
 n76117 , n76118 , n76119 , n76120 , n76121 , n76122 , n76123 , n76124 , n76125 , n76126 , 
 n76127 , n76128 , n76129 , n76130 , n76131 , n76132 , n76133 , n76134 , n76135 , n76136 , 
 n76137 , n76138 , n76139 , n76140 , n76141 , n76142 , n76143 , n76144 , n76145 , n76146 , 
 n76147 , n76148 , n76149 , n76150 , n76151 , n76152 , n76153 , n76154 , n76155 , n76156 , 
 n76157 , n76158 , n76159 , n76160 , n76161 , n76162 , n76163 , n76164 , n76165 , n76166 , 
 n76167 , n76168 , n76169 , n76170 , n76171 , n76172 , n76173 , n76174 , n76175 , n76176 , 
 n76177 , n76178 , n76179 , n76180 , n76181 , n76182 , n76183 , n76184 , n76185 , n76186 , 
 n76187 , n76188 , n76189 , n76190 , n76191 , n76192 , n76193 , n76194 , n76195 , n76196 , 
 n76197 , n76198 , n76199 , n76200 , n76201 , n76202 , n76203 , n76204 , n76205 , n76206 , 
 n76207 , n76208 , n76209 , n76210 , n76211 , n76212 , n76213 , n76214 , n76215 , n76216 , 
 n76217 , n76218 , n76219 , n76220 , n76221 , n76222 , n76223 , n76224 , n76225 , n76226 , 
 n76227 , n76228 , n76229 , n76230 , n76231 , n76232 , n76233 , n76234 , n76235 , n76236 , 
 n76237 , n76238 , n76239 , n76240 , n76241 , n76242 , n76243 , n76244 , n76245 , n76246 , 
 n76247 , n76248 , n76249 , n76250 , n76251 , n76252 , n76253 , n76254 , n76255 , n76256 , 
 n76257 , n76258 , n76259 , n76260 , n76261 , n76262 , n76263 , n76264 , n76265 , n76266 , 
 n76267 , n76268 , n76269 , n76270 , n76271 , n76272 , n76273 , n76274 , n76275 , n76276 , 
 n76277 , n76278 , n76279 , n76280 , n76281 , n76282 , n76283 , n76284 , n76285 , n76286 , 
 n76287 , n76288 , n76289 , n76290 , n76291 , n76292 , n76293 , n76294 , n76295 , n76296 , 
 n76297 , n76298 , n76299 , n76300 , n76301 , n76302 , n76303 , n76304 , n76305 , n76306 , 
 n76307 , n76308 , n76309 , n76310 , n76311 , n76312 , n76313 , n76314 , n76315 , n76316 , 
 n76317 , n76318 , n76319 , n76320 , n76321 , n76322 , n76323 , n76324 , n76325 , n76326 , 
 n76327 , n76328 , n76329 , n76330 , n76331 , n76332 , n76333 , n76334 , n76335 , n76336 , 
 n76337 , n76338 , n76339 , n76340 , n76341 , n76342 , n76343 , n76344 , n76345 , n76346 , 
 n76347 , n76348 , n76349 , n76350 , n76351 , n76352 , n76353 , n76354 , n76355 , n76356 , 
 n76357 , n76358 , n76359 , n76360 , n76361 , n76362 , n76363 , n76364 , n76365 , n76366 , 
 n76367 , n76368 , n76369 , n76370 , n76371 , n76372 , n76373 , n76374 , n76375 , n76376 , 
 n76377 , n76378 , n76379 , n76380 , n76381 , n76382 , n76383 , n76384 , n76385 , n76386 , 
 n76387 , n76388 , n76389 , n76390 , n76391 , n76392 , n76393 , n76394 , n76395 , n76396 , 
 n76397 , n76398 , n76399 , n76400 , n76401 , n76402 , n76403 , n76404 , n76405 , n76406 , 
 n76407 , n76408 , n76409 , n76410 , n76411 , n76412 , n76413 , n76414 , n76415 , n76416 , 
 n76417 , n76418 , n76419 , n76420 , n76421 , n76422 , n76423 , n76424 , n76425 , n76426 , 
 n76427 , n76428 , n76429 , n76430 , n76431 , n76432 , n76433 , n76434 , n76435 , n76436 , 
 n76437 , n76438 , n76439 , n76440 , n76441 , n76442 , n76443 , n76444 , n76445 , n76446 , 
 n76447 , n76448 , n76449 , n76450 , n76451 , n76452 , n76453 , n76454 , n76455 , n76456 , 
 n76457 , n76458 , n76459 , n76460 , n76461 , n76462 , n76463 , n76464 , n76465 , n76466 , 
 n76467 , n76468 , n76469 , n76470 , n76471 , n76472 , n76473 , n76474 , n76475 , n76476 , 
 n76477 , n76478 , n76479 , n76480 , n76481 , n76482 , n76483 , n76484 , n76485 , n76486 , 
 n76487 , n76488 , n76489 , n76490 , n76491 , n76492 , n76493 , n76494 , n76495 , n76496 , 
 n76497 , n76498 , n76499 , n76500 , n76501 , n76502 , n76503 , n76504 , n76505 , n76506 , 
 n76507 , n76508 , n76509 , n76510 , n76511 , n76512 , n76513 , n76514 , n76515 , n76516 , 
 n76517 , n76518 , n76519 , n76520 , n76521 , n76522 , n76523 , n76524 , n76525 , n76526 , 
 n76527 , n76528 , n76529 , n76530 , n76531 , n76532 , n76533 , n76534 , n76535 , n76536 , 
 n76537 , n76538 , n76539 , n76540 , n76541 , n76542 , n76543 , n76544 , n76545 , n76546 , 
 n76547 , n76548 , n76549 , n76550 , n76551 , n76552 , n76553 , n76554 , n76555 , n76556 , 
 n76557 , n76558 , n76559 , n76560 , n76561 , n76562 , n76563 , n76564 , n76565 , n76566 , 
 n76567 , n76568 , n76569 , n76570 , n76571 , n76572 , n76573 , n76574 , n76575 , n76576 , 
 n76577 , n76578 , n76579 , n76580 , n76581 , n76582 , n76583 , n76584 , n76585 , n76586 , 
 n76587 , n76588 , n76589 , n76590 , n76591 , n76592 , n76593 , n76594 , n76595 , n76596 , 
 n76597 , n76598 , n76599 , n76600 , n76601 , n76602 , n76603 , n76604 , n76605 , n76606 , 
 n76607 , n76608 , n76609 , n76610 , n76611 , n76612 , n76613 , n76614 , n76615 , n76616 , 
 n76617 , n76618 , n76619 , n76620 , n76621 , n76622 , n76623 , n76624 , n76625 , n76626 , 
 n76627 , n76628 , n76629 , n76630 , n76631 , n76632 , n76633 , n76634 , n76635 , n76636 , 
 n76637 , n76638 , n76639 , n76640 , n76641 , n76642 , n76643 , n76644 , n76645 , n76646 , 
 n76647 , n76648 , n76649 , n76650 , n76651 , n76652 , n76653 , n76654 , n76655 , n76656 , 
 n76657 , n76658 , n76659 , n76660 , n76661 , n76662 , n76663 , n76664 , n76665 , n76666 , 
 n76667 , n76668 , n76669 , n76670 , n76671 , n76672 , n76673 , n76674 , n76675 , n76676 , 
 n76677 , n76678 , n76679 , n76680 , n76681 , n76682 , n76683 , n76684 , n76685 , n76686 , 
 n76687 , n76688 , n76689 , n76690 , n76691 , n76692 , n76693 , n76694 , n76695 , n76696 , 
 n76697 , n76698 , n76699 , n76700 , n76701 , n76702 , n76703 , n76704 , n76705 , n76706 , 
 n76707 , n76708 , n76709 , n76710 , n76711 , n76712 , n76713 , n76714 , n76715 , n76716 , 
 n76717 , n76718 , n76719 , n76720 , n76721 , n76722 , n76723 , n76724 , n76725 , n76726 , 
 n76727 , n76728 , n76729 , n76730 , n76731 , n76732 , n76733 , n76734 , n76735 , n76736 , 
 n76737 , n76738 , n76739 , n76740 , n76741 , n76742 , n76743 , n76744 , n76745 , n76746 , 
 n76747 , n76748 , n76749 , n76750 , n76751 , n76752 , n76753 , n76754 , n76755 , n76756 , 
 n76757 , n76758 , n76759 , n76760 , n76761 , n76762 , n76763 , n76764 , n76765 , n76766 , 
 n76767 , n76768 , n76769 , n76770 , n76771 , n76772 , n76773 , n76774 , n76775 , n76776 , 
 n76777 , n76778 , n76779 , n76780 , n76781 , n76782 , n76783 , n76784 , n76785 , n76786 , 
 n76787 , n76788 , n76789 , n76790 , n76791 , n76792 , n76793 , n76794 , n76795 , n76796 , 
 n76797 , n76798 , n76799 , n76800 , n76801 , n76802 , n76803 , n76804 , n76805 , n76806 , 
 n76807 , n76808 , n76809 , n76810 , n76811 , n76812 , n76813 , n76814 , n76815 , n76816 , 
 n76817 , n76818 , n76819 , n76820 , n76821 , n76822 , n76823 , n76824 , n76825 , n76826 , 
 n76827 , n76828 , n76829 , n76830 , n76831 , n76832 , n76833 , n76834 , n76835 , n76836 , 
 n76837 , n76838 , n76839 , n76840 , n76841 , n76842 , n76843 , n76844 , n76845 , n76846 , 
 n76847 , n76848 , n76849 , n76850 , n76851 , n76852 , n76853 , n76854 , n76855 , n76856 , 
 n76857 , n76858 , n76859 , n76860 , n76861 , n76862 , n76863 , n76864 , n76865 , n76866 , 
 n76867 , n76868 , n76869 , n76870 , n76871 , n76872 , n76873 , n76874 , n76875 , n76876 , 
 n76877 , n76878 , n76879 , n76880 , n76881 , n76882 , n76883 , n76884 , n76885 , n76886 , 
 n76887 , n76888 , n76889 , n76890 , n76891 , n76892 , n76893 , n76894 , n76895 , n76896 , 
 n76897 , n76898 , n76899 , n76900 , n76901 , n76902 , n76903 , n76904 , n76905 , n76906 , 
 n76907 , n76908 , n76909 , n76910 , n76911 , n76912 , n76913 , n76914 , n76915 , n76916 , 
 n76917 , n76918 , n76919 , n76920 , n76921 , n76922 , n76923 , n76924 , n76925 , n76926 , 
 n76927 , n76928 , n76929 , n76930 , n76931 , n76932 , n76933 , n76934 , n76935 , n76936 , 
 n76937 , n76938 , n76939 , n76940 , n76941 , n76942 , n76943 , n76944 , n76945 , n76946 , 
 n76947 , n76948 , n76949 , n76950 , n76951 , n76952 , n76953 , n76954 , n76955 , n76956 , 
 n76957 , n76958 , n76959 , n76960 , n76961 , n76962 , n76963 , n76964 , n76965 , n76966 , 
 n76967 , n76968 , n76969 , n76970 , n76971 , n76972 , n76973 , n76974 , n76975 , n76976 , 
 n76977 , n76978 , n76979 , n76980 , n76981 , n76982 , n76983 , n76984 , n76985 , n76986 , 
 n76987 , n76988 , n76989 , n76990 , n76991 , n76992 , n76993 , n76994 , n76995 , n76996 , 
 n76997 , n76998 , n76999 , n77000 , n77001 , n77002 , n77003 , n77004 , n77005 , n77006 , 
 n77007 , n77008 , n77009 , n77010 , n77011 , n77012 , n77013 , n77014 , n77015 , n77016 , 
 n77017 , n77018 , n77019 , n77020 , n77021 , n77022 , n77023 , n77024 , n77025 , n77026 , 
 n77027 , n77028 , n77029 , n77030 , n77031 , n77032 , n77033 , n77034 , n77035 , n77036 , 
 n77037 , n77038 , n77039 , n77040 , n77041 , n77042 , n77043 , n77044 , n77045 , n77046 , 
 n77047 , n77048 , n77049 , n77050 , n77051 , n77052 , n77053 , n77054 , n77055 , n77056 , 
 n77057 , n77058 , n77059 , n77060 , n77061 , n77062 , n77063 , n77064 , n77065 , n77066 , 
 n77067 , n77068 , n77069 , n77070 , n77071 , n77072 , n77073 , n77074 , n77075 , n77076 , 
 n77077 , n77078 , n77079 , n77080 , n77081 , n77082 , n77083 , n77084 , n77085 , n77086 , 
 n77087 , n77088 , n77089 , n77090 , n77091 , n77092 , n77093 , n77094 , n77095 , n77096 , 
 n77097 , n77098 , n77099 , n77100 , n77101 , n77102 , n77103 , n77104 , n77105 , n77106 , 
 n77107 , n77108 , n77109 , n77110 , n77111 , n77112 , n77113 , n77114 , n77115 , n77116 , 
 n77117 , n77118 , n77119 , n77120 , n77121 , n77122 , n77123 , n77124 , n77125 , n77126 , 
 n77127 , n77128 , n77129 , n77130 , n77131 , n77132 , n77133 , n77134 , n77135 , n77136 , 
 n77137 , n77138 , n77139 , n77140 , n77141 , n77142 , n77143 , n77144 , n77145 , n77146 , 
 n77147 , n77148 , n77149 , n77150 , n77151 , n77152 , n77153 , n77154 , n77155 , n77156 , 
 n77157 , n77158 , n77159 , n77160 , n77161 , n77162 , n77163 , n77164 , n77165 , n77166 , 
 n77167 , n77168 , n77169 , n77170 , n77171 , n77172 , n77173 , n77174 , n77175 , n77176 , 
 n77177 , n77178 , n77179 , n77180 , n77181 , n77182 , n77183 , n77184 , n77185 , n77186 , 
 n77187 , n77188 , n77189 , n77190 , n77191 , n77192 , n77193 , n77194 , n77195 , n77196 , 
 n77197 , n77198 , n77199 , n77200 , n77201 , n77202 , n77203 , n77204 , n77205 , n77206 , 
 n77207 , n77208 , n77209 , n77210 , n77211 , n77212 , n77213 , n77214 , n77215 , n77216 , 
 n77217 , n77218 , n77219 , n77220 , n77221 , n77222 , n77223 , n77224 , n77225 , n77226 , 
 n77227 , n77228 , n77229 , n77230 , n77231 , n77232 , n77233 , n77234 , n77235 , n77236 , 
 n77237 , n77238 , n77239 , n77240 , n77241 , n77242 , n77243 , n77244 , n77245 , n77246 , 
 n77247 , n77248 , n77249 , n77250 , n77251 , n77252 , n77253 , n77254 , n77255 , n77256 , 
 n77257 , n77258 , n77259 , n77260 , n77261 , n77262 , n77263 , n77264 , n77265 , n77266 , 
 n77267 , n77268 , n77269 , n77270 , n77271 , n77272 , n77273 , n77274 , n77275 , n77276 , 
 n77277 , n77278 , n77279 , n77280 , n77281 , n77282 , n77283 , n77284 , n77285 , n77286 , 
 n77287 , n77288 , n77289 , n77290 , n77291 , n77292 , n77293 , n77294 , n77295 , n77296 , 
 n77297 , n77298 , n77299 , n77300 , n77301 , n77302 , n77303 , n77304 , n77305 , n77306 , 
 n77307 , n77308 , n77309 , n77310 , n77311 , n77312 , n77313 , n77314 , n77315 , n77316 , 
 n77317 , n77318 , n77319 , n77320 , n77321 , n77322 , n77323 , n77324 , n77325 , n77326 , 
 n77327 , n77328 , n77329 , n77330 , n77331 , n77332 , n77333 , n77334 , n77335 , n77336 , 
 n77337 , n77338 , n77339 , n77340 , n77341 , n77342 , n77343 , n77344 , n77345 , n77346 , 
 n77347 , n77348 , n77349 , n77350 , n77351 , n77352 , n77353 , n77354 , n77355 , n77356 , 
 n77357 , n77358 , n77359 , n77360 , n77361 , n77362 , n77363 , n77364 , n77365 , n77366 , 
 n77367 , n77368 , n77369 , n77370 , n77371 , n77372 , n77373 , n77374 , n77375 , n77376 , 
 n77377 , n77378 , n77379 , n77380 , n77381 , n77382 , n77383 , n77384 , n77385 , n77386 , 
 n77387 , n77388 , n77389 , n77390 , n77391 , n77392 , n77393 , n77394 , n77395 , n77396 , 
 n77397 , n77398 , n77399 , n77400 , n77401 , n77402 , n77403 , n77404 , n77405 , n77406 , 
 n77407 , n77408 , n77409 , n77410 , n77411 , n77412 , n77413 , n77414 , n77415 , n77416 , 
 n77417 , n77418 , n77419 , n77420 , n77421 , n77422 , n77423 , n77424 , n77425 , n77426 , 
 n77427 , n77428 , n77429 , n77430 , n77431 , n77432 , n77433 , n77434 , n77435 , n77436 , 
 n77437 , n77438 , n77439 , n77440 , n77441 , n77442 , n77443 , n77444 , n77445 , n77446 , 
 n77447 , n77448 , n77449 , n77450 , n77451 , n77452 , n77453 , n77454 , n77455 , n77456 , 
 n77457 , n77458 , n77459 , n77460 , n77461 , n77462 , n77463 , n77464 , n77465 , n77466 , 
 n77467 , n77468 , n77469 , n77470 , n77471 , n77472 , n77473 , n77474 , n77475 , n77476 , 
 n77477 , n77478 , n77479 , n77480 , n77481 , n77482 , n77483 , n77484 , n77485 , n77486 , 
 n77487 , n77488 , n77489 , n77490 , n77491 , n77492 , n77493 , n77494 , n77495 , n77496 , 
 n77497 , n77498 , n77499 , n77500 , n77501 , n77502 , n77503 , n77504 , n77505 , n77506 , 
 n77507 , n77508 , n77509 , n77510 , n77511 , n77512 , n77513 , n77514 , n77515 , n77516 , 
 n77517 , n77518 , n77519 , n77520 , n77521 , n77522 , n77523 , n77524 , n77525 , n77526 , 
 n77527 , n77528 , n77529 , n77530 , n77531 , n77532 , n77533 , n77534 , n77535 , n77536 , 
 n77537 , n77538 , n77539 , n77540 , n77541 , n77542 , n77543 , n77544 , n77545 , n77546 , 
 n77547 , n77548 , n77549 , n77550 , n77551 , n77552 , n77553 , n77554 , n77555 , n77556 , 
 n77557 , n77558 , n77559 , n77560 , n77561 , n77562 , n77563 , n77564 , n77565 , n77566 , 
 n77567 , n77568 , n77569 , n77570 , n77571 , n77572 , n77573 , n77574 , n77575 , n77576 , 
 n77577 , n77578 , n77579 , n77580 , n77581 , n77582 , n77583 , n77584 , n77585 , n77586 , 
 n77587 , n77588 , n77589 , n77590 , n77591 , n77592 , n77593 , n77594 , n77595 , n77596 , 
 n77597 , n77598 , n77599 , n77600 , n77601 , n77602 , n77603 , n77604 , n77605 , n77606 , 
 n77607 , n77608 , n77609 , n77610 , n77611 , n77612 , n77613 , n77614 , n77615 , n77616 , 
 n77617 , n77618 , n77619 , n77620 , n77621 , n77622 , n77623 , n77624 , n77625 , n77626 , 
 n77627 , n77628 , n77629 , n77630 , n77631 , n77632 , n77633 , n77634 , n77635 , n77636 , 
 n77637 , n77638 , n77639 , n77640 , n77641 , n77642 , n77643 , n77644 , n77645 , n77646 , 
 n77647 , n77648 , n77649 , n77650 , n77651 , n77652 , n77653 , n77654 , n77655 , n77656 , 
 n77657 , n77658 , n77659 , n77660 , n77661 , n77662 , n77663 , n77664 , n77665 , n77666 , 
 n77667 , n77668 , n77669 , n77670 , n77671 , n77672 , n77673 , n77674 , n77675 , n77676 , 
 n77677 , n77678 , n77679 , n77680 , n77681 , n77682 , n77683 , n77684 , n77685 , n77686 , 
 n77687 , n77688 , n77689 , n77690 , n77691 , n77692 , n77693 , n77694 , n77695 , n77696 , 
 n77697 , n77698 , n77699 , n77700 , n77701 , n77702 , n77703 , n77704 , n77705 , n77706 , 
 n77707 , n77708 , n77709 , n77710 , n77711 , n77712 , n77713 , n77714 , n77715 , n77716 , 
 n77717 , n77718 , n77719 , n77720 , n77721 , n77722 , n77723 , n77724 , n77725 , n77726 , 
 n77727 , n77728 , n77729 , n77730 , n77731 , n77732 , n77733 , n77734 , n77735 , n77736 , 
 n77737 , n77738 , n77739 , n77740 , n77741 , n77742 , n77743 , n77744 , n77745 , n77746 , 
 n77747 , n77748 , n77749 , n77750 , n77751 , n77752 , n77753 , n77754 , n77755 , n77756 , 
 n77757 , n77758 , n77759 , n77760 , n77761 , n77762 , n77763 , n77764 , n77765 , n77766 , 
 n77767 , n77768 , n77769 , n77770 , n77771 , n77772 , n77773 , n77774 , n77775 , n77776 , 
 n77777 , n77778 , n77779 , n77780 , n77781 , n77782 , n77783 , n77784 , n77785 , n77786 , 
 n77787 , n77788 , n77789 , n77790 , n77791 , n77792 , n77793 , n77794 , n77795 , n77796 , 
 n77797 , n77798 , n77799 , n77800 , n77801 , n77802 , n77803 , n77804 , n77805 , n77806 , 
 n77807 , n77808 , n77809 , n77810 , n77811 , n77812 , n77813 , n77814 , n77815 , n77816 , 
 n77817 , n77818 , n77819 , n77820 , n77821 , n77822 , n77823 , n77824 , n77825 , n77826 , 
 n77827 , n77828 , n77829 , n77830 , n77831 , n77832 , n77833 , n77834 , n77835 , n77836 , 
 n77837 , n77838 , n77839 , n77840 , n77841 , n77842 , n77843 , n77844 , n77845 , n77846 , 
 n77847 , n77848 , n77849 , n77850 , n77851 , n77852 , n77853 , n77854 , n77855 , n77856 , 
 n77857 , n77858 , n77859 , n77860 , n77861 , n77862 , n77863 , n77864 , n77865 , n77866 , 
 n77867 , n77868 , n77869 , n77870 , n77871 , n77872 , n77873 , n77874 , n77875 , n77876 , 
 n77877 , n77878 , n77879 , n77880 , n77881 , n77882 , n77883 , n77884 , n77885 , n77886 , 
 n77887 , n77888 , n77889 , n77890 , n77891 , n77892 , n77893 , n77894 , n77895 , n77896 , 
 n77897 , n77898 , n77899 , n77900 , n77901 , n77902 , n77903 , n77904 , n77905 , n77906 , 
 n77907 , n77908 , n77909 , n77910 , n77911 , n77912 , n77913 , n77914 , n77915 , n77916 , 
 n77917 , n77918 , n77919 , n77920 , n77921 , n77922 , n77923 , n77924 , n77925 , n77926 , 
 n77927 , n77928 , n77929 , n77930 , n77931 , n77932 , n77933 , n77934 , n77935 , n77936 , 
 n77937 , n77938 , n77939 , n77940 , n77941 , n77942 , n77943 , n77944 , n77945 , n77946 , 
 n77947 , n77948 , n77949 , n77950 , n77951 , n77952 , n77953 , n77954 , n77955 , n77956 , 
 n77957 , n77958 , n77959 , n77960 , n77961 , n77962 , n77963 , n77964 , n77965 , n77966 , 
 n77967 , n77968 , n77969 , n77970 , n77971 , n77972 , n77973 , n77974 , n77975 , n77976 , 
 n77977 , n77978 , n77979 , n77980 , n77981 , n77982 , n77983 , n77984 , n77985 , n77986 , 
 n77987 , n77988 , n77989 , n77990 , n77991 , n77992 , n77993 , n77994 , n77995 , n77996 , 
 n77997 , n77998 , n77999 , n78000 , n78001 , n78002 , n78003 , n78004 , n78005 , n78006 , 
 n78007 , n78008 , n78009 , n78010 , n78011 , n78012 , n78013 , n78014 , n78015 , n78016 , 
 n78017 , n78018 , n78019 , n78020 , n78021 , n78022 , n78023 , n78024 , n78025 , n78026 , 
 n78027 , n78028 , n78029 , n78030 , n78031 , n78032 , n78033 , n78034 , n78035 , n78036 , 
 n78037 , n78038 , n78039 , n78040 , n78041 , n78042 , n78043 , n78044 , n78045 , n78046 , 
 n78047 , n78048 , n78049 , n78050 , n78051 , n78052 , n78053 , n78054 , n78055 , n78056 , 
 n78057 , n78058 , n78059 , n78060 , n78061 , n78062 , n78063 , n78064 , n78065 , n78066 , 
 n78067 , n78068 , n78069 , n78070 , n78071 , n78072 , n78073 , n78074 , n78075 , n78076 , 
 n78077 , n78078 , n78079 , n78080 , n78081 , n78082 , n78083 , n78084 , n78085 , n78086 , 
 n78087 , n78088 , n78089 , n78090 , n78091 , n78092 , n78093 , n78094 , n78095 , n78096 , 
 n78097 , n78098 , n78099 , n78100 , n78101 , n78102 , n78103 , n78104 , n78105 , n78106 , 
 n78107 , n78108 , n78109 , n78110 , n78111 , n78112 , n78113 , n78114 , n78115 , n78116 , 
 n78117 , n78118 , n78119 , n78120 , n78121 , n78122 , n78123 , n78124 , n78125 , n78126 , 
 n78127 , n78128 , n78129 , n78130 , n78131 , n78132 , n78133 , n78134 , n78135 , n78136 , 
 n78137 , n78138 , n78139 , n78140 , n78141 , n78142 , n78143 , n78144 , n78145 , n78146 , 
 n78147 , n78148 , n78149 , n78150 , n78151 , n78152 , n78153 , n78154 , n78155 , n78156 , 
 n78157 , n78158 , n78159 , n78160 , n78161 , n78162 , n78163 , n78164 , n78165 , n78166 , 
 n78167 , n78168 , n78169 , n78170 , n78171 , n78172 , n78173 , n78174 , n78175 , n78176 , 
 n78177 , n78178 , n78179 , n78180 , n78181 , n78182 , n78183 , n78184 , n78185 , n78186 , 
 n78187 , n78188 , n78189 , n78190 , n78191 , n78192 , n78193 , n78194 , n78195 , n78196 , 
 n78197 , n78198 , n78199 , n78200 , n78201 , n78202 , n78203 , n78204 , n78205 , n78206 , 
 n78207 , n78208 , n78209 , n78210 , n78211 , n78212 , n78213 , n78214 , n78215 , n78216 , 
 n78217 , n78218 , n78219 , n78220 , n78221 , n78222 , n78223 , n78224 , n78225 , n78226 , 
 n78227 , n78228 , n78229 , n78230 , n78231 , n78232 , n78233 , n78234 , n78235 , n78236 , 
 n78237 , n78238 , n78239 , n78240 , n78241 , n78242 , n78243 , n78244 , n78245 , n78246 , 
 n78247 , n78248 , n78249 , n78250 , n78251 , n78252 , n78253 , n78254 , n78255 , n78256 , 
 n78257 , n78258 , n78259 , n78260 , n78261 , n78262 , n78263 , n78264 , n78265 , n78266 , 
 n78267 , n78268 , n78269 , n78270 , n78271 , n78272 , n78273 , n78274 , n78275 , n78276 , 
 n78277 , n78278 , n78279 , n78280 , n78281 , n78282 , n78283 , n78284 , n78285 , n78286 , 
 n78287 , n78288 , n78289 , n78290 , n78291 , n78292 , n78293 , n78294 , n78295 , n78296 , 
 n78297 , n78298 , n78299 , n78300 , n78301 , n78302 , n78303 , n78304 , n78305 , n78306 , 
 n78307 , n78308 , n78309 , n78310 , n78311 , n78312 , n78313 , n78314 , n78315 , n78316 , 
 n78317 , n78318 , n78319 , n78320 , n78321 , n78322 , n78323 , n78324 , n78325 , n78326 , 
 n78327 , n78328 , n78329 , n78330 , n78331 , n78332 , n78333 , n78334 , n78335 , n78336 , 
 n78337 , n78338 , n78339 , n78340 , n78341 , n78342 , n78343 , n78344 , n78345 , n78346 , 
 n78347 , n78348 , n78349 , n78350 , n78351 , n78352 , n78353 , n78354 , n78355 , n78356 , 
 n78357 , n78358 , n78359 , n78360 , n78361 , n78362 , n78363 , n78364 , n78365 , n78366 , 
 n78367 , n78368 , n78369 , n78370 , n78371 , n78372 , n78373 , n78374 , n78375 , n78376 , 
 n78377 , n78378 , n78379 , n78380 , n78381 , n78382 , n78383 , n78384 , n78385 , n78386 , 
 n78387 , n78388 , n78389 , n78390 , n78391 , n78392 , n78393 , n78394 , n78395 , n78396 , 
 n78397 , n78398 , n78399 , n78400 , n78401 , n78402 , n78403 , n78404 , n78405 , n78406 , 
 n78407 , n78408 , n78409 , n78410 , n78411 , n78412 , n78413 , n78414 , n78415 , n78416 , 
 n78417 , n78418 , n78419 , n78420 , n78421 , n78422 , n78423 , n78424 , n78425 , n78426 , 
 n78427 , n78428 , n78429 , n78430 , n78431 , n78432 , n78433 , n78434 , n78435 , n78436 , 
 n78437 , n78438 , n78439 , n78440 , n78441 , n78442 , n78443 , n78444 , n78445 , n78446 , 
 n78447 , n78448 , n78449 , n78450 , n78451 , n78452 , n78453 , n78454 , n78455 , n78456 , 
 n78457 , n78458 , n78459 , n78460 , n78461 , n78462 , n78463 , n78464 , n78465 , n78466 , 
 n78467 , n78468 , n78469 , n78470 , n78471 , n78472 , n78473 , n78474 , n78475 , n78476 , 
 n78477 , n78478 , n78479 , n78480 , n78481 , n78482 , n78483 , n78484 , n78485 , n78486 , 
 n78487 , n78488 , n78489 , n78490 , n78491 , n78492 , n78493 , n78494 , n78495 , n78496 , 
 n78497 , n78498 , n78499 , n78500 , n78501 , n78502 , n78503 , n78504 , n78505 , n78506 , 
 n78507 , n78508 , n78509 , n78510 , n78511 , n78512 , n78513 , n78514 , n78515 , n78516 , 
 n78517 , n78518 , n78519 , n78520 , n78521 , n78522 , n78523 , n78524 , n78525 , n78526 , 
 n78527 , n78528 , n78529 , n78530 , n78531 , n78532 , n78533 , n78534 , n78535 , n78536 , 
 n78537 , n78538 , n78539 , n78540 , n78541 , n78542 , n78543 , n78544 , n78545 , n78546 , 
 n78547 , n78548 , n78549 , n78550 , n78551 , n78552 , n78553 , n78554 , n78555 , n78556 , 
 n78557 , n78558 , n78559 , n78560 , n78561 , n78562 , n78563 , n78564 , n78565 , n78566 , 
 n78567 , n78568 , n78569 , n78570 , n78571 , n78572 , n78573 , n78574 , n78575 , n78576 , 
 n78577 , n78578 , n78579 , n78580 , n78581 , n78582 , n78583 , n78584 , n78585 , n78586 , 
 n78587 , n78588 , n78589 , n78590 , n78591 , n78592 , n78593 , n78594 , n78595 , n78596 , 
 n78597 , n78598 , n78599 , n78600 , n78601 , n78602 , n78603 , n78604 , n78605 , n78606 , 
 n78607 , n78608 , n78609 , n78610 , n78611 , n78612 , n78613 , n78614 , n78615 , n78616 , 
 n78617 , n78618 , n78619 , n78620 , n78621 , n78622 , n78623 , n78624 , n78625 , n78626 , 
 C0n , C0 ;
buf ( n736 , n6 );
buf ( n737 , n7 );
buf ( n738 , n8 );
buf ( n739 , n9 );
buf ( n740 , n10 );
buf ( n741 , n11 );
buf ( n742 , n12 );
buf ( n743 , n13 );
buf ( n744 , n14 );
buf ( n745 , n15 );
buf ( n746 , n16 );
buf ( n747 , n17 );
buf ( n748 , n18 );
buf ( n749 , n19 );
buf ( n750 , n20 );
buf ( n751 , n21 );
buf ( n752 , n22 );
buf ( n753 , n23 );
buf ( n754 , n24 );
buf ( n755 , n25 );
buf ( n756 , n26 );
buf ( n757 , n27 );
buf ( n758 , n28 );
buf ( n759 , n29 );
buf ( n760 , n30 );
buf ( n761 , n31 );
buf ( n762 , n32 );
buf ( n763 , n33 );
buf ( n764 , n34 );
buf ( n765 , n35 );
buf ( n766 , n36 );
buf ( n767 , n37 );
buf ( n768 , n38 );
buf ( n769 , n39 );
buf ( n770 , n40 );
buf ( n771 , n41 );
buf ( n772 , n42 );
buf ( n773 , n43 );
buf ( n774 , n44 );
buf ( n775 , n45 );
buf ( n776 , n46 );
buf ( n777 , n47 );
buf ( n778 , n48 );
buf ( n779 , n49 );
buf ( n780 , n50 );
buf ( n781 , n51 );
buf ( n782 , n52 );
buf ( n783 , n53 );
buf ( n784 , n54 );
buf ( n785 , n55 );
buf ( n786 , n56 );
buf ( n787 , n57 );
buf ( n788 , n58 );
buf ( n789 , n59 );
buf ( n790 , n60 );
buf ( n791 , n61 );
buf ( n792 , n62 );
buf ( n793 , n63 );
buf ( n794 , n64 );
buf ( n795 , n65 );
buf ( n796 , n66 );
buf ( n797 , n67 );
buf ( n798 , n68 );
buf ( n799 , n69 );
buf ( n800 , n70 );
buf ( n801 , n71 );
buf ( n802 , n72 );
buf ( n803 , n73 );
buf ( n804 , n74 );
buf ( n805 , n75 );
buf ( n806 , n76 );
buf ( n807 , n77 );
buf ( n808 , n78 );
buf ( n809 , n79 );
buf ( n80 , n810 );
buf ( n81 , n811 );
buf ( n82 , n812 );
buf ( n83 , n813 );
buf ( n84 , n814 );
buf ( n85 , n815 );
buf ( n86 , n816 );
buf ( n87 , n817 );
buf ( n88 , n818 );
buf ( n89 , n819 );
buf ( n90 , n820 );
buf ( n91 , n821 );
buf ( n92 , n822 );
buf ( n93 , n823 );
buf ( n94 , n824 );
buf ( n95 , n825 );
buf ( n96 , n826 );
buf ( n97 , n827 );
buf ( n98 , n828 );
buf ( n99 , n829 );
buf ( n100 , n830 );
buf ( n101 , n831 );
buf ( n102 , n832 );
buf ( n103 , n833 );
buf ( n104 , n834 );
buf ( n105 , n835 );
buf ( n106 , n836 );
buf ( n107 , n837 );
buf ( n108 , n838 );
buf ( n109 , n839 );
buf ( n110 , n840 );
buf ( n111 , n841 );
buf ( n112 , n842 );
buf ( n113 , n843 );
buf ( n114 , n844 );
buf ( n115 , n845 );
buf ( n116 , n846 );
buf ( n117 , n847 );
buf ( n118 , n848 );
buf ( n119 , n849 );
buf ( n120 , n850 );
buf ( n121 , n851 );
buf ( n122 , n852 );
buf ( n123 , n853 );
buf ( n124 , n854 );
buf ( n125 , n855 );
buf ( n126 , n856 );
buf ( n127 , n857 );
buf ( n128 , n858 );
buf ( n129 , n859 );
buf ( n130 , n860 );
buf ( n131 , n861 );
buf ( n132 , n862 );
buf ( n133 , n863 );
buf ( n134 , n864 );
buf ( n135 , n865 );
buf ( n136 , n866 );
buf ( n137 , n867 );
buf ( n138 , n868 );
buf ( n139 , n869 );
buf ( n140 , n870 );
buf ( n141 , n871 );
buf ( n142 , n872 );
buf ( n143 , n873 );
buf ( n144 , n874 );
buf ( n145 , n875 );
buf ( n146 , n876 );
buf ( n147 , n877 );
buf ( n148 , n878 );
buf ( n149 , n879 );
buf ( n150 , n880 );
buf ( n151 , n881 );
buf ( n152 , n882 );
buf ( n153 , n883 );
buf ( n154 , n884 );
buf ( n155 , n885 );
buf ( n156 , n886 );
buf ( n157 , n887 );
buf ( n158 , n888 );
buf ( n159 , n889 );
buf ( n160 , n890 );
buf ( n161 , n891 );
buf ( n162 , n892 );
buf ( n163 , n893 );
buf ( n164 , n894 );
buf ( n165 , n895 );
buf ( n166 , n896 );
buf ( n167 , n897 );
buf ( n168 , n898 );
buf ( n169 , n899 );
buf ( n170 , n900 );
buf ( n171 , n901 );
buf ( n172 , n902 );
buf ( n173 , n903 );
buf ( n174 , n904 );
buf ( n175 , n905 );
buf ( n176 , n906 );
buf ( n177 , n907 );
buf ( n178 , n908 );
buf ( n179 , n909 );
buf ( n180 , n910 );
buf ( n181 , n911 );
buf ( n182 , n912 );
buf ( n183 , n913 );
buf ( n184 , n914 );
buf ( n185 , n915 );
buf ( n186 , n916 );
buf ( n187 , n917 );
buf ( n188 , n918 );
buf ( n189 , n919 );
buf ( n190 , n920 );
buf ( n191 , n921 );
buf ( n192 , n922 );
buf ( n193 , n923 );
buf ( n194 , n924 );
buf ( n195 , n925 );
buf ( n196 , n926 );
buf ( n197 , n927 );
buf ( n198 , n928 );
buf ( n199 , n929 );
buf ( n200 , n930 );
buf ( n201 , n931 );
buf ( n202 , n932 );
buf ( n203 , n933 );
buf ( n204 , n934 );
buf ( n205 , n935 );
buf ( n206 , n936 );
buf ( n207 , n937 );
buf ( n208 , n938 );
buf ( n209 , n939 );
buf ( n210 , n940 );
buf ( n211 , n941 );
buf ( n212 , n942 );
buf ( n213 , n943 );
buf ( n214 , n944 );
buf ( n215 , n945 );
buf ( n216 , n946 );
buf ( n217 , n947 );
buf ( n218 , n948 );
buf ( n219 , n949 );
buf ( n220 , n950 );
buf ( n221 , n951 );
buf ( n222 , n952 );
buf ( n223 , n953 );
buf ( n224 , n954 );
buf ( n225 , n955 );
buf ( n226 , n956 );
buf ( n227 , n957 );
buf ( n228 , n958 );
buf ( n229 , n959 );
buf ( n230 , n960 );
buf ( n231 , n961 );
buf ( n232 , n962 );
buf ( n233 , n963 );
buf ( n234 , n964 );
buf ( n235 , n965 );
buf ( n236 , n966 );
buf ( n237 , n967 );
buf ( n238 , n968 );
buf ( n239 , n969 );
buf ( n240 , n970 );
buf ( n241 , n971 );
buf ( n242 , n972 );
buf ( n243 , n973 );
buf ( n244 , n974 );
buf ( n245 , n975 );
buf ( n246 , n976 );
buf ( n247 , n977 );
buf ( n248 , n978 );
buf ( n249 , n979 );
buf ( n250 , n980 );
buf ( n251 , n981 );
buf ( n252 , n982 );
buf ( n253 , n983 );
buf ( n254 , n984 );
buf ( n255 , n985 );
buf ( n256 , n986 );
buf ( n257 , n987 );
buf ( n258 , n988 );
buf ( n259 , n989 );
buf ( n260 , n990 );
buf ( n261 , n991 );
buf ( n262 , n992 );
buf ( n263 , n993 );
buf ( n264 , n994 );
buf ( n265 , n995 );
buf ( n266 , n996 );
buf ( n267 , n997 );
buf ( n268 , n998 );
buf ( n269 , n999 );
buf ( n270 , n1000 );
buf ( n271 , n1001 );
buf ( n272 , n1002 );
buf ( n273 , n1003 );
buf ( n274 , n1004 );
buf ( n275 , n1005 );
buf ( n276 , n1006 );
buf ( n277 , n1007 );
buf ( n278 , n1008 );
buf ( n279 , n1009 );
buf ( n280 , n1010 );
buf ( n281 , n1011 );
buf ( n282 , n1012 );
buf ( n283 , n1013 );
buf ( n284 , n1014 );
buf ( n285 , n1015 );
buf ( n286 , n1016 );
buf ( n287 , n1017 );
buf ( n288 , n1018 );
buf ( n289 , n1019 );
buf ( n290 , n1020 );
buf ( n291 , n1021 );
buf ( n292 , n1022 );
buf ( n293 , n1023 );
buf ( n294 , n1024 );
buf ( n295 , n1025 );
buf ( n296 , n1026 );
buf ( n297 , n1027 );
buf ( n298 , n1028 );
buf ( n299 , n1029 );
buf ( n300 , n1030 );
buf ( n301 , n1031 );
buf ( n302 , n1032 );
buf ( n303 , n1033 );
buf ( n304 , n1034 );
buf ( n305 , n1035 );
buf ( n306 , n1036 );
buf ( n307 , n1037 );
buf ( n308 , n1038 );
buf ( n309 , n1039 );
buf ( n310 , n1040 );
buf ( n311 , n1041 );
buf ( n312 , n1042 );
buf ( n313 , n1043 );
buf ( n314 , n1044 );
buf ( n315 , n1045 );
buf ( n316 , n1046 );
buf ( n317 , n1047 );
buf ( n318 , n1048 );
buf ( n319 , n1049 );
buf ( n320 , n1050 );
buf ( n321 , n1051 );
buf ( n322 , n1052 );
buf ( n323 , n1053 );
buf ( n324 , n1054 );
buf ( n325 , n1055 );
buf ( n326 , n1056 );
buf ( n327 , n1057 );
buf ( n328 , n1058 );
buf ( n329 , n1059 );
buf ( n330 , n1060 );
buf ( n331 , n1061 );
buf ( n332 , n1062 );
buf ( n333 , n1063 );
buf ( n334 , n1064 );
buf ( n335 , n1065 );
buf ( n336 , n1066 );
buf ( n337 , n1067 );
buf ( n338 , n1068 );
buf ( n339 , n1069 );
buf ( n340 , n1070 );
buf ( n341 , n1071 );
buf ( n342 , n1072 );
buf ( n343 , n1073 );
buf ( n344 , n1074 );
buf ( n345 , n1075 );
buf ( n346 , n1076 );
buf ( n347 , n1077 );
buf ( n348 , n1078 );
buf ( n349 , n1079 );
buf ( n350 , n1080 );
buf ( n351 , n1081 );
buf ( n352 , n1082 );
buf ( n353 , n1083 );
buf ( n354 , n1084 );
buf ( n355 , n1085 );
buf ( n356 , n1086 );
buf ( n357 , n1087 );
buf ( n358 , n1088 );
buf ( n359 , n1089 );
buf ( n360 , n1090 );
buf ( n361 , n1091 );
buf ( n362 , n1092 );
buf ( n363 , n1093 );
buf ( n364 , n1094 );
buf ( n365 , n1095 );
buf ( n366 , n1096 );
buf ( n367 , n1097 );
buf ( n810 , n20184 );
buf ( n811 , n20187 );
buf ( n812 , n20190 );
buf ( n813 , n20193 );
buf ( n814 , n20196 );
buf ( n815 , n20199 );
buf ( n816 , n20202 );
buf ( n817 , n20205 );
buf ( n818 , n20208 );
buf ( n819 , n20211 );
buf ( n820 , n20214 );
buf ( n821 , n20217 );
buf ( n822 , n20220 );
buf ( n823 , n20223 );
buf ( n824 , n20226 );
buf ( n825 , n20229 );
buf ( n826 , n20232 );
buf ( n827 , n20235 );
buf ( n828 , n20238 );
buf ( n829 , n20241 );
buf ( n830 , n20244 );
buf ( n831 , n20247 );
buf ( n832 , n20252 );
buf ( n833 , n20257 );
buf ( n834 , n20262 );
buf ( n835 , n20267 );
buf ( n836 , n20270 );
buf ( n837 , n20273 );
buf ( n838 , n20276 );
buf ( n839 , n20279 );
buf ( n840 , n10629 );
buf ( n841 , n10921 );
buf ( n842 , n45689 );
buf ( n843 , n45667 );
buf ( n844 , n45696 );
buf ( n845 , n45725 );
buf ( n846 , n45766 );
buf ( n847 , n45797 );
buf ( n848 , n45847 );
buf ( n849 , n45911 );
buf ( n850 , n45984 );
buf ( n851 , n46058 );
buf ( n852 , n46103 );
buf ( n853 , n46172 );
buf ( n854 , n46268 );
buf ( n855 , n46349 );
buf ( n856 , n46478 );
buf ( n857 , n46533 );
buf ( n858 , n46630 );
buf ( n859 , n46754 );
buf ( n860 , n46902 );
buf ( n861 , n46973 );
buf ( n862 , n47093 );
buf ( n863 , n47220 );
buf ( n864 , n47355 );
buf ( n865 , n47546 );
buf ( n866 , n47691 );
buf ( n867 , n47782 );
buf ( n868 , n48017 );
buf ( n869 , n48193 );
buf ( n870 , n48275 );
buf ( n871 , n48437 );
buf ( n872 , n48690 );
buf ( n873 , n48802 );
buf ( n874 , n48992 );
buf ( n875 , n49178 );
buf ( n876 , n49480 );
buf ( n877 , n49573 );
buf ( n878 , n49784 );
buf ( n879 , n49980 );
buf ( n880 , n50273 );
buf ( n881 , n50488 );
buf ( n882 , n50628 );
buf ( n883 , n50845 );
buf ( n884 , n51081 );
buf ( n885 , n51302 );
buf ( n886 , n51670 );
buf ( n887 , n51832 );
buf ( n888 , n52086 );
buf ( n889 , n52460 );
buf ( n890 , n52615 );
buf ( n891 , n52873 );
buf ( n892 , n53146 );
buf ( n893 , n53423 );
buf ( n894 , n53846 );
buf ( n895 , n54158 );
buf ( n896 , n54312 );
buf ( n897 , n54607 );
buf ( n898 , n54946 );
buf ( n899 , n55255 );
buf ( n900 , n55578 );
buf ( n901 , n55931 );
buf ( n902 , n56396 );
buf ( n903 , n56577 );
buf ( n904 , n57079 );
buf ( n905 , n57273 );
buf ( n906 , n57603 );
buf ( n907 , n57944 );
buf ( n908 , n58287 );
buf ( n909 , n58623 );
buf ( n910 , n58988 );
buf ( n911 , n59360 );
buf ( n912 , n59723 );
buf ( n913 , n60092 );
buf ( n914 , n60617 );
buf ( n915 , n60816 );
buf ( n916 , n61181 );
buf ( n917 , n61579 );
buf ( n918 , n62009 );
buf ( n919 , n62369 );
buf ( n920 , n62703 );
buf ( n921 , n63100 );
buf ( n922 , n63487 );
buf ( n923 , n63850 );
buf ( n924 , n64217 );
buf ( n925 , n64640 );
buf ( n926 , n65021 );
buf ( n927 , n65414 );
buf ( n928 , n65832 );
buf ( n929 , n66229 );
buf ( n930 , n66715 );
buf ( n931 , n67179 );
buf ( n932 , n67554 );
buf ( n933 , n67993 );
buf ( n934 , n68432 );
buf ( n935 , n68887 );
buf ( n936 , n69296 );
buf ( n937 , n69788 );
buf ( n938 , n70236 );
buf ( n939 , n70660 );
buf ( n940 , n71035 );
buf ( n941 , n71465 );
buf ( n942 , n71858 );
buf ( n943 , n72239 );
buf ( n944 , n72610 );
buf ( n945 , n72998 );
buf ( n946 , n73342 );
buf ( n947 , n73690 );
buf ( n948 , n74082 );
buf ( n949 , n74396 );
buf ( n950 , n74705 );
buf ( n951 , n74998 );
buf ( n952 , n75295 );
buf ( n953 , n75570 );
buf ( n954 , n75839 );
buf ( n955 , n76082 );
buf ( n956 , n76310 );
buf ( n957 , n76698 );
buf ( n958 , n76754 );
buf ( n959 , n76937 );
buf ( n960 , n77108 );
buf ( n961 , n77300 );
buf ( n962 , n77463 );
buf ( n963 , n77616 );
buf ( n964 , n77736 );
buf ( n965 , n77832 );
buf ( n966 , n77985 );
buf ( n967 , n78007 );
buf ( n968 , n78073 );
buf ( n969 , n78103 );
buf ( n970 , n78370 );
buf ( n971 , n78372 );
buf ( n972 , n78374 );
buf ( n973 , n78376 );
buf ( n974 , n78378 );
buf ( n975 , n78380 );
buf ( n976 , n78382 );
buf ( n977 , n78384 );
buf ( n978 , n78386 );
buf ( n979 , n78388 );
buf ( n980 , n78390 );
buf ( n981 , n78392 );
buf ( n982 , n78394 );
buf ( n983 , n78396 );
buf ( n984 , n78398 );
buf ( n985 , n78400 );
buf ( n986 , n78402 );
buf ( n987 , n78404 );
buf ( n988 , n78406 );
buf ( n989 , n78408 );
buf ( n990 , n78410 );
buf ( n991 , n78412 );
buf ( n992 , n78414 );
buf ( n993 , n78416 );
buf ( n994 , n78418 );
buf ( n995 , n78420 );
buf ( n996 , n78422 );
buf ( n997 , n78424 );
buf ( n998 , n78426 );
buf ( n999 , n78428 );
buf ( n1000 , n78430 );
buf ( n1001 , n78432 );
buf ( n1002 , n78434 );
buf ( n1003 , n78436 );
buf ( n1004 , n78438 );
buf ( n1005 , n78440 );
buf ( n1006 , n78442 );
buf ( n1007 , n78444 );
buf ( n1008 , n78446 );
buf ( n1009 , n78448 );
buf ( n1010 , n78450 );
buf ( n1011 , n78452 );
buf ( n1012 , n78454 );
buf ( n1013 , n78456 );
buf ( n1014 , n78458 );
buf ( n1015 , n78460 );
buf ( n1016 , n78462 );
buf ( n1017 , n78464 );
buf ( n1018 , n78466 );
buf ( n1019 , n78468 );
buf ( n1020 , n78470 );
buf ( n1021 , n78472 );
buf ( n1022 , n78474 );
buf ( n1023 , n78476 );
buf ( n1024 , n78478 );
buf ( n1025 , n78480 );
buf ( n1026 , n78482 );
buf ( n1027 , n78484 );
buf ( n1028 , n78486 );
buf ( n1029 , n78488 );
buf ( n1030 , n78490 );
buf ( n1031 , n78492 );
buf ( n1032 , n78494 );
buf ( n1033 , n78496 );
buf ( n1034 , n78498 );
buf ( n1035 , n78500 );
buf ( n1036 , n78502 );
buf ( n1037 , n78504 );
buf ( n1038 , n78506 );
buf ( n1039 , n78508 );
buf ( n1040 , n78510 );
buf ( n1041 , n78512 );
buf ( n1042 , n78514 );
buf ( n1043 , n78516 );
buf ( n1044 , n78518 );
buf ( n1045 , n78520 );
buf ( n1046 , n78522 );
buf ( n1047 , n78524 );
buf ( n1048 , n78526 );
buf ( n1049 , n78528 );
buf ( n1050 , n78530 );
buf ( n1051 , n78532 );
buf ( n1052 , n78534 );
buf ( n1053 , n78536 );
buf ( n1054 , n78538 );
buf ( n1055 , n78540 );
buf ( n1056 , n78542 );
buf ( n1057 , n78544 );
buf ( n1058 , n78546 );
buf ( n1059 , n78548 );
buf ( n1060 , n78550 );
buf ( n1061 , n78552 );
buf ( n1062 , n78554 );
buf ( n1063 , n78556 );
buf ( n1064 , n78558 );
buf ( n1065 , n78560 );
buf ( n1066 , n78562 );
buf ( n1067 , n78564 );
buf ( n1068 , n78566 );
buf ( n1069 , n78568 );
buf ( n1070 , n78570 );
buf ( n1071 , n78572 );
buf ( n1072 , n78574 );
buf ( n1073 , n78576 );
buf ( n1074 , n78578 );
buf ( n1075 , n78580 );
buf ( n1076 , n78582 );
buf ( n1077 , n78584 );
buf ( n1078 , n78586 );
buf ( n1079 , n78588 );
buf ( n1080 , n78590 );
buf ( n1081 , n78592 );
buf ( n1082 , n78594 );
buf ( n1083 , n78596 );
buf ( n1084 , n78598 );
buf ( n1085 , n78600 );
buf ( n1086 , n78602 );
buf ( n1087 , n78604 );
buf ( n1088 , n78606 );
buf ( n1089 , n78608 );
buf ( n1090 , n78610 );
buf ( n1091 , n78612 );
buf ( n1092 , n78614 );
buf ( n1093 , n78616 );
buf ( n1094 , n78618 );
buf ( n1095 , n78620 );
buf ( n1096 , n78622 );
buf ( n1097 , n78626 );
buf ( n1098 , n742 );
buf ( n1099 , n1098 );
buf ( n1100 , n1099 );
buf ( n1101 , n1100 );
buf ( n1102 , n1101 );
buf ( n1103 , n1102 );
buf ( n1104 , n1103 );
buf ( n1105 , n1104 );
buf ( n1106 , n1105 );
buf ( n1107 , n736 );
buf ( n1108 , n737 );
buf ( n1109 , n738 );
buf ( n1110 , n739 );
buf ( n1111 , n740 );
buf ( n1112 , n741 );
buf ( n1113 , n742 );
buf ( n1114 , n746 );
and ( n1115 , n1113 , n1114 );
buf ( n1116 , n743 );
buf ( n1117 , n747 );
and ( n1118 , n1116 , n1117 );
buf ( n1119 , n744 );
buf ( n1120 , n748 );
and ( n1121 , n1119 , n1120 );
buf ( n1122 , n745 );
buf ( n1123 , n749 );
and ( n1124 , n1122 , n1123 );
and ( n1125 , n1120 , n1124 );
and ( n1126 , n1119 , n1124 );
or ( n1127 , n1121 , n1125 , n1126 );
and ( n1128 , n1117 , n1127 );
and ( n1129 , n1116 , n1127 );
or ( n1130 , n1118 , n1128 , n1129 );
and ( n1131 , n1114 , n1130 );
and ( n1132 , n1113 , n1130 );
or ( n1133 , n1115 , n1131 , n1132 );
and ( n1134 , n1112 , n1133 );
and ( n1135 , n1111 , n1134 );
and ( n1136 , n1110 , n1135 );
and ( n1137 , n1109 , n1136 );
and ( n1138 , n1108 , n1137 );
xor ( n1139 , n1107 , n1138 );
buf ( n1140 , n1139 );
buf ( n1141 , n1140 );
xor ( n1142 , n1108 , n1137 );
buf ( n1143 , n1142 );
buf ( n1144 , n1143 );
xor ( n1145 , n1109 , n1136 );
buf ( n1146 , n1145 );
buf ( n1147 , n1146 );
xor ( n1148 , n1110 , n1135 );
buf ( n1149 , n1148 );
buf ( n1150 , n1149 );
xor ( n1151 , n1111 , n1134 );
buf ( n1152 , n1151 );
buf ( n1153 , n1152 );
xor ( n1154 , n1112 , n1133 );
buf ( n1155 , n1154 );
buf ( n1156 , n1155 );
xor ( n1157 , n1113 , n1114 );
xor ( n1158 , n1157 , n1130 );
buf ( n1159 , n1158 );
buf ( n1160 , n1159 );
xor ( n1161 , n1116 , n1117 );
xor ( n1162 , n1161 , n1127 );
buf ( n1163 , n1162 );
buf ( n1164 , n1163 );
xor ( n1165 , n1119 , n1120 );
xor ( n1166 , n1165 , n1124 );
buf ( n1167 , n1166 );
buf ( n1168 , n1167 );
xor ( n1169 , n1122 , n1123 );
buf ( n1170 , n1169 );
buf ( n1171 , n1170 );
buf ( n1172 , n750 );
buf ( n1173 , n1172 );
buf ( n1174 , n1173 );
buf ( n1175 , n1174 );
buf ( n1176 , n751 );
buf ( n1177 , n1176 );
buf ( n1178 , n1177 );
buf ( n1179 , n1178 );
buf ( n1180 , n752 );
buf ( n1181 , n1180 );
buf ( n1182 , n1181 );
buf ( n1183 , n1182 );
buf ( n1184 , n753 );
buf ( n1185 , n1184 );
buf ( n1186 , n1185 );
buf ( n1187 , n1186 );
buf ( n1188 , n754 );
buf ( n1189 , n1188 );
buf ( n1190 , n1189 );
buf ( n1191 , n1190 );
buf ( n1192 , n755 );
buf ( n1193 , n1192 );
buf ( n1194 , n1193 );
buf ( n1195 , n1194 );
buf ( n1196 , n756 );
buf ( n1197 , n1196 );
buf ( n1198 , n1197 );
buf ( n1199 , n1198 );
buf ( n1200 , n762 );
and ( n1201 , n1199 , n1200 );
buf ( n1202 , n757 );
buf ( n1203 , n1202 );
buf ( n1204 , n1203 );
buf ( n1205 , n1204 );
buf ( n1206 , n763 );
and ( n1207 , n1205 , n1206 );
buf ( n1208 , n758 );
buf ( n1209 , n1208 );
buf ( n1210 , n1209 );
buf ( n1211 , n1210 );
buf ( n1212 , n764 );
and ( n1213 , n1211 , n1212 );
buf ( n1214 , n759 );
buf ( n1215 , n1214 );
buf ( n1216 , n1215 );
buf ( n1217 , n1216 );
buf ( n1218 , n765 );
and ( n1219 , n1217 , n1218 );
buf ( n1220 , n760 );
buf ( n1221 , n1220 );
buf ( n1222 , n1221 );
buf ( n1223 , n1222 );
buf ( n1224 , n766 );
and ( n1225 , n1223 , n1224 );
buf ( n1226 , n761 );
buf ( n1227 , n1226 );
buf ( n1228 , n1227 );
buf ( n1229 , n1228 );
buf ( n1230 , n767 );
and ( n1231 , n1229 , n1230 );
and ( n1232 , n1224 , n1231 );
and ( n1233 , n1223 , n1231 );
or ( n1234 , n1225 , n1232 , n1233 );
and ( n1235 , n1218 , n1234 );
and ( n1236 , n1217 , n1234 );
or ( n1237 , n1219 , n1235 , n1236 );
and ( n1238 , n1212 , n1237 );
and ( n1239 , n1211 , n1237 );
or ( n1240 , n1213 , n1238 , n1239 );
and ( n1241 , n1206 , n1240 );
and ( n1242 , n1205 , n1240 );
or ( n1243 , n1207 , n1241 , n1242 );
and ( n1244 , n1200 , n1243 );
and ( n1245 , n1199 , n1243 );
or ( n1246 , n1201 , n1244 , n1245 );
and ( n1247 , n1195 , n1246 );
and ( n1248 , n1191 , n1247 );
and ( n1249 , n1187 , n1248 );
and ( n1250 , n1183 , n1249 );
and ( n1251 , n1179 , n1250 );
and ( n1252 , n1175 , n1251 );
and ( n1253 , n1171 , n1252 );
and ( n1254 , n1168 , n1253 );
and ( n1255 , n1164 , n1254 );
and ( n1256 , n1160 , n1255 );
and ( n1257 , n1156 , n1256 );
and ( n1258 , n1153 , n1257 );
and ( n1259 , n1150 , n1258 );
and ( n1260 , n1147 , n1259 );
and ( n1261 , n1144 , n1260 );
xor ( n1262 , n1141 , n1261 );
buf ( n1263 , n1262 );
buf ( n1264 , n1263 );
buf ( n1265 , n1264 );
buf ( n1266 , n1265 );
xnor ( n1267 , n1106 , n1266 );
buf ( n1268 , n743 );
buf ( n1269 , n1268 );
buf ( n1270 , n1269 );
buf ( n1271 , n1270 );
buf ( n1272 , n1271 );
buf ( n1273 , n1272 );
buf ( n1274 , n1273 );
buf ( n1275 , n1274 );
not ( n1276 , n1275 );
buf ( n1277 , n1103 );
buf ( n1278 , n1277 );
not ( n1279 , n1278 );
and ( n1280 , n1279 , n1275 );
nor ( n1281 , n1276 , n1280 );
xor ( n1282 , n1147 , n1259 );
buf ( n1283 , n1282 );
buf ( n1284 , n1283 );
buf ( n1285 , n1284 );
buf ( n1286 , n1263 );
buf ( n1287 , n1286 );
and ( n1288 , n1285 , n1287 );
and ( n1289 , n1281 , n1288 );
and ( n1290 , n1267 , n1289 );
not ( n1291 , n1105 );
buf ( n1292 , n1273 );
buf ( n1293 , n1292 );
and ( n1294 , n1291 , n1293 );
not ( n1295 , n1293 );
nor ( n1296 , n1294 , n1295 );
buf ( n1297 , n1296 );
xor ( n1298 , n1144 , n1260 );
buf ( n1299 , n1298 );
buf ( n1300 , n1299 );
buf ( n1301 , n1300 );
and ( n1302 , n1301 , n1287 );
xor ( n1303 , n1297 , n1302 );
not ( n1304 , n1296 );
buf ( n1305 , n744 );
buf ( n1306 , n1305 );
buf ( n1307 , n1306 );
buf ( n1308 , n1307 );
buf ( n1309 , n1308 );
buf ( n1310 , n1309 );
buf ( n1311 , n1310 );
buf ( n1312 , n1311 );
and ( n1313 , n1291 , n1312 );
not ( n1314 , n1312 );
nor ( n1315 , n1313 , n1314 );
buf ( n1316 , n1310 );
buf ( n1317 , n1316 );
not ( n1318 , n1317 );
and ( n1319 , n1279 , n1317 );
nor ( n1320 , n1318 , n1319 );
and ( n1321 , n1315 , n1320 );
and ( n1322 , n1304 , n1321 );
xor ( n1323 , n1281 , n1288 );
and ( n1324 , n1321 , n1323 );
and ( n1325 , n1304 , n1323 );
or ( n1326 , n1322 , n1324 , n1325 );
and ( n1327 , n1303 , n1326 );
xor ( n1328 , n1267 , n1289 );
and ( n1329 , n1326 , n1328 );
and ( n1330 , n1303 , n1328 );
or ( n1331 , n1327 , n1329 , n1330 );
xor ( n1332 , n1290 , n1331 );
or ( n1333 , n1106 , n1266 );
and ( n1334 , n1297 , n1302 );
xor ( n1335 , n1333 , n1334 );
xor ( n1336 , n1332 , n1335 );
buf ( n1337 , n1275 );
buf ( n1338 , n1301 );
and ( n1339 , n1337 , n1338 );
xor ( n1340 , n1337 , n1338 );
buf ( n1341 , n745 );
buf ( n1342 , n1341 );
buf ( n1343 , n1342 );
buf ( n1344 , n1343 );
buf ( n1345 , n1344 );
buf ( n1346 , n1345 );
buf ( n1347 , n1346 );
buf ( n1348 , n1347 );
and ( n1349 , n1291 , n1348 );
not ( n1350 , n1348 );
nor ( n1351 , n1349 , n1350 );
buf ( n1352 , n1346 );
buf ( n1353 , n1352 );
not ( n1354 , n1353 );
and ( n1355 , n1279 , n1353 );
nor ( n1356 , n1354 , n1355 );
and ( n1357 , n1351 , n1356 );
and ( n1358 , n1340 , n1357 );
buf ( n1359 , n1299 );
buf ( n1360 , n1359 );
and ( n1361 , n1285 , n1360 );
and ( n1362 , n1357 , n1361 );
and ( n1363 , n1340 , n1361 );
or ( n1364 , n1358 , n1362 , n1363 );
and ( n1365 , n1339 , n1364 );
and ( n1366 , n1275 , n1312 );
buf ( n1367 , n1366 );
xor ( n1368 , n1150 , n1258 );
buf ( n1369 , n1368 );
buf ( n1370 , n1369 );
buf ( n1371 , n1370 );
and ( n1372 , n1371 , n1287 );
or ( n1373 , n1367 , n1372 );
and ( n1374 , n1364 , n1373 );
and ( n1375 , n1339 , n1373 );
or ( n1376 , n1365 , n1374 , n1375 );
xor ( n1377 , n1303 , n1326 );
xor ( n1378 , n1377 , n1328 );
and ( n1379 , n1376 , n1378 );
xor ( n1380 , n1315 , n1320 );
and ( n1381 , n1317 , n1293 );
xor ( n1382 , n1153 , n1257 );
buf ( n1383 , n1382 );
buf ( n1384 , n1383 );
buf ( n1385 , n1384 );
and ( n1386 , n1385 , n1287 );
and ( n1387 , n1381 , n1386 );
and ( n1388 , n1380 , n1387 );
xor ( n1389 , n1304 , n1321 );
xor ( n1390 , n1389 , n1323 );
and ( n1391 , n1388 , n1390 );
xor ( n1392 , n1339 , n1364 );
xor ( n1393 , n1392 , n1373 );
and ( n1394 , n1390 , n1393 );
and ( n1395 , n1388 , n1393 );
or ( n1396 , n1391 , n1394 , n1395 );
and ( n1397 , n1378 , n1396 );
and ( n1398 , n1376 , n1396 );
or ( n1399 , n1379 , n1397 , n1398 );
xnor ( n1400 , n1336 , n1399 );
xor ( n1401 , n1340 , n1357 );
xor ( n1402 , n1401 , n1361 );
xnor ( n1403 , n1367 , n1372 );
and ( n1404 , n1402 , n1403 );
buf ( n1405 , n1317 );
buf ( n1406 , n1285 );
and ( n1407 , n1405 , n1406 );
and ( n1408 , n1275 , n1348 );
buf ( n1409 , n1408 );
and ( n1410 , n1407 , n1409 );
and ( n1411 , n1371 , n1360 );
and ( n1412 , n1409 , n1411 );
and ( n1413 , n1407 , n1411 );
or ( n1414 , n1410 , n1412 , n1413 );
and ( n1415 , n1403 , n1414 );
and ( n1416 , n1402 , n1414 );
or ( n1417 , n1404 , n1415 , n1416 );
not ( n1418 , n1366 );
xor ( n1419 , n1351 , n1356 );
and ( n1420 , n1418 , n1419 );
and ( n1421 , n1353 , n1293 );
and ( n1422 , n1385 , n1360 );
and ( n1423 , n1421 , n1422 );
and ( n1424 , n1419 , n1423 );
and ( n1425 , n1418 , n1423 );
or ( n1426 , n1420 , n1424 , n1425 );
xor ( n1427 , n1380 , n1387 );
and ( n1428 , n1426 , n1427 );
xor ( n1429 , n1381 , n1386 );
xor ( n1430 , n1407 , n1409 );
xor ( n1431 , n1430 , n1411 );
and ( n1432 , n1429 , n1431 );
xor ( n1433 , n1405 , n1406 );
and ( n1434 , n1317 , n1348 );
and ( n1435 , n1353 , n1312 );
and ( n1436 , n1434 , n1435 );
and ( n1437 , n1433 , n1436 );
xor ( n1438 , n1156 , n1256 );
buf ( n1439 , n1438 );
buf ( n1440 , n1439 );
buf ( n1441 , n1440 );
and ( n1442 , n1441 , n1287 );
and ( n1443 , n1436 , n1442 );
and ( n1444 , n1433 , n1442 );
or ( n1445 , n1437 , n1443 , n1444 );
and ( n1446 , n1431 , n1445 );
and ( n1447 , n1429 , n1445 );
or ( n1448 , n1432 , n1446 , n1447 );
and ( n1449 , n1427 , n1448 );
and ( n1450 , n1426 , n1448 );
or ( n1451 , n1428 , n1449 , n1450 );
and ( n1452 , n1417 , n1451 );
xor ( n1453 , n1388 , n1390 );
xor ( n1454 , n1453 , n1393 );
and ( n1455 , n1451 , n1454 );
and ( n1456 , n1417 , n1454 );
or ( n1457 , n1452 , n1455 , n1456 );
xor ( n1458 , n1376 , n1378 );
xor ( n1459 , n1458 , n1396 );
and ( n1460 , n1457 , n1459 );
xor ( n1461 , n1457 , n1459 );
xor ( n1462 , n1402 , n1403 );
xor ( n1463 , n1462 , n1414 );
buf ( n1464 , n1283 );
buf ( n1465 , n1464 );
and ( n1466 , n1371 , n1465 );
not ( n1467 , n1408 );
and ( n1468 , n1466 , n1467 );
xor ( n1469 , n1160 , n1255 );
buf ( n1470 , n1469 );
buf ( n1471 , n1470 );
buf ( n1472 , n1471 );
and ( n1473 , n1472 , n1287 );
and ( n1474 , n1385 , n1465 );
and ( n1475 , n1473 , n1474 );
and ( n1476 , n1467 , n1475 );
and ( n1477 , n1466 , n1475 );
or ( n1478 , n1468 , n1476 , n1477 );
xor ( n1479 , n1418 , n1419 );
xor ( n1480 , n1479 , n1423 );
and ( n1481 , n1478 , n1480 );
xor ( n1482 , n1421 , n1422 );
xor ( n1483 , n1433 , n1436 );
xor ( n1484 , n1483 , n1442 );
and ( n1485 , n1482 , n1484 );
buf ( n1486 , n1353 );
buf ( n1487 , n1371 );
and ( n1488 , n1486 , n1487 );
and ( n1489 , n1441 , n1360 );
or ( n1490 , n1488 , n1489 );
and ( n1491 , n1484 , n1490 );
and ( n1492 , n1482 , n1490 );
or ( n1493 , n1485 , n1491 , n1492 );
and ( n1494 , n1480 , n1493 );
and ( n1495 , n1478 , n1493 );
or ( n1496 , n1481 , n1494 , n1495 );
and ( n1497 , n1463 , n1496 );
xor ( n1498 , n1426 , n1427 );
xor ( n1499 , n1498 , n1448 );
and ( n1500 , n1496 , n1499 );
and ( n1501 , n1463 , n1499 );
or ( n1502 , n1497 , n1500 , n1501 );
xor ( n1503 , n1417 , n1451 );
xor ( n1504 , n1503 , n1454 );
and ( n1505 , n1502 , n1504 );
xor ( n1506 , n1502 , n1504 );
xor ( n1507 , n1429 , n1431 );
xor ( n1508 , n1507 , n1445 );
xor ( n1509 , n1434 , n1435 );
and ( n1510 , n1472 , n1360 );
and ( n1511 , n1441 , n1465 );
and ( n1512 , n1510 , n1511 );
and ( n1513 , n1509 , n1512 );
xor ( n1514 , n1473 , n1474 );
and ( n1515 , n1512 , n1514 );
and ( n1516 , n1509 , n1514 );
or ( n1517 , n1513 , n1515 , n1516 );
xor ( n1518 , n1466 , n1467 );
xor ( n1519 , n1518 , n1475 );
and ( n1520 , n1517 , n1519 );
xnor ( n1521 , n1488 , n1489 );
xor ( n1522 , n1486 , n1487 );
xor ( n1523 , n1164 , n1254 );
buf ( n1524 , n1523 );
buf ( n1525 , n1524 );
buf ( n1526 , n1525 );
and ( n1527 , n1526 , n1287 );
and ( n1528 , n1522 , n1527 );
buf ( n1529 , n1369 );
buf ( n1530 , n1529 );
and ( n1531 , n1385 , n1530 );
and ( n1532 , n1527 , n1531 );
and ( n1533 , n1522 , n1531 );
or ( n1534 , n1528 , n1532 , n1533 );
and ( n1535 , n1521 , n1534 );
xor ( n1536 , n1509 , n1512 );
xor ( n1537 , n1536 , n1514 );
and ( n1538 , n1534 , n1537 );
and ( n1539 , n1521 , n1537 );
or ( n1540 , n1535 , n1538 , n1539 );
and ( n1541 , n1519 , n1540 );
and ( n1542 , n1517 , n1540 );
or ( n1543 , n1520 , n1541 , n1542 );
and ( n1544 , n1508 , n1543 );
xor ( n1545 , n1478 , n1480 );
xor ( n1546 , n1545 , n1493 );
and ( n1547 , n1543 , n1546 );
and ( n1548 , n1508 , n1546 );
or ( n1549 , n1544 , n1547 , n1548 );
xor ( n1550 , n1463 , n1496 );
xor ( n1551 , n1550 , n1499 );
and ( n1552 , n1549 , n1551 );
xor ( n1553 , n1549 , n1551 );
xor ( n1554 , n1508 , n1543 );
xor ( n1555 , n1554 , n1546 );
xor ( n1556 , n1482 , n1484 );
xor ( n1557 , n1556 , n1490 );
xor ( n1558 , n1517 , n1519 );
xor ( n1559 , n1558 , n1540 );
and ( n1560 , n1557 , n1559 );
xor ( n1561 , n1168 , n1253 );
buf ( n1562 , n1561 );
buf ( n1563 , n1562 );
buf ( n1564 , n1563 );
and ( n1565 , n1564 , n1287 );
and ( n1566 , n1472 , n1465 );
and ( n1567 , n1565 , n1566 );
and ( n1568 , n1441 , n1530 );
and ( n1569 , n1566 , n1568 );
and ( n1570 , n1565 , n1568 );
or ( n1571 , n1567 , n1569 , n1570 );
xor ( n1572 , n1510 , n1511 );
and ( n1573 , n1571 , n1572 );
buf ( n1574 , n746 );
buf ( n1575 , n1574 );
buf ( n1576 , n1575 );
buf ( n1577 , n1576 );
buf ( n1578 , n747 );
buf ( n1579 , n1578 );
buf ( n1580 , n1579 );
buf ( n1581 , n1580 );
buf ( n1582 , n748 );
buf ( n1583 , n1582 );
buf ( n1584 , n1583 );
buf ( n1585 , n1584 );
buf ( n1586 , n749 );
buf ( n1587 , n1586 );
buf ( n1588 , n1587 );
buf ( n1589 , n1588 );
buf ( n1590 , n750 );
buf ( n1591 , n1590 );
buf ( n1592 , n1591 );
buf ( n1593 , n1592 );
buf ( n1594 , n751 );
buf ( n1595 , n1594 );
buf ( n1596 , n1595 );
buf ( n1597 , n1596 );
buf ( n1598 , n752 );
buf ( n1599 , n1598 );
buf ( n1600 , n1599 );
buf ( n1601 , n1600 );
buf ( n1602 , n753 );
buf ( n1603 , n1602 );
buf ( n1604 , n1603 );
buf ( n1605 , n1604 );
buf ( n1606 , n762 );
and ( n1607 , n1605 , n1606 );
buf ( n1608 , n754 );
buf ( n1609 , n1608 );
buf ( n1610 , n1609 );
buf ( n1611 , n1610 );
buf ( n1612 , n763 );
and ( n1613 , n1611 , n1612 );
buf ( n1614 , n755 );
buf ( n1615 , n1614 );
buf ( n1616 , n1615 );
buf ( n1617 , n1616 );
buf ( n1618 , n764 );
and ( n1619 , n1617 , n1618 );
buf ( n1620 , n756 );
buf ( n1621 , n1620 );
buf ( n1622 , n1621 );
buf ( n1623 , n1622 );
buf ( n1624 , n765 );
and ( n1625 , n1623 , n1624 );
buf ( n1626 , n757 );
buf ( n1627 , n1626 );
buf ( n1628 , n1627 );
buf ( n1629 , n1628 );
buf ( n1630 , n766 );
and ( n1631 , n1629 , n1630 );
buf ( n1632 , n758 );
buf ( n1633 , n1632 );
buf ( n1634 , n1633 );
buf ( n1635 , n1634 );
buf ( n1636 , n767 );
and ( n1637 , n1635 , n1636 );
buf ( n1638 , n759 );
buf ( n1639 , n1638 );
buf ( n1640 , n1639 );
buf ( n1641 , n1640 );
buf ( n1642 , n768 );
and ( n1643 , n1641 , n1642 );
buf ( n1644 , n760 );
buf ( n1645 , n1644 );
buf ( n1646 , n1645 );
buf ( n1647 , n1646 );
buf ( n1648 , n769 );
and ( n1649 , n1647 , n1648 );
buf ( n1650 , n761 );
buf ( n1651 , n1650 );
buf ( n1652 , n1651 );
buf ( n1653 , n1652 );
buf ( n1654 , n770 );
and ( n1655 , n1653 , n1654 );
and ( n1656 , n1648 , n1655 );
and ( n1657 , n1647 , n1655 );
or ( n1658 , n1649 , n1656 , n1657 );
and ( n1659 , n1642 , n1658 );
and ( n1660 , n1641 , n1658 );
or ( n1661 , n1643 , n1659 , n1660 );
and ( n1662 , n1636 , n1661 );
and ( n1663 , n1635 , n1661 );
or ( n1664 , n1637 , n1662 , n1663 );
and ( n1665 , n1630 , n1664 );
and ( n1666 , n1629 , n1664 );
or ( n1667 , n1631 , n1665 , n1666 );
and ( n1668 , n1624 , n1667 );
and ( n1669 , n1623 , n1667 );
or ( n1670 , n1625 , n1668 , n1669 );
and ( n1671 , n1618 , n1670 );
and ( n1672 , n1617 , n1670 );
or ( n1673 , n1619 , n1671 , n1672 );
and ( n1674 , n1612 , n1673 );
and ( n1675 , n1611 , n1673 );
or ( n1676 , n1613 , n1674 , n1675 );
and ( n1677 , n1606 , n1676 );
and ( n1678 , n1605 , n1676 );
or ( n1679 , n1607 , n1677 , n1678 );
and ( n1680 , n1601 , n1679 );
and ( n1681 , n1597 , n1680 );
and ( n1682 , n1593 , n1681 );
and ( n1683 , n1589 , n1682 );
and ( n1684 , n1585 , n1683 );
and ( n1685 , n1581 , n1684 );
and ( n1686 , n1577 , n1685 );
buf ( n1687 , n1686 );
buf ( n1688 , n1687 );
buf ( n1689 , n1688 );
and ( n1690 , n1291 , n1689 );
not ( n1691 , n1689 );
nor ( n1692 , n1690 , n1691 );
buf ( n1693 , n1687 );
buf ( n1694 , n1693 );
not ( n1695 , n1694 );
and ( n1696 , n1279 , n1694 );
nor ( n1697 , n1695 , n1696 );
and ( n1698 , n1692 , n1697 );
and ( n1699 , n1526 , n1360 );
or ( n1700 , n1698 , n1699 );
and ( n1701 , n1572 , n1700 );
and ( n1702 , n1571 , n1700 );
or ( n1703 , n1573 , n1701 , n1702 );
xor ( n1704 , n1521 , n1534 );
xor ( n1705 , n1704 , n1537 );
and ( n1706 , n1703 , n1705 );
and ( n1707 , n1564 , n1360 );
and ( n1708 , n1526 , n1465 );
and ( n1709 , n1707 , n1708 );
buf ( n1710 , n1383 );
buf ( n1711 , n1710 );
and ( n1712 , n1441 , n1711 );
and ( n1713 , n1708 , n1712 );
and ( n1714 , n1707 , n1712 );
or ( n1715 , n1709 , n1713 , n1714 );
xor ( n1716 , n1577 , n1685 );
buf ( n1717 , n1716 );
buf ( n1718 , n1717 );
buf ( n1719 , n1718 );
and ( n1720 , n1291 , n1719 );
not ( n1721 , n1719 );
nor ( n1722 , n1720 , n1721 );
buf ( n1723 , n1717 );
buf ( n1724 , n1723 );
not ( n1725 , n1724 );
and ( n1726 , n1279 , n1724 );
nor ( n1727 , n1725 , n1726 );
and ( n1728 , n1722 , n1727 );
xor ( n1729 , n1171 , n1252 );
buf ( n1730 , n1729 );
buf ( n1731 , n1730 );
buf ( n1732 , n1731 );
and ( n1733 , n1732 , n1287 );
and ( n1734 , n1728 , n1733 );
and ( n1735 , n1472 , n1530 );
and ( n1736 , n1733 , n1735 );
and ( n1737 , n1728 , n1735 );
or ( n1738 , n1734 , n1736 , n1737 );
and ( n1739 , n1715 , n1738 );
and ( n1740 , n1275 , n1689 );
and ( n1741 , n1694 , n1293 );
and ( n1742 , n1740 , n1741 );
buf ( n1743 , n1385 );
or ( n1744 , n1742 , n1743 );
and ( n1745 , n1738 , n1744 );
and ( n1746 , n1715 , n1744 );
or ( n1747 , n1739 , n1745 , n1746 );
xor ( n1748 , n1522 , n1527 );
xor ( n1749 , n1748 , n1531 );
or ( n1750 , n1747 , n1749 );
and ( n1751 , n1705 , n1750 );
and ( n1752 , n1703 , n1750 );
or ( n1753 , n1706 , n1751 , n1752 );
and ( n1754 , n1559 , n1753 );
and ( n1755 , n1557 , n1753 );
or ( n1756 , n1560 , n1754 , n1755 );
and ( n1757 , n1555 , n1756 );
xor ( n1758 , n1555 , n1756 );
xor ( n1759 , n1557 , n1559 );
xor ( n1760 , n1759 , n1753 );
xor ( n1761 , n1571 , n1572 );
xor ( n1762 , n1761 , n1700 );
xnor ( n1763 , n1747 , n1749 );
and ( n1764 , n1762 , n1763 );
xnor ( n1765 , n1698 , n1699 );
xnor ( n1766 , n1742 , n1743 );
and ( n1767 , n1564 , n1465 );
and ( n1768 , n1526 , n1530 );
and ( n1769 , n1767 , n1768 );
and ( n1770 , n1472 , n1711 );
and ( n1771 , n1768 , n1770 );
and ( n1772 , n1767 , n1770 );
or ( n1773 , n1769 , n1771 , n1772 );
and ( n1774 , n1766 , n1773 );
xor ( n1775 , n1581 , n1684 );
buf ( n1776 , n1775 );
buf ( n1777 , n1776 );
buf ( n1778 , n1777 );
not ( n1779 , n1778 );
and ( n1780 , n1279 , n1778 );
nor ( n1781 , n1779 , n1780 );
and ( n1782 , n1724 , n1293 );
and ( n1783 , n1781 , n1782 );
and ( n1784 , n1694 , n1312 );
and ( n1785 , n1782 , n1784 );
and ( n1786 , n1781 , n1784 );
or ( n1787 , n1783 , n1785 , n1786 );
buf ( n1788 , n1776 );
buf ( n1789 , n1788 );
and ( n1790 , n1291 , n1789 );
not ( n1791 , n1789 );
nor ( n1792 , n1790 , n1791 );
and ( n1793 , n1275 , n1719 );
and ( n1794 , n1792 , n1793 );
and ( n1795 , n1317 , n1689 );
and ( n1796 , n1793 , n1795 );
and ( n1797 , n1792 , n1795 );
or ( n1798 , n1794 , n1796 , n1797 );
and ( n1799 , n1787 , n1798 );
and ( n1800 , n1773 , n1799 );
and ( n1801 , n1766 , n1799 );
or ( n1802 , n1774 , n1800 , n1801 );
and ( n1803 , n1765 , n1802 );
xor ( n1804 , n1565 , n1566 );
xor ( n1805 , n1804 , n1568 );
and ( n1806 , n1802 , n1805 );
and ( n1807 , n1765 , n1805 );
or ( n1808 , n1803 , n1806 , n1807 );
and ( n1809 , n1763 , n1808 );
and ( n1810 , n1762 , n1808 );
or ( n1811 , n1764 , n1809 , n1810 );
xor ( n1812 , n1703 , n1705 );
xor ( n1813 , n1812 , n1750 );
and ( n1814 , n1811 , n1813 );
xor ( n1815 , n1707 , n1708 );
xor ( n1816 , n1815 , n1712 );
xor ( n1817 , n1692 , n1697 );
and ( n1818 , n1816 , n1817 );
xor ( n1819 , n1715 , n1738 );
xor ( n1820 , n1819 , n1744 );
and ( n1821 , n1818 , n1820 );
xor ( n1822 , n1175 , n1251 );
buf ( n1823 , n1822 );
buf ( n1824 , n1823 );
buf ( n1825 , n1824 );
and ( n1826 , n1825 , n1287 );
and ( n1827 , n1732 , n1360 );
and ( n1828 , n1826 , n1827 );
xor ( n1829 , n1728 , n1733 );
xor ( n1830 , n1829 , n1735 );
and ( n1831 , n1828 , n1830 );
xor ( n1832 , n1722 , n1727 );
xor ( n1833 , n1740 , n1741 );
and ( n1834 , n1832 , n1833 );
xor ( n1835 , n1826 , n1827 );
and ( n1836 , n1833 , n1835 );
and ( n1837 , n1832 , n1835 );
or ( n1838 , n1834 , n1836 , n1837 );
and ( n1839 , n1830 , n1838 );
and ( n1840 , n1828 , n1838 );
or ( n1841 , n1831 , n1839 , n1840 );
xor ( n1842 , n1765 , n1802 );
xor ( n1843 , n1842 , n1805 );
and ( n1844 , n1841 , n1843 );
xor ( n1845 , n1816 , n1817 );
xor ( n1846 , n1766 , n1773 );
xor ( n1847 , n1846 , n1799 );
and ( n1848 , n1845 , n1847 );
xor ( n1849 , n1787 , n1798 );
and ( n1850 , n1275 , n1789 );
and ( n1851 , n1778 , n1293 );
and ( n1852 , n1850 , n1851 );
xor ( n1853 , n1179 , n1250 );
buf ( n1854 , n1853 );
buf ( n1855 , n1854 );
buf ( n1856 , n1855 );
and ( n1857 , n1856 , n1287 );
and ( n1858 , n1852 , n1857 );
buf ( n1859 , n1439 );
buf ( n1860 , n1859 );
and ( n1861 , n1472 , n1860 );
and ( n1862 , n1857 , n1861 );
and ( n1863 , n1852 , n1861 );
or ( n1864 , n1858 , n1862 , n1863 );
and ( n1865 , n1849 , n1864 );
xor ( n1866 , n1781 , n1782 );
xor ( n1867 , n1866 , n1784 );
xor ( n1868 , n1792 , n1793 );
xor ( n1869 , n1868 , n1795 );
and ( n1870 , n1867 , n1869 );
and ( n1871 , n1864 , n1870 );
and ( n1872 , n1849 , n1870 );
or ( n1873 , n1865 , n1871 , n1872 );
and ( n1874 , n1847 , n1873 );
and ( n1875 , n1845 , n1873 );
or ( n1876 , n1848 , n1874 , n1875 );
and ( n1877 , n1843 , n1876 );
and ( n1878 , n1841 , n1876 );
or ( n1879 , n1844 , n1877 , n1878 );
and ( n1880 , n1821 , n1879 );
xor ( n1881 , n1762 , n1763 );
xor ( n1882 , n1881 , n1808 );
and ( n1883 , n1879 , n1882 );
and ( n1884 , n1821 , n1882 );
or ( n1885 , n1880 , n1883 , n1884 );
and ( n1886 , n1813 , n1885 );
and ( n1887 , n1811 , n1885 );
or ( n1888 , n1814 , n1886 , n1887 );
and ( n1889 , n1760 , n1888 );
xor ( n1890 , n1760 , n1888 );
xor ( n1891 , n1811 , n1813 );
xor ( n1892 , n1891 , n1885 );
xor ( n1893 , n1818 , n1820 );
xor ( n1894 , n1828 , n1830 );
xor ( n1895 , n1894 , n1838 );
xor ( n1896 , n1832 , n1833 );
xor ( n1897 , n1896 , n1835 );
and ( n1898 , n1825 , n1360 );
and ( n1899 , n1564 , n1530 );
xor ( n1900 , n1898 , n1899 );
and ( n1901 , n1526 , n1711 );
xor ( n1902 , n1900 , n1901 );
xor ( n1903 , n1585 , n1683 );
buf ( n1904 , n1903 );
buf ( n1905 , n1904 );
buf ( n1906 , n1905 );
and ( n1907 , n1291 , n1906 );
not ( n1908 , n1906 );
nor ( n1909 , n1907 , n1908 );
buf ( n1910 , n1904 );
buf ( n1911 , n1910 );
not ( n1912 , n1911 );
and ( n1913 , n1279 , n1911 );
nor ( n1914 , n1912 , n1913 );
and ( n1915 , n1909 , n1914 );
and ( n1916 , n1317 , n1719 );
and ( n1917 , n1724 , n1312 );
and ( n1918 , n1916 , n1917 );
xor ( n1919 , n1915 , n1918 );
and ( n1920 , n1732 , n1465 );
xor ( n1921 , n1919 , n1920 );
and ( n1922 , n1902 , n1921 );
xor ( n1923 , n1852 , n1857 );
xor ( n1924 , n1923 , n1861 );
and ( n1925 , n1921 , n1924 );
and ( n1926 , n1902 , n1924 );
or ( n1927 , n1922 , n1925 , n1926 );
and ( n1928 , n1897 , n1927 );
xor ( n1929 , n1867 , n1869 );
xor ( n1930 , n1909 , n1914 );
xor ( n1931 , n1850 , n1851 );
and ( n1932 , n1930 , n1931 );
and ( n1933 , n1929 , n1932 );
and ( n1934 , n1927 , n1933 );
and ( n1935 , n1897 , n1933 );
or ( n1936 , n1928 , n1934 , n1935 );
and ( n1937 , n1895 , n1936 );
xor ( n1938 , n1845 , n1847 );
xor ( n1939 , n1938 , n1873 );
and ( n1940 , n1936 , n1939 );
and ( n1941 , n1895 , n1939 );
or ( n1942 , n1937 , n1940 , n1941 );
and ( n1943 , n1893 , n1942 );
xor ( n1944 , n1841 , n1843 );
xor ( n1945 , n1944 , n1876 );
and ( n1946 , n1942 , n1945 );
and ( n1947 , n1893 , n1945 );
or ( n1948 , n1943 , n1946 , n1947 );
xor ( n1949 , n1821 , n1879 );
xor ( n1950 , n1949 , n1882 );
and ( n1951 , n1948 , n1950 );
and ( n1952 , n1898 , n1899 );
and ( n1953 , n1899 , n1901 );
and ( n1954 , n1898 , n1901 );
or ( n1955 , n1952 , n1953 , n1954 );
and ( n1956 , n1915 , n1918 );
and ( n1957 , n1918 , n1920 );
and ( n1958 , n1915 , n1920 );
or ( n1959 , n1956 , n1957 , n1958 );
and ( n1960 , n1955 , n1959 );
buf ( n1961 , n1441 );
buf ( n1962 , n1961 );
and ( n1963 , n1959 , n1962 );
and ( n1964 , n1955 , n1962 );
or ( n1965 , n1960 , n1963 , n1964 );
and ( n1966 , n1275 , n1906 );
and ( n1967 , n1911 , n1293 );
and ( n1968 , n1966 , n1967 );
and ( n1969 , n1856 , n1360 );
and ( n1970 , n1968 , n1969 );
and ( n1971 , n1564 , n1711 );
and ( n1972 , n1969 , n1971 );
and ( n1973 , n1968 , n1971 );
or ( n1974 , n1970 , n1972 , n1973 );
and ( n1975 , n1317 , n1789 );
and ( n1976 , n1778 , n1312 );
and ( n1977 , n1975 , n1976 );
and ( n1978 , n1353 , n1719 );
and ( n1979 , n1724 , n1348 );
and ( n1980 , n1978 , n1979 );
and ( n1981 , n1977 , n1980 );
and ( n1982 , n1526 , n1860 );
and ( n1983 , n1980 , n1982 );
and ( n1984 , n1977 , n1982 );
or ( n1985 , n1981 , n1983 , n1984 );
and ( n1986 , n1974 , n1985 );
xor ( n1987 , n1589 , n1682 );
buf ( n1988 , n1987 );
buf ( n1989 , n1988 );
buf ( n1990 , n1989 );
and ( n1991 , n1291 , n1990 );
not ( n1992 , n1990 );
nor ( n1993 , n1991 , n1992 );
buf ( n1994 , n1988 );
buf ( n1995 , n1994 );
not ( n1996 , n1995 );
and ( n1997 , n1279 , n1995 );
nor ( n1998 , n1996 , n1997 );
and ( n1999 , n1993 , n1998 );
and ( n2000 , n1825 , n1465 );
and ( n2001 , n1999 , n2000 );
and ( n2002 , n1732 , n1530 );
and ( n2003 , n2000 , n2002 );
and ( n2004 , n1999 , n2002 );
or ( n2005 , n2001 , n2003 , n2004 );
and ( n2006 , n1985 , n2005 );
and ( n2007 , n1974 , n2005 );
or ( n2008 , n1986 , n2006 , n2007 );
xor ( n2009 , n1183 , n1249 );
buf ( n2010 , n2009 );
buf ( n2011 , n2010 );
buf ( n2012 , n2011 );
and ( n2013 , n2012 , n1287 );
buf ( n2014 , n2013 );
and ( n2015 , n1353 , n1689 );
and ( n2016 , n1694 , n1348 );
and ( n2017 , n2015 , n2016 );
and ( n2018 , n2014 , n2017 );
not ( n2019 , n1961 );
and ( n2020 , n2017 , n2019 );
and ( n2021 , n2014 , n2019 );
or ( n2022 , n2018 , n2020 , n2021 );
and ( n2023 , n2008 , n2022 );
xor ( n2024 , n1767 , n1768 );
xor ( n2025 , n2024 , n1770 );
and ( n2026 , n2022 , n2025 );
and ( n2027 , n2008 , n2025 );
or ( n2028 , n2023 , n2026 , n2027 );
and ( n2029 , n1965 , n2028 );
xor ( n2030 , n1849 , n1864 );
xor ( n2031 , n2030 , n1870 );
xor ( n2032 , n1187 , n1248 );
buf ( n2033 , n2032 );
buf ( n2034 , n2033 );
buf ( n2035 , n2034 );
and ( n2036 , n2035 , n1287 );
and ( n2037 , n1564 , n1860 );
and ( n2038 , n2036 , n2037 );
buf ( n2039 , n1470 );
buf ( n2040 , n2039 );
and ( n2041 , n1526 , n2040 );
and ( n2042 , n2037 , n2041 );
and ( n2043 , n2036 , n2041 );
or ( n2044 , n2038 , n2042 , n2043 );
xor ( n2045 , n1593 , n1681 );
buf ( n2046 , n2045 );
buf ( n2047 , n2046 );
buf ( n2048 , n2047 );
not ( n2049 , n2048 );
and ( n2050 , n1279 , n2048 );
nor ( n2051 , n2049 , n2050 );
and ( n2052 , n1995 , n1293 );
and ( n2053 , n2051 , n2052 );
and ( n2054 , n1778 , n1348 );
and ( n2055 , n2052 , n2054 );
and ( n2056 , n2051 , n2054 );
or ( n2057 , n2053 , n2055 , n2056 );
buf ( n2058 , n2046 );
buf ( n2059 , n2058 );
and ( n2060 , n1291 , n2059 );
not ( n2061 , n2059 );
nor ( n2062 , n2060 , n2061 );
and ( n2063 , n1275 , n1990 );
and ( n2064 , n2062 , n2063 );
and ( n2065 , n1353 , n1789 );
and ( n2066 , n2063 , n2065 );
and ( n2067 , n2062 , n2065 );
or ( n2068 , n2064 , n2066 , n2067 );
and ( n2069 , n2057 , n2068 );
and ( n2070 , n2044 , n2069 );
xor ( n2071 , n1968 , n1969 );
xor ( n2072 , n2071 , n1971 );
and ( n2073 , n2069 , n2072 );
and ( n2074 , n2044 , n2072 );
or ( n2075 , n2070 , n2073 , n2074 );
xor ( n2076 , n1974 , n1985 );
xor ( n2077 , n2076 , n2005 );
and ( n2078 , n2075 , n2077 );
xor ( n2079 , n1902 , n1921 );
xor ( n2080 , n2079 , n1924 );
and ( n2081 , n2077 , n2080 );
and ( n2082 , n2075 , n2080 );
or ( n2083 , n2078 , n2081 , n2082 );
and ( n2084 , n2031 , n2083 );
xor ( n2085 , n1897 , n1927 );
xor ( n2086 , n2085 , n1933 );
and ( n2087 , n2083 , n2086 );
and ( n2088 , n2031 , n2086 );
or ( n2089 , n2084 , n2087 , n2088 );
and ( n2090 , n2028 , n2089 );
and ( n2091 , n1965 , n2089 );
or ( n2092 , n2029 , n2090 , n2091 );
xor ( n2093 , n1893 , n1942 );
xor ( n2094 , n2093 , n1945 );
and ( n2095 , n2092 , n2094 );
xor ( n2096 , n1895 , n1936 );
xor ( n2097 , n2096 , n1939 );
and ( n2098 , n2012 , n1360 );
and ( n2099 , n1856 , n1465 );
and ( n2100 , n2098 , n2099 );
and ( n2101 , n1825 , n1530 );
and ( n2102 , n2099 , n2101 );
and ( n2103 , n2098 , n2101 );
or ( n2104 , n2100 , n2102 , n2103 );
buf ( n2105 , n1472 );
buf ( n2106 , n2105 );
and ( n2107 , n2104 , n2106 );
not ( n2108 , n2013 );
and ( n2109 , n2106 , n2108 );
and ( n2110 , n2104 , n2108 );
or ( n2111 , n2107 , n2109 , n2110 );
and ( n2112 , n1317 , n1906 );
and ( n2113 , n1911 , n1312 );
and ( n2114 , n2112 , n2113 );
and ( n2115 , n1732 , n1711 );
and ( n2116 , n2114 , n2115 );
not ( n2117 , n2105 );
and ( n2118 , n2115 , n2117 );
and ( n2119 , n2114 , n2117 );
or ( n2120 , n2116 , n2118 , n2119 );
xor ( n2121 , n1977 , n1980 );
xor ( n2122 , n2121 , n1982 );
and ( n2123 , n2120 , n2122 );
xor ( n2124 , n1999 , n2000 );
xor ( n2125 , n2124 , n2002 );
and ( n2126 , n2122 , n2125 );
and ( n2127 , n2120 , n2125 );
or ( n2128 , n2123 , n2126 , n2127 );
and ( n2129 , n2111 , n2128 );
xor ( n2130 , n2014 , n2017 );
xor ( n2131 , n2130 , n2019 );
and ( n2132 , n2128 , n2131 );
and ( n2133 , n2111 , n2131 );
or ( n2134 , n2129 , n2132 , n2133 );
xor ( n2135 , n2008 , n2022 );
xor ( n2136 , n2135 , n2025 );
or ( n2137 , n2134 , n2136 );
and ( n2138 , n2097 , n2137 );
xor ( n2139 , n1955 , n1959 );
xor ( n2140 , n2139 , n1962 );
xor ( n2141 , n1916 , n1917 );
xor ( n2142 , n2015 , n2016 );
and ( n2143 , n2141 , n2142 );
xor ( n2144 , n1993 , n1998 );
xor ( n2145 , n1966 , n1967 );
and ( n2146 , n2144 , n2145 );
and ( n2147 , n2142 , n2146 );
and ( n2148 , n2141 , n2146 );
or ( n2149 , n2143 , n2147 , n2148 );
xor ( n2150 , n1929 , n1932 );
and ( n2151 , n2149 , n2150 );
xor ( n2152 , n1930 , n1931 );
xor ( n2153 , n1975 , n1976 );
xor ( n2154 , n1978 , n1979 );
and ( n2155 , n2153 , n2154 );
xor ( n2156 , n2057 , n2068 );
and ( n2157 , n2154 , n2156 );
and ( n2158 , n2153 , n2156 );
or ( n2159 , n2155 , n2157 , n2158 );
and ( n2160 , n2152 , n2159 );
xor ( n2161 , n2141 , n2142 );
xor ( n2162 , n2161 , n2146 );
and ( n2163 , n2159 , n2162 );
and ( n2164 , n2152 , n2162 );
or ( n2165 , n2160 , n2163 , n2164 );
and ( n2166 , n2150 , n2165 );
and ( n2167 , n2149 , n2165 );
or ( n2168 , n2151 , n2166 , n2167 );
and ( n2169 , n2140 , n2168 );
xor ( n2170 , n2031 , n2083 );
xor ( n2171 , n2170 , n2086 );
and ( n2172 , n2168 , n2171 );
and ( n2173 , n2140 , n2171 );
or ( n2174 , n2169 , n2172 , n2173 );
and ( n2175 , n2137 , n2174 );
and ( n2176 , n2097 , n2174 );
or ( n2177 , n2138 , n2175 , n2176 );
and ( n2178 , n2094 , n2177 );
and ( n2179 , n2092 , n2177 );
or ( n2180 , n2095 , n2178 , n2179 );
and ( n2181 , n1950 , n2180 );
and ( n2182 , n1948 , n2180 );
or ( n2183 , n1951 , n2181 , n2182 );
and ( n2184 , n1892 , n2183 );
xor ( n2185 , n1892 , n2183 );
xor ( n2186 , n1948 , n1950 );
xor ( n2187 , n2186 , n2180 );
xor ( n2188 , n1965 , n2028 );
xor ( n2189 , n2188 , n2089 );
xnor ( n2190 , n2134 , n2136 );
and ( n2191 , n2012 , n1465 );
and ( n2192 , n1856 , n1530 );
and ( n2193 , n2191 , n2192 );
and ( n2194 , n1825 , n1711 );
and ( n2195 , n2192 , n2194 );
and ( n2196 , n2191 , n2194 );
or ( n2197 , n2193 , n2195 , n2196 );
and ( n2198 , n2035 , n1360 );
and ( n2199 , n1732 , n1860 );
and ( n2200 , n2198 , n2199 );
and ( n2201 , n1564 , n2040 );
and ( n2202 , n2199 , n2201 );
and ( n2203 , n2198 , n2201 );
or ( n2204 , n2200 , n2202 , n2203 );
and ( n2205 , n2197 , n2204 );
and ( n2206 , n1275 , n2059 );
and ( n2207 , n2048 , n1293 );
and ( n2208 , n2206 , n2207 );
buf ( n2209 , n2208 );
and ( n2210 , n2204 , n2209 );
and ( n2211 , n2197 , n2209 );
or ( n2212 , n2205 , n2210 , n2211 );
xor ( n2213 , n2104 , n2106 );
xor ( n2214 , n2213 , n2108 );
and ( n2215 , n2212 , n2214 );
xor ( n2216 , n2044 , n2069 );
xor ( n2217 , n2216 , n2072 );
and ( n2218 , n2214 , n2217 );
and ( n2219 , n2212 , n2217 );
or ( n2220 , n2215 , n2218 , n2219 );
xor ( n2221 , n2111 , n2128 );
xor ( n2222 , n2221 , n2131 );
and ( n2223 , n2220 , n2222 );
xor ( n2224 , n2075 , n2077 );
xor ( n2225 , n2224 , n2080 );
and ( n2226 , n2222 , n2225 );
and ( n2227 , n2220 , n2225 );
or ( n2228 , n2223 , n2226 , n2227 );
and ( n2229 , n2190 , n2228 );
xor ( n2230 , n2140 , n2168 );
xor ( n2231 , n2230 , n2171 );
and ( n2232 , n2228 , n2231 );
and ( n2233 , n2190 , n2231 );
or ( n2234 , n2229 , n2232 , n2233 );
and ( n2235 , n2189 , n2234 );
xor ( n2236 , n2097 , n2137 );
xor ( n2237 , n2236 , n2174 );
and ( n2238 , n2234 , n2237 );
and ( n2239 , n2189 , n2237 );
or ( n2240 , n2235 , n2238 , n2239 );
xor ( n2241 , n2092 , n2094 );
xor ( n2242 , n2241 , n2177 );
and ( n2243 , n2240 , n2242 );
xor ( n2244 , n2240 , n2242 );
xor ( n2245 , n2189 , n2234 );
xor ( n2246 , n2245 , n2237 );
xor ( n2247 , n1597 , n1680 );
buf ( n2248 , n2247 );
buf ( n2249 , n2248 );
buf ( n2250 , n2249 );
and ( n2251 , n1291 , n2250 );
not ( n2252 , n2250 );
nor ( n2253 , n2251 , n2252 );
buf ( n2254 , n2248 );
buf ( n2255 , n2254 );
not ( n2256 , n2255 );
and ( n2257 , n1279 , n2255 );
nor ( n2258 , n2256 , n2257 );
and ( n2259 , n2253 , n2258 );
and ( n2260 , n1317 , n1990 );
and ( n2261 , n1995 , n1312 );
and ( n2262 , n2260 , n2261 );
and ( n2263 , n2259 , n2262 );
xor ( n2264 , n1191 , n1247 );
buf ( n2265 , n2264 );
buf ( n2266 , n2265 );
buf ( n2267 , n2266 );
and ( n2268 , n2267 , n1287 );
and ( n2269 , n2262 , n2268 );
and ( n2270 , n2259 , n2268 );
or ( n2271 , n2263 , n2269 , n2270 );
xor ( n2272 , n2036 , n2037 );
xor ( n2273 , n2272 , n2041 );
and ( n2274 , n2271 , n2273 );
xor ( n2275 , n2114 , n2115 );
xor ( n2276 , n2275 , n2117 );
and ( n2277 , n2273 , n2276 );
and ( n2278 , n2271 , n2276 );
or ( n2279 , n2274 , n2277 , n2278 );
and ( n2280 , n1353 , n1990 );
and ( n2281 , n1995 , n1348 );
and ( n2282 , n2280 , n2281 );
xor ( n2283 , n1195 , n1246 );
buf ( n2284 , n2283 );
buf ( n2285 , n2284 );
buf ( n2286 , n2285 );
and ( n2287 , n2286 , n1287 );
and ( n2288 , n2282 , n2287 );
and ( n2289 , n1856 , n1711 );
and ( n2290 , n2287 , n2289 );
and ( n2291 , n2282 , n2289 );
or ( n2292 , n2288 , n2290 , n2291 );
and ( n2293 , n2267 , n1360 );
and ( n2294 , n1825 , n1860 );
and ( n2295 , n2293 , n2294 );
and ( n2296 , n1732 , n2040 );
and ( n2297 , n2294 , n2296 );
and ( n2298 , n2293 , n2296 );
or ( n2299 , n2295 , n2297 , n2298 );
and ( n2300 , n2292 , n2299 );
xor ( n2301 , n1601 , n1679 );
buf ( n2302 , n2301 );
buf ( n2303 , n2302 );
buf ( n2304 , n2303 );
and ( n2305 , n1291 , n2304 );
not ( n2306 , n2304 );
nor ( n2307 , n2305 , n2306 );
buf ( n2308 , n2302 );
buf ( n2309 , n2308 );
not ( n2310 , n2309 );
and ( n2311 , n1279 , n2309 );
nor ( n2312 , n2310 , n2311 );
and ( n2313 , n2307 , n2312 );
and ( n2314 , n2035 , n1465 );
and ( n2315 , n2313 , n2314 );
and ( n2316 , n2012 , n1530 );
and ( n2317 , n2314 , n2316 );
and ( n2318 , n2313 , n2316 );
or ( n2319 , n2315 , n2317 , n2318 );
and ( n2320 , n2299 , n2319 );
and ( n2321 , n2292 , n2319 );
or ( n2322 , n2300 , n2320 , n2321 );
xor ( n2323 , n2051 , n2052 );
xor ( n2324 , n2323 , n2054 );
xor ( n2325 , n2062 , n2063 );
xor ( n2326 , n2325 , n2065 );
and ( n2327 , n2324 , n2326 );
and ( n2328 , n2322 , n2327 );
xor ( n2329 , n2098 , n2099 );
xor ( n2330 , n2329 , n2101 );
and ( n2331 , n2327 , n2330 );
and ( n2332 , n2322 , n2330 );
or ( n2333 , n2328 , n2331 , n2332 );
and ( n2334 , n2279 , n2333 );
xor ( n2335 , n2120 , n2122 );
xor ( n2336 , n2335 , n2125 );
and ( n2337 , n2333 , n2336 );
and ( n2338 , n2279 , n2336 );
or ( n2339 , n2334 , n2337 , n2338 );
and ( n2340 , n1275 , n2250 );
and ( n2341 , n2255 , n1293 );
and ( n2342 , n2340 , n2341 );
buf ( n2343 , n1526 );
or ( n2344 , n2342 , n2343 );
not ( n2345 , n2208 );
and ( n2346 , n2344 , n2345 );
and ( n2347 , n1353 , n1906 );
and ( n2348 , n1911 , n1348 );
and ( n2349 , n2347 , n2348 );
and ( n2350 , n2345 , n2349 );
and ( n2351 , n2344 , n2349 );
or ( n2352 , n2346 , n2350 , n2351 );
xor ( n2353 , n2191 , n2192 );
xor ( n2354 , n2353 , n2194 );
xor ( n2355 , n2198 , n2199 );
xor ( n2356 , n2355 , n2201 );
and ( n2357 , n2354 , n2356 );
xor ( n2358 , n2259 , n2262 );
xor ( n2359 , n2358 , n2268 );
and ( n2360 , n2356 , n2359 );
and ( n2361 , n2354 , n2359 );
or ( n2362 , n2357 , n2360 , n2361 );
and ( n2363 , n2352 , n2362 );
xor ( n2364 , n2197 , n2204 );
xor ( n2365 , n2364 , n2209 );
and ( n2366 , n2362 , n2365 );
and ( n2367 , n2352 , n2365 );
or ( n2368 , n2363 , n2366 , n2367 );
xor ( n2369 , n2212 , n2214 );
xor ( n2370 , n2369 , n2217 );
and ( n2371 , n2368 , n2370 );
xor ( n2372 , n2279 , n2333 );
xor ( n2373 , n2372 , n2336 );
and ( n2374 , n2370 , n2373 );
and ( n2375 , n2368 , n2373 );
or ( n2376 , n2371 , n2374 , n2375 );
and ( n2377 , n2339 , n2376 );
xor ( n2378 , n2220 , n2222 );
xor ( n2379 , n2378 , n2225 );
and ( n2380 , n2376 , n2379 );
and ( n2381 , n2339 , n2379 );
or ( n2382 , n2377 , n2380 , n2381 );
xor ( n2383 , n2190 , n2228 );
xor ( n2384 , n2383 , n2231 );
and ( n2385 , n2382 , n2384 );
xor ( n2386 , n2149 , n2150 );
xor ( n2387 , n2386 , n2165 );
xor ( n2388 , n2144 , n2145 );
xor ( n2389 , n2271 , n2273 );
xor ( n2390 , n2389 , n2276 );
and ( n2391 , n2388 , n2390 );
xor ( n2392 , n2112 , n2113 );
xor ( n2393 , n2324 , n2326 );
and ( n2394 , n2392 , n2393 );
and ( n2395 , n2390 , n2394 );
and ( n2396 , n2388 , n2394 );
or ( n2397 , n2391 , n2395 , n2396 );
xor ( n2398 , n2152 , n2159 );
xor ( n2399 , n2398 , n2162 );
and ( n2400 , n2397 , n2399 );
xor ( n2401 , n2153 , n2154 );
xor ( n2402 , n2401 , n2156 );
xor ( n2403 , n2322 , n2327 );
xor ( n2404 , n2403 , n2330 );
and ( n2405 , n2402 , n2404 );
buf ( n2406 , n1524 );
buf ( n2407 , n2406 );
and ( n2408 , n1564 , n2407 );
xor ( n2409 , n2293 , n2294 );
xor ( n2410 , n2409 , n2296 );
and ( n2411 , n2408 , n2410 );
xor ( n2412 , n2253 , n2258 );
xor ( n2413 , n2206 , n2207 );
and ( n2414 , n2412 , n2413 );
xor ( n2415 , n2260 , n2261 );
and ( n2416 , n2413 , n2415 );
and ( n2417 , n2412 , n2415 );
or ( n2418 , n2414 , n2416 , n2417 );
and ( n2419 , n2411 , n2418 );
xor ( n2420 , n2292 , n2299 );
xor ( n2421 , n2420 , n2319 );
and ( n2422 , n2418 , n2421 );
and ( n2423 , n2411 , n2421 );
or ( n2424 , n2419 , n2422 , n2423 );
and ( n2425 , n2404 , n2424 );
and ( n2426 , n2402 , n2424 );
or ( n2427 , n2405 , n2425 , n2426 );
and ( n2428 , n2399 , n2427 );
and ( n2429 , n2397 , n2427 );
or ( n2430 , n2400 , n2428 , n2429 );
and ( n2431 , n2387 , n2430 );
xor ( n2432 , n2339 , n2376 );
xor ( n2433 , n2432 , n2379 );
and ( n2434 , n2430 , n2433 );
and ( n2435 , n2387 , n2433 );
or ( n2436 , n2431 , n2434 , n2435 );
and ( n2437 , n2384 , n2436 );
and ( n2438 , n2382 , n2436 );
or ( n2439 , n2385 , n2437 , n2438 );
and ( n2440 , n2246 , n2439 );
xor ( n2441 , n2246 , n2439 );
xor ( n2442 , n2344 , n2345 );
xor ( n2443 , n2442 , n2349 );
xor ( n2444 , n2354 , n2356 );
xor ( n2445 , n2444 , n2359 );
and ( n2446 , n2443 , n2445 );
xnor ( n2447 , n2342 , n2343 );
and ( n2448 , n1353 , n2059 );
and ( n2449 , n2048 , n1348 );
and ( n2450 , n2448 , n2449 );
and ( n2451 , n2286 , n1360 );
and ( n2452 , n2450 , n2451 );
and ( n2453 , n1732 , n2407 );
and ( n2454 , n2451 , n2453 );
and ( n2455 , n2450 , n2453 );
or ( n2456 , n2452 , n2454 , n2455 );
and ( n2457 , n2447 , n2456 );
and ( n2458 , n1317 , n2250 );
and ( n2459 , n2255 , n1312 );
and ( n2460 , n2458 , n2459 );
and ( n2461 , n2267 , n1465 );
and ( n2462 , n2460 , n2461 );
and ( n2463 , n2035 , n1530 );
and ( n2464 , n2461 , n2463 );
and ( n2465 , n2460 , n2463 );
or ( n2466 , n2462 , n2464 , n2465 );
and ( n2467 , n2456 , n2466 );
and ( n2468 , n2447 , n2466 );
or ( n2469 , n2457 , n2467 , n2468 );
and ( n2470 , n2445 , n2469 );
and ( n2471 , n2443 , n2469 );
or ( n2472 , n2446 , n2470 , n2471 );
xor ( n2473 , n1199 , n1200 );
xor ( n2474 , n2473 , n1243 );
buf ( n2475 , n2474 );
buf ( n2476 , n2475 );
buf ( n2477 , n2476 );
and ( n2478 , n2477 , n1287 );
and ( n2479 , n2012 , n1711 );
and ( n2480 , n2478 , n2479 );
and ( n2481 , n1825 , n2040 );
and ( n2482 , n2479 , n2481 );
and ( n2483 , n2478 , n2481 );
or ( n2484 , n2480 , n2482 , n2483 );
buf ( n2485 , n1694 );
buf ( n2486 , n1564 );
and ( n2487 , n2485 , n2486 );
xor ( n2488 , n1605 , n1606 );
xor ( n2489 , n2488 , n1676 );
buf ( n2490 , n2489 );
buf ( n2491 , n2490 );
buf ( n2492 , n2491 );
and ( n2493 , n1291 , n2492 );
not ( n2494 , n2492 );
nor ( n2495 , n2493 , n2494 );
buf ( n2496 , n2490 );
buf ( n2497 , n2496 );
not ( n2498 , n2497 );
and ( n2499 , n1279 , n2497 );
nor ( n2500 , n2498 , n2499 );
and ( n2501 , n2495 , n2500 );
and ( n2502 , n2487 , n2501 );
and ( n2503 , n1856 , n1860 );
and ( n2504 , n2501 , n2503 );
and ( n2505 , n2487 , n2503 );
or ( n2506 , n2502 , n2504 , n2505 );
and ( n2507 , n2484 , n2506 );
xor ( n2508 , n2282 , n2287 );
xor ( n2509 , n2508 , n2289 );
and ( n2510 , n2506 , n2509 );
and ( n2511 , n2484 , n2509 );
or ( n2512 , n2507 , n2510 , n2511 );
xor ( n2513 , n2347 , n2348 );
xor ( n2514 , n2313 , n2314 );
xor ( n2515 , n2514 , n2316 );
and ( n2516 , n2513 , n2515 );
and ( n2517 , n1275 , n2304 );
and ( n2518 , n2309 , n1293 );
and ( n2519 , n2517 , n2518 );
and ( n2520 , n1317 , n2059 );
or ( n2521 , n2519 , n2520 );
and ( n2522 , n2515 , n2521 );
and ( n2523 , n2513 , n2521 );
or ( n2524 , n2516 , n2522 , n2523 );
and ( n2525 , n2512 , n2524 );
and ( n2526 , n2048 , n1312 );
xor ( n2527 , n2307 , n2312 );
and ( n2528 , n2526 , n2527 );
xor ( n2529 , n2340 , n2341 );
xor ( n2530 , n2280 , n2281 );
and ( n2531 , n2529 , n2530 );
and ( n2532 , n2286 , n1465 );
and ( n2533 , n2267 , n1530 );
and ( n2534 , n2532 , n2533 );
and ( n2535 , n2530 , n2534 );
and ( n2536 , n2529 , n2534 );
or ( n2537 , n2531 , n2535 , n2536 );
and ( n2538 , n2528 , n2537 );
xor ( n2539 , n2408 , n2410 );
and ( n2540 , n2537 , n2539 );
and ( n2541 , n2528 , n2539 );
or ( n2542 , n2538 , n2540 , n2541 );
and ( n2543 , n2524 , n2542 );
and ( n2544 , n2512 , n2542 );
or ( n2545 , n2525 , n2543 , n2544 );
and ( n2546 , n2472 , n2545 );
xor ( n2547 , n2388 , n2390 );
xor ( n2548 , n2547 , n2394 );
and ( n2549 , n2545 , n2548 );
and ( n2550 , n2472 , n2548 );
or ( n2551 , n2546 , n2549 , n2550 );
xor ( n2552 , n2368 , n2370 );
xor ( n2553 , n2552 , n2373 );
and ( n2554 , n2551 , n2553 );
xor ( n2555 , n2352 , n2362 );
xor ( n2556 , n2555 , n2365 );
xor ( n2557 , n2392 , n2393 );
xor ( n2558 , n2412 , n2413 );
xor ( n2559 , n2558 , n2415 );
xor ( n2560 , n2447 , n2456 );
xor ( n2561 , n2560 , n2466 );
and ( n2562 , n2559 , n2561 );
xor ( n2563 , n2484 , n2506 );
xor ( n2564 , n2563 , n2509 );
and ( n2565 , n2561 , n2564 );
and ( n2566 , n2559 , n2564 );
or ( n2567 , n2562 , n2565 , n2566 );
and ( n2568 , n2557 , n2567 );
and ( n2569 , n1353 , n2250 );
and ( n2570 , n2255 , n1348 );
and ( n2571 , n2569 , n2570 );
and ( n2572 , n1694 , n1719 );
and ( n2573 , n1724 , n1689 );
and ( n2574 , n2572 , n2573 );
and ( n2575 , n2571 , n2574 );
buf ( n2576 , n1562 );
buf ( n2577 , n2576 );
and ( n2578 , n1732 , n2577 );
and ( n2579 , n2574 , n2578 );
and ( n2580 , n2571 , n2578 );
or ( n2581 , n2575 , n2579 , n2580 );
xor ( n2582 , n1611 , n1612 );
xor ( n2583 , n2582 , n1673 );
buf ( n2584 , n2583 );
buf ( n2585 , n2584 );
buf ( n2586 , n2585 );
and ( n2587 , n1291 , n2586 );
not ( n2588 , n2586 );
nor ( n2589 , n2587 , n2588 );
buf ( n2590 , n2584 );
buf ( n2591 , n2590 );
not ( n2592 , n2591 );
and ( n2593 , n1279 , n2591 );
nor ( n2594 , n2592 , n2593 );
and ( n2595 , n2589 , n2594 );
and ( n2596 , n1317 , n2304 );
and ( n2597 , n2309 , n1312 );
and ( n2598 , n2596 , n2597 );
and ( n2599 , n2595 , n2598 );
and ( n2600 , n1825 , n2407 );
and ( n2601 , n2598 , n2600 );
and ( n2602 , n2595 , n2600 );
or ( n2603 , n2599 , n2601 , n2602 );
and ( n2604 , n2581 , n2603 );
and ( n2605 , n2477 , n1360 );
and ( n2606 , n2012 , n1860 );
and ( n2607 , n2605 , n2606 );
and ( n2608 , n1856 , n2040 );
and ( n2609 , n2606 , n2608 );
and ( n2610 , n2605 , n2608 );
or ( n2611 , n2607 , n2609 , n2610 );
and ( n2612 , n2603 , n2611 );
and ( n2613 , n2581 , n2611 );
or ( n2614 , n2604 , n2612 , n2613 );
xor ( n2615 , n2478 , n2479 );
xor ( n2616 , n2615 , n2481 );
xor ( n2617 , n2450 , n2451 );
xor ( n2618 , n2617 , n2453 );
and ( n2619 , n2616 , n2618 );
xor ( n2620 , n2487 , n2501 );
xor ( n2621 , n2620 , n2503 );
and ( n2622 , n2618 , n2621 );
and ( n2623 , n2616 , n2621 );
or ( n2624 , n2619 , n2622 , n2623 );
and ( n2625 , n2614 , n2624 );
xnor ( n2626 , n2519 , n2520 );
and ( n2627 , n1275 , n2492 );
and ( n2628 , n2497 , n1293 );
and ( n2629 , n2627 , n2628 );
xor ( n2630 , n1205 , n1206 );
xor ( n2631 , n2630 , n1240 );
buf ( n2632 , n2631 );
buf ( n2633 , n2632 );
buf ( n2634 , n2633 );
and ( n2635 , n2634 , n1287 );
and ( n2636 , n2629 , n2635 );
and ( n2637 , n2035 , n1711 );
and ( n2638 , n2635 , n2637 );
and ( n2639 , n2629 , n2637 );
or ( n2640 , n2636 , n2638 , n2639 );
and ( n2641 , n2626 , n2640 );
xor ( n2642 , n2605 , n2606 );
xor ( n2643 , n2642 , n2608 );
xor ( n2644 , n2495 , n2500 );
and ( n2645 , n2643 , n2644 );
xor ( n2646 , n2517 , n2518 );
and ( n2647 , n2644 , n2646 );
and ( n2648 , n2643 , n2646 );
or ( n2649 , n2645 , n2647 , n2648 );
and ( n2650 , n2640 , n2649 );
and ( n2651 , n2626 , n2649 );
or ( n2652 , n2641 , n2650 , n2651 );
and ( n2653 , n2624 , n2652 );
and ( n2654 , n2614 , n2652 );
or ( n2655 , n2625 , n2653 , n2654 );
and ( n2656 , n2567 , n2655 );
and ( n2657 , n2557 , n2655 );
or ( n2658 , n2568 , n2656 , n2657 );
and ( n2659 , n2556 , n2658 );
xor ( n2660 , n2458 , n2459 );
xor ( n2661 , n2448 , n2449 );
and ( n2662 , n2660 , n2661 );
xor ( n2663 , n2532 , n2533 );
and ( n2664 , n2661 , n2663 );
and ( n2665 , n2660 , n2663 );
or ( n2666 , n2662 , n2664 , n2665 );
xor ( n2667 , n2526 , n2527 );
and ( n2668 , n2666 , n2667 );
xor ( n2669 , n2529 , n2530 );
xor ( n2670 , n2669 , n2534 );
and ( n2671 , n2667 , n2670 );
and ( n2672 , n2666 , n2670 );
or ( n2673 , n2668 , n2671 , n2672 );
xor ( n2674 , n2513 , n2515 );
xor ( n2675 , n2674 , n2521 );
and ( n2676 , n2673 , n2675 );
xor ( n2677 , n2528 , n2537 );
xor ( n2678 , n2677 , n2539 );
and ( n2679 , n2675 , n2678 );
and ( n2680 , n2673 , n2678 );
or ( n2681 , n2676 , n2679 , n2680 );
xor ( n2682 , n2411 , n2418 );
xor ( n2683 , n2682 , n2421 );
and ( n2684 , n2681 , n2683 );
xor ( n2685 , n2443 , n2445 );
xor ( n2686 , n2685 , n2469 );
and ( n2687 , n2683 , n2686 );
and ( n2688 , n2681 , n2686 );
or ( n2689 , n2684 , n2687 , n2688 );
and ( n2690 , n2658 , n2689 );
and ( n2691 , n2556 , n2689 );
or ( n2692 , n2659 , n2690 , n2691 );
and ( n2693 , n2553 , n2692 );
and ( n2694 , n2551 , n2692 );
or ( n2695 , n2554 , n2693 , n2694 );
xor ( n2696 , n2397 , n2399 );
xor ( n2697 , n2696 , n2427 );
xor ( n2698 , n2402 , n2404 );
xor ( n2699 , n2698 , n2424 );
xor ( n2700 , n2472 , n2545 );
xor ( n2701 , n2700 , n2548 );
and ( n2702 , n2699 , n2701 );
xor ( n2703 , n2512 , n2524 );
xor ( n2704 , n2703 , n2542 );
and ( n2705 , n1317 , n2492 );
and ( n2706 , n2497 , n1312 );
and ( n2707 , n2705 , n2706 );
and ( n2708 , n2634 , n1360 );
and ( n2709 , n2707 , n2708 );
and ( n2710 , n2477 , n1465 );
and ( n2711 , n2708 , n2710 );
and ( n2712 , n2707 , n2710 );
or ( n2713 , n2709 , n2711 , n2712 );
xor ( n2714 , n1617 , n1618 );
xor ( n2715 , n2714 , n1670 );
buf ( n2716 , n2715 );
buf ( n2717 , n2716 );
buf ( n2718 , n2717 );
and ( n2719 , n1291 , n2718 );
not ( n2720 , n2718 );
nor ( n2721 , n2719 , n2720 );
buf ( n2722 , n2716 );
buf ( n2723 , n2722 );
not ( n2724 , n2723 );
and ( n2725 , n1279 , n2723 );
nor ( n2726 , n2724 , n2725 );
and ( n2727 , n2721 , n2726 );
and ( n2728 , n1353 , n2304 );
and ( n2729 , n2309 , n1348 );
and ( n2730 , n2728 , n2729 );
and ( n2731 , n2727 , n2730 );
and ( n2732 , n2012 , n2040 );
and ( n2733 , n2730 , n2732 );
and ( n2734 , n2727 , n2732 );
or ( n2735 , n2731 , n2733 , n2734 );
and ( n2736 , n2713 , n2735 );
and ( n2737 , n1275 , n2586 );
and ( n2738 , n2591 , n1293 );
and ( n2739 , n2737 , n2738 );
and ( n2740 , n1694 , n1789 );
and ( n2741 , n1778 , n1689 );
and ( n2742 , n2740 , n2741 );
and ( n2743 , n2739 , n2742 );
and ( n2744 , n1856 , n2407 );
and ( n2745 , n2742 , n2744 );
and ( n2746 , n2739 , n2744 );
or ( n2747 , n2743 , n2745 , n2746 );
and ( n2748 , n2735 , n2747 );
and ( n2749 , n2713 , n2747 );
or ( n2750 , n2736 , n2748 , n2749 );
xor ( n2751 , n2485 , n2486 );
and ( n2752 , n2267 , n1711 );
and ( n2753 , n2035 , n1860 );
and ( n2754 , n2752 , n2753 );
and ( n2755 , n1825 , n2577 );
and ( n2756 , n2753 , n2755 );
and ( n2757 , n2752 , n2755 );
or ( n2758 , n2754 , n2756 , n2757 );
and ( n2759 , n2751 , n2758 );
xor ( n2760 , n1211 , n1212 );
xor ( n2761 , n2760 , n1237 );
buf ( n2762 , n2761 );
buf ( n2763 , n2762 );
buf ( n2764 , n2763 );
and ( n2765 , n2764 , n1287 );
buf ( n2766 , n2765 );
and ( n2767 , n2758 , n2766 );
and ( n2768 , n2751 , n2766 );
or ( n2769 , n2759 , n2767 , n2768 );
and ( n2770 , n2750 , n2769 );
xor ( n2771 , n2460 , n2461 );
xor ( n2772 , n2771 , n2463 );
and ( n2773 , n2769 , n2772 );
and ( n2774 , n2750 , n2772 );
or ( n2775 , n2770 , n2773 , n2774 );
xor ( n2776 , n2581 , n2603 );
xor ( n2777 , n2776 , n2611 );
xor ( n2778 , n2595 , n2598 );
xor ( n2779 , n2778 , n2600 );
xor ( n2780 , n2589 , n2594 );
xor ( n2781 , n2627 , n2628 );
and ( n2782 , n2780 , n2781 );
and ( n2783 , n2779 , n2782 );
xor ( n2784 , n2596 , n2597 );
xor ( n2785 , n2569 , n2570 );
and ( n2786 , n2784 , n2785 );
xor ( n2787 , n2572 , n2573 );
and ( n2788 , n2785 , n2787 );
and ( n2789 , n2784 , n2787 );
or ( n2790 , n2786 , n2788 , n2789 );
and ( n2791 , n2782 , n2790 );
and ( n2792 , n2779 , n2790 );
or ( n2793 , n2783 , n2791 , n2792 );
and ( n2794 , n2777 , n2793 );
xor ( n2795 , n2626 , n2640 );
xor ( n2796 , n2795 , n2649 );
and ( n2797 , n2793 , n2796 );
and ( n2798 , n2777 , n2796 );
or ( n2799 , n2794 , n2797 , n2798 );
and ( n2800 , n2775 , n2799 );
xor ( n2801 , n2559 , n2561 );
xor ( n2802 , n2801 , n2564 );
and ( n2803 , n2799 , n2802 );
and ( n2804 , n2775 , n2802 );
or ( n2805 , n2800 , n2803 , n2804 );
and ( n2806 , n2704 , n2805 );
xor ( n2807 , n2557 , n2567 );
xor ( n2808 , n2807 , n2655 );
and ( n2809 , n2805 , n2808 );
and ( n2810 , n2704 , n2808 );
or ( n2811 , n2806 , n2809 , n2810 );
and ( n2812 , n2701 , n2811 );
and ( n2813 , n2699 , n2811 );
or ( n2814 , n2702 , n2812 , n2813 );
and ( n2815 , n2697 , n2814 );
xor ( n2816 , n2551 , n2553 );
xor ( n2817 , n2816 , n2692 );
and ( n2818 , n2814 , n2817 );
and ( n2819 , n2697 , n2817 );
or ( n2820 , n2815 , n2818 , n2819 );
and ( n2821 , n2695 , n2820 );
xor ( n2822 , n2387 , n2430 );
xor ( n2823 , n2822 , n2433 );
and ( n2824 , n2820 , n2823 );
and ( n2825 , n2695 , n2823 );
or ( n2826 , n2821 , n2824 , n2825 );
xor ( n2827 , n2382 , n2384 );
xor ( n2828 , n2827 , n2436 );
and ( n2829 , n2826 , n2828 );
xor ( n2830 , n2826 , n2828 );
xor ( n2831 , n2695 , n2820 );
xor ( n2832 , n2831 , n2823 );
xor ( n2833 , n2556 , n2658 );
xor ( n2834 , n2833 , n2689 );
xor ( n2835 , n2681 , n2683 );
xor ( n2836 , n2835 , n2686 );
xor ( n2837 , n2614 , n2624 );
xor ( n2838 , n2837 , n2652 );
xor ( n2839 , n2673 , n2675 );
xor ( n2840 , n2839 , n2678 );
and ( n2841 , n2838 , n2840 );
buf ( n2842 , n1724 );
buf ( n2843 , n1732 );
and ( n2844 , n2842 , n2843 );
not ( n2845 , n2765 );
and ( n2846 , n2844 , n2845 );
and ( n2847 , n2286 , n1530 );
and ( n2848 , n2845 , n2847 );
and ( n2849 , n2844 , n2847 );
or ( n2850 , n2846 , n2848 , n2849 );
xor ( n2851 , n2571 , n2574 );
xor ( n2852 , n2851 , n2578 );
and ( n2853 , n2850 , n2852 );
xor ( n2854 , n2629 , n2635 );
xor ( n2855 , n2854 , n2637 );
and ( n2856 , n2852 , n2855 );
and ( n2857 , n2850 , n2855 );
or ( n2858 , n2853 , n2856 , n2857 );
xor ( n2859 , n2616 , n2618 );
xor ( n2860 , n2859 , n2621 );
and ( n2861 , n2858 , n2860 );
xor ( n2862 , n2750 , n2769 );
xor ( n2863 , n2862 , n2772 );
and ( n2864 , n2860 , n2863 );
and ( n2865 , n2858 , n2863 );
or ( n2866 , n2861 , n2864 , n2865 );
and ( n2867 , n2840 , n2866 );
and ( n2868 , n2838 , n2866 );
or ( n2869 , n2841 , n2867 , n2868 );
and ( n2870 , n2836 , n2869 );
xor ( n2871 , n2704 , n2805 );
xor ( n2872 , n2871 , n2808 );
and ( n2873 , n2869 , n2872 );
and ( n2874 , n2836 , n2872 );
or ( n2875 , n2870 , n2873 , n2874 );
and ( n2876 , n2834 , n2875 );
xor ( n2877 , n2699 , n2701 );
xor ( n2878 , n2877 , n2811 );
and ( n2879 , n2875 , n2878 );
and ( n2880 , n2834 , n2878 );
or ( n2881 , n2876 , n2879 , n2880 );
xor ( n2882 , n2697 , n2814 );
xor ( n2883 , n2882 , n2817 );
and ( n2884 , n2881 , n2883 );
xor ( n2885 , n2881 , n2883 );
xor ( n2886 , n2834 , n2875 );
xor ( n2887 , n2886 , n2878 );
xor ( n2888 , n2666 , n2667 );
xor ( n2889 , n2888 , n2670 );
and ( n2890 , n1275 , n2718 );
and ( n2891 , n2723 , n1293 );
and ( n2892 , n2890 , n2891 );
and ( n2893 , n1694 , n1906 );
and ( n2894 , n1911 , n1689 );
and ( n2895 , n2893 , n2894 );
and ( n2896 , n2892 , n2895 );
and ( n2897 , n2286 , n1711 );
and ( n2898 , n2895 , n2897 );
and ( n2899 , n2892 , n2897 );
or ( n2900 , n2896 , n2898 , n2899 );
and ( n2901 , n1724 , n1789 );
and ( n2902 , n1778 , n1719 );
and ( n2903 , n2901 , n2902 );
and ( n2904 , n2634 , n1465 );
and ( n2905 , n2903 , n2904 );
and ( n2906 , n2035 , n2040 );
and ( n2907 , n2904 , n2906 );
and ( n2908 , n2903 , n2906 );
or ( n2909 , n2905 , n2907 , n2908 );
and ( n2910 , n2900 , n2909 );
and ( n2911 , n1317 , n2586 );
and ( n2912 , n2591 , n1312 );
and ( n2913 , n2911 , n2912 );
and ( n2914 , n2764 , n1360 );
or ( n2915 , n2913 , n2914 );
and ( n2916 , n2909 , n2915 );
and ( n2917 , n2900 , n2915 );
or ( n2918 , n2910 , n2916 , n2917 );
xor ( n2919 , n1623 , n1624 );
xor ( n2920 , n2919 , n1667 );
buf ( n2921 , n2920 );
buf ( n2922 , n2921 );
buf ( n2923 , n2922 );
and ( n2924 , n1291 , n2923 );
not ( n2925 , n2923 );
nor ( n2926 , n2924 , n2925 );
buf ( n2927 , n2921 );
buf ( n2928 , n2927 );
not ( n2929 , n2928 );
and ( n2930 , n1279 , n2928 );
nor ( n2931 , n2929 , n2930 );
and ( n2932 , n2926 , n2931 );
xor ( n2933 , n1217 , n1218 );
xor ( n2934 , n2933 , n1234 );
buf ( n2935 , n2934 );
buf ( n2936 , n2935 );
buf ( n2937 , n2936 );
and ( n2938 , n2937 , n1287 );
and ( n2939 , n2932 , n2938 );
and ( n2940 , n1856 , n2577 );
and ( n2941 , n2938 , n2940 );
and ( n2942 , n2932 , n2940 );
or ( n2943 , n2939 , n2941 , n2942 );
and ( n2944 , n2477 , n1530 );
and ( n2945 , n2012 , n2407 );
and ( n2946 , n2944 , n2945 );
buf ( n2947 , n1730 );
buf ( n2948 , n2947 );
and ( n2949 , n1825 , n2948 );
and ( n2950 , n2945 , n2949 );
and ( n2951 , n2944 , n2949 );
or ( n2952 , n2946 , n2950 , n2951 );
and ( n2953 , n2943 , n2952 );
xor ( n2954 , n2842 , n2843 );
and ( n2955 , n1353 , n2492 );
and ( n2956 , n2497 , n1348 );
and ( n2957 , n2955 , n2956 );
and ( n2958 , n2954 , n2957 );
and ( n2959 , n2267 , n1860 );
and ( n2960 , n2957 , n2959 );
and ( n2961 , n2954 , n2959 );
or ( n2962 , n2958 , n2960 , n2961 );
and ( n2963 , n2952 , n2962 );
and ( n2964 , n2943 , n2962 );
or ( n2965 , n2953 , n2963 , n2964 );
and ( n2966 , n2918 , n2965 );
xor ( n2967 , n2751 , n2758 );
xor ( n2968 , n2967 , n2766 );
and ( n2969 , n2965 , n2968 );
and ( n2970 , n2918 , n2968 );
or ( n2971 , n2966 , n2969 , n2970 );
and ( n2972 , n2889 , n2971 );
xor ( n2973 , n2707 , n2708 );
xor ( n2974 , n2973 , n2710 );
xor ( n2975 , n2727 , n2730 );
xor ( n2976 , n2975 , n2732 );
and ( n2977 , n2974 , n2976 );
xor ( n2978 , n2739 , n2742 );
xor ( n2979 , n2978 , n2744 );
and ( n2980 , n2976 , n2979 );
and ( n2981 , n2974 , n2979 );
or ( n2982 , n2977 , n2980 , n2981 );
xor ( n2983 , n2713 , n2735 );
xor ( n2984 , n2983 , n2747 );
or ( n2985 , n2982 , n2984 );
and ( n2986 , n2971 , n2985 );
and ( n2987 , n2889 , n2985 );
or ( n2988 , n2972 , n2986 , n2987 );
xor ( n2989 , n2775 , n2799 );
xor ( n2990 , n2989 , n2802 );
and ( n2991 , n2988 , n2990 );
xor ( n2992 , n2643 , n2644 );
xor ( n2993 , n2992 , n2646 );
xor ( n2994 , n2660 , n2661 );
xor ( n2995 , n2994 , n2663 );
and ( n2996 , n2993 , n2995 );
xor ( n2997 , n2721 , n2726 );
xor ( n2998 , n2737 , n2738 );
and ( n2999 , n2997 , n2998 );
xor ( n3000 , n2705 , n2706 );
xor ( n3001 , n2728 , n2729 );
and ( n3002 , n3000 , n3001 );
xor ( n3003 , n2740 , n2741 );
and ( n3004 , n3001 , n3003 );
and ( n3005 , n3000 , n3003 );
or ( n3006 , n3002 , n3004 , n3005 );
and ( n3007 , n2999 , n3006 );
xor ( n3008 , n2780 , n2781 );
and ( n3009 , n3006 , n3008 );
and ( n3010 , n2999 , n3008 );
or ( n3011 , n3007 , n3009 , n3010 );
and ( n3012 , n2995 , n3011 );
and ( n3013 , n2993 , n3011 );
or ( n3014 , n2996 , n3012 , n3013 );
xor ( n3015 , n2777 , n2793 );
xor ( n3016 , n3015 , n2796 );
and ( n3017 , n3014 , n3016 );
xor ( n3018 , n2858 , n2860 );
xor ( n3019 , n3018 , n2863 );
and ( n3020 , n3016 , n3019 );
and ( n3021 , n3014 , n3019 );
or ( n3022 , n3017 , n3020 , n3021 );
and ( n3023 , n2990 , n3022 );
and ( n3024 , n2988 , n3022 );
or ( n3025 , n2991 , n3023 , n3024 );
xor ( n3026 , n2836 , n2869 );
xor ( n3027 , n3026 , n2872 );
and ( n3028 , n3025 , n3027 );
xor ( n3029 , n2779 , n2782 );
xor ( n3030 , n3029 , n2790 );
xor ( n3031 , n2918 , n2965 );
xor ( n3032 , n3031 , n2968 );
and ( n3033 , n3030 , n3032 );
xnor ( n3034 , n2982 , n2984 );
and ( n3035 , n3032 , n3034 );
and ( n3036 , n3030 , n3034 );
or ( n3037 , n3033 , n3035 , n3036 );
xor ( n3038 , n2932 , n2938 );
xor ( n3039 , n3038 , n2940 );
xor ( n3040 , n2892 , n2895 );
xor ( n3041 , n3040 , n2897 );
and ( n3042 , n3039 , n3041 );
xor ( n3043 , n2954 , n2957 );
xor ( n3044 , n3043 , n2959 );
and ( n3045 , n3041 , n3044 );
and ( n3046 , n3039 , n3044 );
or ( n3047 , n3042 , n3045 , n3046 );
xor ( n3048 , n2943 , n2952 );
xor ( n3049 , n3048 , n2962 );
and ( n3050 , n3047 , n3049 );
xor ( n3051 , n2974 , n2976 );
xor ( n3052 , n3051 , n2979 );
and ( n3053 , n3049 , n3052 );
and ( n3054 , n3047 , n3052 );
or ( n3055 , n3050 , n3053 , n3054 );
xor ( n3056 , n2784 , n2785 );
xor ( n3057 , n3056 , n2787 );
xor ( n3058 , n2926 , n2931 );
xor ( n3059 , n2890 , n2891 );
and ( n3060 , n3058 , n3059 );
xor ( n3061 , n2911 , n2912 );
xor ( n3062 , n2955 , n2956 );
and ( n3063 , n3061 , n3062 );
xor ( n3064 , n2893 , n2894 );
and ( n3065 , n3062 , n3064 );
and ( n3066 , n3061 , n3064 );
or ( n3067 , n3063 , n3065 , n3066 );
and ( n3068 , n3060 , n3067 );
xor ( n3069 , n2997 , n2998 );
and ( n3070 , n3067 , n3069 );
and ( n3071 , n3060 , n3069 );
or ( n3072 , n3068 , n3070 , n3071 );
and ( n3073 , n3057 , n3072 );
xor ( n3074 , n2999 , n3006 );
xor ( n3075 , n3074 , n3008 );
and ( n3076 , n3072 , n3075 );
and ( n3077 , n3057 , n3075 );
or ( n3078 , n3073 , n3076 , n3077 );
and ( n3079 , n3055 , n3078 );
xor ( n3080 , n2993 , n2995 );
xor ( n3081 , n3080 , n3011 );
and ( n3082 , n3078 , n3081 );
and ( n3083 , n3055 , n3081 );
or ( n3084 , n3079 , n3082 , n3083 );
and ( n3085 , n3037 , n3084 );
xor ( n3086 , n2889 , n2971 );
xor ( n3087 , n3086 , n2985 );
and ( n3088 , n3084 , n3087 );
and ( n3089 , n3037 , n3087 );
or ( n3090 , n3085 , n3088 , n3089 );
xor ( n3091 , n2838 , n2840 );
xor ( n3092 , n3091 , n2866 );
and ( n3093 , n3090 , n3092 );
and ( n3094 , n1353 , n2586 );
and ( n3095 , n2591 , n1348 );
and ( n3096 , n3094 , n3095 );
and ( n3097 , n1724 , n1906 );
and ( n3098 , n1911 , n1719 );
and ( n3099 , n3097 , n3098 );
and ( n3100 , n3096 , n3099 );
and ( n3101 , n2267 , n2040 );
and ( n3102 , n3099 , n3101 );
and ( n3103 , n3096 , n3101 );
or ( n3104 , n3100 , n3102 , n3103 );
and ( n3105 , n1317 , n2718 );
and ( n3106 , n2723 , n1312 );
and ( n3107 , n3105 , n3106 );
and ( n3108 , n2937 , n1360 );
and ( n3109 , n3107 , n3108 );
and ( n3110 , n2286 , n1860 );
and ( n3111 , n3108 , n3110 );
and ( n3112 , n3107 , n3110 );
or ( n3113 , n3109 , n3111 , n3112 );
and ( n3114 , n3104 , n3113 );
and ( n3115 , n1275 , n2923 );
and ( n3116 , n2928 , n1293 );
and ( n3117 , n3115 , n3116 );
and ( n3118 , n2764 , n1465 );
and ( n3119 , n3117 , n3118 );
and ( n3120 , n2035 , n2407 );
and ( n3121 , n3118 , n3120 );
and ( n3122 , n3117 , n3120 );
or ( n3123 , n3119 , n3121 , n3122 );
and ( n3124 , n3113 , n3123 );
and ( n3125 , n3104 , n3123 );
or ( n3126 , n3114 , n3124 , n3125 );
xor ( n3127 , n2752 , n2753 );
xor ( n3128 , n3127 , n2755 );
and ( n3129 , n3126 , n3128 );
xor ( n3130 , n2844 , n2845 );
xor ( n3131 , n3130 , n2847 );
and ( n3132 , n3128 , n3131 );
and ( n3133 , n3126 , n3131 );
or ( n3134 , n3129 , n3132 , n3133 );
and ( n3135 , n2477 , n1711 );
and ( n3136 , n2012 , n2577 );
and ( n3137 , n3135 , n3136 );
and ( n3138 , n1856 , n2948 );
and ( n3139 , n3136 , n3138 );
and ( n3140 , n3135 , n3138 );
or ( n3141 , n3137 , n3139 , n3140 );
xor ( n3142 , n1629 , n1630 );
xor ( n3143 , n3142 , n1664 );
buf ( n3144 , n3143 );
buf ( n3145 , n3144 );
buf ( n3146 , n3145 );
and ( n3147 , n1291 , n3146 );
not ( n3148 , n3146 );
nor ( n3149 , n3147 , n3148 );
buf ( n3150 , n3144 );
buf ( n3151 , n3150 );
not ( n3152 , n3151 );
and ( n3153 , n1279 , n3151 );
nor ( n3154 , n3152 , n3153 );
and ( n3155 , n3149 , n3154 );
and ( n3156 , n1694 , n1990 );
and ( n3157 , n1995 , n1689 );
and ( n3158 , n3156 , n3157 );
and ( n3159 , n3155 , n3158 );
and ( n3160 , n2634 , n1530 );
and ( n3161 , n3158 , n3160 );
and ( n3162 , n3155 , n3160 );
or ( n3163 , n3159 , n3161 , n3162 );
and ( n3164 , n3141 , n3163 );
xor ( n3165 , n1223 , n1224 );
xor ( n3166 , n3165 , n1231 );
buf ( n3167 , n3166 );
buf ( n3168 , n3167 );
buf ( n3169 , n3168 );
and ( n3170 , n3169 , n1287 );
buf ( n3171 , n3170 );
and ( n3172 , n3163 , n3171 );
and ( n3173 , n3141 , n3171 );
or ( n3174 , n3164 , n3172 , n3173 );
xnor ( n3175 , n2913 , n2914 );
xor ( n3176 , n2944 , n2945 );
xor ( n3177 , n3176 , n2949 );
and ( n3178 , n3175 , n3177 );
xor ( n3179 , n2903 , n2904 );
xor ( n3180 , n3179 , n2906 );
and ( n3181 , n3177 , n3180 );
and ( n3182 , n3175 , n3180 );
or ( n3183 , n3178 , n3181 , n3182 );
and ( n3184 , n3174 , n3183 );
xor ( n3185 , n2900 , n2909 );
xor ( n3186 , n3185 , n2915 );
and ( n3187 , n3183 , n3186 );
and ( n3188 , n3174 , n3186 );
or ( n3189 , n3184 , n3187 , n3188 );
and ( n3190 , n3134 , n3189 );
xor ( n3191 , n2850 , n2852 );
xor ( n3192 , n3191 , n2855 );
and ( n3193 , n3189 , n3192 );
and ( n3194 , n3134 , n3192 );
or ( n3195 , n3190 , n3193 , n3194 );
xor ( n3196 , n3014 , n3016 );
xor ( n3197 , n3196 , n3019 );
and ( n3198 , n3195 , n3197 );
xor ( n3199 , n3037 , n3084 );
xor ( n3200 , n3199 , n3087 );
and ( n3201 , n3197 , n3200 );
and ( n3202 , n3195 , n3200 );
or ( n3203 , n3198 , n3201 , n3202 );
and ( n3204 , n3092 , n3203 );
and ( n3205 , n3090 , n3203 );
or ( n3206 , n3093 , n3204 , n3205 );
and ( n3207 , n3027 , n3206 );
and ( n3208 , n3025 , n3206 );
or ( n3209 , n3028 , n3207 , n3208 );
and ( n3210 , n2887 , n3209 );
xor ( n3211 , n2887 , n3209 );
xor ( n3212 , n3025 , n3027 );
xor ( n3213 , n3212 , n3206 );
xor ( n3214 , n2988 , n2990 );
xor ( n3215 , n3214 , n3022 );
xor ( n3216 , n3090 , n3092 );
xor ( n3217 , n3216 , n3203 );
and ( n3218 , n3215 , n3217 );
xor ( n3219 , n3195 , n3197 );
xor ( n3220 , n3219 , n3200 );
and ( n3221 , n1275 , n3146 );
and ( n3222 , n3151 , n1293 );
and ( n3223 , n3221 , n3222 );
and ( n3224 , n2764 , n1530 );
and ( n3225 , n3223 , n3224 );
and ( n3226 , n2267 , n2407 );
and ( n3227 , n3224 , n3226 );
and ( n3228 , n3223 , n3226 );
or ( n3229 , n3225 , n3227 , n3228 );
and ( n3230 , n1353 , n2718 );
and ( n3231 , n2723 , n1348 );
and ( n3232 , n3230 , n3231 );
and ( n3233 , n2634 , n1711 );
and ( n3234 , n3232 , n3233 );
and ( n3235 , n2035 , n2577 );
and ( n3236 , n3233 , n3235 );
and ( n3237 , n3232 , n3235 );
or ( n3238 , n3234 , n3236 , n3237 );
and ( n3239 , n3229 , n3238 );
and ( n3240 , n1694 , n2059 );
and ( n3241 , n2048 , n1689 );
and ( n3242 , n3240 , n3241 );
xor ( n3243 , n1229 , n1230 );
buf ( n3244 , n3243 );
buf ( n3245 , n3244 );
buf ( n3246 , n3245 );
and ( n3247 , n3246 , n1287 );
and ( n3248 , n3242 , n3247 );
and ( n3249 , n2937 , n1465 );
and ( n3250 , n3247 , n3249 );
and ( n3251 , n3242 , n3249 );
or ( n3252 , n3248 , n3250 , n3251 );
and ( n3253 , n3238 , n3252 );
and ( n3254 , n3229 , n3252 );
or ( n3255 , n3239 , n3253 , n3254 );
buf ( n3256 , n1778 );
buf ( n3257 , n1825 );
and ( n3258 , n3256 , n3257 );
and ( n3259 , n1317 , n2923 );
and ( n3260 , n2928 , n1312 );
and ( n3261 , n3259 , n3260 );
and ( n3262 , n3169 , n1360 );
or ( n3263 , n3261 , n3262 );
and ( n3264 , n3258 , n3263 );
not ( n3265 , n3170 );
and ( n3266 , n3263 , n3265 );
and ( n3267 , n3258 , n3265 );
or ( n3268 , n3264 , n3266 , n3267 );
and ( n3269 , n3255 , n3268 );
xor ( n3270 , n3104 , n3113 );
xor ( n3271 , n3270 , n3123 );
and ( n3272 , n3268 , n3271 );
and ( n3273 , n3255 , n3271 );
or ( n3274 , n3269 , n3272 , n3273 );
and ( n3275 , n1778 , n1906 );
and ( n3276 , n1911 , n1789 );
and ( n3277 , n3275 , n3276 );
and ( n3278 , n2477 , n1860 );
and ( n3279 , n3277 , n3278 );
and ( n3280 , n2286 , n2040 );
and ( n3281 , n3278 , n3280 );
and ( n3282 , n3277 , n3280 );
or ( n3283 , n3279 , n3281 , n3282 );
xor ( n3284 , n1635 , n1636 );
xor ( n3285 , n3284 , n1661 );
buf ( n3286 , n3285 );
buf ( n3287 , n3286 );
buf ( n3288 , n3287 );
and ( n3289 , n1291 , n3288 );
not ( n3290 , n3288 );
nor ( n3291 , n3289 , n3290 );
buf ( n3292 , n3286 );
buf ( n3293 , n3292 );
not ( n3294 , n3293 );
and ( n3295 , n1279 , n3293 );
nor ( n3296 , n3294 , n3295 );
and ( n3297 , n3291 , n3296 );
and ( n3298 , n2012 , n2948 );
and ( n3299 , n3297 , n3298 );
buf ( n3300 , n1823 );
buf ( n3301 , n3300 );
and ( n3302 , n1856 , n3301 );
and ( n3303 , n3298 , n3302 );
and ( n3304 , n3297 , n3302 );
or ( n3305 , n3299 , n3303 , n3304 );
and ( n3306 , n3283 , n3305 );
xor ( n3307 , n3135 , n3136 );
xor ( n3308 , n3307 , n3138 );
and ( n3309 , n3305 , n3308 );
and ( n3310 , n3283 , n3308 );
or ( n3311 , n3306 , n3309 , n3310 );
xor ( n3312 , n3107 , n3108 );
xor ( n3313 , n3312 , n3110 );
xor ( n3314 , n3155 , n3158 );
xor ( n3315 , n3314 , n3160 );
and ( n3316 , n3313 , n3315 );
xor ( n3317 , n3117 , n3118 );
xor ( n3318 , n3317 , n3120 );
and ( n3319 , n3315 , n3318 );
and ( n3320 , n3313 , n3318 );
or ( n3321 , n3316 , n3319 , n3320 );
and ( n3322 , n3311 , n3321 );
xor ( n3323 , n3141 , n3163 );
xor ( n3324 , n3323 , n3171 );
and ( n3325 , n3321 , n3324 );
and ( n3326 , n3311 , n3324 );
or ( n3327 , n3322 , n3325 , n3326 );
and ( n3328 , n3274 , n3327 );
xor ( n3329 , n3126 , n3128 );
xor ( n3330 , n3329 , n3131 );
and ( n3331 , n3327 , n3330 );
and ( n3332 , n3274 , n3330 );
or ( n3333 , n3328 , n3331 , n3332 );
xor ( n3334 , n3256 , n3257 );
buf ( n3335 , n768 );
buf ( n3336 , n3335 );
buf ( n3337 , n3336 );
buf ( n3338 , n3337 );
buf ( n3339 , n3338 );
and ( n3340 , n3339 , n1287 );
buf ( n3341 , n3340 );
and ( n3342 , n3334 , n3341 );
and ( n3343 , n1724 , n1990 );
and ( n3344 , n1995 , n1719 );
and ( n3345 , n3343 , n3344 );
and ( n3346 , n3341 , n3345 );
and ( n3347 , n3334 , n3345 );
or ( n3348 , n3342 , n3346 , n3347 );
xor ( n3349 , n3096 , n3099 );
xor ( n3350 , n3349 , n3101 );
and ( n3351 , n3348 , n3350 );
xor ( n3352 , n3258 , n3263 );
xor ( n3353 , n3352 , n3265 );
and ( n3354 , n3350 , n3353 );
and ( n3355 , n3348 , n3353 );
or ( n3356 , n3351 , n3354 , n3355 );
xor ( n3357 , n3039 , n3041 );
xor ( n3358 , n3357 , n3044 );
and ( n3359 , n3356 , n3358 );
xor ( n3360 , n3175 , n3177 );
xor ( n3361 , n3360 , n3180 );
and ( n3362 , n3358 , n3361 );
and ( n3363 , n3356 , n3361 );
or ( n3364 , n3359 , n3362 , n3363 );
xor ( n3365 , n3174 , n3183 );
xor ( n3366 , n3365 , n3186 );
and ( n3367 , n3364 , n3366 );
xor ( n3368 , n3047 , n3049 );
xor ( n3369 , n3368 , n3052 );
and ( n3370 , n3366 , n3369 );
and ( n3371 , n3364 , n3369 );
or ( n3372 , n3367 , n3370 , n3371 );
and ( n3373 , n3333 , n3372 );
xor ( n3374 , n3134 , n3189 );
xor ( n3375 , n3374 , n3192 );
and ( n3376 , n3372 , n3375 );
and ( n3377 , n3333 , n3375 );
or ( n3378 , n3373 , n3376 , n3377 );
and ( n3379 , n3220 , n3378 );
xor ( n3380 , n3030 , n3032 );
xor ( n3381 , n3380 , n3034 );
xor ( n3382 , n3055 , n3078 );
xor ( n3383 , n3382 , n3081 );
and ( n3384 , n3381 , n3383 );
xor ( n3385 , n3000 , n3001 );
xor ( n3386 , n3385 , n3003 );
xor ( n3387 , n2901 , n2902 );
xor ( n3388 , n3149 , n3154 );
xor ( n3389 , n3115 , n3116 );
and ( n3390 , n3388 , n3389 );
and ( n3391 , n3387 , n3390 );
xor ( n3392 , n3105 , n3106 );
xor ( n3393 , n3094 , n3095 );
and ( n3394 , n3392 , n3393 );
xor ( n3395 , n3156 , n3157 );
and ( n3396 , n3393 , n3395 );
and ( n3397 , n3392 , n3395 );
or ( n3398 , n3394 , n3396 , n3397 );
and ( n3399 , n3390 , n3398 );
and ( n3400 , n3387 , n3398 );
or ( n3401 , n3391 , n3399 , n3400 );
and ( n3402 , n3386 , n3401 );
xor ( n3403 , n3060 , n3067 );
xor ( n3404 , n3403 , n3069 );
and ( n3405 , n3401 , n3404 );
and ( n3406 , n3386 , n3404 );
or ( n3407 , n3402 , n3405 , n3406 );
xor ( n3408 , n3057 , n3072 );
xor ( n3409 , n3408 , n3075 );
and ( n3410 , n3407 , n3409 );
xor ( n3411 , n3058 , n3059 );
xor ( n3412 , n3061 , n3062 );
xor ( n3413 , n3412 , n3064 );
and ( n3414 , n3411 , n3413 );
xor ( n3415 , n3097 , n3098 );
xor ( n3416 , n3291 , n3296 );
xor ( n3417 , n3221 , n3222 );
and ( n3418 , n3416 , n3417 );
and ( n3419 , n3415 , n3418 );
xor ( n3420 , n3259 , n3260 );
xor ( n3421 , n3230 , n3231 );
and ( n3422 , n3420 , n3421 );
xor ( n3423 , n3240 , n3241 );
and ( n3424 , n3421 , n3423 );
and ( n3425 , n3420 , n3423 );
or ( n3426 , n3422 , n3424 , n3425 );
and ( n3427 , n3418 , n3426 );
and ( n3428 , n3415 , n3426 );
or ( n3429 , n3419 , n3427 , n3428 );
and ( n3430 , n3413 , n3429 );
and ( n3431 , n3411 , n3429 );
or ( n3432 , n3414 , n3430 , n3431 );
xor ( n3433 , n3386 , n3401 );
xor ( n3434 , n3433 , n3404 );
and ( n3435 , n3432 , n3434 );
xor ( n3436 , n3387 , n3390 );
xor ( n3437 , n3436 , n3398 );
xor ( n3438 , n3388 , n3389 );
xor ( n3439 , n3392 , n3393 );
xor ( n3440 , n3439 , n3395 );
and ( n3441 , n3438 , n3440 );
xor ( n3442 , n3343 , n3344 );
xor ( n3443 , n3275 , n3276 );
and ( n3444 , n3442 , n3443 );
xor ( n3445 , n1641 , n1642 );
xor ( n3446 , n3445 , n1658 );
buf ( n3447 , n3446 );
buf ( n3448 , n3447 );
buf ( n3449 , n3448 );
and ( n3450 , n1291 , n3449 );
not ( n3451 , n3449 );
nor ( n3452 , n3450 , n3451 );
buf ( n3453 , n3447 );
buf ( n3454 , n3453 );
not ( n3455 , n3454 );
and ( n3456 , n1279 , n3454 );
nor ( n3457 , n3455 , n3456 );
xor ( n3458 , n3452 , n3457 );
and ( n3459 , n1275 , n3288 );
and ( n3460 , n3293 , n1293 );
xor ( n3461 , n3459 , n3460 );
and ( n3462 , n3458 , n3461 );
and ( n3463 , n3443 , n3462 );
and ( n3464 , n3442 , n3462 );
or ( n3465 , n3444 , n3463 , n3464 );
and ( n3466 , n3440 , n3465 );
and ( n3467 , n3438 , n3465 );
or ( n3468 , n3441 , n3466 , n3467 );
and ( n3469 , n3437 , n3468 );
xor ( n3470 , n3411 , n3413 );
xor ( n3471 , n3470 , n3429 );
and ( n3472 , n3468 , n3471 );
and ( n3473 , n3437 , n3471 );
or ( n3474 , n3469 , n3472 , n3473 );
and ( n3475 , n3434 , n3474 );
and ( n3476 , n3432 , n3474 );
or ( n3477 , n3435 , n3475 , n3476 );
and ( n3478 , n3409 , n3477 );
and ( n3479 , n3407 , n3477 );
or ( n3480 , n3410 , n3478 , n3479 );
and ( n3481 , n3383 , n3480 );
and ( n3482 , n3381 , n3480 );
or ( n3483 , n3384 , n3481 , n3482 );
and ( n3484 , n3378 , n3483 );
and ( n3485 , n3220 , n3483 );
or ( n3486 , n3379 , n3484 , n3485 );
and ( n3487 , n3217 , n3486 );
and ( n3488 , n3215 , n3486 );
or ( n3489 , n3218 , n3487 , n3488 );
and ( n3490 , n3213 , n3489 );
xor ( n3491 , n3213 , n3489 );
xor ( n3492 , n3215 , n3217 );
xor ( n3493 , n3492 , n3486 );
xor ( n3494 , n3333 , n3372 );
xor ( n3495 , n3494 , n3375 );
and ( n3496 , n3246 , n1360 );
and ( n3497 , n2477 , n2040 );
and ( n3498 , n3496 , n3497 );
and ( n3499 , n2286 , n2407 );
and ( n3500 , n3497 , n3499 );
and ( n3501 , n3496 , n3499 );
or ( n3502 , n3498 , n3500 , n3501 );
and ( n3503 , n3169 , n1465 );
and ( n3504 , n2634 , n1860 );
and ( n3505 , n3503 , n3504 );
and ( n3506 , n2267 , n2577 );
and ( n3507 , n3504 , n3506 );
and ( n3508 , n3503 , n3506 );
or ( n3509 , n3505 , n3507 , n3508 );
and ( n3510 , n3502 , n3509 );
and ( n3511 , n3452 , n3457 );
and ( n3512 , n1317 , n3146 );
and ( n3513 , n3151 , n1312 );
and ( n3514 , n3512 , n3513 );
and ( n3515 , n3511 , n3514 );
and ( n3516 , n2012 , n3301 );
and ( n3517 , n3514 , n3516 );
and ( n3518 , n3511 , n3516 );
or ( n3519 , n3515 , n3517 , n3518 );
and ( n3520 , n3509 , n3519 );
and ( n3521 , n3502 , n3519 );
or ( n3522 , n3510 , n3520 , n3521 );
buf ( n3523 , n1911 );
buf ( n3524 , n1856 );
and ( n3525 , n3523 , n3524 );
and ( n3526 , n1353 , n2923 );
and ( n3527 , n2928 , n1348 );
and ( n3528 , n3526 , n3527 );
and ( n3529 , n3525 , n3528 );
and ( n3530 , n1724 , n2059 );
and ( n3531 , n2048 , n1719 );
and ( n3532 , n3530 , n3531 );
and ( n3533 , n3528 , n3532 );
and ( n3534 , n3525 , n3532 );
or ( n3535 , n3529 , n3533 , n3534 );
xor ( n3536 , n3223 , n3224 );
xor ( n3537 , n3536 , n3226 );
and ( n3538 , n3535 , n3537 );
xor ( n3539 , n3232 , n3233 );
xor ( n3540 , n3539 , n3235 );
and ( n3541 , n3537 , n3540 );
and ( n3542 , n3535 , n3540 );
or ( n3543 , n3538 , n3541 , n3542 );
and ( n3544 , n3522 , n3543 );
xnor ( n3545 , n3261 , n3262 );
xor ( n3546 , n3297 , n3298 );
xor ( n3547 , n3546 , n3302 );
and ( n3548 , n3545 , n3547 );
xor ( n3549 , n3242 , n3247 );
xor ( n3550 , n3549 , n3249 );
and ( n3551 , n3547 , n3550 );
and ( n3552 , n3545 , n3550 );
or ( n3553 , n3548 , n3551 , n3552 );
and ( n3554 , n3543 , n3553 );
and ( n3555 , n3522 , n3553 );
or ( n3556 , n3544 , n3554 , n3555 );
and ( n3557 , n3459 , n3460 );
and ( n3558 , n1694 , n2250 );
and ( n3559 , n2255 , n1689 );
and ( n3560 , n3558 , n3559 );
and ( n3561 , n3557 , n3560 );
and ( n3562 , n2764 , n1711 );
and ( n3563 , n3560 , n3562 );
and ( n3564 , n3557 , n3562 );
or ( n3565 , n3561 , n3563 , n3564 );
and ( n3566 , n1778 , n1990 );
and ( n3567 , n1995 , n1789 );
and ( n3568 , n3566 , n3567 );
and ( n3569 , n2937 , n1530 );
and ( n3570 , n3568 , n3569 );
and ( n3571 , n2035 , n2948 );
and ( n3572 , n3569 , n3571 );
and ( n3573 , n3568 , n3571 );
or ( n3574 , n3570 , n3572 , n3573 );
and ( n3575 , n3565 , n3574 );
xor ( n3576 , n3277 , n3278 );
xor ( n3577 , n3576 , n3280 );
and ( n3578 , n3574 , n3577 );
and ( n3579 , n3565 , n3577 );
or ( n3580 , n3575 , n3578 , n3579 );
xor ( n3581 , n3229 , n3238 );
xor ( n3582 , n3581 , n3252 );
and ( n3583 , n3580 , n3582 );
xor ( n3584 , n3283 , n3305 );
xor ( n3585 , n3584 , n3308 );
and ( n3586 , n3582 , n3585 );
and ( n3587 , n3580 , n3585 );
or ( n3588 , n3583 , n3586 , n3587 );
and ( n3589 , n3556 , n3588 );
xor ( n3590 , n3255 , n3268 );
xor ( n3591 , n3590 , n3271 );
and ( n3592 , n3588 , n3591 );
and ( n3593 , n3556 , n3591 );
or ( n3594 , n3589 , n3592 , n3593 );
xor ( n3595 , n3274 , n3327 );
xor ( n3596 , n3595 , n3330 );
and ( n3597 , n3594 , n3596 );
xor ( n3598 , n3364 , n3366 );
xor ( n3599 , n3598 , n3369 );
and ( n3600 , n3596 , n3599 );
and ( n3601 , n3594 , n3599 );
or ( n3602 , n3597 , n3600 , n3601 );
and ( n3603 , n3495 , n3602 );
xor ( n3604 , n3381 , n3383 );
xor ( n3605 , n3604 , n3480 );
and ( n3606 , n3602 , n3605 );
and ( n3607 , n3495 , n3605 );
or ( n3608 , n3603 , n3606 , n3607 );
xor ( n3609 , n3220 , n3378 );
xor ( n3610 , n3609 , n3483 );
and ( n3611 , n3608 , n3610 );
and ( n3612 , n1275 , n3449 );
and ( n3613 , n3454 , n1293 );
and ( n3614 , n3612 , n3613 );
and ( n3615 , n1694 , n2304 );
and ( n3616 , n2309 , n1689 );
and ( n3617 , n3615 , n3616 );
and ( n3618 , n3614 , n3617 );
and ( n3619 , n3339 , n1360 );
and ( n3620 , n3617 , n3619 );
and ( n3621 , n3614 , n3619 );
or ( n3622 , n3618 , n3620 , n3621 );
and ( n3623 , n2764 , n1860 );
and ( n3624 , n2634 , n2040 );
and ( n3625 , n3623 , n3624 );
buf ( n3626 , n1854 );
buf ( n3627 , n3626 );
and ( n3628 , n2012 , n3627 );
and ( n3629 , n3624 , n3628 );
and ( n3630 , n3623 , n3628 );
or ( n3631 , n3625 , n3629 , n3630 );
and ( n3632 , n3622 , n3631 );
and ( n3633 , n1317 , n3288 );
and ( n3634 , n3293 , n1312 );
and ( n3635 , n3633 , n3634 );
and ( n3636 , n2477 , n2407 );
or ( n3637 , n3635 , n3636 );
and ( n3638 , n3631 , n3637 );
and ( n3639 , n3622 , n3637 );
or ( n3640 , n3632 , n3638 , n3639 );
buf ( n3641 , n769 );
buf ( n3642 , n3641 );
buf ( n3643 , n3642 );
buf ( n3644 , n3643 );
buf ( n3645 , n3644 );
and ( n3646 , n3645 , n1287 );
and ( n3647 , n3246 , n1465 );
and ( n3648 , n3646 , n3647 );
and ( n3649 , n2035 , n3301 );
and ( n3650 , n3647 , n3649 );
and ( n3651 , n3646 , n3649 );
or ( n3652 , n3648 , n3650 , n3651 );
and ( n3653 , n1353 , n3146 );
and ( n3654 , n3151 , n1348 );
and ( n3655 , n3653 , n3654 );
and ( n3656 , n1724 , n2250 );
and ( n3657 , n2255 , n1719 );
and ( n3658 , n3656 , n3657 );
and ( n3659 , n3655 , n3658 );
and ( n3660 , n3169 , n1530 );
and ( n3661 , n3658 , n3660 );
and ( n3662 , n3655 , n3660 );
or ( n3663 , n3659 , n3661 , n3662 );
and ( n3664 , n3652 , n3663 );
not ( n3665 , n3340 );
and ( n3666 , n3663 , n3665 );
and ( n3667 , n3652 , n3665 );
or ( n3668 , n3664 , n3666 , n3667 );
and ( n3669 , n3640 , n3668 );
xor ( n3670 , n3334 , n3341 );
xor ( n3671 , n3670 , n3345 );
and ( n3672 , n3668 , n3671 );
and ( n3673 , n3640 , n3671 );
or ( n3674 , n3669 , n3672 , n3673 );
xor ( n3675 , n3313 , n3315 );
xor ( n3676 , n3675 , n3318 );
and ( n3677 , n3674 , n3676 );
xor ( n3678 , n3348 , n3350 );
xor ( n3679 , n3678 , n3353 );
and ( n3680 , n3676 , n3679 );
and ( n3681 , n3674 , n3679 );
or ( n3682 , n3677 , n3680 , n3681 );
xor ( n3683 , n3311 , n3321 );
xor ( n3684 , n3683 , n3324 );
and ( n3685 , n3682 , n3684 );
xor ( n3686 , n3356 , n3358 );
xor ( n3687 , n3686 , n3361 );
and ( n3688 , n3684 , n3687 );
and ( n3689 , n3682 , n3687 );
or ( n3690 , n3685 , n3688 , n3689 );
xor ( n3691 , n3496 , n3497 );
xor ( n3692 , n3691 , n3499 );
xor ( n3693 , n3557 , n3560 );
xor ( n3694 , n3693 , n3562 );
and ( n3695 , n3692 , n3694 );
xor ( n3696 , n3568 , n3569 );
xor ( n3697 , n3696 , n3571 );
and ( n3698 , n3694 , n3697 );
and ( n3699 , n3692 , n3697 );
or ( n3700 , n3695 , n3698 , n3699 );
xor ( n3701 , n3502 , n3509 );
xor ( n3702 , n3701 , n3519 );
and ( n3703 , n3700 , n3702 );
xor ( n3704 , n3565 , n3574 );
xor ( n3705 , n3704 , n3577 );
and ( n3706 , n3702 , n3705 );
and ( n3707 , n3700 , n3705 );
or ( n3708 , n3703 , n3706 , n3707 );
xor ( n3709 , n3522 , n3543 );
xor ( n3710 , n3709 , n3553 );
and ( n3711 , n3708 , n3710 );
xor ( n3712 , n3580 , n3582 );
xor ( n3713 , n3712 , n3585 );
and ( n3714 , n3710 , n3713 );
and ( n3715 , n3708 , n3713 );
or ( n3716 , n3711 , n3714 , n3715 );
and ( n3717 , n2937 , n1711 );
and ( n3718 , n2286 , n2577 );
and ( n3719 , n3717 , n3718 );
and ( n3720 , n2267 , n2948 );
and ( n3721 , n3718 , n3720 );
and ( n3722 , n3717 , n3720 );
or ( n3723 , n3719 , n3721 , n3722 );
xor ( n3724 , n1647 , n1648 );
xor ( n3725 , n3724 , n1655 );
buf ( n3726 , n3725 );
buf ( n3727 , n3726 );
buf ( n3728 , n3727 );
not ( n3729 , n3728 );
and ( n3730 , n1279 , n3728 );
nor ( n3731 , n3729 , n3730 );
and ( n3732 , n2048 , n1789 );
and ( n3733 , n3731 , n3732 );
and ( n3734 , n1995 , n1906 );
and ( n3735 , n3732 , n3734 );
and ( n3736 , n3731 , n3734 );
or ( n3737 , n3733 , n3735 , n3736 );
buf ( n3738 , n3726 );
buf ( n3739 , n3738 );
and ( n3740 , n1291 , n3739 );
not ( n3741 , n3739 );
nor ( n3742 , n3740 , n3741 );
and ( n3743 , n1778 , n2059 );
and ( n3744 , n3742 , n3743 );
and ( n3745 , n1911 , n1990 );
and ( n3746 , n3743 , n3745 );
and ( n3747 , n3742 , n3745 );
or ( n3748 , n3744 , n3746 , n3747 );
and ( n3749 , n3737 , n3748 );
and ( n3750 , n3723 , n3749 );
xor ( n3751 , n3503 , n3504 );
xor ( n3752 , n3751 , n3506 );
and ( n3753 , n3749 , n3752 );
and ( n3754 , n3723 , n3752 );
or ( n3755 , n3750 , n3753 , n3754 );
xor ( n3756 , n3535 , n3537 );
xor ( n3757 , n3756 , n3540 );
and ( n3758 , n3755 , n3757 );
xor ( n3759 , n3545 , n3547 );
xor ( n3760 , n3759 , n3550 );
and ( n3761 , n3757 , n3760 );
and ( n3762 , n3755 , n3760 );
or ( n3763 , n3758 , n3761 , n3762 );
xnor ( n3764 , n3635 , n3636 );
and ( n3765 , n1778 , n2250 );
and ( n3766 , n2255 , n1789 );
and ( n3767 , n3765 , n3766 );
and ( n3768 , n2286 , n2948 );
and ( n3769 , n3767 , n3768 );
and ( n3770 , n2267 , n3301 );
and ( n3771 , n3768 , n3770 );
and ( n3772 , n3767 , n3770 );
or ( n3773 , n3769 , n3771 , n3772 );
and ( n3774 , n3764 , n3773 );
and ( n3775 , n3728 , n1293 );
and ( n3776 , n2497 , n1689 );
and ( n3777 , n3775 , n3776 );
and ( n3778 , n2048 , n1906 );
and ( n3779 , n3776 , n3778 );
and ( n3780 , n3775 , n3778 );
or ( n3781 , n3777 , n3779 , n3780 );
and ( n3782 , n1275 , n3739 );
and ( n3783 , n1694 , n2492 );
and ( n3784 , n3782 , n3783 );
and ( n3785 , n1911 , n2059 );
and ( n3786 , n3783 , n3785 );
and ( n3787 , n3782 , n3785 );
or ( n3788 , n3784 , n3786 , n3787 );
and ( n3789 , n3781 , n3788 );
and ( n3790 , n3773 , n3789 );
and ( n3791 , n3764 , n3789 );
or ( n3792 , n3774 , n3790 , n3791 );
xor ( n3793 , n3646 , n3647 );
xor ( n3794 , n3793 , n3649 );
xor ( n3795 , n3614 , n3617 );
xor ( n3796 , n3795 , n3619 );
and ( n3797 , n3794 , n3796 );
xor ( n3798 , n3623 , n3624 );
xor ( n3799 , n3798 , n3628 );
and ( n3800 , n3796 , n3799 );
and ( n3801 , n3794 , n3799 );
or ( n3802 , n3797 , n3800 , n3801 );
and ( n3803 , n3792 , n3802 );
xor ( n3804 , n3731 , n3732 );
xor ( n3805 , n3804 , n3734 );
xor ( n3806 , n3742 , n3743 );
xor ( n3807 , n3806 , n3745 );
and ( n3808 , n3805 , n3807 );
xor ( n3809 , n3655 , n3658 );
xor ( n3810 , n3809 , n3660 );
and ( n3811 , n3808 , n3810 );
xor ( n3812 , n3717 , n3718 );
xor ( n3813 , n3812 , n3720 );
and ( n3814 , n3810 , n3813 );
and ( n3815 , n3808 , n3813 );
or ( n3816 , n3811 , n3814 , n3815 );
and ( n3817 , n3802 , n3816 );
and ( n3818 , n3792 , n3816 );
or ( n3819 , n3803 , n3817 , n3818 );
xor ( n3820 , n3523 , n3524 );
and ( n3821 , n3246 , n1530 );
and ( n3822 , n2764 , n2040 );
and ( n3823 , n3821 , n3822 );
and ( n3824 , n2634 , n2407 );
and ( n3825 , n3822 , n3824 );
and ( n3826 , n3821 , n3824 );
or ( n3827 , n3823 , n3825 , n3826 );
and ( n3828 , n3820 , n3827 );
buf ( n3829 , n770 );
buf ( n3830 , n3829 );
buf ( n3831 , n3830 );
buf ( n3832 , n3831 );
buf ( n3833 , n3832 );
and ( n3834 , n3833 , n1287 );
buf ( n3835 , n3834 );
and ( n3836 , n3827 , n3835 );
and ( n3837 , n3820 , n3835 );
or ( n3838 , n3828 , n3836 , n3837 );
xor ( n3839 , n3525 , n3528 );
xor ( n3840 , n3839 , n3532 );
and ( n3841 , n3838 , n3840 );
xor ( n3842 , n3511 , n3514 );
xor ( n3843 , n3842 , n3516 );
and ( n3844 , n3840 , n3843 );
and ( n3845 , n3838 , n3843 );
or ( n3846 , n3841 , n3844 , n3845 );
and ( n3847 , n3819 , n3846 );
xor ( n3848 , n3640 , n3668 );
xor ( n3849 , n3848 , n3671 );
and ( n3850 , n3846 , n3849 );
and ( n3851 , n3819 , n3849 );
or ( n3852 , n3847 , n3850 , n3851 );
and ( n3853 , n3763 , n3852 );
xor ( n3854 , n3674 , n3676 );
xor ( n3855 , n3854 , n3679 );
and ( n3856 , n3852 , n3855 );
and ( n3857 , n3763 , n3855 );
or ( n3858 , n3853 , n3856 , n3857 );
and ( n3859 , n3716 , n3858 );
xor ( n3860 , n3556 , n3588 );
xor ( n3861 , n3860 , n3591 );
and ( n3862 , n3858 , n3861 );
and ( n3863 , n3716 , n3861 );
or ( n3864 , n3859 , n3862 , n3863 );
and ( n3865 , n3690 , n3864 );
xor ( n3866 , n3594 , n3596 );
xor ( n3867 , n3866 , n3599 );
and ( n3868 , n3864 , n3867 );
and ( n3869 , n3690 , n3867 );
or ( n3870 , n3865 , n3868 , n3869 );
xor ( n3871 , n3495 , n3602 );
xor ( n3872 , n3871 , n3605 );
and ( n3873 , n3870 , n3872 );
and ( n3874 , n3645 , n1360 );
and ( n3875 , n3169 , n1711 );
and ( n3876 , n3874 , n3875 );
and ( n3877 , n2477 , n2577 );
and ( n3878 , n3875 , n3877 );
and ( n3879 , n3874 , n3877 );
or ( n3880 , n3876 , n3878 , n3879 );
and ( n3881 , n3339 , n1465 );
and ( n3882 , n2937 , n1860 );
and ( n3883 , n3881 , n3882 );
and ( n3884 , n2035 , n3627 );
and ( n3885 , n3882 , n3884 );
and ( n3886 , n3881 , n3884 );
or ( n3887 , n3883 , n3885 , n3886 );
and ( n3888 , n3880 , n3887 );
xor ( n3889 , n1653 , n1654 );
buf ( n3890 , n3889 );
buf ( n3891 , n3890 );
buf ( n3892 , n3891 );
not ( n3893 , n3892 );
and ( n3894 , n1279 , n3892 );
nor ( n3895 , n3893 , n3894 );
and ( n3896 , n3454 , n1312 );
and ( n3897 , n3895 , n3896 );
and ( n3898 , n3293 , n1348 );
and ( n3899 , n3896 , n3898 );
and ( n3900 , n3895 , n3898 );
or ( n3901 , n3897 , n3899 , n3900 );
buf ( n3902 , n3890 );
buf ( n3903 , n3902 );
and ( n3904 , n1291 , n3903 );
not ( n3905 , n3903 );
nor ( n3906 , n3904 , n3905 );
and ( n3907 , n1317 , n3449 );
and ( n3908 , n3906 , n3907 );
and ( n3909 , n1353 , n3288 );
and ( n3910 , n3907 , n3909 );
and ( n3911 , n3906 , n3909 );
or ( n3912 , n3908 , n3910 , n3911 );
and ( n3913 , n3901 , n3912 );
and ( n3914 , n3887 , n3913 );
and ( n3915 , n3880 , n3913 );
or ( n3916 , n3888 , n3914 , n3915 );
xor ( n3917 , n3652 , n3663 );
xor ( n3918 , n3917 , n3665 );
and ( n3919 , n3916 , n3918 );
xor ( n3920 , n3723 , n3749 );
xor ( n3921 , n3920 , n3752 );
and ( n3922 , n3918 , n3921 );
and ( n3923 , n3916 , n3921 );
or ( n3924 , n3919 , n3922 , n3923 );
and ( n3925 , n3246 , n1711 );
and ( n3926 , n2764 , n2407 );
and ( n3927 , n3925 , n3926 );
buf ( n3928 , n2010 );
buf ( n3929 , n3928 );
and ( n3930 , n2035 , n3929 );
and ( n3931 , n3926 , n3930 );
and ( n3932 , n3925 , n3930 );
or ( n3933 , n3927 , n3931 , n3932 );
and ( n3934 , n1778 , n2304 );
and ( n3935 , n2309 , n1789 );
and ( n3936 , n3934 , n3935 );
and ( n3937 , n3339 , n1530 );
and ( n3938 , n3936 , n3937 );
and ( n3939 , n2477 , n2948 );
and ( n3940 , n3937 , n3939 );
and ( n3941 , n3936 , n3939 );
or ( n3942 , n3938 , n3940 , n3941 );
and ( n3943 , n3933 , n3942 );
and ( n3944 , n1995 , n2059 );
and ( n3945 , n2048 , n1990 );
and ( n3946 , n3944 , n3945 );
and ( n3947 , n2937 , n2040 );
or ( n3948 , n3946 , n3947 );
and ( n3949 , n3942 , n3948 );
and ( n3950 , n3933 , n3948 );
or ( n3951 , n3943 , n3949 , n3950 );
buf ( n3952 , n1995 );
buf ( n3953 , n2012 );
and ( n3954 , n3952 , n3953 );
and ( n3955 , n1724 , n2304 );
and ( n3956 , n2309 , n1719 );
and ( n3957 , n3955 , n3956 );
and ( n3958 , n3954 , n3957 );
not ( n3959 , n3834 );
and ( n3960 , n3957 , n3959 );
and ( n3961 , n3954 , n3959 );
or ( n3962 , n3958 , n3960 , n3961 );
and ( n3963 , n3951 , n3962 );
xor ( n3964 , n3820 , n3827 );
xor ( n3965 , n3964 , n3835 );
and ( n3966 , n3962 , n3965 );
and ( n3967 , n3951 , n3965 );
or ( n3968 , n3963 , n3966 , n3967 );
xor ( n3969 , n3622 , n3631 );
xor ( n3970 , n3969 , n3637 );
and ( n3971 , n3968 , n3970 );
xor ( n3972 , n3692 , n3694 );
xor ( n3973 , n3972 , n3697 );
and ( n3974 , n3970 , n3973 );
and ( n3975 , n3968 , n3973 );
or ( n3976 , n3971 , n3974 , n3975 );
and ( n3977 , n3924 , n3976 );
xor ( n3978 , n3700 , n3702 );
xor ( n3979 , n3978 , n3705 );
and ( n3980 , n3976 , n3979 );
and ( n3981 , n3924 , n3979 );
or ( n3982 , n3977 , n3980 , n3981 );
xor ( n3983 , n3708 , n3710 );
xor ( n3984 , n3983 , n3713 );
and ( n3985 , n3982 , n3984 );
xor ( n3986 , n3763 , n3852 );
xor ( n3987 , n3986 , n3855 );
and ( n3988 , n3984 , n3987 );
and ( n3989 , n3982 , n3987 );
or ( n3990 , n3985 , n3988 , n3989 );
xor ( n3991 , n3682 , n3684 );
xor ( n3992 , n3991 , n3687 );
and ( n3993 , n3990 , n3992 );
xor ( n3994 , n3716 , n3858 );
xor ( n3995 , n3994 , n3861 );
and ( n3996 , n3992 , n3995 );
and ( n3997 , n3990 , n3995 );
or ( n3998 , n3993 , n3996 , n3997 );
xor ( n3999 , n3690 , n3864 );
xor ( n4000 , n3999 , n3867 );
and ( n4001 , n3998 , n4000 );
and ( n4002 , n3872 , n4001 );
and ( n4003 , n3870 , n4001 );
or ( n4004 , n3873 , n4002 , n4003 );
and ( n4005 , n3610 , n4004 );
and ( n4006 , n3608 , n4004 );
or ( n4007 , n3611 , n4005 , n4006 );
and ( n4008 , n3493 , n4007 );
xor ( n4009 , n3493 , n4007 );
xor ( n4010 , n3608 , n3610 );
xor ( n4011 , n4010 , n4004 );
xor ( n4012 , n3407 , n3409 );
xor ( n4013 , n4012 , n3477 );
xor ( n4014 , n3998 , n4000 );
and ( n4015 , n4013 , n4014 );
xor ( n4016 , n3432 , n3434 );
xor ( n4017 , n4016 , n3474 );
xor ( n4018 , n3512 , n3513 );
xor ( n4019 , n3526 , n3527 );
and ( n4020 , n4018 , n4019 );
xor ( n4021 , n3558 , n3559 );
and ( n4022 , n4019 , n4021 );
and ( n4023 , n4018 , n4021 );
or ( n4024 , n4020 , n4022 , n4023 );
xor ( n4025 , n3416 , n3417 );
and ( n4026 , n4024 , n4025 );
xor ( n4027 , n3420 , n3421 );
xor ( n4028 , n4027 , n3423 );
and ( n4029 , n4025 , n4028 );
and ( n4030 , n4024 , n4028 );
or ( n4031 , n4026 , n4029 , n4030 );
xor ( n4032 , n3415 , n3418 );
xor ( n4033 , n4032 , n3426 );
and ( n4034 , n4031 , n4033 );
xor ( n4035 , n3530 , n3531 );
xor ( n4036 , n3566 , n3567 );
and ( n4037 , n4035 , n4036 );
xor ( n4038 , n3737 , n3748 );
and ( n4039 , n4036 , n4038 );
and ( n4040 , n4035 , n4038 );
or ( n4041 , n4037 , n4039 , n4040 );
xor ( n4042 , n3612 , n3613 );
xor ( n4043 , n3633 , n3634 );
and ( n4044 , n4042 , n4043 );
xor ( n4045 , n3653 , n3654 );
xor ( n4046 , n3615 , n3616 );
and ( n4047 , n4045 , n4046 );
xor ( n4048 , n3656 , n3657 );
and ( n4049 , n4046 , n4048 );
and ( n4050 , n4045 , n4048 );
or ( n4051 , n4047 , n4049 , n4050 );
and ( n4052 , n4044 , n4051 );
xor ( n4053 , n3458 , n3461 );
and ( n4054 , n4051 , n4053 );
and ( n4055 , n4044 , n4053 );
or ( n4056 , n4052 , n4054 , n4055 );
and ( n4057 , n4041 , n4056 );
xor ( n4058 , n3442 , n3443 );
xor ( n4059 , n4058 , n3462 );
and ( n4060 , n4056 , n4059 );
and ( n4061 , n4041 , n4059 );
or ( n4062 , n4057 , n4060 , n4061 );
and ( n4063 , n4033 , n4062 );
and ( n4064 , n4031 , n4062 );
or ( n4065 , n4034 , n4063 , n4064 );
xor ( n4066 , n3437 , n3468 );
xor ( n4067 , n4066 , n3471 );
and ( n4068 , n4065 , n4067 );
xor ( n4069 , n3438 , n3440 );
xor ( n4070 , n4069 , n3465 );
xor ( n4071 , n4024 , n4025 );
xor ( n4072 , n4071 , n4028 );
xor ( n4073 , n4018 , n4019 );
xor ( n4074 , n4073 , n4021 );
xor ( n4075 , n3901 , n3912 );
xor ( n4076 , n3781 , n3788 );
and ( n4077 , n4075 , n4076 );
xor ( n4078 , n3805 , n3807 );
and ( n4079 , n4076 , n4078 );
and ( n4080 , n4075 , n4078 );
or ( n4081 , n4077 , n4079 , n4080 );
and ( n4082 , n4074 , n4081 );
xor ( n4083 , n3955 , n3956 );
xor ( n4084 , n3765 , n3766 );
and ( n4085 , n4083 , n4084 );
xor ( n4086 , n4042 , n4043 );
and ( n4087 , n4085 , n4086 );
xor ( n4088 , n4045 , n4046 );
xor ( n4089 , n4088 , n4048 );
and ( n4090 , n4086 , n4089 );
and ( n4091 , n4085 , n4089 );
or ( n4092 , n4087 , n4090 , n4091 );
and ( n4093 , n4081 , n4092 );
and ( n4094 , n4074 , n4092 );
or ( n4095 , n4082 , n4093 , n4094 );
and ( n4096 , n4072 , n4095 );
xor ( n4097 , n4041 , n4056 );
xor ( n4098 , n4097 , n4059 );
and ( n4099 , n4095 , n4098 );
and ( n4100 , n4072 , n4098 );
or ( n4101 , n4096 , n4099 , n4100 );
and ( n4102 , n4070 , n4101 );
xor ( n4103 , n4031 , n4033 );
xor ( n4104 , n4103 , n4062 );
and ( n4105 , n4101 , n4104 );
and ( n4106 , n4070 , n4104 );
or ( n4107 , n4102 , n4105 , n4106 );
and ( n4108 , n4067 , n4107 );
and ( n4109 , n4065 , n4107 );
or ( n4110 , n4068 , n4108 , n4109 );
and ( n4111 , n4017 , n4110 );
xor ( n4112 , n3990 , n3992 );
xor ( n4113 , n4112 , n3995 );
and ( n4114 , n4110 , n4113 );
and ( n4115 , n4017 , n4113 );
or ( n4116 , n4111 , n4114 , n4115 );
and ( n4117 , n4014 , n4116 );
and ( n4118 , n4013 , n4116 );
or ( n4119 , n4015 , n4117 , n4118 );
xor ( n4120 , n3870 , n3872 );
xor ( n4121 , n4120 , n4001 );
and ( n4122 , n4119 , n4121 );
xor ( n4123 , n4119 , n4121 );
and ( n4124 , n3645 , n1465 );
and ( n4125 , n3169 , n1860 );
and ( n4126 , n4124 , n4125 );
and ( n4127 , n2286 , n3301 );
and ( n4128 , n4125 , n4127 );
and ( n4129 , n4124 , n4127 );
or ( n4130 , n4126 , n4128 , n4129 );
and ( n4131 , n1275 , n3903 );
and ( n4132 , n3892 , n1293 );
and ( n4133 , n4131 , n4132 );
buf ( n4134 , n771 );
buf ( n4135 , n4134 );
buf ( n4136 , n4135 );
buf ( n4137 , n4136 );
buf ( n4138 , n4137 );
and ( n4139 , n4138 , n1287 );
and ( n4140 , n4133 , n4139 );
and ( n4141 , n3833 , n1360 );
and ( n4142 , n4139 , n4141 );
and ( n4143 , n4133 , n4141 );
or ( n4144 , n4140 , n4142 , n4143 );
and ( n4145 , n4130 , n4144 );
buf ( n4146 , n771 );
buf ( n4147 , n4146 );
buf ( n4148 , n4147 );
buf ( n4149 , n4148 );
buf ( n4150 , n4149 );
not ( n4151 , n4150 );
and ( n4152 , n1279 , n4150 );
nor ( n4153 , n4151 , n4152 );
and ( n4154 , n2591 , n1689 );
and ( n4155 , n4153 , n4154 );
and ( n4156 , n2255 , n1906 );
and ( n4157 , n4154 , n4156 );
and ( n4158 , n4153 , n4156 );
or ( n4159 , n4155 , n4157 , n4158 );
buf ( n4160 , n4148 );
buf ( n4161 , n4160 );
and ( n4162 , n1291 , n4161 );
not ( n4163 , n4161 );
nor ( n4164 , n4162 , n4163 );
and ( n4165 , n1694 , n2586 );
and ( n4166 , n4164 , n4165 );
and ( n4167 , n1911 , n2250 );
and ( n4168 , n4165 , n4167 );
and ( n4169 , n4164 , n4167 );
or ( n4170 , n4166 , n4168 , n4169 );
and ( n4171 , n4159 , n4170 );
and ( n4172 , n4144 , n4171 );
and ( n4173 , n4130 , n4171 );
or ( n4174 , n4145 , n4172 , n4173 );
and ( n4175 , n1317 , n3739 );
and ( n4176 , n3728 , n1312 );
and ( n4177 , n4175 , n4176 );
and ( n4178 , n2634 , n2577 );
and ( n4179 , n4177 , n4178 );
and ( n4180 , n2267 , n3627 );
and ( n4181 , n4178 , n4180 );
and ( n4182 , n4177 , n4180 );
or ( n4183 , n4179 , n4181 , n4182 );
xor ( n4184 , n3895 , n3896 );
xor ( n4185 , n4184 , n3898 );
xor ( n4186 , n3906 , n3907 );
xor ( n4187 , n4186 , n3909 );
and ( n4188 , n4185 , n4187 );
and ( n4189 , n4183 , n4188 );
xor ( n4190 , n3874 , n3875 );
xor ( n4191 , n4190 , n3877 );
and ( n4192 , n4188 , n4191 );
and ( n4193 , n4183 , n4191 );
or ( n4194 , n4189 , n4192 , n4193 );
and ( n4195 , n4174 , n4194 );
xor ( n4196 , n3764 , n3773 );
xor ( n4197 , n4196 , n3789 );
and ( n4198 , n4194 , n4197 );
and ( n4199 , n4174 , n4197 );
or ( n4200 , n4195 , n4198 , n4199 );
xor ( n4201 , n3838 , n3840 );
xor ( n4202 , n4201 , n3843 );
and ( n4203 , n4200 , n4202 );
xor ( n4204 , n3916 , n3918 );
xor ( n4205 , n4204 , n3921 );
and ( n4206 , n4202 , n4205 );
and ( n4207 , n4200 , n4205 );
or ( n4208 , n4203 , n4206 , n4207 );
xor ( n4209 , n3755 , n3757 );
xor ( n4210 , n4209 , n3760 );
and ( n4211 , n4208 , n4210 );
xor ( n4212 , n3819 , n3846 );
xor ( n4213 , n4212 , n3849 );
and ( n4214 , n4210 , n4213 );
and ( n4215 , n4208 , n4213 );
or ( n4216 , n4211 , n4214 , n4215 );
xor ( n4217 , n3952 , n3953 );
and ( n4218 , n1353 , n3449 );
and ( n4219 , n3454 , n1348 );
and ( n4220 , n4218 , n4219 );
and ( n4221 , n4217 , n4220 );
and ( n4222 , n1724 , n2492 );
and ( n4223 , n2497 , n1719 );
and ( n4224 , n4222 , n4223 );
and ( n4225 , n4220 , n4224 );
and ( n4226 , n4217 , n4224 );
or ( n4227 , n4221 , n4225 , n4226 );
xor ( n4228 , n3767 , n3768 );
xor ( n4229 , n4228 , n3770 );
and ( n4230 , n4227 , n4229 );
xor ( n4231 , n3954 , n3957 );
xor ( n4232 , n4231 , n3959 );
and ( n4233 , n4229 , n4232 );
and ( n4234 , n4227 , n4232 );
or ( n4235 , n4230 , n4233 , n4234 );
xor ( n4236 , n3775 , n3776 );
xor ( n4237 , n4236 , n3778 );
xor ( n4238 , n3782 , n3783 );
xor ( n4239 , n4238 , n3785 );
and ( n4240 , n4237 , n4239 );
xor ( n4241 , n3881 , n3882 );
xor ( n4242 , n4241 , n3884 );
and ( n4243 , n4240 , n4242 );
xor ( n4244 , n3821 , n3822 );
xor ( n4245 , n4244 , n3824 );
and ( n4246 , n4242 , n4245 );
and ( n4247 , n4240 , n4245 );
or ( n4248 , n4243 , n4246 , n4247 );
and ( n4249 , n4235 , n4248 );
xor ( n4250 , n3880 , n3887 );
xor ( n4251 , n4250 , n3913 );
and ( n4252 , n4248 , n4251 );
and ( n4253 , n4235 , n4251 );
or ( n4254 , n4249 , n4252 , n4253 );
xor ( n4255 , n3792 , n3802 );
xor ( n4256 , n4255 , n3816 );
and ( n4257 , n4254 , n4256 );
xor ( n4258 , n3968 , n3970 );
xor ( n4259 , n4258 , n3973 );
and ( n4260 , n4256 , n4259 );
and ( n4261 , n4254 , n4259 );
or ( n4262 , n4257 , n4260 , n4261 );
and ( n4263 , n1911 , n2304 );
and ( n4264 , n2309 , n1906 );
and ( n4265 , n4263 , n4264 );
and ( n4266 , n3169 , n2040 );
and ( n4267 , n4265 , n4266 );
and ( n4268 , n2286 , n3627 );
and ( n4269 , n4266 , n4268 );
and ( n4270 , n4265 , n4268 );
or ( n4271 , n4267 , n4269 , n4270 );
and ( n4272 , n1694 , n2718 );
and ( n4273 , n2723 , n1689 );
and ( n4274 , n4272 , n4273 );
and ( n4275 , n3833 , n1465 );
and ( n4276 , n4274 , n4275 );
and ( n4277 , n2267 , n3929 );
and ( n4278 , n4275 , n4277 );
and ( n4279 , n4274 , n4277 );
or ( n4280 , n4276 , n4278 , n4279 );
and ( n4281 , n4271 , n4280 );
and ( n4282 , n1778 , n2492 );
and ( n4283 , n2497 , n1789 );
and ( n4284 , n4282 , n4283 );
and ( n4285 , n3246 , n1860 );
and ( n4286 , n4284 , n4285 );
and ( n4287 , n2634 , n2948 );
and ( n4288 , n4285 , n4287 );
and ( n4289 , n4284 , n4287 );
or ( n4290 , n4286 , n4288 , n4289 );
and ( n4291 , n4280 , n4290 );
and ( n4292 , n4271 , n4290 );
or ( n4293 , n4281 , n4291 , n4292 );
and ( n4294 , n4138 , n1360 );
and ( n4295 , n3339 , n1711 );
and ( n4296 , n4294 , n4295 );
and ( n4297 , n2764 , n2577 );
and ( n4298 , n4295 , n4297 );
and ( n4299 , n4294 , n4297 );
or ( n4300 , n4296 , n4298 , n4299 );
and ( n4301 , n1275 , n4161 );
buf ( n4302 , n4301 );
buf ( n4303 , n4302 );
and ( n4304 , n4300 , n4303 );
and ( n4305 , n3892 , n1312 );
and ( n4306 , n3728 , n1348 );
and ( n4307 , n4305 , n4306 );
and ( n4308 , n2591 , n1719 );
and ( n4309 , n4306 , n4308 );
and ( n4310 , n4305 , n4308 );
or ( n4311 , n4307 , n4309 , n4310 );
and ( n4312 , n1317 , n3903 );
and ( n4313 , n1353 , n3739 );
and ( n4314 , n4312 , n4313 );
and ( n4315 , n1724 , n2586 );
and ( n4316 , n4313 , n4315 );
and ( n4317 , n4312 , n4315 );
or ( n4318 , n4314 , n4316 , n4317 );
and ( n4319 , n4311 , n4318 );
and ( n4320 , n4303 , n4319 );
and ( n4321 , n4300 , n4319 );
or ( n4322 , n4304 , n4320 , n4321 );
and ( n4323 , n4293 , n4322 );
xor ( n4324 , n4153 , n4154 );
xor ( n4325 , n4324 , n4156 );
xor ( n4326 , n4164 , n4165 );
xor ( n4327 , n4326 , n4167 );
and ( n4328 , n4325 , n4327 );
xor ( n4329 , n3936 , n3937 );
xor ( n4330 , n4329 , n3939 );
and ( n4331 , n4328 , n4330 );
xor ( n4332 , n4133 , n4139 );
xor ( n4333 , n4332 , n4141 );
and ( n4334 , n4330 , n4333 );
and ( n4335 , n4328 , n4333 );
or ( n4336 , n4331 , n4334 , n4335 );
and ( n4337 , n4322 , n4336 );
and ( n4338 , n4293 , n4336 );
or ( n4339 , n4323 , n4337 , n4338 );
xnor ( n4340 , n3946 , n3947 );
xor ( n4341 , n4124 , n4125 );
xor ( n4342 , n4341 , n4127 );
and ( n4343 , n4340 , n4342 );
xor ( n4344 , n4217 , n4220 );
xor ( n4345 , n4344 , n4224 );
and ( n4346 , n4342 , n4345 );
and ( n4347 , n4340 , n4345 );
or ( n4348 , n4343 , n4346 , n4347 );
xor ( n4349 , n4130 , n4144 );
xor ( n4350 , n4349 , n4171 );
and ( n4351 , n4348 , n4350 );
xor ( n4352 , n3933 , n3942 );
xor ( n4353 , n4352 , n3948 );
and ( n4354 , n4350 , n4353 );
and ( n4355 , n4348 , n4353 );
or ( n4356 , n4351 , n4354 , n4355 );
and ( n4357 , n4339 , n4356 );
buf ( n4358 , n772 );
buf ( n4359 , n4358 );
buf ( n4360 , n4359 );
buf ( n4361 , n4360 );
buf ( n4362 , n4361 );
and ( n4363 , n1291 , n4362 );
not ( n4364 , n4362 );
nor ( n4365 , n4363 , n4364 );
buf ( n4366 , n4360 );
buf ( n4367 , n4366 );
not ( n4368 , n4367 );
and ( n4369 , n1279 , n4367 );
nor ( n4370 , n4368 , n4369 );
and ( n4371 , n4365 , n4370 );
and ( n4372 , n3645 , n1530 );
and ( n4373 , n4371 , n4372 );
and ( n4374 , n2477 , n3301 );
and ( n4375 , n4372 , n4374 );
and ( n4376 , n4371 , n4374 );
or ( n4377 , n4373 , n4375 , n4376 );
and ( n4378 , n1995 , n2250 );
and ( n4379 , n2255 , n1990 );
and ( n4380 , n4378 , n4379 );
buf ( n4381 , n772 );
buf ( n4382 , n4381 );
buf ( n4383 , n4382 );
buf ( n4384 , n4383 );
buf ( n4385 , n4384 );
and ( n4386 , n4385 , n1287 );
and ( n4387 , n4380 , n4386 );
and ( n4388 , n2937 , n2407 );
and ( n4389 , n4386 , n4388 );
and ( n4390 , n4380 , n4388 );
or ( n4391 , n4387 , n4389 , n4390 );
and ( n4392 , n4377 , n4391 );
xor ( n4393 , n4177 , n4178 );
xor ( n4394 , n4393 , n4180 );
and ( n4395 , n4391 , n4394 );
and ( n4396 , n4377 , n4394 );
or ( n4397 , n4392 , n4395 , n4396 );
xor ( n4398 , n4227 , n4229 );
xor ( n4399 , n4398 , n4232 );
and ( n4400 , n4397 , n4399 );
xor ( n4401 , n4240 , n4242 );
xor ( n4402 , n4401 , n4245 );
and ( n4403 , n4399 , n4402 );
and ( n4404 , n4397 , n4402 );
or ( n4405 , n4400 , n4403 , n4404 );
and ( n4406 , n4356 , n4405 );
and ( n4407 , n4339 , n4405 );
or ( n4408 , n4357 , n4406 , n4407 );
xor ( n4409 , n3794 , n3796 );
xor ( n4410 , n4409 , n3799 );
xor ( n4411 , n3808 , n3810 );
xor ( n4412 , n4411 , n3813 );
and ( n4413 , n4410 , n4412 );
xor ( n4414 , n3951 , n3962 );
xor ( n4415 , n4414 , n3965 );
and ( n4416 , n4412 , n4415 );
and ( n4417 , n4410 , n4415 );
or ( n4418 , n4413 , n4416 , n4417 );
and ( n4419 , n4408 , n4418 );
xor ( n4420 , n4200 , n4202 );
xor ( n4421 , n4420 , n4205 );
and ( n4422 , n4418 , n4421 );
and ( n4423 , n4408 , n4421 );
or ( n4424 , n4419 , n4422 , n4423 );
and ( n4425 , n4262 , n4424 );
xor ( n4426 , n3924 , n3976 );
xor ( n4427 , n4426 , n3979 );
and ( n4428 , n4424 , n4427 );
and ( n4429 , n4262 , n4427 );
or ( n4430 , n4425 , n4428 , n4429 );
and ( n4431 , n4216 , n4430 );
xor ( n4432 , n3982 , n3984 );
xor ( n4433 , n4432 , n3987 );
and ( n4434 , n4430 , n4433 );
and ( n4435 , n4216 , n4433 );
or ( n4436 , n4431 , n4434 , n4435 );
xor ( n4437 , n4065 , n4067 );
xor ( n4438 , n4437 , n4107 );
xor ( n4439 , n4216 , n4430 );
xor ( n4440 , n4439 , n4433 );
and ( n4441 , n4438 , n4440 );
xor ( n4442 , n4208 , n4210 );
xor ( n4443 , n4442 , n4213 );
xor ( n4444 , n4262 , n4424 );
xor ( n4445 , n4444 , n4427 );
and ( n4446 , n4443 , n4445 );
and ( n4447 , n4440 , n4446 );
and ( n4448 , n4438 , n4446 );
or ( n4449 , n4441 , n4447 , n4448 );
and ( n4450 , n4436 , n4449 );
xor ( n4451 , n4017 , n4110 );
xor ( n4452 , n4451 , n4113 );
and ( n4453 , n4449 , n4452 );
and ( n4454 , n4436 , n4452 );
or ( n4455 , n4450 , n4453 , n4454 );
xor ( n4456 , n4013 , n4014 );
xor ( n4457 , n4456 , n4116 );
and ( n4458 , n4455 , n4457 );
xor ( n4459 , n4455 , n4457 );
xor ( n4460 , n4070 , n4101 );
xor ( n4461 , n4460 , n4104 );
xor ( n4462 , n4035 , n4036 );
xor ( n4463 , n4462 , n4038 );
xor ( n4464 , n4044 , n4051 );
xor ( n4465 , n4464 , n4053 );
and ( n4466 , n4463 , n4465 );
xor ( n4467 , n4159 , n4170 );
xor ( n4468 , n4185 , n4187 );
and ( n4469 , n4467 , n4468 );
xor ( n4470 , n4237 , n4239 );
and ( n4471 , n4468 , n4470 );
and ( n4472 , n4467 , n4470 );
or ( n4473 , n4469 , n4471 , n4472 );
xor ( n4474 , n4294 , n4295 );
xor ( n4475 , n4474 , n4297 );
xor ( n4476 , n4131 , n4132 );
and ( n4477 , n4475 , n4476 );
xor ( n4478 , n4175 , n4176 );
xor ( n4479 , n4218 , n4219 );
and ( n4480 , n4478 , n4479 );
xor ( n4481 , n4222 , n4223 );
and ( n4482 , n4479 , n4481 );
and ( n4483 , n4478 , n4481 );
or ( n4484 , n4480 , n4482 , n4483 );
and ( n4485 , n4477 , n4484 );
xor ( n4486 , n3934 , n3935 );
xor ( n4487 , n3944 , n3945 );
and ( n4488 , n4486 , n4487 );
and ( n4489 , n4150 , n1293 );
and ( n4490 , n3169 , n2407 );
and ( n4491 , n4489 , n4490 );
and ( n4492 , n4487 , n4491 );
and ( n4493 , n4486 , n4491 );
or ( n4494 , n4488 , n4492 , n4493 );
and ( n4495 , n4484 , n4494 );
and ( n4496 , n4477 , n4494 );
or ( n4497 , n4485 , n4495 , n4496 );
and ( n4498 , n4473 , n4497 );
xor ( n4499 , n4075 , n4076 );
xor ( n4500 , n4499 , n4078 );
and ( n4501 , n4497 , n4500 );
and ( n4502 , n4473 , n4500 );
or ( n4503 , n4498 , n4501 , n4502 );
and ( n4504 , n4465 , n4503 );
and ( n4505 , n4463 , n4503 );
or ( n4506 , n4466 , n4504 , n4505 );
xor ( n4507 , n4072 , n4095 );
xor ( n4508 , n4507 , n4098 );
and ( n4509 , n4506 , n4508 );
xor ( n4510 , n4254 , n4256 );
xor ( n4511 , n4510 , n4259 );
and ( n4512 , n4508 , n4511 );
and ( n4513 , n4506 , n4511 );
or ( n4514 , n4509 , n4512 , n4513 );
and ( n4515 , n4461 , n4514 );
and ( n4516 , n1995 , n2304 );
and ( n4517 , n2309 , n1990 );
and ( n4518 , n4516 , n4517 );
and ( n4519 , n2937 , n2577 );
and ( n4520 , n4518 , n4519 );
buf ( n4521 , n2033 );
buf ( n4522 , n4521 );
and ( n4523 , n2267 , n4522 );
and ( n4524 , n4519 , n4523 );
and ( n4525 , n4518 , n4523 );
or ( n4526 , n4520 , n4524 , n4525 );
and ( n4527 , n1353 , n3903 );
and ( n4528 , n3892 , n1348 );
and ( n4529 , n4527 , n4528 );
and ( n4530 , n4385 , n1360 );
and ( n4531 , n4529 , n4530 );
and ( n4532 , n3339 , n1860 );
and ( n4533 , n4530 , n4532 );
and ( n4534 , n4529 , n4532 );
or ( n4535 , n4531 , n4533 , n4534 );
and ( n4536 , n4526 , n4535 );
and ( n4537 , n1778 , n2586 );
and ( n4538 , n2591 , n1789 );
and ( n4539 , n4537 , n4538 );
and ( n4540 , n4138 , n1465 );
and ( n4541 , n4539 , n4540 );
and ( n4542 , n2286 , n3929 );
and ( n4543 , n4540 , n4542 );
and ( n4544 , n4539 , n4542 );
or ( n4545 , n4541 , n4543 , n4544 );
and ( n4546 , n4535 , n4545 );
and ( n4547 , n4526 , n4545 );
or ( n4548 , n4536 , n4546 , n4547 );
and ( n4549 , n2048 , n2250 );
and ( n4550 , n2255 , n2059 );
and ( n4551 , n4549 , n4550 );
and ( n4552 , n3833 , n1530 );
and ( n4553 , n4551 , n4552 );
and ( n4554 , n2764 , n2948 );
and ( n4555 , n4552 , n4554 );
and ( n4556 , n4551 , n4554 );
or ( n4557 , n4553 , n4555 , n4556 );
buf ( n4558 , n2048 );
buf ( n4559 , n2035 );
and ( n4560 , n4558 , n4559 );
and ( n4561 , n4557 , n4560 );
not ( n4562 , n4302 );
and ( n4563 , n4560 , n4562 );
and ( n4564 , n4557 , n4562 );
or ( n4565 , n4561 , n4563 , n4564 );
and ( n4566 , n4548 , n4565 );
xor ( n4567 , n3925 , n3926 );
xor ( n4568 , n4567 , n3930 );
and ( n4569 , n4565 , n4568 );
and ( n4570 , n4548 , n4568 );
or ( n4571 , n4566 , n4569 , n4570 );
and ( n4572 , n1275 , n4362 );
and ( n4573 , n4367 , n1293 );
and ( n4574 , n4572 , n4573 );
buf ( n4575 , n773 );
buf ( n4576 , n4575 );
buf ( n4577 , n4576 );
buf ( n4578 , n4577 );
buf ( n4579 , n4578 );
and ( n4580 , n4579 , n1287 );
and ( n4581 , n4574 , n4580 );
and ( n4582 , n3645 , n1711 );
and ( n4583 , n4580 , n4582 );
and ( n4584 , n4574 , n4582 );
or ( n4585 , n4581 , n4583 , n4584 );
and ( n4586 , n1694 , n2923 );
and ( n4587 , n2928 , n1689 );
and ( n4588 , n4586 , n4587 );
and ( n4589 , n1911 , n2492 );
and ( n4590 , n2497 , n1906 );
and ( n4591 , n4589 , n4590 );
and ( n4592 , n4588 , n4591 );
and ( n4593 , n2634 , n3301 );
and ( n4594 , n4591 , n4593 );
and ( n4595 , n4588 , n4593 );
or ( n4596 , n4592 , n4594 , n4595 );
and ( n4597 , n4585 , n4596 );
and ( n4598 , n1317 , n4161 );
and ( n4599 , n4150 , n1312 );
and ( n4600 , n4598 , n4599 );
and ( n4601 , n3246 , n2040 );
and ( n4602 , n4600 , n4601 );
and ( n4603 , n2477 , n3627 );
and ( n4604 , n4601 , n4603 );
and ( n4605 , n4600 , n4603 );
or ( n4606 , n4602 , n4604 , n4605 );
and ( n4607 , n4596 , n4606 );
and ( n4608 , n4585 , n4606 );
or ( n4609 , n4597 , n4607 , n4608 );
xor ( n4610 , n4271 , n4280 );
xor ( n4611 , n4610 , n4290 );
and ( n4612 , n4609 , n4611 );
xor ( n4613 , n4377 , n4391 );
xor ( n4614 , n4613 , n4394 );
and ( n4615 , n4611 , n4614 );
and ( n4616 , n4609 , n4614 );
or ( n4617 , n4612 , n4615 , n4616 );
and ( n4618 , n4571 , n4617 );
xor ( n4619 , n4183 , n4188 );
xor ( n4620 , n4619 , n4191 );
and ( n4621 , n4617 , n4620 );
and ( n4622 , n4571 , n4620 );
or ( n4623 , n4618 , n4621 , n4622 );
xor ( n4624 , n4174 , n4194 );
xor ( n4625 , n4624 , n4197 );
and ( n4626 , n4623 , n4625 );
xor ( n4627 , n4235 , n4248 );
xor ( n4628 , n4627 , n4251 );
and ( n4629 , n4625 , n4628 );
and ( n4630 , n4623 , n4628 );
or ( n4631 , n4626 , n4629 , n4630 );
xor ( n4632 , n4074 , n4081 );
xor ( n4633 , n4632 , n4092 );
xor ( n4634 , n4410 , n4412 );
xor ( n4635 , n4634 , n4415 );
and ( n4636 , n4633 , n4635 );
xor ( n4637 , n4085 , n4086 );
xor ( n4638 , n4637 , n4089 );
xor ( n4639 , n4348 , n4350 );
xor ( n4640 , n4639 , n4353 );
and ( n4641 , n4638 , n4640 );
xor ( n4642 , n4397 , n4399 );
xor ( n4643 , n4642 , n4402 );
and ( n4644 , n4640 , n4643 );
and ( n4645 , n4638 , n4643 );
or ( n4646 , n4641 , n4644 , n4645 );
and ( n4647 , n4635 , n4646 );
and ( n4648 , n4633 , n4646 );
or ( n4649 , n4636 , n4647 , n4648 );
and ( n4650 , n4631 , n4649 );
xor ( n4651 , n4408 , n4418 );
xor ( n4652 , n4651 , n4421 );
and ( n4653 , n4649 , n4652 );
and ( n4654 , n4631 , n4652 );
or ( n4655 , n4650 , n4653 , n4654 );
and ( n4656 , n4514 , n4655 );
and ( n4657 , n4461 , n4655 );
or ( n4658 , n4515 , n4656 , n4657 );
xor ( n4659 , n4083 , n4084 );
xor ( n4660 , n4328 , n4330 );
xor ( n4661 , n4660 , n4333 );
and ( n4662 , n4659 , n4661 );
xor ( n4663 , n4340 , n4342 );
xor ( n4664 , n4663 , n4345 );
and ( n4665 , n4661 , n4664 );
and ( n4666 , n4659 , n4664 );
or ( n4667 , n4662 , n4665 , n4666 );
xor ( n4668 , n4284 , n4285 );
xor ( n4669 , n4668 , n4287 );
xor ( n4670 , n4371 , n4372 );
xor ( n4671 , n4670 , n4374 );
and ( n4672 , n4669 , n4671 );
xor ( n4673 , n4380 , n4386 );
xor ( n4674 , n4673 , n4388 );
and ( n4675 , n4671 , n4674 );
and ( n4676 , n4669 , n4674 );
or ( n4677 , n4672 , n4675 , n4676 );
xor ( n4678 , n4265 , n4266 );
xor ( n4679 , n4678 , n4268 );
xor ( n4680 , n4274 , n4275 );
xor ( n4681 , n4680 , n4277 );
and ( n4682 , n4679 , n4681 );
xor ( n4683 , n4311 , n4318 );
and ( n4684 , n4681 , n4683 );
and ( n4685 , n4679 , n4683 );
or ( n4686 , n4682 , n4684 , n4685 );
and ( n4687 , n4677 , n4686 );
xor ( n4688 , n4325 , n4327 );
xor ( n4689 , n4305 , n4306 );
xor ( n4690 , n4689 , n4308 );
xor ( n4691 , n4312 , n4313 );
xor ( n4692 , n4691 , n4315 );
and ( n4693 , n4690 , n4692 );
and ( n4694 , n4688 , n4693 );
xor ( n4695 , n4558 , n4559 );
not ( n4696 , n4301 );
and ( n4697 , n4695 , n4696 );
xor ( n4698 , n4365 , n4370 );
and ( n4699 , n4696 , n4698 );
and ( n4700 , n4695 , n4698 );
or ( n4701 , n4697 , n4699 , n4700 );
and ( n4702 , n4693 , n4701 );
and ( n4703 , n4688 , n4701 );
or ( n4704 , n4694 , n4702 , n4703 );
and ( n4705 , n4686 , n4704 );
and ( n4706 , n4677 , n4704 );
or ( n4707 , n4687 , n4705 , n4706 );
and ( n4708 , n4667 , n4707 );
xor ( n4709 , n4272 , n4273 );
xor ( n4710 , n4282 , n4283 );
and ( n4711 , n4709 , n4710 );
xor ( n4712 , n4263 , n4264 );
and ( n4713 , n4710 , n4712 );
and ( n4714 , n4709 , n4712 );
or ( n4715 , n4711 , n4713 , n4714 );
xor ( n4716 , n4378 , n4379 );
buf ( n4717 , n774 );
buf ( n4718 , n4717 );
buf ( n4719 , n4718 );
buf ( n4720 , n4719 );
buf ( n4721 , n4720 );
and ( n4722 , n4721 , n1287 );
and ( n4723 , n2477 , n3929 );
and ( n4724 , n4722 , n4723 );
and ( n4725 , n2286 , n4522 );
and ( n4726 , n4723 , n4725 );
and ( n4727 , n4722 , n4725 );
or ( n4728 , n4724 , n4726 , n4727 );
and ( n4729 , n4716 , n4728 );
buf ( n4730 , n773 );
buf ( n4731 , n4730 );
buf ( n4732 , n4731 );
buf ( n4733 , n4732 );
buf ( n4734 , n4733 );
and ( n4735 , n1291 , n4734 );
not ( n4736 , n4734 );
nor ( n4737 , n4735 , n4736 );
buf ( n4738 , n4732 );
buf ( n4739 , n4738 );
not ( n4740 , n4739 );
and ( n4741 , n1279 , n4739 );
nor ( n4742 , n4740 , n4741 );
and ( n4743 , n4737 , n4742 );
and ( n4744 , n4728 , n4743 );
and ( n4745 , n4716 , n4743 );
or ( n4746 , n4729 , n4744 , n4745 );
and ( n4747 , n4715 , n4746 );
xor ( n4748 , n4475 , n4476 );
and ( n4749 , n4746 , n4748 );
and ( n4750 , n4715 , n4748 );
or ( n4751 , n4747 , n4749 , n4750 );
xor ( n4752 , n4467 , n4468 );
xor ( n4753 , n4752 , n4470 );
and ( n4754 , n4751 , n4753 );
xor ( n4755 , n4477 , n4484 );
xor ( n4756 , n4755 , n4494 );
and ( n4757 , n4753 , n4756 );
and ( n4758 , n4751 , n4756 );
or ( n4759 , n4754 , n4757 , n4758 );
and ( n4760 , n4707 , n4759 );
and ( n4761 , n4667 , n4759 );
or ( n4762 , n4708 , n4760 , n4761 );
xor ( n4763 , n4463 , n4465 );
xor ( n4764 , n4763 , n4503 );
and ( n4765 , n4762 , n4764 );
xor ( n4766 , n4339 , n4356 );
xor ( n4767 , n4766 , n4405 );
and ( n4768 , n4764 , n4767 );
and ( n4769 , n4762 , n4767 );
or ( n4770 , n4765 , n4768 , n4769 );
xor ( n4771 , n4623 , n4625 );
xor ( n4772 , n4771 , n4628 );
xor ( n4773 , n4473 , n4497 );
xor ( n4774 , n4773 , n4500 );
xor ( n4775 , n4293 , n4322 );
xor ( n4776 , n4775 , n4336 );
and ( n4777 , n4774 , n4776 );
xor ( n4778 , n4571 , n4617 );
xor ( n4779 , n4778 , n4620 );
and ( n4780 , n4776 , n4779 );
and ( n4781 , n4774 , n4779 );
or ( n4782 , n4777 , n4780 , n4781 );
and ( n4783 , n4772 , n4782 );
xor ( n4784 , n4300 , n4303 );
xor ( n4785 , n4784 , n4319 );
xor ( n4786 , n4548 , n4565 );
xor ( n4787 , n4786 , n4568 );
and ( n4788 , n4785 , n4787 );
xor ( n4789 , n4609 , n4611 );
xor ( n4790 , n4789 , n4614 );
and ( n4791 , n4787 , n4790 );
and ( n4792 , n4785 , n4790 );
or ( n4793 , n4788 , n4791 , n4792 );
xor ( n4794 , n4478 , n4479 );
xor ( n4795 , n4794 , n4481 );
xor ( n4796 , n4486 , n4487 );
xor ( n4797 , n4796 , n4491 );
and ( n4798 , n4795 , n4797 );
xor ( n4799 , n4585 , n4596 );
xor ( n4800 , n4799 , n4606 );
and ( n4801 , n4797 , n4800 );
and ( n4802 , n4795 , n4800 );
or ( n4803 , n4798 , n4801 , n4802 );
xor ( n4804 , n4526 , n4535 );
xor ( n4805 , n4804 , n4545 );
xor ( n4806 , n4557 , n4560 );
xor ( n4807 , n4806 , n4562 );
and ( n4808 , n4805 , n4807 );
xor ( n4809 , n4669 , n4671 );
xor ( n4810 , n4809 , n4674 );
and ( n4811 , n4807 , n4810 );
and ( n4812 , n4805 , n4810 );
or ( n4813 , n4808 , n4811 , n4812 );
and ( n4814 , n4803 , n4813 );
and ( n4815 , n4138 , n1530 );
and ( n4816 , n3246 , n2407 );
and ( n4817 , n4815 , n4816 );
and ( n4818 , n2634 , n3627 );
and ( n4819 , n4816 , n4818 );
and ( n4820 , n4815 , n4818 );
or ( n4821 , n4817 , n4819 , n4820 );
and ( n4822 , n1778 , n2718 );
and ( n4823 , n2723 , n1789 );
and ( n4824 , n4822 , n4823 );
and ( n4825 , n3833 , n1711 );
and ( n4826 , n4824 , n4825 );
and ( n4827 , n3169 , n2577 );
and ( n4828 , n4825 , n4827 );
and ( n4829 , n4824 , n4827 );
or ( n4830 , n4826 , n4828 , n4829 );
and ( n4831 , n4821 , n4830 );
and ( n4832 , n1694 , n3146 );
and ( n4833 , n3151 , n1689 );
and ( n4834 , n4832 , n4833 );
and ( n4835 , n4579 , n1360 );
and ( n4836 , n4834 , n4835 );
and ( n4837 , n2937 , n2948 );
and ( n4838 , n4835 , n4837 );
and ( n4839 , n4834 , n4837 );
or ( n4840 , n4836 , n4838 , n4839 );
and ( n4841 , n4830 , n4840 );
and ( n4842 , n4821 , n4840 );
or ( n4843 , n4831 , n4841 , n4842 );
xor ( n4844 , n4518 , n4519 );
xor ( n4845 , n4844 , n4523 );
xor ( n4846 , n4529 , n4530 );
xor ( n4847 , n4846 , n4532 );
and ( n4848 , n4845 , n4847 );
xor ( n4849 , n4539 , n4540 );
xor ( n4850 , n4849 , n4542 );
and ( n4851 , n4847 , n4850 );
and ( n4852 , n4845 , n4850 );
or ( n4853 , n4848 , n4851 , n4852 );
and ( n4854 , n4843 , n4853 );
xor ( n4855 , n4574 , n4580 );
xor ( n4856 , n4855 , n4582 );
xor ( n4857 , n4588 , n4591 );
xor ( n4858 , n4857 , n4593 );
and ( n4859 , n4856 , n4858 );
xor ( n4860 , n4551 , n4552 );
xor ( n4861 , n4860 , n4554 );
and ( n4862 , n4858 , n4861 );
and ( n4863 , n4856 , n4861 );
or ( n4864 , n4859 , n4862 , n4863 );
and ( n4865 , n4853 , n4864 );
and ( n4866 , n4843 , n4864 );
or ( n4867 , n4854 , n4865 , n4866 );
and ( n4868 , n4813 , n4867 );
and ( n4869 , n4803 , n4867 );
or ( n4870 , n4814 , n4868 , n4869 );
and ( n4871 , n4793 , n4870 );
and ( n4872 , n2723 , n1719 );
and ( n4873 , n4385 , n1465 );
and ( n4874 , n4872 , n4873 );
xor ( n4875 , n4489 , n4490 );
and ( n4876 , n4874 , n4875 );
xor ( n4877 , n4600 , n4601 );
xor ( n4878 , n4877 , n4603 );
and ( n4879 , n4875 , n4878 );
and ( n4880 , n4874 , n4878 );
or ( n4881 , n4876 , n4879 , n4880 );
xor ( n4882 , n4690 , n4692 );
buf ( n4883 , n2255 );
buf ( n4884 , n2267 );
and ( n4885 , n4883 , n4884 );
and ( n4886 , n1353 , n4161 );
and ( n4887 , n4150 , n1348 );
and ( n4888 , n4886 , n4887 );
and ( n4889 , n4885 , n4888 );
and ( n4890 , n1724 , n2923 );
and ( n4891 , n2928 , n1719 );
and ( n4892 , n4890 , n4891 );
and ( n4893 , n4888 , n4892 );
and ( n4894 , n4885 , n4892 );
or ( n4895 , n4889 , n4893 , n4894 );
and ( n4896 , n4882 , n4895 );
and ( n4897 , n1911 , n2586 );
and ( n4898 , n2591 , n1906 );
and ( n4899 , n4897 , n4898 );
and ( n4900 , n3645 , n1860 );
and ( n4901 , n4899 , n4900 );
and ( n4902 , n2764 , n3301 );
and ( n4903 , n4900 , n4902 );
and ( n4904 , n4899 , n4902 );
or ( n4905 , n4901 , n4903 , n4904 );
and ( n4906 , n4895 , n4905 );
and ( n4907 , n4882 , n4905 );
or ( n4908 , n4896 , n4906 , n4907 );
and ( n4909 , n4881 , n4908 );
and ( n4910 , n1995 , n2492 );
and ( n4911 , n2497 , n1990 );
and ( n4912 , n4910 , n4911 );
and ( n4913 , n2048 , n2304 );
and ( n4914 , n2309 , n2059 );
and ( n4915 , n4913 , n4914 );
and ( n4916 , n4912 , n4915 );
and ( n4917 , n3339 , n2040 );
and ( n4918 , n4915 , n4917 );
and ( n4919 , n4912 , n4917 );
or ( n4920 , n4916 , n4918 , n4919 );
and ( n4921 , n1275 , n4734 );
and ( n4922 , n4739 , n1293 );
and ( n4923 , n4921 , n4922 );
and ( n4924 , n1724 , n2718 );
or ( n4925 , n4923 , n4924 );
and ( n4926 , n4920 , n4925 );
xor ( n4927 , n4722 , n4723 );
xor ( n4928 , n4927 , n4725 );
xor ( n4929 , n4737 , n4742 );
and ( n4930 , n4928 , n4929 );
xor ( n4931 , n4572 , n4573 );
and ( n4932 , n4929 , n4931 );
and ( n4933 , n4928 , n4931 );
or ( n4934 , n4930 , n4932 , n4933 );
and ( n4935 , n4925 , n4934 );
and ( n4936 , n4920 , n4934 );
or ( n4937 , n4926 , n4935 , n4936 );
and ( n4938 , n4908 , n4937 );
and ( n4939 , n4881 , n4937 );
or ( n4940 , n4909 , n4938 , n4939 );
xor ( n4941 , n4598 , n4599 );
xor ( n4942 , n4527 , n4528 );
and ( n4943 , n4941 , n4942 );
xor ( n4944 , n4586 , n4587 );
and ( n4945 , n4942 , n4944 );
and ( n4946 , n4941 , n4944 );
or ( n4947 , n4943 , n4945 , n4946 );
xor ( n4948 , n4537 , n4538 );
xor ( n4949 , n4589 , n4590 );
and ( n4950 , n4948 , n4949 );
xor ( n4951 , n4516 , n4517 );
and ( n4952 , n4949 , n4951 );
and ( n4953 , n4948 , n4951 );
or ( n4954 , n4950 , n4952 , n4953 );
and ( n4955 , n4947 , n4954 );
xor ( n4956 , n4549 , n4550 );
and ( n4957 , n3833 , n1860 );
and ( n4958 , n3645 , n2040 );
and ( n4959 , n4957 , n4958 );
and ( n4960 , n3246 , n2577 );
and ( n4961 , n4958 , n4960 );
and ( n4962 , n4957 , n4960 );
or ( n4963 , n4959 , n4961 , n4962 );
and ( n4964 , n4956 , n4963 );
and ( n4965 , n4385 , n1530 );
and ( n4966 , n4138 , n1711 );
and ( n4967 , n4965 , n4966 );
and ( n4968 , n3339 , n2407 );
and ( n4969 , n4966 , n4968 );
and ( n4970 , n4965 , n4968 );
or ( n4971 , n4967 , n4969 , n4970 );
and ( n4972 , n4963 , n4971 );
and ( n4973 , n4956 , n4971 );
or ( n4974 , n4964 , n4972 , n4973 );
and ( n4975 , n4954 , n4974 );
and ( n4976 , n4947 , n4974 );
or ( n4977 , n4955 , n4975 , n4976 );
buf ( n4978 , n774 );
buf ( n4979 , n4978 );
buf ( n4980 , n4979 );
buf ( n4981 , n4980 );
buf ( n4982 , n4981 );
and ( n4983 , n1291 , n4982 );
not ( n4984 , n4982 );
nor ( n4985 , n4983 , n4984 );
and ( n4986 , n1317 , n4362 );
or ( n4987 , n4985 , n4986 );
buf ( n4988 , n4980 );
buf ( n4989 , n4988 );
not ( n4990 , n4989 );
and ( n4991 , n1279 , n4989 );
nor ( n4992 , n4990 , n4991 );
and ( n4993 , n4367 , n1312 );
and ( n4994 , n4992 , n4993 );
and ( n4995 , n4987 , n4994 );
xor ( n4996 , n4872 , n4873 );
and ( n4997 , n4994 , n4996 );
and ( n4998 , n4987 , n4996 );
or ( n4999 , n4995 , n4997 , n4998 );
xor ( n5000 , n4695 , n4696 );
xor ( n5001 , n5000 , n4698 );
and ( n5002 , n4999 , n5001 );
xor ( n5003 , n4709 , n4710 );
xor ( n5004 , n5003 , n4712 );
and ( n5005 , n5001 , n5004 );
and ( n5006 , n4999 , n5004 );
or ( n5007 , n5002 , n5005 , n5006 );
and ( n5008 , n4977 , n5007 );
xor ( n5009 , n4679 , n4681 );
xor ( n5010 , n5009 , n4683 );
and ( n5011 , n5007 , n5010 );
and ( n5012 , n4977 , n5010 );
or ( n5013 , n5008 , n5011 , n5012 );
and ( n5014 , n4940 , n5013 );
xor ( n5015 , n4659 , n4661 );
xor ( n5016 , n5015 , n4664 );
and ( n5017 , n5013 , n5016 );
and ( n5018 , n4940 , n5016 );
or ( n5019 , n5014 , n5017 , n5018 );
and ( n5020 , n4870 , n5019 );
and ( n5021 , n4793 , n5019 );
or ( n5022 , n4871 , n5020 , n5021 );
and ( n5023 , n4782 , n5022 );
and ( n5024 , n4772 , n5022 );
or ( n5025 , n4783 , n5023 , n5024 );
and ( n5026 , n4770 , n5025 );
xor ( n5027 , n4506 , n4508 );
xor ( n5028 , n5027 , n4511 );
and ( n5029 , n5025 , n5028 );
and ( n5030 , n4770 , n5028 );
or ( n5031 , n5026 , n5029 , n5030 );
xor ( n5032 , n4443 , n4445 );
and ( n5033 , n5031 , n5032 );
xor ( n5034 , n4633 , n4635 );
xor ( n5035 , n5034 , n4646 );
xor ( n5036 , n4638 , n4640 );
xor ( n5037 , n5036 , n4643 );
xor ( n5038 , n4667 , n4707 );
xor ( n5039 , n5038 , n4759 );
and ( n5040 , n5037 , n5039 );
xor ( n5041 , n4677 , n4686 );
xor ( n5042 , n5041 , n4704 );
xor ( n5043 , n4751 , n4753 );
xor ( n5044 , n5043 , n4756 );
and ( n5045 , n5042 , n5044 );
xor ( n5046 , n4688 , n4693 );
xor ( n5047 , n5046 , n4701 );
xor ( n5048 , n4715 , n4746 );
xor ( n5049 , n5048 , n4748 );
and ( n5050 , n5047 , n5049 );
xor ( n5051 , n4716 , n4728 );
xor ( n5052 , n5051 , n4743 );
xor ( n5053 , n4821 , n4830 );
xor ( n5054 , n5053 , n4840 );
and ( n5055 , n5052 , n5054 );
xor ( n5056 , n4845 , n4847 );
xor ( n5057 , n5056 , n4850 );
and ( n5058 , n5054 , n5057 );
and ( n5059 , n5052 , n5057 );
or ( n5060 , n5055 , n5058 , n5059 );
and ( n5061 , n5049 , n5060 );
and ( n5062 , n5047 , n5060 );
or ( n5063 , n5050 , n5061 , n5062 );
and ( n5064 , n5044 , n5063 );
and ( n5065 , n5042 , n5063 );
or ( n5066 , n5045 , n5064 , n5065 );
and ( n5067 , n5039 , n5066 );
and ( n5068 , n5037 , n5066 );
or ( n5069 , n5040 , n5067 , n5068 );
and ( n5070 , n5035 , n5069 );
xor ( n5071 , n4856 , n4858 );
xor ( n5072 , n5071 , n4861 );
and ( n5073 , n4721 , n1360 );
and ( n5074 , n2634 , n3929 );
and ( n5075 , n5073 , n5074 );
buf ( n5076 , n2265 );
buf ( n5077 , n5076 );
and ( n5078 , n2286 , n5077 );
and ( n5079 , n5074 , n5078 );
and ( n5080 , n5073 , n5078 );
or ( n5081 , n5075 , n5079 , n5080 );
buf ( n5082 , n775 );
buf ( n5083 , n5082 );
buf ( n5084 , n5083 );
buf ( n5085 , n5084 );
buf ( n5086 , n5085 );
and ( n5087 , n1291 , n5086 );
not ( n5088 , n5086 );
nor ( n5089 , n5087 , n5088 );
buf ( n5090 , n5084 );
buf ( n5091 , n5090 );
not ( n5092 , n5091 );
and ( n5093 , n1279 , n5091 );
nor ( n5094 , n5092 , n5093 );
and ( n5095 , n5089 , n5094 );
and ( n5096 , n1911 , n2718 );
and ( n5097 , n2723 , n1906 );
and ( n5098 , n5096 , n5097 );
and ( n5099 , n5095 , n5098 );
and ( n5100 , n4579 , n1465 );
and ( n5101 , n5098 , n5100 );
and ( n5102 , n5095 , n5100 );
or ( n5103 , n5099 , n5101 , n5102 );
and ( n5104 , n5081 , n5103 );
and ( n5105 , n1317 , n4734 );
and ( n5106 , n4739 , n1312 );
and ( n5107 , n5105 , n5106 );
and ( n5108 , n1778 , n2923 );
and ( n5109 , n2928 , n1789 );
and ( n5110 , n5108 , n5109 );
and ( n5111 , n5107 , n5110 );
and ( n5112 , n2477 , n4522 );
and ( n5113 , n5110 , n5112 );
and ( n5114 , n5107 , n5112 );
or ( n5115 , n5111 , n5113 , n5114 );
and ( n5116 , n5103 , n5115 );
and ( n5117 , n5081 , n5115 );
or ( n5118 , n5104 , n5116 , n5117 );
and ( n5119 , n5072 , n5118 );
and ( n5120 , n1694 , n3288 );
and ( n5121 , n3293 , n1689 );
and ( n5122 , n5120 , n5121 );
and ( n5123 , n3169 , n2948 );
and ( n5124 , n5122 , n5123 );
and ( n5125 , n2937 , n3301 );
and ( n5126 , n5123 , n5125 );
and ( n5127 , n5122 , n5125 );
or ( n5128 , n5124 , n5126 , n5127 );
xor ( n5129 , n4885 , n4888 );
xor ( n5130 , n5129 , n4892 );
and ( n5131 , n5128 , n5130 );
xor ( n5132 , n4815 , n4816 );
xor ( n5133 , n5132 , n4818 );
and ( n5134 , n5130 , n5133 );
and ( n5135 , n5128 , n5133 );
or ( n5136 , n5131 , n5134 , n5135 );
and ( n5137 , n5118 , n5136 );
and ( n5138 , n5072 , n5136 );
or ( n5139 , n5119 , n5137 , n5138 );
xor ( n5140 , n4899 , n4900 );
xor ( n5141 , n5140 , n4902 );
xor ( n5142 , n4912 , n4915 );
xor ( n5143 , n5142 , n4917 );
and ( n5144 , n5141 , n5143 );
xor ( n5145 , n4834 , n4835 );
xor ( n5146 , n5145 , n4837 );
and ( n5147 , n5143 , n5146 );
and ( n5148 , n5141 , n5146 );
or ( n5149 , n5144 , n5147 , n5148 );
xor ( n5150 , n4824 , n4825 );
xor ( n5151 , n5150 , n4827 );
xnor ( n5152 , n4923 , n4924 );
and ( n5153 , n5151 , n5152 );
and ( n5154 , n4367 , n1348 );
and ( n5155 , n3151 , n1719 );
and ( n5156 , n5154 , n5155 );
and ( n5157 , n2309 , n2250 );
and ( n5158 , n5155 , n5157 );
and ( n5159 , n5154 , n5157 );
or ( n5160 , n5156 , n5158 , n5159 );
and ( n5161 , n1353 , n4362 );
and ( n5162 , n1724 , n3146 );
and ( n5163 , n5161 , n5162 );
and ( n5164 , n2255 , n2304 );
and ( n5165 , n5162 , n5164 );
and ( n5166 , n5161 , n5164 );
or ( n5167 , n5163 , n5165 , n5166 );
and ( n5168 , n5160 , n5167 );
and ( n5169 , n5152 , n5168 );
and ( n5170 , n5151 , n5168 );
or ( n5171 , n5153 , n5169 , n5170 );
and ( n5172 , n5149 , n5171 );
buf ( n5173 , n775 );
buf ( n5174 , n5173 );
buf ( n5175 , n5174 );
buf ( n5176 , n5175 );
buf ( n5177 , n5176 );
and ( n5178 , n5177 , n1287 );
and ( n5179 , n2764 , n3627 );
and ( n5180 , n5178 , n5179 );
xor ( n5181 , n4957 , n4958 );
xor ( n5182 , n5181 , n4960 );
and ( n5183 , n5179 , n5182 );
and ( n5184 , n5178 , n5182 );
or ( n5185 , n5180 , n5183 , n5184 );
xor ( n5186 , n5073 , n5074 );
xor ( n5187 , n5186 , n5078 );
xnor ( n5188 , n4985 , n4986 );
and ( n5189 , n5187 , n5188 );
xor ( n5190 , n4883 , n4884 );
and ( n5191 , n5188 , n5190 );
and ( n5192 , n5187 , n5190 );
or ( n5193 , n5189 , n5191 , n5192 );
and ( n5194 , n5185 , n5193 );
xor ( n5195 , n4921 , n4922 );
xor ( n5196 , n4886 , n4887 );
and ( n5197 , n5195 , n5196 );
xor ( n5198 , n4832 , n4833 );
and ( n5199 , n5196 , n5198 );
and ( n5200 , n5195 , n5198 );
or ( n5201 , n5197 , n5199 , n5200 );
and ( n5202 , n5193 , n5201 );
and ( n5203 , n5185 , n5201 );
or ( n5204 , n5194 , n5202 , n5203 );
and ( n5205 , n5171 , n5204 );
and ( n5206 , n5149 , n5204 );
or ( n5207 , n5172 , n5205 , n5206 );
and ( n5208 , n5139 , n5207 );
xor ( n5209 , n4890 , n4891 );
xor ( n5210 , n4822 , n4823 );
and ( n5211 , n5209 , n5210 );
xor ( n5212 , n4897 , n4898 );
and ( n5213 , n5210 , n5212 );
and ( n5214 , n5209 , n5212 );
or ( n5215 , n5211 , n5213 , n5214 );
xor ( n5216 , n4910 , n4911 );
xor ( n5217 , n4913 , n4914 );
and ( n5218 , n5216 , n5217 );
and ( n5219 , n1275 , n4982 );
and ( n5220 , n1995 , n2586 );
or ( n5221 , n5219 , n5220 );
and ( n5222 , n5217 , n5221 );
and ( n5223 , n5216 , n5221 );
or ( n5224 , n5218 , n5222 , n5223 );
and ( n5225 , n5215 , n5224 );
and ( n5226 , n2048 , n2492 );
and ( n5227 , n2497 , n2059 );
and ( n5228 , n5226 , n5227 );
and ( n5229 , n4989 , n1293 );
and ( n5230 , n2591 , n1990 );
and ( n5231 , n5229 , n5230 );
buf ( n5232 , n2716 );
buf ( n5233 , n5232 );
buf ( n5234 , n2010 );
buf ( n5235 , n5234 );
buf ( n5236 , n2033 );
buf ( n5237 , n5236 );
xor ( n5238 , n5235 , n5237 );
buf ( n5239 , n2265 );
buf ( n5240 , n5239 );
xor ( n5241 , n5237 , n5240 );
not ( n5242 , n5241 );
and ( n5243 , n5238 , n5242 );
and ( n5244 , n5233 , n5243 );
buf ( n5245 , n2584 );
buf ( n5246 , n5245 );
and ( n5247 , n5246 , n5241 );
nor ( n5248 , n5244 , n5247 );
and ( n5249 , n5237 , n5240 );
not ( n5250 , n5249 );
and ( n5251 , n5235 , n5250 );
xnor ( n5252 , n5248 , n5251 );
buf ( n5253 , n3144 );
buf ( n5254 , n5253 );
buf ( n5255 , n1823 );
buf ( n5256 , n5255 );
buf ( n5257 , n1854 );
buf ( n5258 , n5257 );
xor ( n5259 , n5256 , n5258 );
xor ( n5260 , n5258 , n5235 );
not ( n5261 , n5260 );
and ( n5262 , n5259 , n5261 );
and ( n5263 , n5254 , n5262 );
buf ( n5264 , n2921 );
buf ( n5265 , n5264 );
and ( n5266 , n5265 , n5260 );
nor ( n5267 , n5263 , n5266 );
and ( n5268 , n5258 , n5235 );
not ( n5269 , n5268 );
and ( n5270 , n5256 , n5269 );
xnor ( n5271 , n5267 , n5270 );
and ( n5272 , n5252 , n5271 );
buf ( n5273 , n3447 );
buf ( n5274 , n5273 );
buf ( n5275 , n1562 );
buf ( n5276 , n5275 );
buf ( n5277 , n1730 );
buf ( n5278 , n5277 );
xor ( n5279 , n5276 , n5278 );
xor ( n5280 , n5278 , n5256 );
not ( n5281 , n5280 );
and ( n5282 , n5279 , n5281 );
and ( n5283 , n5274 , n5282 );
buf ( n5284 , n3286 );
buf ( n5285 , n5284 );
and ( n5286 , n5285 , n5280 );
nor ( n5287 , n5283 , n5286 );
and ( n5288 , n5278 , n5256 );
not ( n5289 , n5288 );
and ( n5290 , n5276 , n5289 );
xnor ( n5291 , n5287 , n5290 );
and ( n5292 , n5271 , n5291 );
and ( n5293 , n5252 , n5291 );
or ( n5294 , n5272 , n5292 , n5293 );
buf ( n5295 , n1776 );
buf ( n5296 , n5295 );
buf ( n5297 , n3167 );
buf ( n5298 , n5297 );
buf ( n5299 , n3244 );
buf ( n5300 , n5299 );
xor ( n5301 , n5298 , n5300 );
buf ( n5302 , n3337 );
buf ( n5303 , n5302 );
xor ( n5304 , n5300 , n5303 );
not ( n5305 , n5304 );
and ( n5306 , n5301 , n5305 );
and ( n5307 , n5296 , n5306 );
buf ( n5308 , n1717 );
buf ( n5309 , n5308 );
and ( n5310 , n5309 , n5304 );
nor ( n5311 , n5307 , n5310 );
and ( n5312 , n5300 , n5303 );
not ( n5313 , n5312 );
and ( n5314 , n5298 , n5313 );
xnor ( n5315 , n5311 , n5314 );
buf ( n5316 , n2490 );
buf ( n5317 , n5316 );
buf ( n5318 , n2284 );
buf ( n5319 , n5318 );
xor ( n5320 , n5240 , n5319 );
buf ( n5321 , n2475 );
buf ( n5322 , n5321 );
xor ( n5323 , n5319 , n5322 );
not ( n5324 , n5323 );
and ( n5325 , n5320 , n5324 );
and ( n5326 , n5317 , n5325 );
buf ( n5327 , n2302 );
buf ( n5328 , n5327 );
and ( n5329 , n5328 , n5323 );
nor ( n5330 , n5326 , n5329 );
and ( n5331 , n5319 , n5322 );
not ( n5332 , n5331 );
and ( n5333 , n5240 , n5332 );
xnor ( n5334 , n5330 , n5333 );
and ( n5335 , n5315 , n5334 );
buf ( n5336 , n777 );
buf ( n5337 , n5336 );
buf ( n5338 , n5337 );
buf ( n5339 , n5338 );
buf ( n5340 , n5339 );
buf ( n5341 , n1263 );
buf ( n5342 , n5341 );
and ( n5343 , n5340 , n5342 );
and ( n5344 , n5334 , n5343 );
and ( n5345 , n5315 , n5343 );
or ( n5346 , n5335 , n5344 , n5345 );
xor ( n5347 , n5294 , n5346 );
and ( n5348 , n5328 , n5325 );
buf ( n5349 , n2248 );
buf ( n5350 , n5349 );
and ( n5351 , n5350 , n5323 );
nor ( n5352 , n5348 , n5351 );
xnor ( n5353 , n5352 , n5333 );
buf ( n5354 , n4148 );
buf ( n5355 , n5354 );
buf ( n5356 , n1383 );
buf ( n5357 , n5356 );
buf ( n5358 , n1439 );
buf ( n5359 , n5358 );
xor ( n5360 , n5357 , n5359 );
buf ( n5361 , n1470 );
buf ( n5362 , n5361 );
xor ( n5363 , n5359 , n5362 );
not ( n5364 , n5363 );
and ( n5365 , n5360 , n5364 );
and ( n5366 , n5355 , n5365 );
buf ( n5367 , n3890 );
buf ( n5368 , n5367 );
and ( n5369 , n5368 , n5363 );
nor ( n5370 , n5366 , n5369 );
and ( n5371 , n5359 , n5362 );
not ( n5372 , n5371 );
and ( n5373 , n5357 , n5372 );
xnor ( n5374 , n5370 , n5373 );
xor ( n5375 , n5353 , n5374 );
buf ( n5376 , n1273 );
buf ( n5377 , n5376 );
buf ( n5378 , n776 );
buf ( n5379 , n5378 );
buf ( n5380 , n5379 );
buf ( n5381 , n5380 );
buf ( n5382 , n5381 );
buf ( n5383 , n777 );
buf ( n5384 , n5383 );
buf ( n5385 , n5384 );
buf ( n5386 , n5385 );
buf ( n5387 , n5386 );
xor ( n5388 , n5382 , n5387 );
not ( n5389 , n5387 );
and ( n5390 , n5388 , n5389 );
and ( n5391 , n5377 , n5390 );
buf ( n5392 , n1103 );
buf ( n5393 , n5392 );
and ( n5394 , n5393 , n5387 );
nor ( n5395 , n5391 , n5394 );
xnor ( n5396 , n5395 , n5382 );
buf ( n5397 , n4383 );
buf ( n5398 , n5397 );
buf ( n5399 , n4577 );
buf ( n5400 , n5399 );
buf ( n5401 , n4719 );
buf ( n5402 , n5401 );
and ( n5403 , n5400 , n5402 );
not ( n5404 , n5403 );
and ( n5405 , n5398 , n5404 );
and ( n5406 , n5396 , n5405 );
buf ( n5407 , n1310 );
buf ( n5408 , n5407 );
buf ( n5409 , n5175 );
buf ( n5410 , n5409 );
xor ( n5411 , n5402 , n5410 );
xor ( n5412 , n5410 , n5382 );
not ( n5413 , n5412 );
and ( n5414 , n5411 , n5413 );
and ( n5415 , n5408 , n5414 );
and ( n5416 , n5377 , n5412 );
nor ( n5417 , n5415 , n5416 );
and ( n5418 , n5410 , n5382 );
not ( n5419 , n5418 );
and ( n5420 , n5402 , n5419 );
xnor ( n5421 , n5417 , n5420 );
and ( n5422 , n5406 , n5421 );
buf ( n5423 , n3831 );
buf ( n5424 , n5423 );
buf ( n5425 , n4136 );
buf ( n5426 , n5425 );
and ( n5427 , n5426 , n5398 );
not ( n5428 , n5427 );
and ( n5429 , n5424 , n5428 );
and ( n5430 , n5421 , n5429 );
and ( n5431 , n5406 , n5429 );
or ( n5432 , n5422 , n5430 , n5431 );
and ( n5433 , n5393 , n5390 );
not ( n5434 , n5433 );
xnor ( n5435 , n5434 , n5382 );
buf ( n5436 , n1346 );
buf ( n5437 , n5436 );
xor ( n5438 , n5400 , n5402 );
and ( n5439 , n5437 , n5438 );
not ( n5440 , n5439 );
xnor ( n5441 , n5440 , n5405 );
xor ( n5442 , n5435 , n5441 );
xor ( n5443 , n5396 , n5405 );
and ( n5444 , n5437 , n5414 );
and ( n5445 , n5408 , n5412 );
nor ( n5446 , n5444 , n5445 );
xnor ( n5447 , n5446 , n5420 );
and ( n5448 , n5443 , n5447 );
and ( n5449 , n5447 , n5429 );
and ( n5450 , n5443 , n5429 );
or ( n5451 , n5448 , n5449 , n5450 );
and ( n5452 , n5442 , n5451 );
xor ( n5453 , n5406 , n5421 );
xor ( n5454 , n5453 , n5429 );
and ( n5455 , n5451 , n5454 );
and ( n5456 , n5442 , n5454 );
or ( n5457 , n5452 , n5455 , n5456 );
xor ( n5458 , n5432 , n5457 );
and ( n5459 , n5435 , n5441 );
and ( n5460 , n5377 , n5414 );
and ( n5461 , n5393 , n5412 );
nor ( n5462 , n5460 , n5461 );
xnor ( n5463 , n5462 , n5420 );
not ( n5464 , n5463 );
xor ( n5465 , n5459 , n5464 );
xor ( n5466 , n5398 , n5400 );
not ( n5467 , n5438 );
and ( n5468 , n5466 , n5467 );
and ( n5469 , n5437 , n5468 );
and ( n5470 , n5408 , n5438 );
nor ( n5471 , n5469 , n5470 );
xnor ( n5472 , n5471 , n5405 );
xor ( n5473 , n5472 , n5429 );
buf ( n5474 , n3643 );
buf ( n5475 , n5474 );
and ( n5476 , n5475 , n5424 );
not ( n5477 , n5476 );
and ( n5478 , n5303 , n5477 );
xor ( n5479 , n5473 , n5478 );
xor ( n5480 , n5465 , n5479 );
xor ( n5481 , n5458 , n5480 );
xor ( n5482 , n5375 , n5481 );
xor ( n5483 , n5347 , n5482 );
xor ( n5484 , n5303 , n5475 );
xor ( n5485 , n5475 , n5424 );
not ( n5486 , n5485 );
and ( n5487 , n5484 , n5486 );
and ( n5488 , n5296 , n5487 );
and ( n5489 , n5309 , n5485 );
nor ( n5490 , n5488 , n5489 );
xnor ( n5491 , n5490 , n5478 );
buf ( n5492 , n2632 );
buf ( n5493 , n5492 );
xor ( n5494 , n5322 , n5493 );
buf ( n5495 , n2762 );
buf ( n5496 , n5495 );
xor ( n5497 , n5493 , n5496 );
not ( n5498 , n5497 );
and ( n5499 , n5494 , n5498 );
and ( n5500 , n5317 , n5499 );
and ( n5501 , n5328 , n5497 );
nor ( n5502 , n5500 , n5501 );
and ( n5503 , n5493 , n5496 );
not ( n5504 , n5503 );
and ( n5505 , n5322 , n5504 );
xnor ( n5506 , n5502 , n5505 );
xor ( n5507 , n5491 , n5506 );
buf ( n5508 , n1299 );
buf ( n5509 , n5508 );
buf ( n5510 , n1283 );
buf ( n5511 , n5510 );
xor ( n5512 , n5509 , n5511 );
and ( n5513 , n5340 , n5512 );
xor ( n5514 , n5507 , n5513 );
and ( n5515 , n5437 , n5390 );
and ( n5516 , n5408 , n5387 );
nor ( n5517 , n5515 , n5516 );
xnor ( n5518 , n5517 , n5382 );
and ( n5519 , n5518 , n5420 );
and ( n5520 , n5420 , n5405 );
and ( n5521 , n5518 , n5405 );
or ( n5522 , n5519 , n5520 , n5521 );
and ( n5523 , n5514 , n5522 );
and ( n5524 , n5285 , n5243 );
and ( n5525 , n5254 , n5241 );
nor ( n5526 , n5524 , n5525 );
xnor ( n5527 , n5526 , n5251 );
buf ( n5528 , n3726 );
buf ( n5529 , n5528 );
and ( n5530 , n5529 , n5262 );
and ( n5531 , n5274 , n5260 );
nor ( n5532 , n5530 , n5531 );
xnor ( n5533 , n5532 , n5270 );
and ( n5534 , n5527 , n5533 );
buf ( n5535 , n4732 );
buf ( n5536 , n5535 );
buf ( n5537 , n1524 );
buf ( n5538 , n5537 );
xor ( n5539 , n5362 , n5538 );
xor ( n5540 , n5538 , n5276 );
not ( n5541 , n5540 );
and ( n5542 , n5539 , n5541 );
and ( n5543 , n5536 , n5542 );
buf ( n5544 , n4360 );
buf ( n5545 , n5544 );
and ( n5546 , n5545 , n5540 );
nor ( n5547 , n5543 , n5546 );
and ( n5548 , n5538 , n5276 );
not ( n5549 , n5548 );
and ( n5550 , n5362 , n5549 );
xnor ( n5551 , n5547 , n5550 );
and ( n5552 , n5533 , n5551 );
and ( n5553 , n5527 , n5551 );
or ( n5554 , n5534 , n5552 , n5553 );
and ( n5555 , n5522 , n5554 );
and ( n5556 , n5514 , n5554 );
or ( n5557 , n5523 , n5555 , n5556 );
not ( n5558 , n5513 );
and ( n5559 , n5509 , n5511 );
not ( n5560 , n5559 );
and ( n5561 , n5342 , n5560 );
and ( n5562 , n5558 , n5561 );
buf ( n5563 , n778 );
buf ( n5564 , n5563 );
buf ( n5565 , n5564 );
buf ( n5566 , n779 );
buf ( n5567 , n5566 );
and ( n5568 , n5564 , n5567 );
buf ( n5569 , n779 );
buf ( n5570 , n5569 );
buf ( n5571 , n778 );
buf ( n5572 , n5571 );
and ( n5573 , n5570 , n5572 );
and ( n5574 , n5568 , n5573 );
and ( n5575 , n5565 , n5574 );
xor ( n5576 , n5568 , n5573 );
buf ( n5577 , n780 );
buf ( n5578 , n5577 );
and ( n5579 , n5564 , n5578 );
buf ( n5580 , n780 );
buf ( n5581 , n5580 );
and ( n5582 , n5581 , n5572 );
and ( n5583 , n5579 , n5582 );
and ( n5584 , n5576 , n5583 );
buf ( n5585 , n5570 );
xor ( n5586 , n5579 , n5582 );
and ( n5587 , n5585 , n5586 );
buf ( n5588 , n781 );
buf ( n5589 , n5588 );
and ( n5590 , n5564 , n5589 );
buf ( n5591 , n781 );
buf ( n5592 , n5591 );
and ( n5593 , n5592 , n5572 );
and ( n5594 , n5590 , n5593 );
and ( n5595 , n5586 , n5594 );
and ( n5596 , n5585 , n5594 );
or ( n5597 , n5587 , n5595 , n5596 );
and ( n5598 , n5583 , n5597 );
and ( n5599 , n5576 , n5597 );
or ( n5600 , n5584 , n5598 , n5599 );
and ( n5601 , n5574 , n5600 );
and ( n5602 , n5565 , n5600 );
or ( n5603 , n5575 , n5601 , n5602 );
xor ( n5604 , n5565 , n5574 );
xor ( n5605 , n5604 , n5600 );
buf ( n5606 , n782 );
buf ( n5607 , n5606 );
and ( n5608 , n5607 , n5572 );
and ( n5609 , n5592 , n5567 );
or ( n5610 , n5608 , n5609 );
buf ( n5611 , n782 );
buf ( n5612 , n5611 );
and ( n5613 , n5564 , n5612 );
and ( n5614 , n5570 , n5589 );
or ( n5615 , n5613 , n5614 );
and ( n5616 , n5610 , n5615 );
and ( n5617 , n5581 , n5567 );
and ( n5618 , n5570 , n5578 );
and ( n5619 , n5617 , n5618 );
xor ( n5620 , n5590 , n5593 );
and ( n5621 , n5618 , n5620 );
and ( n5622 , n5617 , n5620 );
or ( n5623 , n5619 , n5621 , n5622 );
and ( n5624 , n5616 , n5623 );
xor ( n5625 , n5585 , n5586 );
xor ( n5626 , n5625 , n5594 );
and ( n5627 , n5623 , n5626 );
and ( n5628 , n5616 , n5626 );
or ( n5629 , n5624 , n5627 , n5628 );
xor ( n5630 , n5576 , n5583 );
xor ( n5631 , n5630 , n5597 );
and ( n5632 , n5629 , n5631 );
xor ( n5633 , n5610 , n5615 );
xnor ( n5634 , n5608 , n5609 );
xnor ( n5635 , n5613 , n5614 );
and ( n5636 , n5634 , n5635 );
and ( n5637 , n5633 , n5636 );
buf ( n5638 , n5581 );
buf ( n5639 , n783 );
buf ( n5640 , n5639 );
and ( n5641 , n5564 , n5640 );
buf ( n5642 , n783 );
buf ( n5643 , n5642 );
and ( n5644 , n5643 , n5572 );
and ( n5645 , n5641 , n5644 );
and ( n5646 , n5638 , n5645 );
and ( n5647 , n5570 , n5612 );
and ( n5648 , n5607 , n5567 );
and ( n5649 , n5647 , n5648 );
and ( n5650 , n5645 , n5649 );
and ( n5651 , n5638 , n5649 );
or ( n5652 , n5646 , n5650 , n5651 );
and ( n5653 , n5636 , n5652 );
and ( n5654 , n5633 , n5652 );
or ( n5655 , n5637 , n5653 , n5654 );
xor ( n5656 , n5616 , n5623 );
xor ( n5657 , n5656 , n5626 );
and ( n5658 , n5655 , n5657 );
xor ( n5659 , n5617 , n5618 );
xor ( n5660 , n5659 , n5620 );
and ( n5661 , n5581 , n5589 );
and ( n5662 , n5592 , n5578 );
and ( n5663 , n5661 , n5662 );
xor ( n5664 , n5634 , n5635 );
and ( n5665 , n5663 , n5664 );
buf ( n5666 , n784 );
buf ( n5667 , n5666 );
and ( n5668 , n5667 , n5572 );
and ( n5669 , n5643 , n5567 );
and ( n5670 , n5668 , n5669 );
and ( n5671 , n5607 , n5578 );
and ( n5672 , n5669 , n5671 );
and ( n5673 , n5668 , n5671 );
or ( n5674 , n5670 , n5672 , n5673 );
buf ( n5675 , n784 );
buf ( n5676 , n5675 );
and ( n5677 , n5564 , n5676 );
and ( n5678 , n5570 , n5640 );
and ( n5679 , n5677 , n5678 );
and ( n5680 , n5581 , n5612 );
and ( n5681 , n5678 , n5680 );
and ( n5682 , n5677 , n5680 );
or ( n5683 , n5679 , n5681 , n5682 );
and ( n5684 , n5674 , n5683 );
and ( n5685 , n5664 , n5684 );
and ( n5686 , n5663 , n5684 );
or ( n5687 , n5665 , n5685 , n5686 );
and ( n5688 , n5660 , n5687 );
xor ( n5689 , n5633 , n5636 );
xor ( n5690 , n5689 , n5652 );
and ( n5691 , n5687 , n5690 );
and ( n5692 , n5660 , n5690 );
or ( n5693 , n5688 , n5691 , n5692 );
and ( n5694 , n5657 , n5693 );
and ( n5695 , n5655 , n5693 );
or ( n5696 , n5658 , n5694 , n5695 );
and ( n5697 , n5631 , n5696 );
and ( n5698 , n5629 , n5696 );
or ( n5699 , n5632 , n5697 , n5698 );
and ( n5700 , n5605 , n5699 );
xor ( n5701 , n5629 , n5631 );
xor ( n5702 , n5701 , n5696 );
xor ( n5703 , n5655 , n5657 );
xor ( n5704 , n5703 , n5693 );
xor ( n5705 , n5641 , n5644 );
xor ( n5706 , n5647 , n5648 );
and ( n5707 , n5705 , n5706 );
xor ( n5708 , n5661 , n5662 );
and ( n5709 , n5706 , n5708 );
and ( n5710 , n5705 , n5708 );
or ( n5711 , n5707 , n5709 , n5710 );
xor ( n5712 , n5638 , n5645 );
xor ( n5713 , n5712 , n5649 );
and ( n5714 , n5711 , n5713 );
xor ( n5715 , n5674 , n5683 );
xor ( n5716 , n5668 , n5669 );
xor ( n5717 , n5716 , n5671 );
xor ( n5718 , n5677 , n5678 );
xor ( n5719 , n5718 , n5680 );
and ( n5720 , n5717 , n5719 );
and ( n5721 , n5715 , n5720 );
xor ( n5722 , n5705 , n5706 );
xor ( n5723 , n5722 , n5708 );
and ( n5724 , n5720 , n5723 );
and ( n5725 , n5715 , n5723 );
or ( n5726 , n5721 , n5724 , n5725 );
and ( n5727 , n5713 , n5726 );
and ( n5728 , n5711 , n5726 );
or ( n5729 , n5714 , n5727 , n5728 );
xor ( n5730 , n5660 , n5687 );
xor ( n5731 , n5730 , n5690 );
and ( n5732 , n5729 , n5731 );
xor ( n5733 , n5663 , n5664 );
xor ( n5734 , n5733 , n5684 );
buf ( n5735 , n786 );
buf ( n5736 , n5735 );
and ( n5737 , n5564 , n5736 );
and ( n5738 , n5581 , n5676 );
and ( n5739 , n5737 , n5738 );
and ( n5740 , n5592 , n5640 );
and ( n5741 , n5738 , n5740 );
and ( n5742 , n5737 , n5740 );
or ( n5743 , n5739 , n5741 , n5742 );
buf ( n5744 , n785 );
buf ( n5745 , n5744 );
and ( n5746 , n5745 , n5572 );
and ( n5747 , n5743 , n5746 );
and ( n5748 , n5643 , n5578 );
and ( n5749 , n5746 , n5748 );
and ( n5750 , n5743 , n5748 );
or ( n5751 , n5747 , n5749 , n5750 );
buf ( n5752 , n786 );
buf ( n5753 , n5752 );
and ( n5754 , n5753 , n5572 );
and ( n5755 , n5667 , n5578 );
and ( n5756 , n5754 , n5755 );
and ( n5757 , n5643 , n5589 );
and ( n5758 , n5755 , n5757 );
and ( n5759 , n5754 , n5757 );
or ( n5760 , n5756 , n5758 , n5759 );
buf ( n5761 , n785 );
buf ( n5762 , n5761 );
and ( n5763 , n5564 , n5762 );
and ( n5764 , n5760 , n5763 );
and ( n5765 , n5581 , n5640 );
and ( n5766 , n5763 , n5765 );
and ( n5767 , n5760 , n5765 );
or ( n5768 , n5764 , n5766 , n5767 );
and ( n5769 , n5751 , n5768 );
buf ( n5770 , n5592 );
and ( n5771 , n5570 , n5676 );
and ( n5772 , n5667 , n5567 );
and ( n5773 , n5771 , n5772 );
and ( n5774 , n5770 , n5773 );
xor ( n5775 , n5717 , n5719 );
and ( n5776 , n5773 , n5775 );
and ( n5777 , n5770 , n5775 );
or ( n5778 , n5774 , n5776 , n5777 );
and ( n5779 , n5769 , n5778 );
xor ( n5780 , n5715 , n5720 );
xor ( n5781 , n5780 , n5723 );
and ( n5782 , n5778 , n5781 );
and ( n5783 , n5769 , n5781 );
or ( n5784 , n5779 , n5782 , n5783 );
and ( n5785 , n5734 , n5784 );
xor ( n5786 , n5711 , n5713 );
xor ( n5787 , n5786 , n5726 );
and ( n5788 , n5784 , n5787 );
and ( n5789 , n5734 , n5787 );
or ( n5790 , n5785 , n5788 , n5789 );
and ( n5791 , n5731 , n5790 );
and ( n5792 , n5729 , n5790 );
or ( n5793 , n5732 , n5791 , n5792 );
and ( n5794 , n5704 , n5793 );
xor ( n5795 , n5729 , n5731 );
xor ( n5796 , n5795 , n5790 );
xor ( n5797 , n5734 , n5784 );
xor ( n5798 , n5797 , n5787 );
and ( n5799 , n5607 , n5589 );
and ( n5800 , n5592 , n5612 );
and ( n5801 , n5799 , n5800 );
xor ( n5802 , n5771 , n5772 );
and ( n5803 , n5800 , n5802 );
and ( n5804 , n5799 , n5802 );
or ( n5805 , n5801 , n5803 , n5804 );
xor ( n5806 , n5751 , n5768 );
and ( n5807 , n5805 , n5806 );
xor ( n5808 , n5743 , n5746 );
xor ( n5809 , n5808 , n5748 );
xor ( n5810 , n5760 , n5763 );
xor ( n5811 , n5810 , n5765 );
and ( n5812 , n5809 , n5811 );
and ( n5813 , n5806 , n5812 );
and ( n5814 , n5805 , n5812 );
or ( n5815 , n5807 , n5813 , n5814 );
xor ( n5816 , n5769 , n5778 );
xor ( n5817 , n5816 , n5781 );
and ( n5818 , n5815 , n5817 );
and ( n5819 , n5570 , n5762 );
and ( n5820 , n5745 , n5567 );
and ( n5821 , n5819 , n5820 );
and ( n5822 , n5753 , n5567 );
and ( n5823 , n5667 , n5589 );
or ( n5824 , n5822 , n5823 );
and ( n5825 , n5570 , n5736 );
and ( n5826 , n5592 , n5676 );
or ( n5827 , n5825 , n5826 );
and ( n5828 , n5824 , n5827 );
and ( n5829 , n5821 , n5828 );
xor ( n5830 , n5754 , n5755 );
xor ( n5831 , n5830 , n5757 );
xor ( n5832 , n5737 , n5738 );
xor ( n5833 , n5832 , n5740 );
and ( n5834 , n5831 , n5833 );
and ( n5835 , n5828 , n5834 );
and ( n5836 , n5821 , n5834 );
or ( n5837 , n5829 , n5835 , n5836 );
xor ( n5838 , n5770 , n5773 );
xor ( n5839 , n5838 , n5775 );
and ( n5840 , n5837 , n5839 );
buf ( n5841 , n5607 );
xor ( n5842 , n5819 , n5820 );
and ( n5843 , n5841 , n5842 );
and ( n5844 , n5581 , n5762 );
and ( n5845 , n5745 , n5578 );
and ( n5846 , n5844 , n5845 );
and ( n5847 , n5842 , n5846 );
and ( n5848 , n5841 , n5846 );
or ( n5849 , n5843 , n5847 , n5848 );
xor ( n5850 , n5799 , n5800 );
xor ( n5851 , n5850 , n5802 );
and ( n5852 , n5849 , n5851 );
xor ( n5853 , n5809 , n5811 );
and ( n5854 , n5851 , n5853 );
and ( n5855 , n5849 , n5853 );
or ( n5856 , n5852 , n5854 , n5855 );
and ( n5857 , n5839 , n5856 );
and ( n5858 , n5837 , n5856 );
or ( n5859 , n5840 , n5857 , n5858 );
and ( n5860 , n5817 , n5859 );
and ( n5861 , n5815 , n5859 );
or ( n5862 , n5818 , n5860 , n5861 );
and ( n5863 , n5798 , n5862 );
buf ( n5864 , n787 );
buf ( n5865 , n5864 );
and ( n5866 , n5865 , n5572 );
not ( n5867 , n5866 );
xnor ( n5868 , n5825 , n5826 );
and ( n5869 , n5867 , n5868 );
buf ( n5870 , n787 );
buf ( n5871 , n5870 );
and ( n5872 , n5564 , n5871 );
not ( n5873 , n5872 );
xnor ( n5874 , n5822 , n5823 );
and ( n5875 , n5873 , n5874 );
and ( n5876 , n5869 , n5875 );
buf ( n5877 , n5866 );
buf ( n5878 , n5872 );
and ( n5879 , n5877 , n5878 );
and ( n5880 , n5876 , n5879 );
xor ( n5881 , n5824 , n5827 );
xor ( n5882 , n5831 , n5833 );
and ( n5883 , n5881 , n5882 );
and ( n5884 , n5865 , n5567 );
and ( n5885 , n5745 , n5589 );
and ( n5886 , n5884 , n5885 );
and ( n5887 , n5667 , n5612 );
and ( n5888 , n5885 , n5887 );
and ( n5889 , n5884 , n5887 );
or ( n5890 , n5886 , n5888 , n5889 );
and ( n5891 , n5570 , n5871 );
and ( n5892 , n5592 , n5762 );
and ( n5893 , n5891 , n5892 );
and ( n5894 , n5607 , n5676 );
and ( n5895 , n5892 , n5894 );
and ( n5896 , n5891 , n5894 );
or ( n5897 , n5893 , n5895 , n5896 );
and ( n5898 , n5890 , n5897 );
and ( n5899 , n5882 , n5898 );
and ( n5900 , n5881 , n5898 );
or ( n5901 , n5883 , n5899 , n5900 );
and ( n5902 , n5879 , n5901 );
and ( n5903 , n5876 , n5901 );
or ( n5904 , n5880 , n5902 , n5903 );
xor ( n5905 , n5805 , n5806 );
xor ( n5906 , n5905 , n5812 );
and ( n5907 , n5904 , n5906 );
xor ( n5908 , n5821 , n5828 );
xor ( n5909 , n5908 , n5834 );
and ( n5910 , n5643 , n5612 );
and ( n5911 , n5607 , n5640 );
and ( n5912 , n5910 , n5911 );
xor ( n5913 , n5844 , n5845 );
and ( n5914 , n5911 , n5913 );
and ( n5915 , n5910 , n5913 );
or ( n5916 , n5912 , n5914 , n5915 );
xor ( n5917 , n5841 , n5842 );
xor ( n5918 , n5917 , n5846 );
and ( n5919 , n5916 , n5918 );
xor ( n5920 , n5869 , n5875 );
and ( n5921 , n5918 , n5920 );
and ( n5922 , n5916 , n5920 );
or ( n5923 , n5919 , n5921 , n5922 );
and ( n5924 , n5909 , n5923 );
xor ( n5925 , n5877 , n5878 );
buf ( n5926 , n788 );
buf ( n5927 , n5926 );
and ( n5928 , n5570 , n5927 );
and ( n5929 , n5581 , n5871 );
and ( n5930 , n5928 , n5929 );
and ( n5931 , n5607 , n5762 );
and ( n5932 , n5929 , n5931 );
and ( n5933 , n5928 , n5931 );
or ( n5934 , n5930 , n5932 , n5933 );
buf ( n5935 , n788 );
buf ( n5936 , n5935 );
and ( n5937 , n5936 , n5572 );
and ( n5938 , n5934 , n5937 );
and ( n5939 , n5753 , n5578 );
and ( n5940 , n5937 , n5939 );
and ( n5941 , n5934 , n5939 );
or ( n5942 , n5938 , n5940 , n5941 );
and ( n5943 , n5936 , n5567 );
and ( n5944 , n5865 , n5578 );
and ( n5945 , n5943 , n5944 );
and ( n5946 , n5745 , n5612 );
and ( n5947 , n5944 , n5946 );
and ( n5948 , n5943 , n5946 );
or ( n5949 , n5945 , n5947 , n5948 );
and ( n5950 , n5564 , n5927 );
and ( n5951 , n5949 , n5950 );
and ( n5952 , n5581 , n5736 );
and ( n5953 , n5950 , n5952 );
and ( n5954 , n5949 , n5952 );
or ( n5955 , n5951 , n5953 , n5954 );
and ( n5956 , n5942 , n5955 );
and ( n5957 , n5925 , n5956 );
xor ( n5958 , n5867 , n5868 );
xor ( n5959 , n5873 , n5874 );
and ( n5960 , n5958 , n5959 );
and ( n5961 , n5956 , n5960 );
and ( n5962 , n5925 , n5960 );
or ( n5963 , n5957 , n5961 , n5962 );
and ( n5964 , n5923 , n5963 );
and ( n5965 , n5909 , n5963 );
or ( n5966 , n5924 , n5964 , n5965 );
and ( n5967 , n5906 , n5966 );
and ( n5968 , n5904 , n5966 );
or ( n5969 , n5907 , n5967 , n5968 );
xor ( n5970 , n5815 , n5817 );
xor ( n5971 , n5970 , n5859 );
and ( n5972 , n5969 , n5971 );
xor ( n5973 , n5837 , n5839 );
xor ( n5974 , n5973 , n5856 );
xor ( n5975 , n5849 , n5851 );
xor ( n5976 , n5975 , n5853 );
xor ( n5977 , n5876 , n5879 );
xor ( n5978 , n5977 , n5901 );
and ( n5979 , n5976 , n5978 );
xor ( n5980 , n5890 , n5897 );
xor ( n5981 , n5884 , n5885 );
xor ( n5982 , n5981 , n5887 );
xor ( n5983 , n5891 , n5892 );
xor ( n5984 , n5983 , n5894 );
and ( n5985 , n5982 , n5984 );
and ( n5986 , n5980 , n5985 );
buf ( n5987 , n5643 );
buf ( n5988 , n789 );
buf ( n5989 , n5988 );
and ( n5990 , n5564 , n5989 );
buf ( n5991 , n789 );
buf ( n5992 , n5991 );
and ( n5993 , n5992 , n5572 );
and ( n5994 , n5990 , n5993 );
and ( n5995 , n5987 , n5994 );
and ( n5996 , n5592 , n5736 );
and ( n5997 , n5753 , n5589 );
and ( n5998 , n5996 , n5997 );
and ( n5999 , n5994 , n5998 );
and ( n6000 , n5987 , n5998 );
or ( n6001 , n5995 , n5999 , n6000 );
and ( n6002 , n5985 , n6001 );
and ( n6003 , n5980 , n6001 );
or ( n6004 , n5986 , n6002 , n6003 );
xor ( n6005 , n5881 , n5882 );
xor ( n6006 , n6005 , n5898 );
and ( n6007 , n6004 , n6006 );
xor ( n6008 , n5910 , n5911 );
xor ( n6009 , n6008 , n5913 );
xor ( n6010 , n5942 , n5955 );
and ( n6011 , n6009 , n6010 );
xor ( n6012 , n5958 , n5959 );
and ( n6013 , n6010 , n6012 );
and ( n6014 , n6009 , n6012 );
or ( n6015 , n6011 , n6013 , n6014 );
and ( n6016 , n6006 , n6015 );
and ( n6017 , n6004 , n6015 );
or ( n6018 , n6007 , n6016 , n6017 );
and ( n6019 , n5978 , n6018 );
and ( n6020 , n5976 , n6018 );
or ( n6021 , n5979 , n6019 , n6020 );
and ( n6022 , n5974 , n6021 );
xor ( n6023 , n5904 , n5906 );
xor ( n6024 , n6023 , n5966 );
and ( n6025 , n6021 , n6024 );
and ( n6026 , n5974 , n6024 );
or ( n6027 , n6022 , n6025 , n6026 );
and ( n6028 , n5971 , n6027 );
and ( n6029 , n5969 , n6027 );
or ( n6030 , n5972 , n6028 , n6029 );
and ( n6031 , n5862 , n6030 );
and ( n6032 , n5798 , n6030 );
or ( n6033 , n5863 , n6031 , n6032 );
and ( n6034 , n5796 , n6033 );
xor ( n6035 , n5798 , n5862 );
xor ( n6036 , n6035 , n6030 );
xor ( n6037 , n5969 , n5971 );
xor ( n6038 , n6037 , n6027 );
xor ( n6039 , n5934 , n5937 );
xor ( n6040 , n6039 , n5939 );
xor ( n6041 , n5949 , n5950 );
xor ( n6042 , n6041 , n5952 );
and ( n6043 , n6040 , n6042 );
and ( n6044 , n5643 , n5676 );
and ( n6045 , n5667 , n5640 );
and ( n6046 , n6044 , n6045 );
xor ( n6047 , n5982 , n5984 );
and ( n6048 , n6046 , n6047 );
and ( n6049 , n5936 , n5578 );
and ( n6050 , n5753 , n5612 );
or ( n6051 , n6049 , n6050 );
and ( n6052 , n5581 , n5927 );
and ( n6053 , n5607 , n5736 );
or ( n6054 , n6052 , n6053 );
and ( n6055 , n6051 , n6054 );
and ( n6056 , n6047 , n6055 );
and ( n6057 , n6046 , n6055 );
or ( n6058 , n6048 , n6056 , n6057 );
and ( n6059 , n6043 , n6058 );
and ( n6060 , n5992 , n5567 );
and ( n6061 , n5865 , n5589 );
or ( n6062 , n6060 , n6061 );
and ( n6063 , n5570 , n5989 );
and ( n6064 , n5592 , n5871 );
or ( n6065 , n6063 , n6064 );
and ( n6066 , n6062 , n6065 );
xor ( n6067 , n5943 , n5944 );
xor ( n6068 , n6067 , n5946 );
xor ( n6069 , n5928 , n5929 );
xor ( n6070 , n6069 , n5931 );
and ( n6071 , n6068 , n6070 );
and ( n6072 , n6066 , n6071 );
xor ( n6073 , n5990 , n5993 );
xor ( n6074 , n5996 , n5997 );
and ( n6075 , n6073 , n6074 );
xor ( n6076 , n6044 , n6045 );
and ( n6077 , n6074 , n6076 );
and ( n6078 , n6073 , n6076 );
or ( n6079 , n6075 , n6077 , n6078 );
and ( n6080 , n6071 , n6079 );
and ( n6081 , n6066 , n6079 );
or ( n6082 , n6072 , n6080 , n6081 );
and ( n6083 , n6058 , n6082 );
and ( n6084 , n6043 , n6082 );
or ( n6085 , n6059 , n6083 , n6084 );
xor ( n6086 , n5916 , n5918 );
xor ( n6087 , n6086 , n5920 );
and ( n6088 , n6085 , n6087 );
xor ( n6089 , n5925 , n5956 );
xor ( n6090 , n6089 , n5960 );
and ( n6091 , n6087 , n6090 );
and ( n6092 , n6085 , n6090 );
or ( n6093 , n6088 , n6091 , n6092 );
xor ( n6094 , n5909 , n5923 );
xor ( n6095 , n6094 , n5963 );
and ( n6096 , n6093 , n6095 );
xor ( n6097 , n5980 , n5985 );
xor ( n6098 , n6097 , n6001 );
xor ( n6099 , n5987 , n5994 );
xor ( n6100 , n6099 , n5998 );
xor ( n6101 , n6040 , n6042 );
and ( n6102 , n6100 , n6101 );
and ( n6103 , n5745 , n5640 );
xnor ( n6104 , n6052 , n6053 );
or ( n6105 , n6103 , n6104 );
and ( n6106 , n5643 , n5762 );
xnor ( n6107 , n6049 , n6050 );
or ( n6108 , n6106 , n6107 );
and ( n6109 , n6105 , n6108 );
and ( n6110 , n6101 , n6109 );
and ( n6111 , n6100 , n6109 );
or ( n6112 , n6102 , n6110 , n6111 );
and ( n6113 , n6098 , n6112 );
buf ( n6114 , n790 );
buf ( n6115 , n6114 );
and ( n6116 , n6115 , n5572 );
xnor ( n6117 , n6063 , n6064 );
or ( n6118 , n6116 , n6117 );
buf ( n6119 , n790 );
buf ( n6120 , n6119 );
and ( n6121 , n5564 , n6120 );
xnor ( n6122 , n6060 , n6061 );
or ( n6123 , n6121 , n6122 );
and ( n6124 , n6118 , n6123 );
xor ( n6125 , n6051 , n6054 );
xor ( n6126 , n6062 , n6065 );
and ( n6127 , n6125 , n6126 );
xor ( n6128 , n6068 , n6070 );
and ( n6129 , n6126 , n6128 );
and ( n6130 , n6125 , n6128 );
or ( n6131 , n6127 , n6129 , n6130 );
and ( n6132 , n6124 , n6131 );
buf ( n6133 , n791 );
buf ( n6134 , n6133 );
and ( n6135 , n6134 , n5572 );
and ( n6136 , n5936 , n5589 );
and ( n6137 , n6135 , n6136 );
and ( n6138 , n5753 , n5640 );
and ( n6139 , n6136 , n6138 );
and ( n6140 , n6135 , n6138 );
or ( n6141 , n6137 , n6139 , n6140 );
buf ( n6142 , n791 );
buf ( n6143 , n6142 );
and ( n6144 , n5564 , n6143 );
and ( n6145 , n5592 , n5927 );
and ( n6146 , n6144 , n6145 );
and ( n6147 , n5643 , n5736 );
and ( n6148 , n6145 , n6147 );
and ( n6149 , n6144 , n6147 );
or ( n6150 , n6146 , n6148 , n6149 );
and ( n6151 , n6141 , n6150 );
and ( n6152 , n6115 , n5567 );
and ( n6153 , n5992 , n5578 );
or ( n6154 , n6152 , n6153 );
and ( n6155 , n5570 , n6120 );
and ( n6156 , n5581 , n5989 );
or ( n6157 , n6155 , n6156 );
and ( n6158 , n6154 , n6157 );
and ( n6159 , n6151 , n6158 );
xor ( n6160 , n6073 , n6074 );
xor ( n6161 , n6160 , n6076 );
and ( n6162 , n6158 , n6161 );
and ( n6163 , n6151 , n6161 );
or ( n6164 , n6159 , n6162 , n6163 );
and ( n6165 , n6131 , n6164 );
and ( n6166 , n6124 , n6164 );
or ( n6167 , n6132 , n6165 , n6166 );
and ( n6168 , n6112 , n6167 );
and ( n6169 , n6098 , n6167 );
or ( n6170 , n6113 , n6168 , n6169 );
xor ( n6171 , n6004 , n6006 );
xor ( n6172 , n6171 , n6015 );
and ( n6173 , n6170 , n6172 );
xor ( n6174 , n6085 , n6087 );
xor ( n6175 , n6174 , n6090 );
and ( n6176 , n6172 , n6175 );
and ( n6177 , n6170 , n6175 );
or ( n6178 , n6173 , n6176 , n6177 );
and ( n6179 , n6095 , n6178 );
and ( n6180 , n6093 , n6178 );
or ( n6181 , n6096 , n6179 , n6180 );
xor ( n6182 , n5974 , n6021 );
xor ( n6183 , n6182 , n6024 );
and ( n6184 , n6181 , n6183 );
xor ( n6185 , n5976 , n5978 );
xor ( n6186 , n6185 , n6018 );
xor ( n6187 , n6093 , n6095 );
xor ( n6188 , n6187 , n6178 );
and ( n6189 , n6186 , n6188 );
xor ( n6190 , n6009 , n6010 );
xor ( n6191 , n6190 , n6012 );
xor ( n6192 , n6043 , n6058 );
xor ( n6193 , n6192 , n6082 );
and ( n6194 , n6191 , n6193 );
xor ( n6195 , n6046 , n6047 );
xor ( n6196 , n6195 , n6055 );
xor ( n6197 , n6066 , n6071 );
xor ( n6198 , n6197 , n6079 );
and ( n6199 , n6196 , n6198 );
xor ( n6200 , n6105 , n6108 );
xor ( n6201 , n6118 , n6123 );
and ( n6202 , n6200 , n6201 );
xnor ( n6203 , n6103 , n6104 );
xnor ( n6204 , n6106 , n6107 );
and ( n6205 , n6203 , n6204 );
and ( n6206 , n6201 , n6205 );
and ( n6207 , n6200 , n6205 );
or ( n6208 , n6202 , n6206 , n6207 );
and ( n6209 , n6198 , n6208 );
and ( n6210 , n6196 , n6208 );
or ( n6211 , n6199 , n6209 , n6210 );
and ( n6212 , n6193 , n6211 );
and ( n6213 , n6191 , n6211 );
or ( n6214 , n6194 , n6212 , n6213 );
xor ( n6215 , n6170 , n6172 );
xor ( n6216 , n6215 , n6175 );
and ( n6217 , n6214 , n6216 );
xnor ( n6218 , n6116 , n6117 );
xnor ( n6219 , n6121 , n6122 );
and ( n6220 , n6218 , n6219 );
buf ( n6221 , n5667 );
and ( n6222 , n5607 , n5871 );
and ( n6223 , n5865 , n5612 );
and ( n6224 , n6222 , n6223 );
and ( n6225 , n6221 , n6224 );
xor ( n6226 , n6141 , n6150 );
and ( n6227 , n6224 , n6226 );
and ( n6228 , n6221 , n6226 );
or ( n6229 , n6225 , n6227 , n6228 );
and ( n6230 , n6220 , n6229 );
xor ( n6231 , n6154 , n6157 );
and ( n6232 , n5865 , n5640 );
and ( n6233 , n5753 , n5676 );
or ( n6234 , n6232 , n6233 );
and ( n6235 , n5643 , n5871 );
and ( n6236 , n5667 , n5736 );
or ( n6237 , n6235 , n6236 );
and ( n6238 , n6234 , n6237 );
and ( n6239 , n6231 , n6238 );
xor ( n6240 , n6135 , n6136 );
xor ( n6241 , n6240 , n6138 );
xor ( n6242 , n6144 , n6145 );
xor ( n6243 , n6242 , n6147 );
and ( n6244 , n6241 , n6243 );
and ( n6245 , n6238 , n6244 );
and ( n6246 , n6231 , n6244 );
or ( n6247 , n6239 , n6245 , n6246 );
and ( n6248 , n6229 , n6247 );
and ( n6249 , n6220 , n6247 );
or ( n6250 , n6230 , n6248 , n6249 );
xnor ( n6251 , n6152 , n6153 );
xnor ( n6252 , n6155 , n6156 );
and ( n6253 , n6251 , n6252 );
and ( n6254 , n5745 , n5676 );
and ( n6255 , n5667 , n5762 );
and ( n6256 , n6254 , n6255 );
xor ( n6257 , n6222 , n6223 );
and ( n6258 , n6255 , n6257 );
and ( n6259 , n6254 , n6257 );
or ( n6260 , n6256 , n6258 , n6259 );
and ( n6261 , n6253 , n6260 );
and ( n6262 , n5570 , n6143 );
and ( n6263 , n6134 , n5567 );
and ( n6264 , n6262 , n6263 );
and ( n6265 , n5581 , n6120 );
and ( n6266 , n6115 , n5578 );
and ( n6267 , n6265 , n6266 );
and ( n6268 , n6264 , n6267 );
and ( n6269 , n5592 , n5989 );
and ( n6270 , n5992 , n5589 );
and ( n6271 , n6269 , n6270 );
and ( n6272 , n6267 , n6271 );
and ( n6273 , n6264 , n6271 );
or ( n6274 , n6268 , n6272 , n6273 );
and ( n6275 , n6260 , n6274 );
and ( n6276 , n6253 , n6274 );
or ( n6277 , n6261 , n6275 , n6276 );
xor ( n6278 , n6125 , n6126 );
xor ( n6279 , n6278 , n6128 );
and ( n6280 , n6277 , n6279 );
xor ( n6281 , n6151 , n6158 );
xor ( n6282 , n6281 , n6161 );
and ( n6283 , n6279 , n6282 );
and ( n6284 , n6277 , n6282 );
or ( n6285 , n6280 , n6283 , n6284 );
and ( n6286 , n6250 , n6285 );
xor ( n6287 , n6100 , n6101 );
xor ( n6288 , n6287 , n6109 );
and ( n6289 , n6285 , n6288 );
and ( n6290 , n6250 , n6288 );
or ( n6291 , n6286 , n6289 , n6290 );
xor ( n6292 , n6098 , n6112 );
xor ( n6293 , n6292 , n6167 );
and ( n6294 , n6291 , n6293 );
xor ( n6295 , n6124 , n6131 );
xor ( n6296 , n6295 , n6164 );
xor ( n6297 , n6203 , n6204 );
xor ( n6298 , n6218 , n6219 );
and ( n6299 , n6297 , n6298 );
and ( n6300 , n5607 , n5927 );
and ( n6301 , n5936 , n5612 );
and ( n6302 , n6300 , n6301 );
xor ( n6303 , n6234 , n6237 );
and ( n6304 , n6302 , n6303 );
xor ( n6305 , n6241 , n6243 );
and ( n6306 , n6303 , n6305 );
and ( n6307 , n6302 , n6305 );
or ( n6308 , n6304 , n6306 , n6307 );
and ( n6309 , n6298 , n6308 );
and ( n6310 , n6297 , n6308 );
or ( n6311 , n6299 , n6309 , n6310 );
xor ( n6312 , n6251 , n6252 );
buf ( n6313 , n793 );
buf ( n6314 , n6313 );
and ( n6315 , n6314 , n5572 );
buf ( n6316 , n792 );
buf ( n6317 , n6316 );
and ( n6318 , n6317 , n5567 );
and ( n6319 , n6315 , n6318 );
and ( n6320 , n5936 , n5640 );
and ( n6321 , n6318 , n6320 );
and ( n6322 , n6315 , n6320 );
or ( n6323 , n6319 , n6321 , n6322 );
and ( n6324 , n5745 , n5736 );
and ( n6325 , n5753 , n5762 );
and ( n6326 , n6324 , n6325 );
and ( n6327 , n6323 , n6326 );
buf ( n6328 , n792 );
buf ( n6329 , n6328 );
and ( n6330 , n5564 , n6329 );
and ( n6331 , n6326 , n6330 );
and ( n6332 , n6323 , n6330 );
or ( n6333 , n6327 , n6331 , n6332 );
and ( n6334 , n6312 , n6333 );
xnor ( n6335 , n6232 , n6233 );
xnor ( n6336 , n6235 , n6236 );
and ( n6337 , n6335 , n6336 );
and ( n6338 , n6333 , n6337 );
and ( n6339 , n6312 , n6337 );
or ( n6340 , n6334 , n6338 , n6339 );
and ( n6341 , n6317 , n5572 );
buf ( n6342 , n5745 );
and ( n6343 , n6341 , n6342 );
xor ( n6344 , n6262 , n6263 );
and ( n6345 , n6342 , n6344 );
and ( n6346 , n6341 , n6344 );
or ( n6347 , n6343 , n6345 , n6346 );
xor ( n6348 , n6265 , n6266 );
xor ( n6349 , n6269 , n6270 );
and ( n6350 , n6348 , n6349 );
xor ( n6351 , n6300 , n6301 );
and ( n6352 , n6349 , n6351 );
and ( n6353 , n6348 , n6351 );
or ( n6354 , n6350 , n6352 , n6353 );
and ( n6355 , n6347 , n6354 );
buf ( n6356 , n793 );
buf ( n6357 , n6356 );
and ( n6358 , n5564 , n6357 );
and ( n6359 , n5570 , n6329 );
and ( n6360 , n6358 , n6359 );
and ( n6361 , n5643 , n5927 );
and ( n6362 , n6359 , n6361 );
and ( n6363 , n6358 , n6361 );
or ( n6364 , n6360 , n6362 , n6363 );
and ( n6365 , n5581 , n6143 );
and ( n6366 , n6134 , n5578 );
and ( n6367 , n6365 , n6366 );
and ( n6368 , n6364 , n6367 );
and ( n6369 , n5592 , n6120 );
and ( n6370 , n6115 , n5589 );
and ( n6371 , n6369 , n6370 );
and ( n6372 , n6367 , n6371 );
and ( n6373 , n6364 , n6371 );
or ( n6374 , n6368 , n6372 , n6373 );
and ( n6375 , n6354 , n6374 );
and ( n6376 , n6347 , n6374 );
or ( n6377 , n6355 , n6375 , n6376 );
and ( n6378 , n6340 , n6377 );
xor ( n6379 , n6221 , n6224 );
xor ( n6380 , n6379 , n6226 );
and ( n6381 , n6377 , n6380 );
and ( n6382 , n6340 , n6380 );
or ( n6383 , n6378 , n6381 , n6382 );
and ( n6384 , n6311 , n6383 );
xor ( n6385 , n6200 , n6201 );
xor ( n6386 , n6385 , n6205 );
and ( n6387 , n6383 , n6386 );
and ( n6388 , n6311 , n6386 );
or ( n6389 , n6384 , n6387 , n6388 );
and ( n6390 , n6296 , n6389 );
xor ( n6391 , n6196 , n6198 );
xor ( n6392 , n6391 , n6208 );
and ( n6393 , n6389 , n6392 );
and ( n6394 , n6296 , n6392 );
or ( n6395 , n6390 , n6393 , n6394 );
and ( n6396 , n6293 , n6395 );
and ( n6397 , n6291 , n6395 );
or ( n6398 , n6294 , n6396 , n6397 );
and ( n6399 , n6216 , n6398 );
and ( n6400 , n6214 , n6398 );
or ( n6401 , n6217 , n6399 , n6400 );
and ( n6402 , n6188 , n6401 );
and ( n6403 , n6186 , n6401 );
or ( n6404 , n6189 , n6402 , n6403 );
and ( n6405 , n6183 , n6404 );
and ( n6406 , n6181 , n6404 );
or ( n6407 , n6184 , n6405 , n6406 );
or ( n6408 , n6038 , n6407 );
or ( n6409 , n6036 , n6408 );
and ( n6410 , n6033 , n6409 );
and ( n6411 , n5796 , n6409 );
or ( n6412 , n6034 , n6410 , n6411 );
and ( n6413 , n5793 , n6412 );
and ( n6414 , n5704 , n6412 );
or ( n6415 , n5794 , n6413 , n6414 );
or ( n6416 , n5702 , n6415 );
and ( n6417 , n5699 , n6416 );
and ( n6418 , n5605 , n6416 );
or ( n6419 , n5700 , n6417 , n6418 );
xnor ( n6420 , n5603 , n6419 );
xor ( n6421 , n5605 , n5699 );
xor ( n6422 , n6421 , n6416 );
not ( n6423 , n6422 );
xnor ( n6424 , n5702 , n6415 );
xor ( n6425 , n5704 , n5793 );
xor ( n6426 , n6425 , n6412 );
not ( n6427 , n6426 );
xor ( n6428 , n5796 , n6033 );
xor ( n6429 , n6428 , n6409 );
xnor ( n6430 , n6036 , n6408 );
xnor ( n6431 , n6038 , n6407 );
xor ( n6432 , n6181 , n6183 );
xor ( n6433 , n6432 , n6404 );
not ( n6434 , n6433 );
xor ( n6435 , n6186 , n6188 );
xor ( n6436 , n6435 , n6401 );
xor ( n6437 , n6191 , n6193 );
xor ( n6438 , n6437 , n6211 );
xor ( n6439 , n6250 , n6285 );
xor ( n6440 , n6439 , n6288 );
xor ( n6441 , n6220 , n6229 );
xor ( n6442 , n6441 , n6247 );
xor ( n6443 , n6277 , n6279 );
xor ( n6444 , n6443 , n6282 );
and ( n6445 , n6442 , n6444 );
xor ( n6446 , n6231 , n6238 );
xor ( n6447 , n6446 , n6244 );
xor ( n6448 , n6253 , n6260 );
xor ( n6449 , n6448 , n6274 );
and ( n6450 , n6447 , n6449 );
xor ( n6451 , n6254 , n6255 );
xor ( n6452 , n6451 , n6257 );
xor ( n6453 , n6264 , n6267 );
xor ( n6454 , n6453 , n6271 );
and ( n6455 , n6452 , n6454 );
and ( n6456 , n5607 , n5989 );
and ( n6457 , n5992 , n5612 );
and ( n6458 , n6456 , n6457 );
and ( n6459 , n5667 , n5871 );
and ( n6460 , n5865 , n5676 );
and ( n6461 , n6459 , n6460 );
and ( n6462 , n6458 , n6461 );
xor ( n6463 , n6323 , n6326 );
xor ( n6464 , n6463 , n6330 );
and ( n6465 , n6461 , n6464 );
and ( n6466 , n6458 , n6464 );
or ( n6467 , n6462 , n6465 , n6466 );
and ( n6468 , n6454 , n6467 );
and ( n6469 , n6452 , n6467 );
or ( n6470 , n6455 , n6468 , n6469 );
and ( n6471 , n6449 , n6470 );
and ( n6472 , n6447 , n6470 );
or ( n6473 , n6450 , n6471 , n6472 );
and ( n6474 , n6444 , n6473 );
and ( n6475 , n6442 , n6473 );
or ( n6476 , n6445 , n6474 , n6475 );
and ( n6477 , n6440 , n6476 );
xor ( n6478 , n6296 , n6389 );
xor ( n6479 , n6478 , n6392 );
and ( n6480 , n6476 , n6479 );
and ( n6481 , n6440 , n6479 );
or ( n6482 , n6477 , n6480 , n6481 );
and ( n6483 , n6438 , n6482 );
xor ( n6484 , n6291 , n6293 );
xor ( n6485 , n6484 , n6395 );
and ( n6486 , n6482 , n6485 );
and ( n6487 , n6438 , n6485 );
or ( n6488 , n6483 , n6486 , n6487 );
xor ( n6489 , n6214 , n6216 );
xor ( n6490 , n6489 , n6398 );
and ( n6491 , n6488 , n6490 );
xor ( n6492 , n6438 , n6482 );
xor ( n6493 , n6492 , n6485 );
xor ( n6494 , n6335 , n6336 );
and ( n6495 , n6134 , n5589 );
and ( n6496 , n6115 , n5612 );
and ( n6497 , n6495 , n6496 );
and ( n6498 , n5992 , n5640 );
and ( n6499 , n6496 , n6498 );
and ( n6500 , n6495 , n6498 );
or ( n6501 , n6497 , n6499 , n6500 );
and ( n6502 , n5592 , n6143 );
and ( n6503 , n5607 , n6120 );
and ( n6504 , n6502 , n6503 );
and ( n6505 , n5643 , n5989 );
and ( n6506 , n6503 , n6505 );
and ( n6507 , n6502 , n6505 );
or ( n6508 , n6504 , n6506 , n6507 );
and ( n6509 , n6501 , n6508 );
and ( n6510 , n6494 , n6509 );
and ( n6511 , n6314 , n5567 );
and ( n6512 , n6317 , n5578 );
or ( n6513 , n6511 , n6512 );
and ( n6514 , n5570 , n6357 );
and ( n6515 , n5581 , n6329 );
or ( n6516 , n6514 , n6515 );
and ( n6517 , n6513 , n6516 );
and ( n6518 , n6509 , n6517 );
and ( n6519 , n6494 , n6517 );
or ( n6520 , n6510 , n6518 , n6519 );
and ( n6521 , n5936 , n5676 );
not ( n6522 , n6521 );
and ( n6523 , n5865 , n5762 );
and ( n6524 , n6522 , n6523 );
and ( n6525 , n5667 , n5927 );
not ( n6526 , n6525 );
and ( n6527 , n5745 , n5871 );
and ( n6528 , n6526 , n6527 );
and ( n6529 , n6524 , n6528 );
buf ( n6530 , n6521 );
buf ( n6531 , n6525 );
and ( n6532 , n6530 , n6531 );
and ( n6533 , n6529 , n6532 );
xor ( n6534 , n6315 , n6318 );
xor ( n6535 , n6534 , n6320 );
xor ( n6536 , n6358 , n6359 );
xor ( n6537 , n6536 , n6361 );
and ( n6538 , n6535 , n6537 );
and ( n6539 , n6532 , n6538 );
and ( n6540 , n6529 , n6538 );
or ( n6541 , n6533 , n6539 , n6540 );
and ( n6542 , n6520 , n6541 );
xor ( n6543 , n6365 , n6366 );
xor ( n6544 , n6369 , n6370 );
and ( n6545 , n6543 , n6544 );
xor ( n6546 , n6456 , n6457 );
and ( n6547 , n6544 , n6546 );
and ( n6548 , n6543 , n6546 );
or ( n6549 , n6545 , n6547 , n6548 );
xor ( n6550 , n6341 , n6342 );
xor ( n6551 , n6550 , n6344 );
and ( n6552 , n6549 , n6551 );
xor ( n6553 , n6348 , n6349 );
xor ( n6554 , n6553 , n6351 );
and ( n6555 , n6551 , n6554 );
and ( n6556 , n6549 , n6554 );
or ( n6557 , n6552 , n6555 , n6556 );
and ( n6558 , n6541 , n6557 );
and ( n6559 , n6520 , n6557 );
or ( n6560 , n6542 , n6558 , n6559 );
xor ( n6561 , n6302 , n6303 );
xor ( n6562 , n6561 , n6305 );
xor ( n6563 , n6312 , n6333 );
xor ( n6564 , n6563 , n6337 );
and ( n6565 , n6562 , n6564 );
xor ( n6566 , n6347 , n6354 );
xor ( n6567 , n6566 , n6374 );
and ( n6568 , n6564 , n6567 );
and ( n6569 , n6562 , n6567 );
or ( n6570 , n6565 , n6568 , n6569 );
and ( n6571 , n6560 , n6570 );
xor ( n6572 , n6297 , n6298 );
xor ( n6573 , n6572 , n6308 );
and ( n6574 , n6570 , n6573 );
and ( n6575 , n6560 , n6573 );
or ( n6576 , n6571 , n6574 , n6575 );
xor ( n6577 , n6311 , n6383 );
xor ( n6578 , n6577 , n6386 );
and ( n6579 , n6576 , n6578 );
xor ( n6580 , n6340 , n6377 );
xor ( n6581 , n6580 , n6380 );
xor ( n6582 , n6364 , n6367 );
xor ( n6583 , n6582 , n6371 );
xnor ( n6584 , n6514 , n6515 );
not ( n6585 , n6584 );
xor ( n6586 , n6526 , n6527 );
and ( n6587 , n6585 , n6586 );
xnor ( n6588 , n6511 , n6512 );
not ( n6589 , n6588 );
xor ( n6590 , n6522 , n6523 );
and ( n6591 , n6589 , n6590 );
and ( n6592 , n6587 , n6591 );
and ( n6593 , n6583 , n6592 );
buf ( n6594 , n6584 );
buf ( n6595 , n6588 );
and ( n6596 , n6594 , n6595 );
and ( n6597 , n6592 , n6596 );
and ( n6598 , n6583 , n6596 );
or ( n6599 , n6593 , n6597 , n6598 );
xor ( n6600 , n6459 , n6460 );
xor ( n6601 , n6324 , n6325 );
and ( n6602 , n6600 , n6601 );
xor ( n6603 , n6501 , n6508 );
and ( n6604 , n6601 , n6603 );
and ( n6605 , n6600 , n6603 );
or ( n6606 , n6602 , n6604 , n6605 );
xor ( n6607 , n6513 , n6516 );
xor ( n6608 , n6524 , n6528 );
and ( n6609 , n6607 , n6608 );
xor ( n6610 , n6530 , n6531 );
and ( n6611 , n6608 , n6610 );
and ( n6612 , n6607 , n6610 );
or ( n6613 , n6609 , n6611 , n6612 );
and ( n6614 , n6606 , n6613 );
xor ( n6615 , n6535 , n6537 );
and ( n6616 , n6317 , n5589 );
and ( n6617 , n6134 , n5612 );
and ( n6618 , n6616 , n6617 );
and ( n6619 , n5936 , n5762 );
and ( n6620 , n6617 , n6619 );
and ( n6621 , n6616 , n6619 );
or ( n6622 , n6618 , n6620 , n6621 );
and ( n6623 , n6314 , n5578 );
and ( n6624 , n6115 , n5640 );
and ( n6625 , n6623 , n6624 );
and ( n6626 , n5992 , n5676 );
and ( n6627 , n6624 , n6626 );
and ( n6628 , n6623 , n6626 );
or ( n6629 , n6625 , n6627 , n6628 );
and ( n6630 , n6622 , n6629 );
and ( n6631 , n5753 , n5871 );
and ( n6632 , n5865 , n5736 );
and ( n6633 , n6631 , n6632 );
and ( n6634 , n6629 , n6633 );
and ( n6635 , n6622 , n6633 );
or ( n6636 , n6630 , n6634 , n6635 );
and ( n6637 , n6615 , n6636 );
buf ( n6638 , n5753 );
and ( n6639 , n5592 , n6329 );
and ( n6640 , n5607 , n6143 );
and ( n6641 , n6639 , n6640 );
and ( n6642 , n5745 , n5927 );
and ( n6643 , n6640 , n6642 );
and ( n6644 , n6639 , n6642 );
or ( n6645 , n6641 , n6643 , n6644 );
and ( n6646 , n6638 , n6645 );
and ( n6647 , n5581 , n6357 );
and ( n6648 , n5643 , n6120 );
and ( n6649 , n6647 , n6648 );
and ( n6650 , n5667 , n5989 );
and ( n6651 , n6648 , n6650 );
and ( n6652 , n6647 , n6650 );
or ( n6653 , n6649 , n6651 , n6652 );
and ( n6654 , n6645 , n6653 );
and ( n6655 , n6638 , n6653 );
or ( n6656 , n6646 , n6654 , n6655 );
and ( n6657 , n6636 , n6656 );
and ( n6658 , n6615 , n6656 );
or ( n6659 , n6637 , n6657 , n6658 );
and ( n6660 , n6613 , n6659 );
and ( n6661 , n6606 , n6659 );
or ( n6662 , n6614 , n6660 , n6661 );
and ( n6663 , n6599 , n6662 );
xor ( n6664 , n6458 , n6461 );
xor ( n6665 , n6664 , n6464 );
xor ( n6666 , n6494 , n6509 );
xor ( n6667 , n6666 , n6517 );
and ( n6668 , n6665 , n6667 );
xor ( n6669 , n6529 , n6532 );
xor ( n6670 , n6669 , n6538 );
and ( n6671 , n6667 , n6670 );
and ( n6672 , n6665 , n6670 );
or ( n6673 , n6668 , n6671 , n6672 );
and ( n6674 , n6662 , n6673 );
and ( n6675 , n6599 , n6673 );
or ( n6676 , n6663 , n6674 , n6675 );
and ( n6677 , n6581 , n6676 );
xor ( n6678 , n6452 , n6454 );
xor ( n6679 , n6678 , n6467 );
xor ( n6680 , n6520 , n6541 );
xor ( n6681 , n6680 , n6557 );
and ( n6682 , n6679 , n6681 );
xor ( n6683 , n6562 , n6564 );
xor ( n6684 , n6683 , n6567 );
and ( n6685 , n6681 , n6684 );
and ( n6686 , n6679 , n6684 );
or ( n6687 , n6682 , n6685 , n6686 );
and ( n6688 , n6676 , n6687 );
and ( n6689 , n6581 , n6687 );
or ( n6690 , n6677 , n6688 , n6689 );
and ( n6691 , n6578 , n6690 );
and ( n6692 , n6576 , n6690 );
or ( n6693 , n6579 , n6691 , n6692 );
xor ( n6694 , n6440 , n6476 );
xor ( n6695 , n6694 , n6479 );
and ( n6696 , n6693 , n6695 );
xor ( n6697 , n6442 , n6444 );
xor ( n6698 , n6697 , n6473 );
xor ( n6699 , n6447 , n6449 );
xor ( n6700 , n6699 , n6470 );
xor ( n6701 , n6560 , n6570 );
xor ( n6702 , n6701 , n6573 );
and ( n6703 , n6700 , n6702 );
xor ( n6704 , n6549 , n6551 );
xor ( n6705 , n6704 , n6554 );
xor ( n6706 , n6502 , n6503 );
xor ( n6707 , n6706 , n6505 );
not ( n6708 , n6707 );
xor ( n6709 , n6589 , n6590 );
and ( n6710 , n6708 , n6709 );
xor ( n6711 , n6495 , n6496 );
xor ( n6712 , n6711 , n6498 );
not ( n6713 , n6712 );
xor ( n6714 , n6585 , n6586 );
and ( n6715 , n6713 , n6714 );
and ( n6716 , n6710 , n6715 );
and ( n6717 , n6705 , n6716 );
buf ( n6718 , n6707 );
buf ( n6719 , n6712 );
and ( n6720 , n6718 , n6719 );
and ( n6721 , n6716 , n6720 );
and ( n6722 , n6705 , n6720 );
or ( n6723 , n6717 , n6721 , n6722 );
xor ( n6724 , n6543 , n6544 );
xor ( n6725 , n6724 , n6546 );
xor ( n6726 , n6587 , n6591 );
and ( n6727 , n6725 , n6726 );
xor ( n6728 , n6594 , n6595 );
and ( n6729 , n6726 , n6728 );
and ( n6730 , n6725 , n6728 );
or ( n6731 , n6727 , n6729 , n6730 );
xor ( n6732 , n6616 , n6617 );
xor ( n6733 , n6732 , n6619 );
xor ( n6734 , n6623 , n6624 );
xor ( n6735 , n6734 , n6626 );
or ( n6736 , n6733 , n6735 );
and ( n6737 , n6317 , n5612 );
and ( n6738 , n6134 , n5640 );
and ( n6739 , n6737 , n6738 );
and ( n6740 , n6115 , n5676 );
and ( n6741 , n6738 , n6740 );
and ( n6742 , n6737 , n6740 );
or ( n6743 , n6739 , n6741 , n6742 );
and ( n6744 , n5607 , n6329 );
and ( n6745 , n5643 , n6143 );
and ( n6746 , n6744 , n6745 );
and ( n6747 , n5667 , n6120 );
and ( n6748 , n6745 , n6747 );
and ( n6749 , n6744 , n6747 );
or ( n6750 , n6746 , n6748 , n6749 );
and ( n6751 , n6743 , n6750 );
and ( n6752 , n6736 , n6751 );
and ( n6753 , n5992 , n5762 );
and ( n6754 , n5936 , n5736 );
and ( n6755 , n6753 , n6754 );
and ( n6756 , n5745 , n5989 );
and ( n6757 , n5753 , n5927 );
and ( n6758 , n6756 , n6757 );
and ( n6759 , n6755 , n6758 );
and ( n6760 , n6751 , n6759 );
and ( n6761 , n6736 , n6759 );
or ( n6762 , n6752 , n6760 , n6761 );
xor ( n6763 , n6600 , n6601 );
xor ( n6764 , n6763 , n6603 );
and ( n6765 , n6762 , n6764 );
xor ( n6766 , n6607 , n6608 );
xor ( n6767 , n6766 , n6610 );
and ( n6768 , n6764 , n6767 );
and ( n6769 , n6762 , n6767 );
or ( n6770 , n6765 , n6768 , n6769 );
and ( n6771 , n6731 , n6770 );
xor ( n6772 , n6583 , n6592 );
xor ( n6773 , n6772 , n6596 );
and ( n6774 , n6770 , n6773 );
and ( n6775 , n6731 , n6773 );
or ( n6776 , n6771 , n6774 , n6775 );
and ( n6777 , n6723 , n6776 );
xor ( n6778 , n6599 , n6662 );
xor ( n6779 , n6778 , n6673 );
and ( n6780 , n6776 , n6779 );
and ( n6781 , n6723 , n6779 );
or ( n6782 , n6777 , n6780 , n6781 );
and ( n6783 , n6702 , n6782 );
and ( n6784 , n6700 , n6782 );
or ( n6785 , n6703 , n6783 , n6784 );
and ( n6786 , n6698 , n6785 );
xor ( n6787 , n6576 , n6578 );
xor ( n6788 , n6787 , n6690 );
and ( n6789 , n6785 , n6788 );
and ( n6790 , n6698 , n6788 );
or ( n6791 , n6786 , n6789 , n6790 );
and ( n6792 , n6695 , n6791 );
and ( n6793 , n6693 , n6791 );
or ( n6794 , n6696 , n6792 , n6793 );
and ( n6795 , n6493 , n6794 );
xor ( n6796 , n6693 , n6695 );
xor ( n6797 , n6796 , n6791 );
xor ( n6798 , n6581 , n6676 );
xor ( n6799 , n6798 , n6687 );
xor ( n6800 , n6679 , n6681 );
xor ( n6801 , n6800 , n6684 );
xor ( n6802 , n6606 , n6613 );
xor ( n6803 , n6802 , n6659 );
xor ( n6804 , n6665 , n6667 );
xor ( n6805 , n6804 , n6670 );
and ( n6806 , n6803 , n6805 );
xor ( n6807 , n6615 , n6636 );
xor ( n6808 , n6807 , n6656 );
xor ( n6809 , n6710 , n6715 );
and ( n6810 , n6808 , n6809 );
xor ( n6811 , n6718 , n6719 );
and ( n6812 , n6809 , n6811 );
and ( n6813 , n6808 , n6811 );
or ( n6814 , n6810 , n6812 , n6813 );
and ( n6815 , n6805 , n6814 );
and ( n6816 , n6803 , n6814 );
or ( n6817 , n6806 , n6815 , n6816 );
and ( n6818 , n6801 , n6817 );
xor ( n6819 , n6756 , n6757 );
and ( n6820 , n5865 , n5927 );
and ( n6821 , n5936 , n5871 );
and ( n6822 , n6820 , n6821 );
and ( n6823 , n6819 , n6822 );
and ( n6824 , n5592 , n6357 );
and ( n6825 , n6822 , n6824 );
and ( n6826 , n6819 , n6824 );
or ( n6827 , n6823 , n6825 , n6826 );
xor ( n6828 , n6639 , n6640 );
xor ( n6829 , n6828 , n6642 );
and ( n6830 , n6827 , n6829 );
xor ( n6831 , n6647 , n6648 );
xor ( n6832 , n6831 , n6650 );
and ( n6833 , n6829 , n6832 );
and ( n6834 , n6827 , n6832 );
or ( n6835 , n6830 , n6833 , n6834 );
xor ( n6836 , n6622 , n6629 );
xor ( n6837 , n6836 , n6633 );
and ( n6838 , n6835 , n6837 );
xor ( n6839 , n6708 , n6709 );
xor ( n6840 , n6713 , n6714 );
and ( n6841 , n6839 , n6840 );
and ( n6842 , n6838 , n6841 );
xor ( n6843 , n6638 , n6645 );
xor ( n6844 , n6843 , n6653 );
xor ( n6845 , n6631 , n6632 );
xnor ( n6846 , n6733 , n6735 );
and ( n6847 , n6845 , n6846 );
xor ( n6848 , n6743 , n6750 );
and ( n6849 , n6846 , n6848 );
and ( n6850 , n6845 , n6848 );
or ( n6851 , n6847 , n6849 , n6850 );
and ( n6852 , n6844 , n6851 );
xor ( n6853 , n6736 , n6751 );
xor ( n6854 , n6853 , n6759 );
and ( n6855 , n6851 , n6854 );
and ( n6856 , n6844 , n6854 );
or ( n6857 , n6852 , n6855 , n6856 );
and ( n6858 , n6841 , n6857 );
and ( n6859 , n6838 , n6857 );
or ( n6860 , n6842 , n6858 , n6859 );
xor ( n6861 , n6705 , n6716 );
xor ( n6862 , n6861 , n6720 );
and ( n6863 , n6860 , n6862 );
xor ( n6864 , n6731 , n6770 );
xor ( n6865 , n6864 , n6773 );
and ( n6866 , n6862 , n6865 );
and ( n6867 , n6860 , n6865 );
or ( n6868 , n6863 , n6866 , n6867 );
and ( n6869 , n6817 , n6868 );
and ( n6870 , n6801 , n6868 );
or ( n6871 , n6818 , n6869 , n6870 );
and ( n6872 , n6799 , n6871 );
xor ( n6873 , n6700 , n6702 );
xor ( n6874 , n6873 , n6782 );
and ( n6875 , n6871 , n6874 );
and ( n6876 , n6799 , n6874 );
or ( n6877 , n6872 , n6875 , n6876 );
xor ( n6878 , n6698 , n6785 );
xor ( n6879 , n6878 , n6788 );
and ( n6880 , n6877 , n6879 );
xor ( n6881 , n6723 , n6776 );
xor ( n6882 , n6881 , n6779 );
xor ( n6883 , n6725 , n6726 );
xor ( n6884 , n6883 , n6728 );
xor ( n6885 , n6762 , n6764 );
xor ( n6886 , n6885 , n6767 );
and ( n6887 , n6884 , n6886 );
xor ( n6888 , n6835 , n6837 );
xor ( n6889 , n6839 , n6840 );
and ( n6890 , n6888 , n6889 );
and ( n6891 , n5667 , n6143 );
and ( n6892 , n5745 , n6120 );
and ( n6893 , n6891 , n6892 );
and ( n6894 , n5753 , n5989 );
and ( n6895 , n6892 , n6894 );
and ( n6896 , n6891 , n6894 );
or ( n6897 , n6893 , n6895 , n6896 );
and ( n6898 , n6115 , n5736 );
and ( n6899 , n5992 , n5871 );
and ( n6900 , n6898 , n6899 );
and ( n6901 , n5607 , n6357 );
and ( n6902 , n6900 , n6901 );
and ( n6903 , n5643 , n6329 );
and ( n6904 , n6901 , n6903 );
and ( n6905 , n6900 , n6903 );
or ( n6906 , n6902 , n6904 , n6905 );
and ( n6907 , n6897 , n6906 );
xor ( n6908 , n6737 , n6738 );
xor ( n6909 , n6908 , n6740 );
and ( n6910 , n6906 , n6909 );
and ( n6911 , n6897 , n6909 );
or ( n6912 , n6907 , n6910 , n6911 );
and ( n6913 , n6134 , n5676 );
and ( n6914 , n6115 , n5762 );
and ( n6915 , n6913 , n6914 );
and ( n6916 , n5992 , n5736 );
and ( n6917 , n6914 , n6916 );
and ( n6918 , n6913 , n6916 );
or ( n6919 , n6915 , n6917 , n6918 );
and ( n6920 , n5753 , n6120 );
and ( n6921 , n5865 , n5989 );
and ( n6922 , n6920 , n6921 );
and ( n6923 , n6314 , n5612 );
and ( n6924 , n6922 , n6923 );
and ( n6925 , n6317 , n5640 );
and ( n6926 , n6923 , n6925 );
and ( n6927 , n6922 , n6925 );
or ( n6928 , n6924 , n6926 , n6927 );
and ( n6929 , n6919 , n6928 );
xor ( n6930 , n6744 , n6745 );
xor ( n6931 , n6930 , n6747 );
and ( n6932 , n6928 , n6931 );
and ( n6933 , n6919 , n6931 );
or ( n6934 , n6929 , n6932 , n6933 );
and ( n6935 , n6912 , n6934 );
and ( n6936 , n6889 , n6935 );
and ( n6937 , n6888 , n6935 );
or ( n6938 , n6890 , n6936 , n6937 );
and ( n6939 , n6886 , n6938 );
and ( n6940 , n6884 , n6938 );
or ( n6941 , n6887 , n6939 , n6940 );
xor ( n6942 , n6803 , n6805 );
xor ( n6943 , n6942 , n6814 );
and ( n6944 , n6941 , n6943 );
xor ( n6945 , n6860 , n6862 );
xor ( n6946 , n6945 , n6865 );
and ( n6947 , n6943 , n6946 );
and ( n6948 , n6941 , n6946 );
or ( n6949 , n6944 , n6947 , n6948 );
and ( n6950 , n6882 , n6949 );
xor ( n6951 , n6801 , n6817 );
xor ( n6952 , n6951 , n6868 );
and ( n6953 , n6949 , n6952 );
and ( n6954 , n6882 , n6952 );
or ( n6955 , n6950 , n6953 , n6954 );
xor ( n6956 , n6799 , n6871 );
xor ( n6957 , n6956 , n6874 );
and ( n6958 , n6955 , n6957 );
xor ( n6959 , n6882 , n6949 );
xor ( n6960 , n6959 , n6952 );
xor ( n6961 , n6808 , n6809 );
xor ( n6962 , n6961 , n6811 );
xor ( n6963 , n6838 , n6841 );
xor ( n6964 , n6963 , n6857 );
and ( n6965 , n6962 , n6964 );
xor ( n6966 , n6755 , n6758 );
and ( n6967 , n6314 , n5589 );
buf ( n6968 , n5865 );
and ( n6969 , n6967 , n6968 );
xor ( n6970 , n6753 , n6754 );
and ( n6971 , n6968 , n6970 );
and ( n6972 , n6967 , n6970 );
or ( n6973 , n6969 , n6971 , n6972 );
and ( n6974 , n6966 , n6973 );
xor ( n6975 , n6827 , n6829 );
xor ( n6976 , n6975 , n6832 );
and ( n6977 , n6973 , n6976 );
and ( n6978 , n6966 , n6976 );
or ( n6979 , n6974 , n6977 , n6978 );
xor ( n6980 , n6844 , n6851 );
xor ( n6981 , n6980 , n6854 );
and ( n6982 , n6979 , n6981 );
xor ( n6983 , n6819 , n6822 );
xor ( n6984 , n6983 , n6824 );
and ( n6985 , n6314 , n5640 );
and ( n6986 , n6317 , n5676 );
and ( n6987 , n6985 , n6986 );
and ( n6988 , n6134 , n5762 );
and ( n6989 , n6986 , n6988 );
and ( n6990 , n6985 , n6988 );
or ( n6991 , n6987 , n6989 , n6990 );
and ( n6992 , n5643 , n6357 );
and ( n6993 , n5667 , n6329 );
and ( n6994 , n6992 , n6993 );
and ( n6995 , n5745 , n6143 );
and ( n6996 , n6993 , n6995 );
and ( n6997 , n6992 , n6995 );
or ( n6998 , n6994 , n6996 , n6997 );
and ( n6999 , n6991 , n6998 );
and ( n7000 , n6984 , n6999 );
xor ( n7001 , n6913 , n6914 );
xor ( n7002 , n7001 , n6916 );
xor ( n7003 , n6891 , n6892 );
xor ( n7004 , n7003 , n6894 );
and ( n7005 , n7002 , n7004 );
and ( n7006 , n6999 , n7005 );
and ( n7007 , n6984 , n7005 );
or ( n7008 , n7000 , n7006 , n7007 );
xor ( n7009 , n6845 , n6846 );
xor ( n7010 , n7009 , n6848 );
and ( n7011 , n7008 , n7010 );
xor ( n7012 , n6912 , n6934 );
and ( n7013 , n7010 , n7012 );
and ( n7014 , n7008 , n7012 );
or ( n7015 , n7011 , n7013 , n7014 );
and ( n7016 , n6981 , n7015 );
and ( n7017 , n6979 , n7015 );
or ( n7018 , n6982 , n7016 , n7017 );
and ( n7019 , n6964 , n7018 );
and ( n7020 , n6962 , n7018 );
or ( n7021 , n6965 , n7019 , n7020 );
xor ( n7022 , n6941 , n6943 );
xor ( n7023 , n7022 , n6946 );
and ( n7024 , n7021 , n7023 );
xor ( n7025 , n6884 , n6886 );
xor ( n7026 , n7025 , n6938 );
xor ( n7027 , n6897 , n6906 );
xor ( n7028 , n7027 , n6909 );
xor ( n7029 , n6919 , n6928 );
xor ( n7030 , n7029 , n6931 );
and ( n7031 , n7028 , n7030 );
xor ( n7032 , n6967 , n6968 );
xor ( n7033 , n7032 , n6970 );
xor ( n7034 , n6920 , n6921 );
and ( n7035 , n6317 , n5762 );
and ( n7036 , n6134 , n5736 );
and ( n7037 , n7035 , n7036 );
and ( n7038 , n6115 , n5871 );
and ( n7039 , n7036 , n7038 );
and ( n7040 , n7035 , n7038 );
or ( n7041 , n7037 , n7039 , n7040 );
and ( n7042 , n7034 , n7041 );
and ( n7043 , n5936 , n5989 );
and ( n7044 , n5992 , n5927 );
and ( n7045 , n7043 , n7044 );
and ( n7046 , n7041 , n7045 );
and ( n7047 , n7034 , n7045 );
or ( n7048 , n7042 , n7046 , n7047 );
xor ( n7049 , n6922 , n6923 );
xor ( n7050 , n7049 , n6925 );
and ( n7051 , n7048 , n7050 );
and ( n7052 , n7033 , n7051 );
xor ( n7053 , n6820 , n6821 );
xor ( n7054 , n6900 , n6901 );
xor ( n7055 , n7054 , n6903 );
and ( n7056 , n7053 , n7055 );
xor ( n7057 , n6991 , n6998 );
and ( n7058 , n7055 , n7057 );
and ( n7059 , n7053 , n7057 );
or ( n7060 , n7056 , n7058 , n7059 );
and ( n7061 , n7051 , n7060 );
and ( n7062 , n7033 , n7060 );
or ( n7063 , n7052 , n7061 , n7062 );
and ( n7064 , n7031 , n7063 );
xor ( n7065 , n6966 , n6973 );
xor ( n7066 , n7065 , n6976 );
and ( n7067 , n7063 , n7066 );
and ( n7068 , n7031 , n7066 );
or ( n7069 , n7064 , n7067 , n7068 );
xor ( n7070 , n6888 , n6889 );
xor ( n7071 , n7070 , n6935 );
and ( n7072 , n7069 , n7071 );
xor ( n7073 , n7002 , n7004 );
xor ( n7074 , n6985 , n6986 );
xor ( n7075 , n7074 , n6988 );
xor ( n7076 , n6992 , n6993 );
xor ( n7077 , n7076 , n6995 );
and ( n7078 , n7075 , n7077 );
and ( n7079 , n7073 , n7078 );
buf ( n7080 , n5936 );
xor ( n7081 , n6898 , n6899 );
and ( n7082 , n7080 , n7081 );
and ( n7083 , n5745 , n6329 );
and ( n7084 , n5753 , n6143 );
and ( n7085 , n7083 , n7084 );
and ( n7086 , n5865 , n6120 );
and ( n7087 , n7084 , n7086 );
and ( n7088 , n7083 , n7086 );
or ( n7089 , n7085 , n7087 , n7088 );
and ( n7090 , n7081 , n7089 );
and ( n7091 , n7080 , n7089 );
or ( n7092 , n7082 , n7090 , n7091 );
and ( n7093 , n7078 , n7092 );
and ( n7094 , n7073 , n7092 );
or ( n7095 , n7079 , n7093 , n7094 );
xor ( n7096 , n6984 , n6999 );
xor ( n7097 , n7096 , n7005 );
and ( n7098 , n7095 , n7097 );
xor ( n7099 , n7028 , n7030 );
and ( n7100 , n7097 , n7099 );
and ( n7101 , n7095 , n7099 );
or ( n7102 , n7098 , n7100 , n7101 );
xor ( n7103 , n7008 , n7010 );
xor ( n7104 , n7103 , n7012 );
and ( n7105 , n7102 , n7104 );
xor ( n7106 , n7031 , n7063 );
xor ( n7107 , n7106 , n7066 );
and ( n7108 , n7104 , n7107 );
and ( n7109 , n7102 , n7107 );
or ( n7110 , n7105 , n7108 , n7109 );
and ( n7111 , n7071 , n7110 );
and ( n7112 , n7069 , n7110 );
or ( n7113 , n7072 , n7111 , n7112 );
and ( n7114 , n7026 , n7113 );
xor ( n7115 , n6962 , n6964 );
xor ( n7116 , n7115 , n7018 );
and ( n7117 , n7113 , n7116 );
and ( n7118 , n7026 , n7116 );
or ( n7119 , n7114 , n7117 , n7118 );
and ( n7120 , n7023 , n7119 );
and ( n7121 , n7021 , n7119 );
or ( n7122 , n7024 , n7120 , n7121 );
and ( n7123 , n6960 , n7122 );
xor ( n7124 , n7021 , n7023 );
xor ( n7125 , n7124 , n7119 );
xor ( n7126 , n7026 , n7113 );
xor ( n7127 , n7126 , n7116 );
xor ( n7128 , n6979 , n6981 );
xor ( n7129 , n7128 , n7015 );
xor ( n7130 , n7069 , n7071 );
xor ( n7131 , n7130 , n7110 );
and ( n7132 , n7129 , n7131 );
xor ( n7133 , n7048 , n7050 );
and ( n7134 , n5865 , n6143 );
and ( n7135 , n5936 , n6120 );
and ( n7136 , n7134 , n7135 );
and ( n7137 , n6314 , n5676 );
and ( n7138 , n7136 , n7137 );
and ( n7139 , n6134 , n5871 );
and ( n7140 , n6115 , n5927 );
and ( n7141 , n7139 , n7140 );
and ( n7142 , n5667 , n6357 );
and ( n7143 , n7141 , n7142 );
and ( n7144 , n7138 , n7143 );
and ( n7145 , n7133 , n7144 );
xor ( n7146 , n7034 , n7041 );
xor ( n7147 , n7146 , n7045 );
xor ( n7148 , n7075 , n7077 );
and ( n7149 , n7147 , n7148 );
xor ( n7150 , n7083 , n7084 );
xor ( n7151 , n7150 , n7086 );
xor ( n7152 , n7043 , n7044 );
and ( n7153 , n7151 , n7152 );
and ( n7154 , n6314 , n5762 );
and ( n7155 , n6317 , n5736 );
and ( n7156 , n7154 , n7155 );
and ( n7157 , n7152 , n7156 );
and ( n7158 , n7151 , n7156 );
or ( n7159 , n7153 , n7157 , n7158 );
and ( n7160 , n7148 , n7159 );
and ( n7161 , n7147 , n7159 );
or ( n7162 , n7149 , n7160 , n7161 );
and ( n7163 , n7144 , n7162 );
and ( n7164 , n7133 , n7162 );
or ( n7165 , n7145 , n7163 , n7164 );
xor ( n7166 , n7033 , n7051 );
xor ( n7167 , n7166 , n7060 );
and ( n7168 , n7165 , n7167 );
xor ( n7169 , n7053 , n7055 );
xor ( n7170 , n7169 , n7057 );
xor ( n7171 , n7073 , n7078 );
xor ( n7172 , n7171 , n7092 );
and ( n7173 , n7170 , n7172 );
xor ( n7174 , n7080 , n7081 );
xor ( n7175 , n7174 , n7089 );
xor ( n7176 , n7138 , n7143 );
and ( n7177 , n7175 , n7176 );
and ( n7178 , n5992 , n6120 );
and ( n7179 , n6115 , n5989 );
and ( n7180 , n7178 , n7179 );
and ( n7181 , n5745 , n6357 );
and ( n7182 , n7180 , n7181 );
and ( n7183 , n5753 , n6329 );
and ( n7184 , n7181 , n7183 );
and ( n7185 , n7180 , n7183 );
or ( n7186 , n7182 , n7184 , n7185 );
xor ( n7187 , n7035 , n7036 );
xor ( n7188 , n7187 , n7038 );
and ( n7189 , n7186 , n7188 );
and ( n7190 , n7176 , n7189 );
and ( n7191 , n7175 , n7189 );
or ( n7192 , n7177 , n7190 , n7191 );
and ( n7193 , n7172 , n7192 );
and ( n7194 , n7170 , n7192 );
or ( n7195 , n7173 , n7193 , n7194 );
and ( n7196 , n7167 , n7195 );
and ( n7197 , n7165 , n7195 );
or ( n7198 , n7168 , n7196 , n7197 );
xor ( n7199 , n7102 , n7104 );
xor ( n7200 , n7199 , n7107 );
and ( n7201 , n7198 , n7200 );
xor ( n7202 , n7095 , n7097 );
xor ( n7203 , n7202 , n7099 );
xor ( n7204 , n7133 , n7144 );
xor ( n7205 , n7204 , n7162 );
xor ( n7206 , n7136 , n7137 );
xor ( n7207 , n7141 , n7142 );
and ( n7208 , n7206 , n7207 );
xor ( n7209 , n7147 , n7148 );
xor ( n7210 , n7209 , n7159 );
and ( n7211 , n7208 , n7210 );
and ( n7212 , n5753 , n6357 );
and ( n7213 , n5865 , n6329 );
and ( n7214 , n7212 , n7213 );
and ( n7215 , n5936 , n6143 );
and ( n7216 , n7213 , n7215 );
and ( n7217 , n7212 , n7215 );
or ( n7218 , n7214 , n7216 , n7217 );
xor ( n7219 , n7139 , n7140 );
and ( n7220 , n7218 , n7219 );
xor ( n7221 , n7151 , n7152 );
xor ( n7222 , n7221 , n7156 );
and ( n7223 , n7220 , n7222 );
xor ( n7224 , n7186 , n7188 );
and ( n7225 , n7222 , n7224 );
and ( n7226 , n7220 , n7224 );
or ( n7227 , n7223 , n7225 , n7226 );
and ( n7228 , n7210 , n7227 );
and ( n7229 , n7208 , n7227 );
or ( n7230 , n7211 , n7228 , n7229 );
and ( n7231 , n7205 , n7230 );
xor ( n7232 , n7170 , n7172 );
xor ( n7233 , n7232 , n7192 );
and ( n7234 , n7230 , n7233 );
and ( n7235 , n7205 , n7233 );
or ( n7236 , n7231 , n7234 , n7235 );
and ( n7237 , n7203 , n7236 );
xor ( n7238 , n7165 , n7167 );
xor ( n7239 , n7238 , n7195 );
and ( n7240 , n7236 , n7239 );
and ( n7241 , n7203 , n7239 );
or ( n7242 , n7237 , n7240 , n7241 );
and ( n7243 , n7200 , n7242 );
and ( n7244 , n7198 , n7242 );
or ( n7245 , n7201 , n7243 , n7244 );
and ( n7246 , n7131 , n7245 );
and ( n7247 , n7129 , n7245 );
or ( n7248 , n7132 , n7246 , n7247 );
or ( n7249 , n7127 , n7248 );
or ( n7250 , n7125 , n7249 );
and ( n7251 , n7122 , n7250 );
and ( n7252 , n6960 , n7250 );
or ( n7253 , n7123 , n7251 , n7252 );
and ( n7254 , n6957 , n7253 );
and ( n7255 , n6955 , n7253 );
or ( n7256 , n6958 , n7254 , n7255 );
and ( n7257 , n6879 , n7256 );
and ( n7258 , n6877 , n7256 );
or ( n7259 , n6880 , n7257 , n7258 );
or ( n7260 , n6797 , n7259 );
and ( n7261 , n6794 , n7260 );
and ( n7262 , n6493 , n7260 );
or ( n7263 , n6795 , n7261 , n7262 );
and ( n7264 , n6490 , n7263 );
and ( n7265 , n6488 , n7263 );
or ( n7266 , n6491 , n7264 , n7265 );
and ( n7267 , n6436 , n7266 );
xor ( n7268 , n6436 , n7266 );
xor ( n7269 , n6488 , n6490 );
xor ( n7270 , n7269 , n7263 );
not ( n7271 , n7270 );
xor ( n7272 , n6493 , n6794 );
xor ( n7273 , n7272 , n7260 );
xnor ( n7274 , n6797 , n7259 );
xor ( n7275 , n6877 , n6879 );
xor ( n7276 , n7275 , n7256 );
xor ( n7277 , n6955 , n6957 );
xor ( n7278 , n7277 , n7253 );
not ( n7279 , n7278 );
xor ( n7280 , n6960 , n7122 );
xor ( n7281 , n7280 , n7250 );
not ( n7282 , n7281 );
xnor ( n7283 , n7125 , n7249 );
xnor ( n7284 , n7127 , n7248 );
xor ( n7285 , n7129 , n7131 );
xor ( n7286 , n7285 , n7245 );
not ( n7287 , n7286 );
xor ( n7288 , n7198 , n7200 );
xor ( n7289 , n7288 , n7242 );
xor ( n7290 , n7203 , n7236 );
xor ( n7291 , n7290 , n7239 );
xor ( n7292 , n7206 , n7207 );
xor ( n7293 , n7134 , n7135 );
and ( n7294 , n6314 , n5736 );
and ( n7295 , n6317 , n5871 );
and ( n7296 , n7294 , n7295 );
and ( n7297 , n6134 , n5927 );
and ( n7298 , n7295 , n7297 );
and ( n7299 , n7294 , n7297 );
or ( n7300 , n7296 , n7298 , n7299 );
and ( n7301 , n7293 , n7300 );
xor ( n7302 , n7180 , n7181 );
xor ( n7303 , n7302 , n7183 );
and ( n7304 , n7300 , n7303 );
and ( n7305 , n7293 , n7303 );
or ( n7306 , n7301 , n7304 , n7305 );
and ( n7307 , n7292 , n7306 );
buf ( n7308 , n5992 );
xor ( n7309 , n7154 , n7155 );
and ( n7310 , n7308 , n7309 );
xor ( n7311 , n7218 , n7219 );
and ( n7312 , n7309 , n7311 );
and ( n7313 , n7308 , n7311 );
or ( n7314 , n7310 , n7312 , n7313 );
and ( n7315 , n7306 , n7314 );
and ( n7316 , n7292 , n7314 );
or ( n7317 , n7307 , n7315 , n7316 );
xor ( n7318 , n7175 , n7176 );
xor ( n7319 , n7318 , n7189 );
and ( n7320 , n7317 , n7319 );
and ( n7321 , n6317 , n5927 );
and ( n7322 , n6134 , n5989 );
and ( n7323 , n7321 , n7322 );
and ( n7324 , n5936 , n6329 );
and ( n7325 , n5992 , n6143 );
and ( n7326 , n7324 , n7325 );
and ( n7327 , n7323 , n7326 );
xor ( n7328 , n7294 , n7295 );
xor ( n7329 , n7328 , n7297 );
xor ( n7330 , n7212 , n7213 );
xor ( n7331 , n7330 , n7215 );
and ( n7332 , n7329 , n7331 );
and ( n7333 , n7327 , n7332 );
xor ( n7334 , n7293 , n7300 );
xor ( n7335 , n7334 , n7303 );
and ( n7336 , n7332 , n7335 );
and ( n7337 , n7327 , n7335 );
or ( n7338 , n7333 , n7336 , n7337 );
xor ( n7339 , n7178 , n7179 );
xor ( n7340 , n7323 , n7326 );
and ( n7341 , n7339 , n7340 );
xor ( n7342 , n7329 , n7331 );
and ( n7343 , n7340 , n7342 );
and ( n7344 , n7339 , n7342 );
or ( n7345 , n7341 , n7343 , n7344 );
xor ( n7346 , n7324 , n7325 );
and ( n7347 , n6115 , n6143 );
and ( n7348 , n6134 , n6120 );
and ( n7349 , n7347 , n7348 );
and ( n7350 , n7346 , n7349 );
and ( n7351 , n5865 , n6357 );
and ( n7352 , n7349 , n7351 );
and ( n7353 , n7346 , n7351 );
or ( n7354 , n7350 , n7352 , n7353 );
and ( n7355 , n6314 , n5927 );
and ( n7356 , n6317 , n5989 );
and ( n7357 , n7355 , n7356 );
and ( n7358 , n5936 , n6357 );
and ( n7359 , n5992 , n6329 );
and ( n7360 , n7358 , n7359 );
and ( n7361 , n7357 , n7360 );
and ( n7362 , n7354 , n7361 );
and ( n7363 , n6314 , n5871 );
buf ( n7364 , n6115 );
and ( n7365 , n7363 , n7364 );
xor ( n7366 , n7321 , n7322 );
and ( n7367 , n7364 , n7366 );
and ( n7368 , n7363 , n7366 );
or ( n7369 , n7365 , n7367 , n7368 );
and ( n7370 , n7361 , n7369 );
and ( n7371 , n7354 , n7369 );
or ( n7372 , n7362 , n7370 , n7371 );
and ( n7373 , n7345 , n7372 );
xor ( n7374 , n7308 , n7309 );
xor ( n7375 , n7374 , n7311 );
and ( n7376 , n7372 , n7375 );
and ( n7377 , n7345 , n7375 );
or ( n7378 , n7373 , n7376 , n7377 );
and ( n7379 , n7338 , n7378 );
xor ( n7380 , n7220 , n7222 );
xor ( n7381 , n7380 , n7224 );
and ( n7382 , n7378 , n7381 );
and ( n7383 , n7338 , n7381 );
or ( n7384 , n7379 , n7382 , n7383 );
and ( n7385 , n7319 , n7384 );
and ( n7386 , n7317 , n7384 );
or ( n7387 , n7320 , n7385 , n7386 );
xor ( n7388 , n7205 , n7230 );
xor ( n7389 , n7388 , n7233 );
and ( n7390 , n7387 , n7389 );
xor ( n7391 , n7208 , n7210 );
xor ( n7392 , n7391 , n7227 );
xor ( n7393 , n7292 , n7306 );
xor ( n7394 , n7393 , n7314 );
xor ( n7395 , n7346 , n7349 );
xor ( n7396 , n7395 , n7351 );
xor ( n7397 , n7357 , n7360 );
and ( n7398 , n7396 , n7397 );
and ( n7399 , n6314 , n5989 );
and ( n7400 , n6317 , n6120 );
and ( n7401 , n7399 , n7400 );
and ( n7402 , n5992 , n6357 );
and ( n7403 , n6115 , n6329 );
and ( n7404 , n7402 , n7403 );
and ( n7405 , n7401 , n7404 );
and ( n7406 , n7397 , n7405 );
and ( n7407 , n7396 , n7405 );
or ( n7408 , n7398 , n7406 , n7407 );
xor ( n7409 , n7339 , n7340 );
xor ( n7410 , n7409 , n7342 );
and ( n7411 , n7408 , n7410 );
xor ( n7412 , n7354 , n7361 );
xor ( n7413 , n7412 , n7369 );
and ( n7414 , n7410 , n7413 );
and ( n7415 , n7408 , n7413 );
or ( n7416 , n7411 , n7414 , n7415 );
xor ( n7417 , n7327 , n7332 );
xor ( n7418 , n7417 , n7335 );
and ( n7419 , n7416 , n7418 );
xor ( n7420 , n7345 , n7372 );
xor ( n7421 , n7420 , n7375 );
and ( n7422 , n7418 , n7421 );
and ( n7423 , n7416 , n7421 );
or ( n7424 , n7419 , n7422 , n7423 );
and ( n7425 , n7394 , n7424 );
xor ( n7426 , n7338 , n7378 );
xor ( n7427 , n7426 , n7381 );
and ( n7428 , n7424 , n7427 );
and ( n7429 , n7394 , n7427 );
or ( n7430 , n7425 , n7428 , n7429 );
and ( n7431 , n7392 , n7430 );
xor ( n7432 , n7317 , n7319 );
xor ( n7433 , n7432 , n7384 );
and ( n7434 , n7430 , n7433 );
and ( n7435 , n7392 , n7433 );
or ( n7436 , n7431 , n7434 , n7435 );
and ( n7437 , n7389 , n7436 );
and ( n7438 , n7387 , n7436 );
or ( n7439 , n7390 , n7437 , n7438 );
and ( n7440 , n7291 , n7439 );
xor ( n7441 , n7387 , n7389 );
xor ( n7442 , n7441 , n7436 );
xor ( n7443 , n7392 , n7430 );
xor ( n7444 , n7443 , n7433 );
xor ( n7445 , n7394 , n7424 );
xor ( n7446 , n7445 , n7427 );
xor ( n7447 , n7416 , n7418 );
xor ( n7448 , n7447 , n7421 );
xor ( n7449 , n7355 , n7356 );
xor ( n7450 , n7358 , n7359 );
and ( n7451 , n7449 , n7450 );
xor ( n7452 , n7363 , n7364 );
xor ( n7453 , n7452 , n7366 );
and ( n7454 , n7451 , n7453 );
xor ( n7455 , n7347 , n7348 );
xor ( n7456 , n7401 , n7404 );
and ( n7457 , n7455 , n7456 );
xor ( n7458 , n7449 , n7450 );
and ( n7459 , n7456 , n7458 );
and ( n7460 , n7455 , n7458 );
or ( n7461 , n7457 , n7459 , n7460 );
and ( n7462 , n7453 , n7461 );
and ( n7463 , n7451 , n7461 );
or ( n7464 , n7454 , n7462 , n7463 );
xor ( n7465 , n7408 , n7410 );
xor ( n7466 , n7465 , n7413 );
and ( n7467 , n7464 , n7466 );
xor ( n7468 , n7396 , n7397 );
xor ( n7469 , n7468 , n7405 );
and ( n7470 , n6115 , n6357 );
and ( n7471 , n6314 , n6120 );
and ( n7472 , n7470 , n7471 );
buf ( n7473 , n6134 );
or ( n7474 , n7472 , n7473 );
xor ( n7475 , n7399 , n7400 );
xor ( n7476 , n7402 , n7403 );
and ( n7477 , n7475 , n7476 );
and ( n7478 , n7474 , n7477 );
and ( n7479 , n6134 , n6329 );
and ( n7480 , n6317 , n6143 );
and ( n7481 , n7479 , n7480 );
xnor ( n7482 , n7472 , n7473 );
or ( n7483 , n7481 , n7482 );
and ( n7484 , n7477 , n7483 );
and ( n7485 , n7474 , n7483 );
or ( n7486 , n7478 , n7484 , n7485 );
and ( n7487 , n7469 , n7486 );
xor ( n7488 , n7451 , n7453 );
xor ( n7489 , n7488 , n7461 );
and ( n7490 , n7486 , n7489 );
and ( n7491 , n7469 , n7489 );
or ( n7492 , n7487 , n7490 , n7491 );
and ( n7493 , n7466 , n7492 );
and ( n7494 , n7464 , n7492 );
or ( n7495 , n7467 , n7493 , n7494 );
and ( n7496 , n7448 , n7495 );
xor ( n7497 , n7455 , n7456 );
xor ( n7498 , n7497 , n7458 );
xor ( n7499 , n7475 , n7476 );
xnor ( n7500 , n7481 , n7482 );
and ( n7501 , n7499 , n7500 );
xor ( n7502 , n7470 , n7471 );
xor ( n7503 , n7479 , n7480 );
and ( n7504 , n7502 , n7503 );
and ( n7505 , n6317 , n6357 );
and ( n7506 , n6314 , n6329 );
and ( n7507 , n7505 , n7506 );
and ( n7508 , n6134 , n6357 );
and ( n7509 , n7507 , n7508 );
and ( n7510 , n7503 , n7509 );
and ( n7511 , n7502 , n7509 );
or ( n7512 , n7504 , n7510 , n7511 );
and ( n7513 , n7500 , n7512 );
and ( n7514 , n7499 , n7512 );
or ( n7515 , n7501 , n7513 , n7514 );
and ( n7516 , n7498 , n7515 );
xor ( n7517 , n7474 , n7477 );
xor ( n7518 , n7517 , n7483 );
and ( n7519 , n7515 , n7518 );
and ( n7520 , n7498 , n7518 );
or ( n7521 , n7516 , n7519 , n7520 );
xor ( n7522 , n7469 , n7486 );
xor ( n7523 , n7522 , n7489 );
or ( n7524 , n7521 , n7523 );
xor ( n7525 , n7464 , n7466 );
xor ( n7526 , n7525 , n7492 );
or ( n7527 , n7524 , n7526 );
and ( n7528 , n7495 , n7527 );
and ( n7529 , n7448 , n7527 );
or ( n7530 , n7496 , n7528 , n7529 );
or ( n7531 , n7446 , n7530 );
or ( n7532 , n7444 , n7531 );
or ( n7533 , n7442 , n7532 );
and ( n7534 , n7439 , n7533 );
and ( n7535 , n7291 , n7533 );
or ( n7536 , n7440 , n7534 , n7535 );
and ( n7537 , n7289 , n7536 );
xor ( n7538 , n7289 , n7536 );
xor ( n7539 , n7291 , n7439 );
xor ( n7540 , n7539 , n7533 );
not ( n7541 , n7540 );
xnor ( n7542 , n7442 , n7532 );
xnor ( n7543 , n7444 , n7531 );
xnor ( n7544 , n7446 , n7530 );
xor ( n7545 , n7448 , n7495 );
xor ( n7546 , n7545 , n7527 );
not ( n7547 , n7546 );
xnor ( n7548 , n7524 , n7526 );
xnor ( n7549 , n7521 , n7523 );
xor ( n7550 , n7498 , n7515 );
xor ( n7551 , n7550 , n7518 );
buf ( n7552 , n6317 );
not ( n7553 , n7552 );
xor ( n7554 , n7507 , n7508 );
and ( n7555 , n7553 , n7554 );
buf ( n7556 , n7552 );
and ( n7557 , n7555 , n7556 );
xor ( n7558 , n7502 , n7503 );
xor ( n7559 , n7558 , n7509 );
and ( n7560 , n7556 , n7559 );
and ( n7561 , n7555 , n7559 );
or ( n7562 , n7557 , n7560 , n7561 );
xor ( n7563 , n7499 , n7500 );
xor ( n7564 , n7563 , n7512 );
and ( n7565 , n7562 , n7564 );
and ( n7566 , n6314 , n6143 );
xor ( n7567 , n7553 , n7554 );
or ( n7568 , n7566 , n7567 );
xor ( n7569 , n7555 , n7556 );
xor ( n7570 , n7569 , n7559 );
or ( n7571 , n7568 , n7570 );
and ( n7572 , n7564 , n7571 );
and ( n7573 , n7562 , n7571 );
or ( n7574 , n7565 , n7572 , n7573 );
and ( n7575 , n7551 , n7574 );
xor ( n7576 , n7551 , n7574 );
xor ( n7577 , n7562 , n7564 );
xor ( n7578 , n7577 , n7571 );
and ( n7579 , n7576 , n7578 );
or ( n7580 , n7575 , n7579 );
and ( n7581 , n7549 , n7580 );
and ( n7582 , n7548 , n7581 );
and ( n7583 , n7547 , n7582 );
or ( n7584 , n7546 , n7583 );
and ( n7585 , n7544 , n7584 );
and ( n7586 , n7543 , n7585 );
and ( n7587 , n7542 , n7586 );
and ( n7588 , n7541 , n7587 );
or ( n7589 , n7540 , n7588 );
and ( n7590 , n7538 , n7589 );
or ( n7591 , n7537 , n7590 );
and ( n7592 , n7287 , n7591 );
or ( n7593 , n7286 , n7592 );
and ( n7594 , n7284 , n7593 );
and ( n7595 , n7283 , n7594 );
and ( n7596 , n7282 , n7595 );
or ( n7597 , n7281 , n7596 );
and ( n7598 , n7279 , n7597 );
or ( n7599 , n7278 , n7598 );
and ( n7600 , n7276 , n7599 );
and ( n7601 , n7274 , n7600 );
and ( n7602 , n7273 , n7601 );
and ( n7603 , n7271 , n7602 );
or ( n7604 , n7270 , n7603 );
and ( n7605 , n7268 , n7604 );
or ( n7606 , n7267 , n7605 );
and ( n7607 , n6434 , n7606 );
or ( n7608 , n6433 , n7607 );
and ( n7609 , n6431 , n7608 );
and ( n7610 , n6430 , n7609 );
and ( n7611 , n6429 , n7610 );
and ( n7612 , n6427 , n7611 );
or ( n7613 , n6426 , n7612 );
and ( n7614 , n6424 , n7613 );
and ( n7615 , n6423 , n7614 );
or ( n7616 , n6422 , n7615 );
xor ( n7617 , n6420 , n7616 );
buf ( n7618 , n7617 );
buf ( n7619 , n7618 );
buf ( n7620 , n7619 );
xor ( n7621 , n5562 , n7620 );
and ( n7622 , n5285 , n5262 );
and ( n7623 , n5254 , n5260 );
nor ( n7624 , n7622 , n7623 );
xnor ( n7625 , n7624 , n5270 );
and ( n7626 , n5529 , n5282 );
and ( n7627 , n5274 , n5280 );
nor ( n7628 , n7626 , n7627 );
xnor ( n7629 , n7628 , n5290 );
xor ( n7630 , n7625 , n7629 );
xor ( n7631 , n5342 , n5509 );
not ( n7632 , n5512 );
and ( n7633 , n7631 , n7632 );
and ( n7634 , n5340 , n7633 );
buf ( n7635 , n776 );
buf ( n7636 , n7635 );
buf ( n7637 , n7636 );
buf ( n7638 , n7637 );
buf ( n7639 , n7638 );
and ( n7640 , n7639 , n5512 );
nor ( n7641 , n7634 , n7640 );
xnor ( n7642 , n7641 , n5561 );
xor ( n7643 , n7630 , n7642 );
xor ( n7644 , n7621 , n7643 );
and ( n7645 , n5557 , n7644 );
buf ( n7646 , n1988 );
buf ( n7647 , n7646 );
and ( n7648 , n7647 , n5306 );
buf ( n7649 , n1904 );
buf ( n7650 , n7649 );
and ( n7651 , n7650 , n5304 );
nor ( n7652 , n7648 , n7651 );
xnor ( n7653 , n7652 , n5314 );
and ( n7654 , n5368 , n5282 );
and ( n7655 , n5529 , n5280 );
nor ( n7656 , n7654 , n7655 );
xnor ( n7657 , n7656 , n5290 );
and ( n7658 , n7653 , n7657 );
buf ( n7659 , n4980 );
buf ( n7660 , n7659 );
and ( n7661 , n7660 , n5365 );
and ( n7662 , n5536 , n5363 );
nor ( n7663 , n7661 , n7662 );
xnor ( n7664 , n7663 , n5373 );
and ( n7665 , n7657 , n7664 );
and ( n7666 , n7653 , n7664 );
or ( n7667 , n7658 , n7665 , n7666 );
and ( n7668 , n5408 , n5390 );
and ( n7669 , n5377 , n5387 );
nor ( n7670 , n7668 , n7669 );
xnor ( n7671 , n7670 , n5382 );
and ( n7672 , n5437 , n5412 );
not ( n7673 , n7672 );
xnor ( n7674 , n7673 , n5420 );
and ( n7675 , n7671 , n7674 );
and ( n7676 , n7674 , n5405 );
and ( n7677 , n7671 , n5405 );
or ( n7678 , n7675 , n7676 , n7677 );
xor ( n7679 , n7667 , n7678 );
and ( n7680 , n5265 , n5243 );
and ( n7681 , n5233 , n5241 );
nor ( n7682 , n7680 , n7681 );
xnor ( n7683 , n7682 , n5251 );
and ( n7684 , n5355 , n5542 );
and ( n7685 , n5368 , n5540 );
nor ( n7686 , n7684 , n7685 );
xnor ( n7687 , n7686 , n5550 );
xor ( n7688 , n7683 , n7687 );
buf ( n7689 , n5084 );
buf ( n7690 , n7689 );
buf ( n7691 , n1369 );
buf ( n7692 , n7691 );
xor ( n7693 , n5511 , n7692 );
xor ( n7694 , n7692 , n5357 );
not ( n7695 , n7694 );
and ( n7696 , n7693 , n7695 );
and ( n7697 , n7690 , n7696 );
and ( n7698 , n7660 , n7694 );
nor ( n7699 , n7697 , n7698 );
and ( n7700 , n7692 , n5357 );
not ( n7701 , n7700 );
and ( n7702 , n5511 , n7701 );
xnor ( n7703 , n7699 , n7702 );
xor ( n7704 , n7688 , n7703 );
xor ( n7705 , n7679 , n7704 );
and ( n7706 , n7644 , n7705 );
and ( n7707 , n5557 , n7705 );
or ( n7708 , n7645 , n7706 , n7707 );
and ( n7709 , n5309 , n5487 );
buf ( n7710 , n1687 );
buf ( n7711 , n7710 );
and ( n7712 , n7711 , n5485 );
nor ( n7713 , n7709 , n7712 );
xnor ( n7714 , n7713 , n5478 );
buf ( n7715 , n2046 );
buf ( n7716 , n7715 );
buf ( n7717 , n2935 );
buf ( n7718 , n7717 );
xor ( n7719 , n5496 , n7718 );
xor ( n7720 , n7718 , n5298 );
not ( n7721 , n7720 );
and ( n7722 , n7719 , n7721 );
and ( n7723 , n7716 , n7722 );
and ( n7724 , n7647 , n7720 );
nor ( n7725 , n7723 , n7724 );
and ( n7726 , n7718 , n5298 );
not ( n7727 , n7726 );
and ( n7728 , n5496 , n7727 );
xnor ( n7729 , n7725 , n7728 );
and ( n7730 , n7714 , n7729 );
and ( n7731 , n5328 , n5499 );
and ( n7732 , n5350 , n5497 );
nor ( n7733 , n7731 , n7732 );
xnor ( n7734 , n7733 , n5505 );
and ( n7735 , n7729 , n7734 );
and ( n7736 , n7714 , n7734 );
or ( n7737 , n7730 , n7735 , n7736 );
and ( n7738 , n7683 , n7687 );
and ( n7739 , n7687 , n7703 );
and ( n7740 , n7683 , n7703 );
or ( n7741 , n7738 , n7739 , n7740 );
xor ( n7742 , n7737 , n7741 );
and ( n7743 , n7625 , n7629 );
and ( n7744 , n7629 , n7642 );
and ( n7745 , n7625 , n7642 );
or ( n7746 , n7743 , n7744 , n7745 );
xor ( n7747 , n5315 , n5334 );
xor ( n7748 , n7747 , n5343 );
xor ( n7749 , n7746 , n7748 );
and ( n7750 , n5368 , n5542 );
and ( n7751 , n5529 , n5540 );
nor ( n7752 , n7750 , n7751 );
xnor ( n7753 , n7752 , n5550 );
and ( n7754 , n7660 , n7696 );
and ( n7755 , n5536 , n7694 );
nor ( n7756 , n7754 , n7755 );
xnor ( n7757 , n7756 , n7702 );
xor ( n7758 , n7753 , n7757 );
and ( n7759 , n7639 , n7633 );
and ( n7760 , n7690 , n5512 );
nor ( n7761 , n7759 , n7760 );
xnor ( n7762 , n7761 , n5561 );
xor ( n7763 , n7758 , n7762 );
xor ( n7764 , n7749 , n7763 );
xor ( n7765 , n7742 , n7764 );
xor ( n7766 , n7708 , n7765 );
and ( n7767 , n7650 , n5306 );
and ( n7768 , n5296 , n5304 );
nor ( n7769 , n7767 , n7768 );
xnor ( n7770 , n7769 , n5314 );
and ( n7771 , n5246 , n5325 );
and ( n7772 , n5317 , n5323 );
nor ( n7773 , n7771 , n7772 );
xnor ( n7774 , n7773 , n5333 );
and ( n7775 , n7770 , n7774 );
and ( n7776 , n5536 , n5365 );
and ( n7777 , n5545 , n5363 );
nor ( n7778 , n7776 , n7777 );
xnor ( n7779 , n7778 , n5373 );
and ( n7780 , n7774 , n7779 );
and ( n7781 , n7770 , n7779 );
or ( n7782 , n7775 , n7780 , n7781 );
and ( n7783 , n7647 , n7722 );
and ( n7784 , n7650 , n7720 );
nor ( n7785 , n7783 , n7784 );
xnor ( n7786 , n7785 , n7728 );
and ( n7787 , n5350 , n5499 );
and ( n7788 , n7716 , n5497 );
nor ( n7789 , n7787 , n7788 );
xnor ( n7790 , n7789 , n5505 );
xor ( n7791 , n7786 , n7790 );
and ( n7792 , n5545 , n5365 );
and ( n7793 , n5355 , n5363 );
nor ( n7794 , n7792 , n7793 );
xnor ( n7795 , n7794 , n5373 );
xor ( n7796 , n7791 , n7795 );
xnor ( n7797 , n7782 , n7796 );
and ( n7798 , n5254 , n5243 );
and ( n7799 , n5265 , n5241 );
nor ( n7800 , n7798 , n7799 );
xnor ( n7801 , n7800 , n5251 );
and ( n7802 , n5274 , n5262 );
and ( n7803 , n5285 , n5260 );
nor ( n7804 , n7802 , n7803 );
xnor ( n7805 , n7804 , n5270 );
and ( n7806 , n7801 , n7805 );
and ( n7807 , n5545 , n5542 );
and ( n7808 , n5355 , n5540 );
nor ( n7809 , n7807 , n7808 );
xnor ( n7810 , n7809 , n5550 );
and ( n7811 , n7805 , n7810 );
and ( n7812 , n7801 , n7810 );
or ( n7813 , n7806 , n7811 , n7812 );
and ( n7814 , n5491 , n5506 );
and ( n7815 , n5506 , n5513 );
and ( n7816 , n5491 , n5513 );
or ( n7817 , n7814 , n7815 , n7816 );
and ( n7818 , n7813 , n7817 );
xor ( n7819 , n7714 , n7729 );
xor ( n7820 , n7819 , n7734 );
and ( n7821 , n7817 , n7820 );
and ( n7822 , n7813 , n7820 );
or ( n7823 , n7818 , n7821 , n7822 );
xor ( n7824 , n7797 , n7823 );
and ( n7825 , n5350 , n7722 );
and ( n7826 , n7716 , n7720 );
nor ( n7827 , n7825 , n7826 );
xnor ( n7828 , n7827 , n7728 );
and ( n7829 , n5233 , n5325 );
and ( n7830 , n5246 , n5323 );
nor ( n7831 , n7829 , n7830 );
xnor ( n7832 , n7831 , n5333 );
and ( n7833 , n7828 , n7832 );
and ( n7834 , n7639 , n7696 );
and ( n7835 , n7690 , n7694 );
nor ( n7836 , n7834 , n7835 );
xnor ( n7837 , n7836 , n7702 );
and ( n7838 , n7832 , n7837 );
and ( n7839 , n7828 , n7837 );
or ( n7840 , n7833 , n7838 , n7839 );
xor ( n7841 , n7770 , n7774 );
xor ( n7842 , n7841 , n7779 );
or ( n7843 , n7840 , n7842 );
xor ( n7844 , n7824 , n7843 );
xor ( n7845 , n7766 , n7844 );
and ( n7846 , n7716 , n5306 );
and ( n7847 , n7647 , n5304 );
nor ( n7848 , n7846 , n7847 );
xnor ( n7849 , n7848 , n5314 );
and ( n7850 , n5328 , n7722 );
and ( n7851 , n5350 , n7720 );
nor ( n7852 , n7850 , n7851 );
xnor ( n7853 , n7852 , n7728 );
and ( n7854 , n7849 , n7853 );
and ( n7855 , n5265 , n5325 );
and ( n7856 , n5233 , n5323 );
nor ( n7857 , n7855 , n7856 );
xnor ( n7858 , n7857 , n5333 );
and ( n7859 , n7853 , n7858 );
and ( n7860 , n7849 , n7858 );
or ( n7861 , n7854 , n7859 , n7860 );
xor ( n7862 , n5424 , n5426 );
xor ( n7863 , n5426 , n5398 );
not ( n7864 , n7863 );
and ( n7865 , n7862 , n7864 );
and ( n7866 , n5309 , n7865 );
and ( n7867 , n7711 , n7863 );
nor ( n7868 , n7866 , n7867 );
xnor ( n7869 , n7868 , n5429 );
and ( n7870 , n5246 , n5499 );
and ( n7871 , n5317 , n5497 );
nor ( n7872 , n7870 , n7871 );
xnor ( n7873 , n7872 , n5505 );
and ( n7874 , n7869 , n7873 );
and ( n7875 , n7690 , n5365 );
and ( n7876 , n7660 , n5363 );
nor ( n7877 , n7875 , n7876 );
xnor ( n7878 , n7877 , n5373 );
and ( n7879 , n7873 , n7878 );
and ( n7880 , n7869 , n7878 );
or ( n7881 , n7874 , n7879 , n7880 );
and ( n7882 , n7861 , n7881 );
and ( n7883 , n7650 , n5487 );
and ( n7884 , n5296 , n5485 );
nor ( n7885 , n7883 , n7884 );
xnor ( n7886 , n7885 , n5478 );
and ( n7887 , n5355 , n5282 );
and ( n7888 , n5368 , n5280 );
nor ( n7889 , n7887 , n7888 );
xnor ( n7890 , n7889 , n5290 );
and ( n7891 , n7886 , n7890 );
and ( n7892 , n5340 , n7696 );
and ( n7893 , n7639 , n7694 );
nor ( n7894 , n7892 , n7893 );
xnor ( n7895 , n7894 , n7702 );
and ( n7896 , n7890 , n7895 );
and ( n7897 , n7886 , n7895 );
or ( n7898 , n7891 , n7896 , n7897 );
and ( n7899 , n7881 , n7898 );
and ( n7900 , n7861 , n7898 );
or ( n7901 , n7882 , n7899 , n7900 );
and ( n7902 , n7711 , n7865 );
not ( n7903 , n7902 );
xnor ( n7904 , n7903 , n5429 );
xor ( n7905 , n6423 , n7614 );
buf ( n7906 , n7905 );
buf ( n7907 , n7906 );
buf ( n7908 , n7907 );
and ( n7909 , n7904 , n7908 );
xor ( n7910 , n7653 , n7657 );
xor ( n7911 , n7910 , n7664 );
and ( n7912 , n7908 , n7911 );
and ( n7913 , n7904 , n7911 );
or ( n7914 , n7909 , n7912 , n7913 );
xor ( n7915 , n7901 , n7914 );
xor ( n7916 , n7828 , n7832 );
xor ( n7917 , n7916 , n7837 );
xor ( n7918 , n7801 , n7805 );
xor ( n7919 , n7918 , n7810 );
and ( n7920 , n7917 , n7919 );
xor ( n7921 , n7671 , n7674 );
xor ( n7922 , n7921 , n5405 );
and ( n7923 , n7919 , n7922 );
and ( n7924 , n7917 , n7922 );
or ( n7925 , n7920 , n7923 , n7924 );
xor ( n7926 , n7915 , n7925 );
xor ( n7927 , n5557 , n7644 );
xor ( n7928 , n7927 , n7705 );
and ( n7929 , n7926 , n7928 );
xor ( n7930 , n7917 , n7919 );
xor ( n7931 , n7930 , n7922 );
xor ( n7932 , n5514 , n5522 );
xor ( n7933 , n7932 , n5554 );
and ( n7934 , n7931 , n7933 );
xor ( n7935 , n5527 , n5533 );
xor ( n7936 , n7935 , n5551 );
and ( n7937 , n5296 , n7865 );
and ( n7938 , n5309 , n7863 );
nor ( n7939 , n7937 , n7938 );
xnor ( n7940 , n7939 , n5429 );
and ( n7941 , n5545 , n5282 );
and ( n7942 , n5355 , n5280 );
nor ( n7943 , n7941 , n7942 );
xnor ( n7944 , n7943 , n5290 );
and ( n7945 , n7940 , n7944 );
and ( n7946 , n7639 , n5365 );
and ( n7947 , n7690 , n5363 );
nor ( n7948 , n7946 , n7947 );
xnor ( n7949 , n7948 , n5373 );
and ( n7950 , n7944 , n7949 );
and ( n7951 , n7940 , n7949 );
or ( n7952 , n7945 , n7950 , n7951 );
and ( n7953 , n7647 , n5487 );
and ( n7954 , n7650 , n5485 );
nor ( n7955 , n7953 , n7954 );
xnor ( n7956 , n7955 , n5478 );
and ( n7957 , n5350 , n5306 );
and ( n7958 , n7716 , n5304 );
nor ( n7959 , n7957 , n7958 );
xnor ( n7960 , n7959 , n5314 );
and ( n7961 , n7956 , n7960 );
and ( n7962 , n5254 , n5325 );
and ( n7963 , n5265 , n5323 );
nor ( n7964 , n7962 , n7963 );
xnor ( n7965 , n7964 , n5333 );
and ( n7966 , n7960 , n7965 );
and ( n7967 , n7956 , n7965 );
or ( n7968 , n7961 , n7966 , n7967 );
xor ( n7969 , n7952 , n7968 );
xor ( n7970 , n7886 , n7890 );
xor ( n7971 , n7970 , n7895 );
xor ( n7972 , n7969 , n7971 );
and ( n7973 , n7936 , n7972 );
xor ( n7974 , n7849 , n7853 );
xor ( n7975 , n7974 , n7858 );
xor ( n7976 , n7869 , n7873 );
xor ( n7977 , n7976 , n7878 );
xnor ( n7978 , n7975 , n7977 );
and ( n7979 , n7972 , n7978 );
and ( n7980 , n7936 , n7978 );
or ( n7981 , n7973 , n7979 , n7980 );
and ( n7982 , n7933 , n7981 );
and ( n7983 , n7931 , n7981 );
or ( n7984 , n7934 , n7982 , n7983 );
and ( n7985 , n7928 , n7984 );
and ( n7986 , n7926 , n7984 );
or ( n7987 , n7929 , n7985 , n7986 );
and ( n7988 , n7845 , n7987 );
and ( n7989 , n5562 , n7620 );
and ( n7990 , n7620 , n7643 );
and ( n7991 , n5562 , n7643 );
or ( n7992 , n7989 , n7990 , n7991 );
and ( n7993 , n7667 , n7678 );
and ( n7994 , n7678 , n7704 );
and ( n7995 , n7667 , n7704 );
or ( n7996 , n7993 , n7994 , n7995 );
xor ( n7997 , n7992 , n7996 );
and ( n7998 , n7711 , n5487 );
not ( n7999 , n7998 );
xnor ( n8000 , n7999 , n5478 );
xor ( n8001 , n5252 , n5271 );
xor ( n8002 , n8001 , n5291 );
xor ( n8003 , n8000 , n8002 );
xor ( n8004 , n7997 , n8003 );
xor ( n8005 , n7861 , n7881 );
xor ( n8006 , n8005 , n7898 );
and ( n8007 , n7952 , n7968 );
and ( n8008 , n7968 , n7971 );
and ( n8009 , n7952 , n7971 );
or ( n8010 , n8007 , n8008 , n8009 );
and ( n8011 , n8006 , n8010 );
or ( n8012 , n7975 , n7977 );
and ( n8013 , n8010 , n8012 );
and ( n8014 , n8006 , n8012 );
or ( n8015 , n8011 , n8013 , n8014 );
and ( n8016 , n5340 , n7694 );
not ( n8017 , n8016 );
and ( n8018 , n8017 , n7702 );
xor ( n8019 , n6424 , n7613 );
buf ( n8020 , n8019 );
buf ( n8021 , n8020 );
buf ( n8022 , n8021 );
and ( n8023 , n8018 , n8022 );
and ( n8024 , n7711 , n5468 );
not ( n8025 , n8024 );
xnor ( n8026 , n8025 , n5405 );
and ( n8027 , n5317 , n7722 );
and ( n8028 , n5328 , n7720 );
nor ( n8029 , n8027 , n8028 );
xnor ( n8030 , n8029 , n7728 );
and ( n8031 , n8026 , n8030 );
and ( n8032 , n8030 , n8016 );
and ( n8033 , n8026 , n8016 );
or ( n8034 , n8031 , n8032 , n8033 );
and ( n8035 , n8022 , n8034 );
and ( n8036 , n8018 , n8034 );
or ( n8037 , n8023 , n8035 , n8036 );
and ( n8038 , n5437 , n5387 );
not ( n8039 , n8038 );
xnor ( n8040 , n8039 , n5382 );
and ( n8041 , n8040 , n5420 );
and ( n8042 , n5233 , n5499 );
and ( n8043 , n5246 , n5497 );
nor ( n8044 , n8042 , n8043 );
xnor ( n8045 , n8044 , n5505 );
and ( n8046 , n5420 , n8045 );
and ( n8047 , n8040 , n8045 );
or ( n8048 , n8041 , n8046 , n8047 );
and ( n8049 , n5274 , n5243 );
and ( n8050 , n5285 , n5241 );
nor ( n8051 , n8049 , n8050 );
xnor ( n8052 , n8051 , n5251 );
and ( n8053 , n5368 , n5262 );
and ( n8054 , n5529 , n5260 );
nor ( n8055 , n8053 , n8054 );
xnor ( n8056 , n8055 , n5270 );
and ( n8057 , n8052 , n8056 );
and ( n8058 , n7660 , n5542 );
and ( n8059 , n5536 , n5540 );
nor ( n8060 , n8058 , n8059 );
xnor ( n8061 , n8060 , n5550 );
and ( n8062 , n8056 , n8061 );
and ( n8063 , n8052 , n8061 );
or ( n8064 , n8057 , n8062 , n8063 );
and ( n8065 , n8048 , n8064 );
xor ( n8066 , n5518 , n5420 );
xor ( n8067 , n8066 , n5405 );
and ( n8068 , n8064 , n8067 );
and ( n8069 , n8048 , n8067 );
or ( n8070 , n8065 , n8068 , n8069 );
and ( n8071 , n8037 , n8070 );
xor ( n8072 , n7904 , n7908 );
xor ( n8073 , n8072 , n7911 );
and ( n8074 , n8070 , n8073 );
and ( n8075 , n8037 , n8073 );
or ( n8076 , n8071 , n8074 , n8075 );
and ( n8077 , n8015 , n8076 );
xor ( n8078 , n5443 , n5447 );
xor ( n8079 , n8078 , n5429 );
xor ( n8080 , n7813 , n7817 );
xor ( n8081 , n8080 , n7820 );
xor ( n8082 , n8079 , n8081 );
xnor ( n8083 , n7840 , n7842 );
xor ( n8084 , n8082 , n8083 );
and ( n8085 , n8076 , n8084 );
and ( n8086 , n8015 , n8084 );
or ( n8087 , n8077 , n8085 , n8086 );
xor ( n8088 , n8004 , n8087 );
xor ( n8089 , n5442 , n5451 );
xor ( n8090 , n8089 , n5454 );
and ( n8091 , n8079 , n8081 );
and ( n8092 , n8081 , n8083 );
and ( n8093 , n8079 , n8083 );
or ( n8094 , n8091 , n8092 , n8093 );
xor ( n8095 , n8090 , n8094 );
and ( n8096 , n7901 , n7914 );
and ( n8097 , n7914 , n7925 );
and ( n8098 , n7901 , n7925 );
or ( n8099 , n8096 , n8097 , n8098 );
xor ( n8100 , n8095 , n8099 );
xor ( n8101 , n8088 , n8100 );
and ( n8102 , n7987 , n8101 );
and ( n8103 , n7845 , n8101 );
or ( n8104 , n7988 , n8102 , n8103 );
xor ( n8105 , n5483 , n8104 );
and ( n8106 , n7797 , n7823 );
and ( n8107 , n7823 , n7843 );
and ( n8108 , n7797 , n7843 );
or ( n8109 , n8106 , n8107 , n8108 );
and ( n8110 , n7992 , n7996 );
and ( n8111 , n7996 , n8003 );
and ( n8112 , n7992 , n8003 );
or ( n8113 , n8110 , n8111 , n8112 );
xor ( n8114 , n8109 , n8113 );
and ( n8115 , n7746 , n7748 );
and ( n8116 , n7748 , n7763 );
and ( n8117 , n7746 , n7763 );
or ( n8118 , n8115 , n8116 , n8117 );
or ( n8119 , n7782 , n7796 );
xor ( n8120 , n8118 , n8119 );
and ( n8121 , n8000 , n8002 );
xor ( n8122 , n8120 , n8121 );
xor ( n8123 , n8114 , n8122 );
and ( n8124 , n8004 , n8087 );
and ( n8125 , n8087 , n8100 );
and ( n8126 , n8004 , n8100 );
or ( n8127 , n8124 , n8125 , n8126 );
xor ( n8128 , n8123 , n8127 );
and ( n8129 , n8090 , n8094 );
and ( n8130 , n8094 , n8099 );
and ( n8131 , n8090 , n8099 );
or ( n8132 , n8129 , n8130 , n8131 );
and ( n8133 , n7708 , n7765 );
and ( n8134 , n7765 , n7844 );
and ( n8135 , n7708 , n7844 );
or ( n8136 , n8133 , n8134 , n8135 );
xor ( n8137 , n8132 , n8136 );
and ( n8138 , n5309 , n5306 );
and ( n8139 , n7711 , n5304 );
nor ( n8140 , n8138 , n8139 );
xnor ( n8141 , n8140 , n5314 );
and ( n8142 , n7650 , n7722 );
and ( n8143 , n5296 , n7720 );
nor ( n8144 , n8142 , n8143 );
xnor ( n8145 , n8144 , n7728 );
xor ( n8146 , n8141 , n8145 );
and ( n8147 , n7716 , n5499 );
and ( n8148 , n7647 , n5497 );
nor ( n8149 , n8147 , n8148 );
xnor ( n8150 , n8149 , n5505 );
xor ( n8151 , n8146 , n8150 );
and ( n8152 , n5246 , n5243 );
and ( n8153 , n5317 , n5241 );
nor ( n8154 , n8152 , n8153 );
xnor ( n8155 , n8154 , n5251 );
and ( n8156 , n5529 , n5542 );
and ( n8157 , n5274 , n5540 );
nor ( n8158 , n8156 , n8157 );
xnor ( n8159 , n8158 , n5550 );
xor ( n8160 , n8155 , n8159 );
and ( n8161 , n7690 , n7633 );
and ( n8162 , n7660 , n5512 );
nor ( n8163 , n8161 , n8162 );
xnor ( n8164 , n8163 , n5561 );
xor ( n8165 , n8160 , n8164 );
xor ( n8166 , n8151 , n8165 );
and ( n8167 , n7786 , n7790 );
and ( n8168 , n7790 , n7795 );
and ( n8169 , n7786 , n7795 );
or ( n8170 , n8167 , n8168 , n8169 );
xor ( n8171 , n8166 , n8170 );
and ( n8172 , n7753 , n7757 );
and ( n8173 , n7757 , n7762 );
and ( n8174 , n7753 , n7762 );
or ( n8175 , n8172 , n8173 , n8174 );
not ( n8176 , n5382 );
and ( n8177 , n5265 , n5262 );
and ( n8178 , n5233 , n5260 );
nor ( n8179 , n8177 , n8178 );
xnor ( n8180 , n8179 , n5270 );
xor ( n8181 , n8176 , n8180 );
and ( n8182 , n5285 , n5282 );
and ( n8183 , n5254 , n5280 );
nor ( n8184 , n8182 , n8183 );
xnor ( n8185 , n8184 , n5290 );
xor ( n8186 , n8181 , n8185 );
xor ( n8187 , n8175 , n8186 );
and ( n8188 , n5536 , n7696 );
and ( n8189 , n5545 , n7694 );
nor ( n8190 , n8188 , n8189 );
xnor ( n8191 , n8190 , n7702 );
and ( n8192 , n7639 , n5342 );
xor ( n8193 , n8191 , n8192 );
xor ( n8194 , n8187 , n8193 );
xor ( n8195 , n8171 , n8194 );
and ( n8196 , n7737 , n7741 );
and ( n8197 , n7741 , n7764 );
and ( n8198 , n7737 , n7764 );
or ( n8199 , n8196 , n8197 , n8198 );
xor ( n8200 , n8195 , n8199 );
xor ( n8201 , n8137 , n8200 );
xor ( n8202 , n8128 , n8201 );
xor ( n8203 , n8105 , n8202 );
and ( n8204 , n5246 , n7722 );
and ( n8205 , n5317 , n7720 );
nor ( n8206 , n8204 , n8205 );
xnor ( n8207 , n8206 , n7728 );
and ( n8208 , n5265 , n5499 );
and ( n8209 , n5233 , n5497 );
nor ( n8210 , n8208 , n8209 );
xnor ( n8211 , n8210 , n5505 );
and ( n8212 , n8207 , n8211 );
and ( n8213 , n5340 , n5365 );
and ( n8214 , n7639 , n5363 );
nor ( n8215 , n8213 , n8214 );
xnor ( n8216 , n8215 , n5373 );
and ( n8217 , n8211 , n8216 );
and ( n8218 , n8207 , n8216 );
or ( n8219 , n8212 , n8217 , n8218 );
and ( n8220 , n5309 , n5468 );
and ( n8221 , n7711 , n5438 );
nor ( n8222 , n8220 , n8221 );
xnor ( n8223 , n8222 , n5405 );
and ( n8224 , n7650 , n7865 );
and ( n8225 , n5296 , n7863 );
nor ( n8226 , n8224 , n8225 );
xnor ( n8227 , n8226 , n5429 );
and ( n8228 , n8223 , n8227 );
and ( n8229 , n5285 , n5325 );
and ( n8230 , n5254 , n5323 );
nor ( n8231 , n8229 , n8230 );
xnor ( n8232 , n8231 , n5333 );
and ( n8233 , n8227 , n8232 );
and ( n8234 , n8223 , n8232 );
or ( n8235 , n8228 , n8233 , n8234 );
and ( n8236 , n8219 , n8235 );
xor ( n8237 , n8026 , n8030 );
xor ( n8238 , n8237 , n8016 );
and ( n8239 , n8235 , n8238 );
and ( n8240 , n8219 , n8238 );
or ( n8241 , n8236 , n8239 , n8240 );
and ( n8242 , n7716 , n5487 );
and ( n8243 , n7647 , n5485 );
nor ( n8244 , n8242 , n8243 );
xnor ( n8245 , n8244 , n5478 );
and ( n8246 , n5355 , n5262 );
and ( n8247 , n5368 , n5260 );
nor ( n8248 , n8246 , n8247 );
xnor ( n8249 , n8248 , n5270 );
and ( n8250 , n8245 , n8249 );
and ( n8251 , n7690 , n5542 );
and ( n8252 , n7660 , n5540 );
nor ( n8253 , n8251 , n8252 );
xnor ( n8254 , n8253 , n5550 );
and ( n8255 , n8249 , n8254 );
and ( n8256 , n8245 , n8254 );
or ( n8257 , n8250 , n8255 , n8256 );
xor ( n8258 , n7956 , n7960 );
xor ( n8259 , n8258 , n7965 );
or ( n8260 , n8257 , n8259 );
and ( n8261 , n8241 , n8260 );
xor ( n8262 , n6427 , n7611 );
buf ( n8263 , n8262 );
buf ( n8264 , n8263 );
buf ( n8265 , n8264 );
xor ( n8266 , n7940 , n7944 );
xor ( n8267 , n8266 , n7949 );
and ( n8268 , n8265 , n8267 );
and ( n8269 , n5382 , n5420 );
and ( n8270 , n5328 , n5306 );
and ( n8271 , n5350 , n5304 );
nor ( n8272 , n8270 , n8271 );
xnor ( n8273 , n8272 , n5314 );
and ( n8274 , n5420 , n8273 );
and ( n8275 , n5382 , n8273 );
or ( n8276 , n8269 , n8274 , n8275 );
and ( n8277 , n8267 , n8276 );
and ( n8278 , n8265 , n8276 );
or ( n8279 , n8268 , n8277 , n8278 );
and ( n8280 , n8260 , n8279 );
and ( n8281 , n8241 , n8279 );
or ( n8282 , n8261 , n8280 , n8281 );
and ( n8283 , n5529 , n5243 );
and ( n8284 , n5274 , n5241 );
nor ( n8285 , n8283 , n8284 );
xnor ( n8286 , n8285 , n5251 );
and ( n8287 , n5536 , n5282 );
and ( n8288 , n5545 , n5280 );
nor ( n8289 , n8287 , n8288 );
xnor ( n8290 , n8289 , n5290 );
and ( n8291 , n8286 , n8290 );
and ( n8292 , n5340 , n5363 );
not ( n8293 , n8292 );
and ( n8294 , n8293 , n5373 );
and ( n8295 , n8290 , n8294 );
and ( n8296 , n8286 , n8294 );
or ( n8297 , n8291 , n8295 , n8296 );
xor ( n8298 , n8040 , n5420 );
xor ( n8299 , n8298 , n8045 );
and ( n8300 , n8297 , n8299 );
xor ( n8301 , n8052 , n8056 );
xor ( n8302 , n8301 , n8061 );
and ( n8303 , n8299 , n8302 );
and ( n8304 , n8297 , n8302 );
or ( n8305 , n8300 , n8303 , n8304 );
xor ( n8306 , n8018 , n8022 );
xor ( n8307 , n8306 , n8034 );
and ( n8308 , n8305 , n8307 );
xor ( n8309 , n8048 , n8064 );
xor ( n8310 , n8309 , n8067 );
and ( n8311 , n8307 , n8310 );
and ( n8312 , n8305 , n8310 );
or ( n8313 , n8308 , n8311 , n8312 );
and ( n8314 , n8282 , n8313 );
xor ( n8315 , n8006 , n8010 );
xor ( n8316 , n8315 , n8012 );
and ( n8317 , n8313 , n8316 );
and ( n8318 , n8282 , n8316 );
or ( n8319 , n8314 , n8317 , n8318 );
xor ( n8320 , n8015 , n8076 );
xor ( n8321 , n8320 , n8084 );
and ( n8322 , n8319 , n8321 );
xor ( n8323 , n8037 , n8070 );
xor ( n8324 , n8323 , n8073 );
xor ( n8325 , n8219 , n8235 );
xor ( n8326 , n8325 , n8238 );
xnor ( n8327 , n8257 , n8259 );
and ( n8328 , n8326 , n8327 );
and ( n8329 , n5296 , n5468 );
and ( n8330 , n5309 , n5438 );
nor ( n8331 , n8329 , n8330 );
xnor ( n8332 , n8331 , n5405 );
and ( n8333 , n7647 , n7865 );
and ( n8334 , n7650 , n7863 );
nor ( n8335 , n8333 , n8334 );
xnor ( n8336 , n8335 , n5429 );
and ( n8337 , n8332 , n8336 );
and ( n8338 , n7639 , n5542 );
and ( n8339 , n7690 , n5540 );
nor ( n8340 , n8338 , n8339 );
xnor ( n8341 , n8340 , n5550 );
and ( n8342 , n8336 , n8341 );
and ( n8343 , n8332 , n8341 );
or ( n8344 , n8337 , n8342 , n8343 );
xor ( n8345 , n8223 , n8227 );
xor ( n8346 , n8345 , n8232 );
or ( n8347 , n8344 , n8346 );
and ( n8348 , n8327 , n8347 );
and ( n8349 , n8326 , n8347 );
or ( n8350 , n8328 , n8348 , n8349 );
xor ( n8351 , n6429 , n7610 );
buf ( n8352 , n8351 );
buf ( n8353 , n8352 );
buf ( n8354 , n8353 );
xor ( n8355 , n8207 , n8211 );
xor ( n8356 , n8355 , n8216 );
and ( n8357 , n8354 , n8356 );
xor ( n8358 , n8245 , n8249 );
xor ( n8359 , n8358 , n8254 );
and ( n8360 , n8356 , n8359 );
and ( n8361 , n8354 , n8359 );
or ( n8362 , n8357 , n8360 , n8361 );
and ( n8363 , n7711 , n5414 );
not ( n8364 , n8363 );
xnor ( n8365 , n8364 , n5420 );
and ( n8366 , n5233 , n7722 );
and ( n8367 , n5246 , n7720 );
nor ( n8368 , n8366 , n8367 );
xnor ( n8369 , n8368 , n7728 );
and ( n8370 , n8365 , n8369 );
and ( n8371 , n8369 , n8292 );
and ( n8372 , n8365 , n8292 );
or ( n8373 , n8370 , n8371 , n8372 );
and ( n8374 , n5317 , n5306 );
and ( n8375 , n5328 , n5304 );
nor ( n8376 , n8374 , n8375 );
xnor ( n8377 , n8376 , n5314 );
and ( n8378 , n5274 , n5325 );
and ( n8379 , n5285 , n5323 );
nor ( n8380 , n8378 , n8379 );
xnor ( n8381 , n8380 , n5333 );
or ( n8382 , n8377 , n8381 );
and ( n8383 , n8373 , n8382 );
and ( n8384 , n5350 , n5487 );
and ( n8385 , n7716 , n5485 );
nor ( n8386 , n8384 , n8385 );
xnor ( n8387 , n8386 , n5478 );
and ( n8388 , n7660 , n5282 );
and ( n8389 , n5536 , n5280 );
nor ( n8390 , n8388 , n8389 );
xnor ( n8391 , n8390 , n5290 );
and ( n8392 , n8387 , n8391 );
and ( n8393 , n8382 , n8392 );
and ( n8394 , n8373 , n8392 );
or ( n8395 , n8383 , n8393 , n8394 );
and ( n8396 , n8362 , n8395 );
and ( n8397 , n5254 , n5499 );
and ( n8398 , n5265 , n5497 );
nor ( n8399 , n8397 , n8398 );
xnor ( n8400 , n8399 , n5505 );
and ( n8401 , n5382 , n8400 );
and ( n8402 , n5368 , n5243 );
and ( n8403 , n5529 , n5241 );
nor ( n8404 , n8402 , n8403 );
xnor ( n8405 , n8404 , n5251 );
and ( n8406 , n8400 , n8405 );
and ( n8407 , n5382 , n8405 );
or ( n8408 , n8401 , n8406 , n8407 );
xor ( n8409 , n5382 , n5420 );
xor ( n8410 , n8409 , n8273 );
and ( n8411 , n8408 , n8410 );
xor ( n8412 , n8286 , n8290 );
xor ( n8413 , n8412 , n8294 );
and ( n8414 , n8410 , n8413 );
and ( n8415 , n8408 , n8413 );
or ( n8416 , n8411 , n8414 , n8415 );
and ( n8417 , n8395 , n8416 );
and ( n8418 , n8362 , n8416 );
or ( n8419 , n8396 , n8417 , n8418 );
and ( n8420 , n8350 , n8419 );
xor ( n8421 , n7936 , n7972 );
xor ( n8422 , n8421 , n7978 );
and ( n8423 , n8419 , n8422 );
and ( n8424 , n8350 , n8422 );
or ( n8425 , n8420 , n8423 , n8424 );
and ( n8426 , n8324 , n8425 );
xor ( n8427 , n7931 , n7933 );
xor ( n8428 , n8427 , n7981 );
and ( n8429 , n8425 , n8428 );
and ( n8430 , n8324 , n8428 );
or ( n8431 , n8426 , n8429 , n8430 );
and ( n8432 , n8321 , n8431 );
and ( n8433 , n8319 , n8431 );
or ( n8434 , n8322 , n8432 , n8433 );
xor ( n8435 , n7845 , n7987 );
xor ( n8436 , n8435 , n8101 );
and ( n8437 , n8434 , n8436 );
xor ( n8438 , n7926 , n7928 );
xor ( n8439 , n8438 , n7984 );
xor ( n8440 , n8282 , n8313 );
xor ( n8441 , n8440 , n8316 );
xor ( n8442 , n8241 , n8260 );
xor ( n8443 , n8442 , n8279 );
xor ( n8444 , n8305 , n8307 );
xor ( n8445 , n8444 , n8310 );
and ( n8446 , n8443 , n8445 );
xor ( n8447 , n8265 , n8267 );
xor ( n8448 , n8447 , n8276 );
xor ( n8449 , n8297 , n8299 );
xor ( n8450 , n8449 , n8302 );
and ( n8451 , n8448 , n8450 );
xnor ( n8452 , n8344 , n8346 );
and ( n8453 , n5545 , n5262 );
and ( n8454 , n5355 , n5260 );
nor ( n8455 , n8453 , n8454 );
xnor ( n8456 , n8455 , n5270 );
xor ( n8457 , n6430 , n7609 );
buf ( n8458 , n8457 );
buf ( n8459 , n8458 );
buf ( n8460 , n8459 );
and ( n8461 , n8456 , n8460 );
xor ( n8462 , n8365 , n8369 );
xor ( n8463 , n8462 , n8292 );
and ( n8464 , n8460 , n8463 );
and ( n8465 , n8456 , n8463 );
or ( n8466 , n8461 , n8464 , n8465 );
and ( n8467 , n8452 , n8466 );
xor ( n8468 , n8332 , n8336 );
xor ( n8469 , n8468 , n8341 );
xnor ( n8470 , n8377 , n8381 );
and ( n8471 , n8469 , n8470 );
xor ( n8472 , n8387 , n8391 );
and ( n8473 , n8470 , n8472 );
and ( n8474 , n8469 , n8472 );
or ( n8475 , n8471 , n8473 , n8474 );
and ( n8476 , n8466 , n8475 );
and ( n8477 , n8452 , n8475 );
or ( n8478 , n8467 , n8476 , n8477 );
and ( n8479 , n8450 , n8478 );
and ( n8480 , n8448 , n8478 );
or ( n8481 , n8451 , n8479 , n8480 );
and ( n8482 , n8445 , n8481 );
and ( n8483 , n8443 , n8481 );
or ( n8484 , n8446 , n8482 , n8483 );
and ( n8485 , n8441 , n8484 );
xor ( n8486 , n8324 , n8425 );
xor ( n8487 , n8486 , n8428 );
and ( n8488 , n8484 , n8487 );
and ( n8489 , n8441 , n8487 );
or ( n8490 , n8485 , n8488 , n8489 );
and ( n8491 , n8439 , n8490 );
xor ( n8492 , n8319 , n8321 );
xor ( n8493 , n8492 , n8431 );
and ( n8494 , n8490 , n8493 );
and ( n8495 , n8439 , n8493 );
or ( n8496 , n8491 , n8494 , n8495 );
and ( n8497 , n8436 , n8496 );
and ( n8498 , n8434 , n8496 );
or ( n8499 , n8437 , n8497 , n8498 );
xnor ( n8500 , n8203 , n8499 );
xor ( n8501 , n8434 , n8436 );
xor ( n8502 , n8501 , n8496 );
xor ( n8503 , n8439 , n8490 );
xor ( n8504 , n8503 , n8493 );
and ( n8505 , n5328 , n5487 );
and ( n8506 , n5350 , n5485 );
nor ( n8507 , n8505 , n8506 );
xnor ( n8508 , n8507 , n5478 );
and ( n8509 , n5529 , n5325 );
and ( n8510 , n5274 , n5323 );
nor ( n8511 , n8509 , n8510 );
xnor ( n8512 , n8511 , n5333 );
and ( n8513 , n8508 , n8512 );
and ( n8514 , n7690 , n5282 );
and ( n8515 , n7660 , n5280 );
nor ( n8516 , n8514 , n8515 );
xnor ( n8517 , n8516 , n5290 );
and ( n8518 , n8512 , n8517 );
and ( n8519 , n8508 , n8517 );
or ( n8520 , n8513 , n8518 , n8519 );
and ( n8521 , n5355 , n5243 );
and ( n8522 , n5368 , n5241 );
nor ( n8523 , n8521 , n8522 );
xnor ( n8524 , n8523 , n5251 );
and ( n8525 , n5536 , n5262 );
and ( n8526 , n5545 , n5260 );
nor ( n8527 , n8525 , n8526 );
xnor ( n8528 , n8527 , n5270 );
and ( n8529 , n8524 , n8528 );
and ( n8530 , n5340 , n5542 );
and ( n8531 , n7639 , n5540 );
nor ( n8532 , n8530 , n8531 );
xnor ( n8533 , n8532 , n5550 );
and ( n8534 , n8528 , n8533 );
and ( n8535 , n8524 , n8533 );
or ( n8536 , n8529 , n8534 , n8535 );
and ( n8537 , n8520 , n8536 );
and ( n8538 , n7650 , n5468 );
and ( n8539 , n5296 , n5438 );
nor ( n8540 , n8538 , n8539 );
xnor ( n8541 , n8540 , n5405 );
and ( n8542 , n5340 , n5540 );
not ( n8543 , n8542 );
and ( n8544 , n8543 , n5550 );
or ( n8545 , n8541 , n8544 );
and ( n8546 , n8536 , n8545 );
and ( n8547 , n8520 , n8545 );
or ( n8548 , n8537 , n8546 , n8547 );
and ( n8549 , n5246 , n5306 );
and ( n8550 , n5317 , n5304 );
nor ( n8551 , n8549 , n8550 );
xnor ( n8552 , n8551 , n5314 );
and ( n8553 , n5265 , n7722 );
and ( n8554 , n5233 , n7720 );
nor ( n8555 , n8553 , n8554 );
xnor ( n8556 , n8555 , n7728 );
or ( n8557 , n8552 , n8556 );
and ( n8558 , n5309 , n5414 );
and ( n8559 , n7711 , n5412 );
nor ( n8560 , n8558 , n8559 );
xnor ( n8561 , n8560 , n5420 );
and ( n8562 , n7716 , n7865 );
and ( n8563 , n7647 , n7863 );
nor ( n8564 , n8562 , n8563 );
xnor ( n8565 , n8564 , n5429 );
or ( n8566 , n8561 , n8565 );
and ( n8567 , n8557 , n8566 );
and ( n8568 , n5285 , n5499 );
and ( n8569 , n5254 , n5497 );
nor ( n8570 , n8568 , n8569 );
xnor ( n8571 , n8570 , n5505 );
and ( n8572 , n5382 , n8571 );
xor ( n8573 , n6431 , n7608 );
buf ( n8574 , n8573 );
buf ( n8575 , n8574 );
buf ( n8576 , n8575 );
and ( n8577 , n8571 , n8576 );
and ( n8578 , n5382 , n8576 );
or ( n8579 , n8572 , n8577 , n8578 );
and ( n8580 , n8566 , n8579 );
and ( n8581 , n8557 , n8579 );
or ( n8582 , n8567 , n8580 , n8581 );
and ( n8583 , n8548 , n8582 );
xor ( n8584 , n8354 , n8356 );
xor ( n8585 , n8584 , n8359 );
and ( n8586 , n8582 , n8585 );
and ( n8587 , n8548 , n8585 );
or ( n8588 , n8583 , n8586 , n8587 );
xor ( n8589 , n8326 , n8327 );
xor ( n8590 , n8589 , n8347 );
and ( n8591 , n8588 , n8590 );
xor ( n8592 , n8362 , n8395 );
xor ( n8593 , n8592 , n8416 );
and ( n8594 , n8590 , n8593 );
and ( n8595 , n8588 , n8593 );
or ( n8596 , n8591 , n8594 , n8595 );
xor ( n8597 , n8350 , n8419 );
xor ( n8598 , n8597 , n8422 );
and ( n8599 , n8596 , n8598 );
xor ( n8600 , n8373 , n8382 );
xor ( n8601 , n8600 , n8392 );
xor ( n8602 , n8408 , n8410 );
xor ( n8603 , n8602 , n8413 );
and ( n8604 , n8601 , n8603 );
xor ( n8605 , n5382 , n8400 );
xor ( n8606 , n8605 , n8405 );
and ( n8607 , n7711 , n5390 );
not ( n8608 , n8607 );
xnor ( n8609 , n8608 , n5382 );
and ( n8610 , n5317 , n5487 );
and ( n8611 , n5328 , n5485 );
nor ( n8612 , n8610 , n8611 );
xnor ( n8613 , n8612 , n5478 );
and ( n8614 , n8609 , n8613 );
and ( n8615 , n8613 , n8542 );
and ( n8616 , n8609 , n8542 );
or ( n8617 , n8614 , n8615 , n8616 );
and ( n8618 , n7647 , n5468 );
and ( n8619 , n7650 , n5438 );
nor ( n8620 , n8618 , n8619 );
xnor ( n8621 , n8620 , n5405 );
and ( n8622 , n5368 , n5325 );
and ( n8623 , n5529 , n5323 );
nor ( n8624 , n8622 , n8623 );
xnor ( n8625 , n8624 , n5333 );
and ( n8626 , n8621 , n8625 );
and ( n8627 , n7639 , n5282 );
and ( n8628 , n7690 , n5280 );
nor ( n8629 , n8627 , n8628 );
xnor ( n8630 , n8629 , n5290 );
and ( n8631 , n8625 , n8630 );
and ( n8632 , n8621 , n8630 );
or ( n8633 , n8626 , n8631 , n8632 );
and ( n8634 , n8617 , n8633 );
and ( n8635 , n8606 , n8634 );
xor ( n8636 , n8508 , n8512 );
xor ( n8637 , n8636 , n8517 );
xor ( n8638 , n8524 , n8528 );
xor ( n8639 , n8638 , n8533 );
and ( n8640 , n8637 , n8639 );
xnor ( n8641 , n8541 , n8544 );
and ( n8642 , n8639 , n8641 );
and ( n8643 , n8637 , n8641 );
or ( n8644 , n8640 , n8642 , n8643 );
and ( n8645 , n8634 , n8644 );
and ( n8646 , n8606 , n8644 );
or ( n8647 , n8635 , n8645 , n8646 );
and ( n8648 , n8603 , n8647 );
and ( n8649 , n8601 , n8647 );
or ( n8650 , n8604 , n8648 , n8649 );
xnor ( n8651 , n8552 , n8556 );
xnor ( n8652 , n8561 , n8565 );
and ( n8653 , n8651 , n8652 );
and ( n8654 , n5296 , n5414 );
and ( n8655 , n5309 , n5412 );
nor ( n8656 , n8654 , n8655 );
xnor ( n8657 , n8656 , n5420 );
and ( n8658 , n5350 , n7865 );
and ( n8659 , n7716 , n7863 );
nor ( n8660 , n8658 , n8659 );
xnor ( n8661 , n8660 , n5429 );
and ( n8662 , n8657 , n8661 );
and ( n8663 , n5233 , n5306 );
and ( n8664 , n5246 , n5304 );
nor ( n8665 , n8663 , n8664 );
xnor ( n8666 , n8665 , n5314 );
and ( n8667 , n8661 , n8666 );
and ( n8668 , n8657 , n8666 );
or ( n8669 , n8662 , n8667 , n8668 );
and ( n8670 , n8652 , n8669 );
and ( n8671 , n8651 , n8669 );
or ( n8672 , n8653 , n8670 , n8671 );
xor ( n8673 , n8456 , n8460 );
xor ( n8674 , n8673 , n8463 );
and ( n8675 , n8672 , n8674 );
xor ( n8676 , n8469 , n8470 );
xor ( n8677 , n8676 , n8472 );
and ( n8678 , n8674 , n8677 );
and ( n8679 , n8672 , n8677 );
or ( n8680 , n8675 , n8678 , n8679 );
xor ( n8681 , n8452 , n8466 );
xor ( n8682 , n8681 , n8475 );
and ( n8683 , n8680 , n8682 );
xor ( n8684 , n8548 , n8582 );
xor ( n8685 , n8684 , n8585 );
and ( n8686 , n8682 , n8685 );
and ( n8687 , n8680 , n8685 );
or ( n8688 , n8683 , n8686 , n8687 );
and ( n8689 , n8650 , n8688 );
xor ( n8690 , n8448 , n8450 );
xor ( n8691 , n8690 , n8478 );
and ( n8692 , n8688 , n8691 );
and ( n8693 , n8650 , n8691 );
or ( n8694 , n8689 , n8692 , n8693 );
and ( n8695 , n8598 , n8694 );
and ( n8696 , n8596 , n8694 );
or ( n8697 , n8599 , n8695 , n8696 );
xor ( n8698 , n8441 , n8484 );
xor ( n8699 , n8698 , n8487 );
and ( n8700 , n8697 , n8699 );
xor ( n8701 , n8443 , n8445 );
xor ( n8702 , n8701 , n8481 );
xor ( n8703 , n8588 , n8590 );
xor ( n8704 , n8703 , n8593 );
xor ( n8705 , n8520 , n8536 );
xor ( n8706 , n8705 , n8545 );
xor ( n8707 , n8557 , n8566 );
xor ( n8708 , n8707 , n8579 );
and ( n8709 , n8706 , n8708 );
and ( n8710 , n5254 , n7722 );
and ( n8711 , n5265 , n7720 );
nor ( n8712 , n8710 , n8711 );
xnor ( n8713 , n8712 , n7728 );
and ( n8714 , n5274 , n5499 );
and ( n8715 , n5285 , n5497 );
nor ( n8716 , n8714 , n8715 );
xnor ( n8717 , n8716 , n5505 );
and ( n8718 , n8713 , n8717 );
and ( n8719 , n5545 , n5243 );
and ( n8720 , n5355 , n5241 );
nor ( n8721 , n8719 , n8720 );
xnor ( n8722 , n8721 , n5251 );
and ( n8723 , n8717 , n8722 );
and ( n8724 , n8713 , n8722 );
or ( n8725 , n8718 , n8723 , n8724 );
xor ( n8726 , n5382 , n8571 );
xor ( n8727 , n8726 , n8576 );
and ( n8728 , n8725 , n8727 );
xor ( n8729 , n8617 , n8633 );
and ( n8730 , n8727 , n8729 );
and ( n8731 , n8725 , n8729 );
or ( n8732 , n8728 , n8730 , n8731 );
and ( n8733 , n8708 , n8732 );
and ( n8734 , n8706 , n8732 );
or ( n8735 , n8709 , n8733 , n8734 );
and ( n8736 , n7660 , n5262 );
and ( n8737 , n5536 , n5260 );
nor ( n8738 , n8736 , n8737 );
xnor ( n8739 , n8738 , n5270 );
xor ( n8740 , n6434 , n7606 );
buf ( n8741 , n8740 );
buf ( n8742 , n8741 );
buf ( n8743 , n8742 );
and ( n8744 , n8739 , n8743 );
xor ( n8745 , n8609 , n8613 );
xor ( n8746 , n8745 , n8542 );
and ( n8747 , n8743 , n8746 );
and ( n8748 , n8739 , n8746 );
or ( n8749 , n8744 , n8747 , n8748 );
xor ( n8750 , n8621 , n8625 );
xor ( n8751 , n8750 , n8630 );
and ( n8752 , n7716 , n5468 );
and ( n8753 , n7647 , n5438 );
nor ( n8754 , n8752 , n8753 );
xnor ( n8755 , n8754 , n5405 );
and ( n8756 , n7690 , n5262 );
and ( n8757 , n7660 , n5260 );
nor ( n8758 , n8756 , n8757 );
xnor ( n8759 , n8758 , n5270 );
and ( n8760 , n8755 , n8759 );
and ( n8761 , n5340 , n5282 );
and ( n8762 , n7639 , n5280 );
nor ( n8763 , n8761 , n8762 );
xnor ( n8764 , n8763 , n5290 );
and ( n8765 , n8759 , n8764 );
and ( n8766 , n8755 , n8764 );
or ( n8767 , n8760 , n8765 , n8766 );
and ( n8768 , n8751 , n8767 );
and ( n8769 , n5309 , n5390 );
and ( n8770 , n7711 , n5387 );
nor ( n8771 , n8769 , n8770 );
xnor ( n8772 , n8771 , n5382 );
and ( n8773 , n7650 , n5414 );
and ( n8774 , n5296 , n5412 );
nor ( n8775 , n8773 , n8774 );
xnor ( n8776 , n8775 , n5420 );
and ( n8777 , n8772 , n8776 );
and ( n8778 , n5328 , n7865 );
and ( n8779 , n5350 , n7863 );
nor ( n8780 , n8778 , n8779 );
xnor ( n8781 , n8780 , n5429 );
and ( n8782 , n8776 , n8781 );
and ( n8783 , n8772 , n8781 );
or ( n8784 , n8777 , n8782 , n8783 );
and ( n8785 , n8767 , n8784 );
and ( n8786 , n8751 , n8784 );
or ( n8787 , n8768 , n8785 , n8786 );
and ( n8788 , n8749 , n8787 );
and ( n8789 , n5246 , n5487 );
and ( n8790 , n5317 , n5485 );
nor ( n8791 , n8789 , n8790 );
xnor ( n8792 , n8791 , n5478 );
and ( n8793 , n5265 , n5306 );
and ( n8794 , n5233 , n5304 );
nor ( n8795 , n8793 , n8794 );
xnor ( n8796 , n8795 , n5314 );
and ( n8797 , n8792 , n8796 );
and ( n8798 , n5285 , n7722 );
and ( n8799 , n5254 , n7720 );
nor ( n8800 , n8798 , n8799 );
xnor ( n8801 , n8800 , n7728 );
and ( n8802 , n8796 , n8801 );
and ( n8803 , n8792 , n8801 );
or ( n8804 , n8797 , n8802 , n8803 );
and ( n8805 , n5529 , n5499 );
and ( n8806 , n5274 , n5497 );
nor ( n8807 , n8805 , n8806 );
xnor ( n8808 , n8807 , n5505 );
and ( n8809 , n5355 , n5325 );
and ( n8810 , n5368 , n5323 );
nor ( n8811 , n8809 , n8810 );
xnor ( n8812 , n8811 , n5333 );
and ( n8813 , n8808 , n8812 );
and ( n8814 , n5536 , n5243 );
and ( n8815 , n5545 , n5241 );
nor ( n8816 , n8814 , n8815 );
xnor ( n8817 , n8816 , n5251 );
and ( n8818 , n8812 , n8817 );
and ( n8819 , n8808 , n8817 );
or ( n8820 , n8813 , n8818 , n8819 );
and ( n8821 , n8804 , n8820 );
xor ( n8822 , n8657 , n8661 );
xor ( n8823 , n8822 , n8666 );
and ( n8824 , n8820 , n8823 );
and ( n8825 , n8804 , n8823 );
or ( n8826 , n8821 , n8824 , n8825 );
and ( n8827 , n8787 , n8826 );
and ( n8828 , n8749 , n8826 );
or ( n8829 , n8788 , n8827 , n8828 );
xor ( n8830 , n8606 , n8634 );
xor ( n8831 , n8830 , n8644 );
and ( n8832 , n8829 , n8831 );
xor ( n8833 , n8672 , n8674 );
xor ( n8834 , n8833 , n8677 );
and ( n8835 , n8831 , n8834 );
and ( n8836 , n8829 , n8834 );
or ( n8837 , n8832 , n8835 , n8836 );
and ( n8838 , n8735 , n8837 );
xor ( n8839 , n8601 , n8603 );
xor ( n8840 , n8839 , n8647 );
and ( n8841 , n8837 , n8840 );
and ( n8842 , n8735 , n8840 );
or ( n8843 , n8838 , n8841 , n8842 );
and ( n8844 , n8704 , n8843 );
xor ( n8845 , n8650 , n8688 );
xor ( n8846 , n8845 , n8691 );
and ( n8847 , n8843 , n8846 );
and ( n8848 , n8704 , n8846 );
or ( n8849 , n8844 , n8847 , n8848 );
and ( n8850 , n8702 , n8849 );
xor ( n8851 , n8596 , n8598 );
xor ( n8852 , n8851 , n8694 );
and ( n8853 , n8849 , n8852 );
and ( n8854 , n8702 , n8852 );
or ( n8855 , n8850 , n8853 , n8854 );
and ( n8856 , n8699 , n8855 );
and ( n8857 , n8697 , n8855 );
or ( n8858 , n8700 , n8856 , n8857 );
and ( n8859 , n8504 , n8858 );
xor ( n8860 , n8504 , n8858 );
xor ( n8861 , n8697 , n8699 );
xor ( n8862 , n8861 , n8855 );
xor ( n8863 , n8702 , n8849 );
xor ( n8864 , n8863 , n8852 );
xor ( n8865 , n8680 , n8682 );
xor ( n8866 , n8865 , n8685 );
xor ( n8867 , n8637 , n8639 );
xor ( n8868 , n8867 , n8641 );
xor ( n8869 , n8651 , n8652 );
xor ( n8870 , n8869 , n8669 );
and ( n8871 , n8868 , n8870 );
xor ( n8872 , n8713 , n8717 );
xor ( n8873 , n8872 , n8722 );
and ( n8874 , n5340 , n5280 );
not ( n8875 , n8874 );
and ( n8876 , n8875 , n5290 );
xor ( n8877 , n7268 , n7604 );
buf ( n8878 , n8877 );
buf ( n8879 , n8878 );
buf ( n8880 , n8879 );
and ( n8881 , n8876 , n8880 );
xor ( n8882 , n8755 , n8759 );
xor ( n8883 , n8882 , n8764 );
and ( n8884 , n8880 , n8883 );
and ( n8885 , n8876 , n8883 );
or ( n8886 , n8881 , n8884 , n8885 );
and ( n8887 , n8873 , n8886 );
and ( n8888 , n5296 , n5390 );
and ( n8889 , n5309 , n5387 );
nor ( n8890 , n8888 , n8889 );
xnor ( n8891 , n8890 , n5382 );
and ( n8892 , n5350 , n5468 );
and ( n8893 , n7716 , n5438 );
nor ( n8894 , n8892 , n8893 );
xnor ( n8895 , n8894 , n5405 );
and ( n8896 , n8891 , n8895 );
and ( n8897 , n5545 , n5325 );
and ( n8898 , n5355 , n5323 );
nor ( n8899 , n8897 , n8898 );
xnor ( n8900 , n8899 , n5333 );
and ( n8901 , n8895 , n8900 );
and ( n8902 , n8891 , n8900 );
or ( n8903 , n8896 , n8901 , n8902 );
and ( n8904 , n7660 , n5243 );
and ( n8905 , n5536 , n5241 );
nor ( n8906 , n8904 , n8905 );
xnor ( n8907 , n8906 , n5251 );
and ( n8908 , n7639 , n5262 );
and ( n8909 , n7690 , n5260 );
nor ( n8910 , n8908 , n8909 );
xnor ( n8911 , n8910 , n5270 );
and ( n8912 , n8907 , n8911 );
and ( n8913 , n8903 , n8912 );
and ( n8914 , n7647 , n5414 );
and ( n8915 , n7650 , n5412 );
nor ( n8916 , n8914 , n8915 );
xnor ( n8917 , n8916 , n5420 );
and ( n8918 , n5317 , n7865 );
and ( n8919 , n5328 , n7863 );
nor ( n8920 , n8918 , n8919 );
xnor ( n8921 , n8920 , n5429 );
and ( n8922 , n8917 , n8921 );
and ( n8923 , n5233 , n5487 );
and ( n8924 , n5246 , n5485 );
nor ( n8925 , n8923 , n8924 );
xnor ( n8926 , n8925 , n5478 );
and ( n8927 , n8921 , n8926 );
and ( n8928 , n8917 , n8926 );
or ( n8929 , n8922 , n8927 , n8928 );
and ( n8930 , n8912 , n8929 );
and ( n8931 , n8903 , n8929 );
or ( n8932 , n8913 , n8930 , n8931 );
and ( n8933 , n8886 , n8932 );
and ( n8934 , n8873 , n8932 );
or ( n8935 , n8887 , n8933 , n8934 );
and ( n8936 , n8870 , n8935 );
and ( n8937 , n8868 , n8935 );
or ( n8938 , n8871 , n8936 , n8937 );
and ( n8939 , n5254 , n5306 );
and ( n8940 , n5265 , n5304 );
nor ( n8941 , n8939 , n8940 );
xnor ( n8942 , n8941 , n5314 );
and ( n8943 , n5274 , n7722 );
and ( n8944 , n5285 , n7720 );
nor ( n8945 , n8943 , n8944 );
xnor ( n8946 , n8945 , n7728 );
and ( n8947 , n8942 , n8946 );
and ( n8948 , n5368 , n5499 );
and ( n8949 , n5529 , n5497 );
nor ( n8950 , n8948 , n8949 );
xnor ( n8951 , n8950 , n5505 );
and ( n8952 , n8946 , n8951 );
and ( n8953 , n8942 , n8951 );
or ( n8954 , n8947 , n8952 , n8953 );
xor ( n8955 , n8772 , n8776 );
xor ( n8956 , n8955 , n8781 );
and ( n8957 , n8954 , n8956 );
xor ( n8958 , n8792 , n8796 );
xor ( n8959 , n8958 , n8801 );
and ( n8960 , n8956 , n8959 );
and ( n8961 , n8954 , n8959 );
or ( n8962 , n8957 , n8960 , n8961 );
xor ( n8963 , n8739 , n8743 );
xor ( n8964 , n8963 , n8746 );
and ( n8965 , n8962 , n8964 );
xor ( n8966 , n8751 , n8767 );
xor ( n8967 , n8966 , n8784 );
and ( n8968 , n8964 , n8967 );
and ( n8969 , n8962 , n8967 );
or ( n8970 , n8965 , n8968 , n8969 );
xor ( n8971 , n8725 , n8727 );
xor ( n8972 , n8971 , n8729 );
and ( n8973 , n8970 , n8972 );
xor ( n8974 , n8749 , n8787 );
xor ( n8975 , n8974 , n8826 );
and ( n8976 , n8972 , n8975 );
and ( n8977 , n8970 , n8975 );
or ( n8978 , n8973 , n8976 , n8977 );
and ( n8979 , n8938 , n8978 );
xor ( n8980 , n8706 , n8708 );
xor ( n8981 , n8980 , n8732 );
and ( n8982 , n8978 , n8981 );
and ( n8983 , n8938 , n8981 );
or ( n8984 , n8979 , n8982 , n8983 );
and ( n8985 , n8866 , n8984 );
xor ( n8986 , n8735 , n8837 );
xor ( n8987 , n8986 , n8840 );
and ( n8988 , n8984 , n8987 );
and ( n8989 , n8866 , n8987 );
or ( n8990 , n8985 , n8988 , n8989 );
xor ( n8991 , n8704 , n8843 );
xor ( n8992 , n8991 , n8846 );
and ( n8993 , n8990 , n8992 );
xor ( n8994 , n8829 , n8831 );
xor ( n8995 , n8994 , n8834 );
xor ( n8996 , n8804 , n8820 );
xor ( n8997 , n8996 , n8823 );
xor ( n8998 , n8808 , n8812 );
xor ( n8999 , n8998 , n8817 );
xor ( n9000 , n7271 , n7602 );
buf ( n9001 , n9000 );
buf ( n9002 , n9001 );
buf ( n9003 , n9002 );
and ( n9004 , n8874 , n9003 );
xor ( n9005 , n8907 , n8911 );
and ( n9006 , n9003 , n9005 );
and ( n9007 , n8874 , n9005 );
or ( n9008 , n9004 , n9006 , n9007 );
and ( n9009 , n8999 , n9008 );
and ( n9010 , n7716 , n5414 );
and ( n9011 , n7647 , n5412 );
nor ( n9012 , n9010 , n9011 );
xnor ( n9013 , n9012 , n5420 );
and ( n9014 , n5328 , n5468 );
and ( n9015 , n5350 , n5438 );
nor ( n9016 , n9014 , n9015 );
xnor ( n9017 , n9016 , n5405 );
and ( n9018 , n9013 , n9017 );
and ( n9019 , n5536 , n5325 );
and ( n9020 , n5545 , n5323 );
nor ( n9021 , n9019 , n9020 );
xnor ( n9022 , n9021 , n5333 );
and ( n9023 , n9017 , n9022 );
and ( n9024 , n9013 , n9022 );
or ( n9025 , n9018 , n9023 , n9024 );
and ( n9026 , n5285 , n5306 );
and ( n9027 , n5254 , n5304 );
nor ( n9028 , n9026 , n9027 );
xnor ( n9029 , n9028 , n5314 );
and ( n9030 , n5529 , n7722 );
and ( n9031 , n5274 , n7720 );
nor ( n9032 , n9030 , n9031 );
xnor ( n9033 , n9032 , n7728 );
and ( n9034 , n9029 , n9033 );
and ( n9035 , n5355 , n5499 );
and ( n9036 , n5368 , n5497 );
nor ( n9037 , n9035 , n9036 );
xnor ( n9038 , n9037 , n5505 );
and ( n9039 , n9033 , n9038 );
and ( n9040 , n9029 , n9038 );
or ( n9041 , n9034 , n9039 , n9040 );
and ( n9042 , n9025 , n9041 );
and ( n9043 , n5265 , n5487 );
and ( n9044 , n5233 , n5485 );
nor ( n9045 , n9043 , n9044 );
xnor ( n9046 , n9045 , n5478 );
and ( n9047 , n7690 , n5243 );
and ( n9048 , n7660 , n5241 );
nor ( n9049 , n9047 , n9048 );
xnor ( n9050 , n9049 , n5251 );
and ( n9051 , n9046 , n9050 );
xor ( n9052 , n7273 , n7601 );
buf ( n9053 , n9052 );
buf ( n9054 , n9053 );
buf ( n9055 , n9054 );
and ( n9056 , n9050 , n9055 );
and ( n9057 , n9046 , n9055 );
or ( n9058 , n9051 , n9056 , n9057 );
and ( n9059 , n9041 , n9058 );
and ( n9060 , n9025 , n9058 );
or ( n9061 , n9042 , n9059 , n9060 );
and ( n9062 , n9008 , n9061 );
and ( n9063 , n8999 , n9061 );
or ( n9064 , n9009 , n9062 , n9063 );
and ( n9065 , n8997 , n9064 );
xor ( n9066 , n8876 , n8880 );
xor ( n9067 , n9066 , n8883 );
xor ( n9068 , n8903 , n8912 );
xor ( n9069 , n9068 , n8929 );
and ( n9070 , n9067 , n9069 );
xor ( n9071 , n8954 , n8956 );
xor ( n9072 , n9071 , n8959 );
and ( n9073 , n9069 , n9072 );
and ( n9074 , n9067 , n9072 );
or ( n9075 , n9070 , n9073 , n9074 );
and ( n9076 , n9064 , n9075 );
and ( n9077 , n8997 , n9075 );
or ( n9078 , n9065 , n9076 , n9077 );
xor ( n9079 , n8868 , n8870 );
xor ( n9080 , n9079 , n8935 );
and ( n9081 , n9078 , n9080 );
xor ( n9082 , n8970 , n8972 );
xor ( n9083 , n9082 , n8975 );
and ( n9084 , n9080 , n9083 );
and ( n9085 , n9078 , n9083 );
or ( n9086 , n9081 , n9084 , n9085 );
and ( n9087 , n8995 , n9086 );
xor ( n9088 , n8938 , n8978 );
xor ( n9089 , n9088 , n8981 );
and ( n9090 , n9086 , n9089 );
and ( n9091 , n8995 , n9089 );
or ( n9092 , n9087 , n9090 , n9091 );
xor ( n9093 , n8866 , n8984 );
xor ( n9094 , n9093 , n8987 );
and ( n9095 , n9092 , n9094 );
xor ( n9096 , n8995 , n9086 );
xor ( n9097 , n9096 , n9089 );
xor ( n9098 , n8873 , n8886 );
xor ( n9099 , n9098 , n8932 );
xor ( n9100 , n8962 , n8964 );
xor ( n9101 , n9100 , n8967 );
and ( n9102 , n9099 , n9101 );
and ( n9103 , n5254 , n5487 );
and ( n9104 , n5265 , n5485 );
nor ( n9105 , n9103 , n9104 );
xnor ( n9106 , n9105 , n5478 );
and ( n9107 , n5368 , n7722 );
and ( n9108 , n5529 , n7720 );
nor ( n9109 , n9107 , n9108 );
xnor ( n9110 , n9109 , n7728 );
and ( n9111 , n9106 , n9110 );
and ( n9112 , n5545 , n5499 );
and ( n9113 , n5355 , n5497 );
nor ( n9114 , n9112 , n9113 );
xnor ( n9115 , n9114 , n5505 );
and ( n9116 , n9110 , n9115 );
and ( n9117 , n9106 , n9115 );
or ( n9118 , n9111 , n9116 , n9117 );
and ( n9119 , n5246 , n7865 );
and ( n9120 , n5317 , n7863 );
nor ( n9121 , n9119 , n9120 );
xnor ( n9122 , n9121 , n5429 );
and ( n9123 , n9118 , n9122 );
and ( n9124 , n5340 , n5260 );
not ( n9125 , n9124 );
and ( n9126 , n9125 , n5270 );
and ( n9127 , n9122 , n9126 );
and ( n9128 , n9118 , n9126 );
or ( n9129 , n9123 , n9127 , n9128 );
and ( n9130 , n7650 , n5390 );
and ( n9131 , n5296 , n5387 );
nor ( n9132 , n9130 , n9131 );
xnor ( n9133 , n9132 , n5382 );
and ( n9134 , n5340 , n5262 );
and ( n9135 , n7639 , n5260 );
nor ( n9136 , n9134 , n9135 );
xnor ( n9137 , n9136 , n5270 );
and ( n9138 , n9133 , n9137 );
xor ( n9139 , n9029 , n9033 );
xor ( n9140 , n9139 , n9038 );
and ( n9141 , n9137 , n9140 );
and ( n9142 , n9133 , n9140 );
or ( n9143 , n9138 , n9141 , n9142 );
and ( n9144 , n9129 , n9143 );
xor ( n9145 , n8891 , n8895 );
xor ( n9146 , n9145 , n8900 );
and ( n9147 , n9143 , n9146 );
and ( n9148 , n9129 , n9146 );
or ( n9149 , n9144 , n9147 , n9148 );
xor ( n9150 , n8917 , n8921 );
xor ( n9151 , n9150 , n8926 );
xor ( n9152 , n8942 , n8946 );
xor ( n9153 , n9152 , n8951 );
and ( n9154 , n9151 , n9153 );
xor ( n9155 , n9013 , n9017 );
xor ( n9156 , n9155 , n9022 );
and ( n9157 , n7660 , n5325 );
and ( n9158 , n5536 , n5323 );
nor ( n9159 , n9157 , n9158 );
xnor ( n9160 , n9159 , n5333 );
and ( n9161 , n7639 , n5243 );
and ( n9162 , n7690 , n5241 );
nor ( n9163 , n9161 , n9162 );
xnor ( n9164 , n9163 , n5251 );
or ( n9165 , n9160 , n9164 );
and ( n9166 , n9156 , n9165 );
and ( n9167 , n5317 , n5468 );
and ( n9168 , n5328 , n5438 );
nor ( n9169 , n9167 , n9168 );
xnor ( n9170 , n9169 , n5405 );
and ( n9171 , n5233 , n7865 );
and ( n9172 , n5246 , n7863 );
nor ( n9173 , n9171 , n9172 );
xnor ( n9174 , n9173 , n5429 );
and ( n9175 , n9170 , n9174 );
and ( n9176 , n5274 , n5306 );
and ( n9177 , n5285 , n5304 );
nor ( n9178 , n9176 , n9177 );
xnor ( n9179 , n9178 , n5314 );
and ( n9180 , n9174 , n9179 );
and ( n9181 , n9170 , n9179 );
or ( n9182 , n9175 , n9180 , n9181 );
and ( n9183 , n9165 , n9182 );
and ( n9184 , n9156 , n9182 );
or ( n9185 , n9166 , n9183 , n9184 );
and ( n9186 , n9153 , n9185 );
and ( n9187 , n9151 , n9185 );
or ( n9188 , n9154 , n9186 , n9187 );
and ( n9189 , n9149 , n9188 );
xor ( n9190 , n8999 , n9008 );
xor ( n9191 , n9190 , n9061 );
and ( n9192 , n9188 , n9191 );
and ( n9193 , n9149 , n9191 );
or ( n9194 , n9189 , n9192 , n9193 );
and ( n9195 , n9101 , n9194 );
and ( n9196 , n9099 , n9194 );
or ( n9197 , n9102 , n9195 , n9196 );
xor ( n9198 , n9078 , n9080 );
xor ( n9199 , n9198 , n9083 );
and ( n9200 , n9197 , n9199 );
xor ( n9201 , n8997 , n9064 );
xor ( n9202 , n9201 , n9075 );
xor ( n9203 , n9067 , n9069 );
xor ( n9204 , n9203 , n9072 );
xor ( n9205 , n8874 , n9003 );
xor ( n9206 , n9205 , n9005 );
xor ( n9207 , n9025 , n9041 );
xor ( n9208 , n9207 , n9058 );
and ( n9209 , n9206 , n9208 );
xor ( n9210 , n9129 , n9143 );
xor ( n9211 , n9210 , n9146 );
and ( n9212 , n9208 , n9211 );
and ( n9213 , n9206 , n9211 );
or ( n9214 , n9209 , n9212 , n9213 );
and ( n9215 , n9204 , n9214 );
xor ( n9216 , n9046 , n9050 );
xor ( n9217 , n9216 , n9055 );
xor ( n9218 , n9118 , n9122 );
xor ( n9219 , n9218 , n9126 );
and ( n9220 , n9217 , n9219 );
xor ( n9221 , n9133 , n9137 );
xor ( n9222 , n9221 , n9140 );
and ( n9223 , n9219 , n9222 );
and ( n9224 , n9217 , n9222 );
or ( n9225 , n9220 , n9223 , n9224 );
and ( n9226 , n7647 , n5390 );
and ( n9227 , n7650 , n5387 );
nor ( n9228 , n9226 , n9227 );
xnor ( n9229 , n9228 , n5382 );
and ( n9230 , n5350 , n5414 );
and ( n9231 , n7716 , n5412 );
nor ( n9232 , n9230 , n9231 );
xnor ( n9233 , n9232 , n5420 );
and ( n9234 , n9229 , n9233 );
xor ( n9235 , n9106 , n9110 );
xor ( n9236 , n9235 , n9115 );
and ( n9237 , n9233 , n9236 );
and ( n9238 , n9229 , n9236 );
or ( n9239 , n9234 , n9237 , n9238 );
xor ( n9240 , n7274 , n7600 );
buf ( n9241 , n9240 );
buf ( n9242 , n9241 );
buf ( n9243 , n9242 );
and ( n9244 , n9124 , n9243 );
xnor ( n9245 , n9160 , n9164 );
and ( n9246 , n9243 , n9245 );
and ( n9247 , n9124 , n9245 );
or ( n9248 , n9244 , n9246 , n9247 );
and ( n9249 , n9239 , n9248 );
and ( n9250 , n5328 , n5414 );
and ( n9251 , n5350 , n5412 );
nor ( n9252 , n9250 , n9251 );
xnor ( n9253 , n9252 , n5420 );
and ( n9254 , n7690 , n5325 );
and ( n9255 , n7660 , n5323 );
nor ( n9256 , n9254 , n9255 );
xnor ( n9257 , n9256 , n5333 );
and ( n9258 , n9253 , n9257 );
and ( n9259 , n5340 , n5243 );
and ( n9260 , n7639 , n5241 );
nor ( n9261 , n9259 , n9260 );
xnor ( n9262 , n9261 , n5251 );
and ( n9263 , n9257 , n9262 );
and ( n9264 , n9253 , n9262 );
or ( n9265 , n9258 , n9263 , n9264 );
and ( n9266 , n5265 , n7865 );
and ( n9267 , n5233 , n7863 );
nor ( n9268 , n9266 , n9267 );
xnor ( n9269 , n9268 , n5429 );
and ( n9270 , n5340 , n5241 );
not ( n9271 , n9270 );
and ( n9272 , n9271 , n5251 );
and ( n9273 , n9269 , n9272 );
and ( n9274 , n9265 , n9273 );
and ( n9275 , n7716 , n5390 );
and ( n9276 , n7647 , n5387 );
nor ( n9277 , n9275 , n9276 );
xnor ( n9278 , n9277 , n5382 );
and ( n9279 , n5246 , n5468 );
and ( n9280 , n5317 , n5438 );
nor ( n9281 , n9279 , n9280 );
xnor ( n9282 , n9281 , n5405 );
and ( n9283 , n9278 , n9282 );
and ( n9284 , n5285 , n5487 );
and ( n9285 , n5254 , n5485 );
nor ( n9286 , n9284 , n9285 );
xnor ( n9287 , n9286 , n5478 );
and ( n9288 , n9282 , n9287 );
and ( n9289 , n9278 , n9287 );
or ( n9290 , n9283 , n9288 , n9289 );
and ( n9291 , n9273 , n9290 );
and ( n9292 , n9265 , n9290 );
or ( n9293 , n9274 , n9291 , n9292 );
and ( n9294 , n9248 , n9293 );
and ( n9295 , n9239 , n9293 );
or ( n9296 , n9249 , n9294 , n9295 );
and ( n9297 , n9225 , n9296 );
xor ( n9298 , n9151 , n9153 );
xor ( n9299 , n9298 , n9185 );
and ( n9300 , n9296 , n9299 );
and ( n9301 , n9225 , n9299 );
or ( n9302 , n9297 , n9300 , n9301 );
and ( n9303 , n9214 , n9302 );
and ( n9304 , n9204 , n9302 );
or ( n9305 , n9215 , n9303 , n9304 );
and ( n9306 , n9202 , n9305 );
xor ( n9307 , n9099 , n9101 );
xor ( n9308 , n9307 , n9194 );
and ( n9309 , n9305 , n9308 );
and ( n9310 , n9202 , n9308 );
or ( n9311 , n9306 , n9309 , n9310 );
and ( n9312 , n9199 , n9311 );
and ( n9313 , n9197 , n9311 );
or ( n9314 , n9200 , n9312 , n9313 );
or ( n9315 , n9097 , n9314 );
and ( n9316 , n9094 , n9315 );
and ( n9317 , n9092 , n9315 );
or ( n9318 , n9095 , n9316 , n9317 );
and ( n9319 , n8992 , n9318 );
and ( n9320 , n8990 , n9318 );
or ( n9321 , n8993 , n9319 , n9320 );
or ( n9322 , n8864 , n9321 );
and ( n9323 , n8862 , n9322 );
xor ( n9324 , n8862 , n9322 );
xnor ( n9325 , n8864 , n9321 );
xor ( n9326 , n8990 , n8992 );
xor ( n9327 , n9326 , n9318 );
not ( n9328 , n9327 );
xor ( n9329 , n9092 , n9094 );
xor ( n9330 , n9329 , n9315 );
not ( n9331 , n9330 );
xnor ( n9332 , n9097 , n9314 );
xor ( n9333 , n9197 , n9199 );
xor ( n9334 , n9333 , n9311 );
xor ( n9335 , n9149 , n9188 );
xor ( n9336 , n9335 , n9191 );
xor ( n9337 , n9156 , n9165 );
xor ( n9338 , n9337 , n9182 );
and ( n9339 , n5529 , n5306 );
and ( n9340 , n5274 , n5304 );
nor ( n9341 , n9339 , n9340 );
xnor ( n9342 , n9341 , n5314 );
and ( n9343 , n5355 , n7722 );
and ( n9344 , n5368 , n7720 );
nor ( n9345 , n9343 , n9344 );
xnor ( n9346 , n9345 , n7728 );
and ( n9347 , n9342 , n9346 );
and ( n9348 , n5536 , n5499 );
and ( n9349 , n5545 , n5497 );
nor ( n9350 , n9348 , n9349 );
xnor ( n9351 , n9350 , n5505 );
and ( n9352 , n9346 , n9351 );
and ( n9353 , n9342 , n9351 );
or ( n9354 , n9347 , n9352 , n9353 );
xor ( n9355 , n9170 , n9174 );
xor ( n9356 , n9355 , n9179 );
and ( n9357 , n9354 , n9356 );
xor ( n9358 , n9229 , n9233 );
xor ( n9359 , n9358 , n9236 );
and ( n9360 , n9356 , n9359 );
and ( n9361 , n9354 , n9359 );
or ( n9362 , n9357 , n9360 , n9361 );
and ( n9363 , n9338 , n9362 );
xor ( n9364 , n7276 , n7599 );
buf ( n9365 , n9364 );
buf ( n9366 , n9365 );
buf ( n9367 , n9366 );
xor ( n9368 , n9253 , n9257 );
xor ( n9369 , n9368 , n9262 );
and ( n9370 , n9367 , n9369 );
xor ( n9371 , n9269 , n9272 );
and ( n9372 , n9369 , n9371 );
and ( n9373 , n9367 , n9371 );
or ( n9374 , n9370 , n9372 , n9373 );
and ( n9375 , n5274 , n5487 );
and ( n9376 , n5285 , n5485 );
nor ( n9377 , n9375 , n9376 );
xnor ( n9378 , n9377 , n5478 );
and ( n9379 , n5368 , n5306 );
and ( n9380 , n5529 , n5304 );
nor ( n9381 , n9379 , n9380 );
xnor ( n9382 , n9381 , n5314 );
and ( n9383 , n9378 , n9382 );
and ( n9384 , n5545 , n7722 );
and ( n9385 , n5355 , n7720 );
nor ( n9386 , n9384 , n9385 );
xnor ( n9387 , n9386 , n7728 );
and ( n9388 , n9382 , n9387 );
and ( n9389 , n9378 , n9387 );
or ( n9390 , n9383 , n9388 , n9389 );
and ( n9391 , n5350 , n5390 );
and ( n9392 , n7716 , n5387 );
nor ( n9393 , n9391 , n9392 );
xnor ( n9394 , n9393 , n5382 );
and ( n9395 , n7639 , n5325 );
and ( n9396 , n7690 , n5323 );
nor ( n9397 , n9395 , n9396 );
xnor ( n9398 , n9397 , n5333 );
and ( n9399 , n9394 , n9398 );
and ( n9400 , n9390 , n9399 );
xor ( n9401 , n9278 , n9282 );
xor ( n9402 , n9401 , n9287 );
and ( n9403 , n9399 , n9402 );
and ( n9404 , n9390 , n9402 );
or ( n9405 , n9400 , n9403 , n9404 );
and ( n9406 , n9374 , n9405 );
xor ( n9407 , n9124 , n9243 );
xor ( n9408 , n9407 , n9245 );
and ( n9409 , n9405 , n9408 );
and ( n9410 , n9374 , n9408 );
or ( n9411 , n9406 , n9409 , n9410 );
and ( n9412 , n9362 , n9411 );
and ( n9413 , n9338 , n9411 );
or ( n9414 , n9363 , n9412 , n9413 );
xor ( n9415 , n9206 , n9208 );
xor ( n9416 , n9415 , n9211 );
and ( n9417 , n9414 , n9416 );
xor ( n9418 , n9225 , n9296 );
xor ( n9419 , n9418 , n9299 );
and ( n9420 , n9416 , n9419 );
and ( n9421 , n9414 , n9419 );
or ( n9422 , n9417 , n9420 , n9421 );
and ( n9423 , n9336 , n9422 );
xor ( n9424 , n9204 , n9214 );
xor ( n9425 , n9424 , n9302 );
and ( n9426 , n9422 , n9425 );
and ( n9427 , n9336 , n9425 );
or ( n9428 , n9423 , n9426 , n9427 );
xor ( n9429 , n9202 , n9305 );
xor ( n9430 , n9429 , n9308 );
and ( n9431 , n9428 , n9430 );
xor ( n9432 , n9336 , n9422 );
xor ( n9433 , n9432 , n9425 );
xor ( n9434 , n9217 , n9219 );
xor ( n9435 , n9434 , n9222 );
xor ( n9436 , n9239 , n9248 );
xor ( n9437 , n9436 , n9293 );
and ( n9438 , n9435 , n9437 );
xor ( n9439 , n9265 , n9273 );
xor ( n9440 , n9439 , n9290 );
xor ( n9441 , n9342 , n9346 );
xor ( n9442 , n9441 , n9351 );
and ( n9443 , n5529 , n5487 );
and ( n9444 , n5274 , n5485 );
nor ( n9445 , n9443 , n9444 );
xnor ( n9446 , n9445 , n5478 );
and ( n9447 , n5355 , n5306 );
and ( n9448 , n5368 , n5304 );
nor ( n9449 , n9447 , n9448 );
xnor ( n9450 , n9449 , n5314 );
and ( n9451 , n9446 , n9450 );
and ( n9452 , n5233 , n5468 );
and ( n9453 , n5246 , n5438 );
nor ( n9454 , n9452 , n9453 );
xnor ( n9455 , n9454 , n5405 );
and ( n9456 , n9451 , n9455 );
and ( n9457 , n7660 , n5499 );
and ( n9458 , n5536 , n5497 );
nor ( n9459 , n9457 , n9458 );
xnor ( n9460 , n9459 , n5505 );
and ( n9461 , n9455 , n9460 );
and ( n9462 , n9451 , n9460 );
or ( n9463 , n9456 , n9461 , n9462 );
and ( n9464 , n9442 , n9463 );
and ( n9465 , n5317 , n5414 );
and ( n9466 , n5328 , n5412 );
nor ( n9467 , n9465 , n9466 );
xnor ( n9468 , n9467 , n5420 );
and ( n9469 , n9468 , n9270 );
xor ( n9470 , n9378 , n9382 );
xor ( n9471 , n9470 , n9387 );
and ( n9472 , n9270 , n9471 );
and ( n9473 , n9468 , n9471 );
or ( n9474 , n9469 , n9472 , n9473 );
and ( n9475 , n9463 , n9474 );
and ( n9476 , n9442 , n9474 );
or ( n9477 , n9464 , n9475 , n9476 );
and ( n9478 , n9440 , n9477 );
and ( n9479 , n5254 , n7865 );
and ( n9480 , n5265 , n7863 );
nor ( n9481 , n9479 , n9480 );
xnor ( n9482 , n9481 , n5429 );
xor ( n9483 , n7279 , n7597 );
buf ( n9484 , n9483 );
buf ( n9485 , n9484 );
buf ( n9486 , n9485 );
and ( n9487 , n9482 , n9486 );
xor ( n9488 , n9394 , n9398 );
and ( n9489 , n9486 , n9488 );
and ( n9490 , n9482 , n9488 );
or ( n9491 , n9487 , n9489 , n9490 );
xor ( n9492 , n9367 , n9369 );
xor ( n9493 , n9492 , n9371 );
and ( n9494 , n9491 , n9493 );
xor ( n9495 , n9390 , n9399 );
xor ( n9496 , n9495 , n9402 );
and ( n9497 , n9493 , n9496 );
and ( n9498 , n9491 , n9496 );
or ( n9499 , n9494 , n9497 , n9498 );
and ( n9500 , n9477 , n9499 );
and ( n9501 , n9440 , n9499 );
or ( n9502 , n9478 , n9500 , n9501 );
and ( n9503 , n9437 , n9502 );
and ( n9504 , n9435 , n9502 );
or ( n9505 , n9438 , n9503 , n9504 );
xor ( n9506 , n9414 , n9416 );
xor ( n9507 , n9506 , n9419 );
and ( n9508 , n9505 , n9507 );
xor ( n9509 , n9338 , n9362 );
xor ( n9510 , n9509 , n9411 );
xor ( n9511 , n9354 , n9356 );
xor ( n9512 , n9511 , n9359 );
xor ( n9513 , n9374 , n9405 );
xor ( n9514 , n9513 , n9408 );
and ( n9515 , n9512 , n9514 );
and ( n9516 , n5328 , n5390 );
and ( n9517 , n5350 , n5387 );
nor ( n9518 , n9516 , n9517 );
xnor ( n9519 , n9518 , n5382 );
and ( n9520 , n5246 , n5414 );
and ( n9521 , n5317 , n5412 );
nor ( n9522 , n9520 , n9521 );
xnor ( n9523 , n9522 , n5420 );
and ( n9524 , n9519 , n9523 );
and ( n9525 , n5265 , n5468 );
and ( n9526 , n5233 , n5438 );
nor ( n9527 , n9525 , n9526 );
xnor ( n9528 , n9527 , n5405 );
and ( n9529 , n9523 , n9528 );
and ( n9530 , n9519 , n9528 );
or ( n9531 , n9524 , n9529 , n9530 );
and ( n9532 , n5536 , n7722 );
and ( n9533 , n5545 , n7720 );
nor ( n9534 , n9532 , n9533 );
xnor ( n9535 , n9534 , n7728 );
and ( n9536 , n5340 , n5325 );
and ( n9537 , n7639 , n5323 );
nor ( n9538 , n9536 , n9537 );
xnor ( n9539 , n9538 , n5333 );
and ( n9540 , n9535 , n9539 );
and ( n9541 , n5340 , n5323 );
not ( n9542 , n9541 );
and ( n9543 , n9542 , n5333 );
and ( n9544 , n9539 , n9543 );
and ( n9545 , n9535 , n9543 );
or ( n9546 , n9540 , n9544 , n9545 );
and ( n9547 , n9531 , n9546 );
xor ( n9548 , n9451 , n9455 );
xor ( n9549 , n9548 , n9460 );
and ( n9550 , n9546 , n9549 );
and ( n9551 , n9531 , n9549 );
or ( n9552 , n9547 , n9550 , n9551 );
xor ( n9553 , n9468 , n9270 );
xor ( n9554 , n9553 , n9471 );
xor ( n9555 , n9446 , n9450 );
and ( n9556 , n5285 , n7865 );
and ( n9557 , n5254 , n7863 );
nor ( n9558 , n9556 , n9557 );
xnor ( n9559 , n9558 , n5429 );
and ( n9560 , n9555 , n9559 );
and ( n9561 , n7690 , n5499 );
and ( n9562 , n7660 , n5497 );
nor ( n9563 , n9561 , n9562 );
xnor ( n9564 , n9563 , n5505 );
and ( n9565 , n9559 , n9564 );
and ( n9566 , n9555 , n9564 );
or ( n9567 , n9560 , n9565 , n9566 );
and ( n9568 , n9554 , n9567 );
xor ( n9569 , n7282 , n7595 );
buf ( n9570 , n9569 );
buf ( n9571 , n9570 );
buf ( n9572 , n9571 );
and ( n9573 , n5368 , n5487 );
and ( n9574 , n5529 , n5485 );
nor ( n9575 , n9573 , n9574 );
xnor ( n9576 , n9575 , n5478 );
not ( n9577 , n9576 );
and ( n9578 , n5545 , n5306 );
and ( n9579 , n5355 , n5304 );
nor ( n9580 , n9578 , n9579 );
xnor ( n9581 , n9580 , n5314 );
and ( n9582 , n9577 , n9581 );
and ( n9583 , n9572 , n9582 );
buf ( n9584 , n9576 );
and ( n9585 , n9582 , n9584 );
and ( n9586 , n9572 , n9584 );
or ( n9587 , n9583 , n9585 , n9586 );
and ( n9588 , n9567 , n9587 );
and ( n9589 , n9554 , n9587 );
or ( n9590 , n9568 , n9588 , n9589 );
and ( n9591 , n9552 , n9590 );
xor ( n9592 , n9442 , n9463 );
xor ( n9593 , n9592 , n9474 );
and ( n9594 , n9590 , n9593 );
and ( n9595 , n9552 , n9593 );
or ( n9596 , n9591 , n9594 , n9595 );
and ( n9597 , n9514 , n9596 );
and ( n9598 , n9512 , n9596 );
or ( n9599 , n9515 , n9597 , n9598 );
and ( n9600 , n9510 , n9599 );
xor ( n9601 , n9435 , n9437 );
xor ( n9602 , n9601 , n9502 );
and ( n9603 , n9599 , n9602 );
and ( n9604 , n9510 , n9602 );
or ( n9605 , n9600 , n9603 , n9604 );
and ( n9606 , n9507 , n9605 );
and ( n9607 , n9505 , n9605 );
or ( n9608 , n9508 , n9606 , n9607 );
and ( n9609 , n9433 , n9608 );
xor ( n9610 , n9505 , n9507 );
xor ( n9611 , n9610 , n9605 );
xor ( n9612 , n9440 , n9477 );
xor ( n9613 , n9612 , n9499 );
xor ( n9614 , n9491 , n9493 );
xor ( n9615 , n9614 , n9496 );
and ( n9616 , n5317 , n5390 );
and ( n9617 , n5328 , n5387 );
nor ( n9618 , n9616 , n9617 );
xnor ( n9619 , n9618 , n5382 );
and ( n9620 , n5233 , n5414 );
and ( n9621 , n5246 , n5412 );
nor ( n9622 , n9620 , n9621 );
xnor ( n9623 , n9622 , n5420 );
and ( n9624 , n9619 , n9623 );
and ( n9625 , n5254 , n5468 );
and ( n9626 , n5265 , n5438 );
nor ( n9627 , n9625 , n9626 );
xnor ( n9628 , n9627 , n5405 );
and ( n9629 , n9623 , n9628 );
and ( n9630 , n9619 , n9628 );
or ( n9631 , n9624 , n9629 , n9630 );
and ( n9632 , n5274 , n7865 );
and ( n9633 , n5285 , n7863 );
nor ( n9634 , n9632 , n9633 );
xnor ( n9635 , n9634 , n5429 );
and ( n9636 , n7660 , n7722 );
and ( n9637 , n5536 , n7720 );
nor ( n9638 , n9636 , n9637 );
xnor ( n9639 , n9638 , n7728 );
and ( n9640 , n9635 , n9639 );
and ( n9641 , n7639 , n5499 );
and ( n9642 , n7690 , n5497 );
nor ( n9643 , n9641 , n9642 );
xnor ( n9644 , n9643 , n5505 );
and ( n9645 , n9639 , n9644 );
and ( n9646 , n9635 , n9644 );
or ( n9647 , n9640 , n9645 , n9646 );
and ( n9648 , n9631 , n9647 );
xor ( n9649 , n9519 , n9523 );
xor ( n9650 , n9649 , n9528 );
and ( n9651 , n9647 , n9650 );
and ( n9652 , n9631 , n9650 );
or ( n9653 , n9648 , n9651 , n9652 );
xor ( n9654 , n9482 , n9486 );
xor ( n9655 , n9654 , n9488 );
and ( n9656 , n9653 , n9655 );
xor ( n9657 , n9535 , n9539 );
xor ( n9658 , n9657 , n9543 );
xor ( n9659 , n9555 , n9559 );
xor ( n9660 , n9659 , n9564 );
and ( n9661 , n9658 , n9660 );
xor ( n9662 , n7283 , n7594 );
buf ( n9663 , n9662 );
buf ( n9664 , n9663 );
buf ( n9665 , n9664 );
and ( n9666 , n9541 , n9665 );
xor ( n9667 , n9577 , n9581 );
and ( n9668 , n9665 , n9667 );
and ( n9669 , n9541 , n9667 );
or ( n9670 , n9666 , n9668 , n9669 );
and ( n9671 , n9660 , n9670 );
and ( n9672 , n9658 , n9670 );
or ( n9673 , n9661 , n9671 , n9672 );
and ( n9674 , n9655 , n9673 );
and ( n9675 , n9653 , n9673 );
or ( n9676 , n9656 , n9674 , n9675 );
and ( n9677 , n9615 , n9676 );
and ( n9678 , n5355 , n5487 );
and ( n9679 , n5368 , n5485 );
nor ( n9680 , n9678 , n9679 );
xnor ( n9681 , n9680 , n5478 );
and ( n9682 , n5536 , n5306 );
and ( n9683 , n5545 , n5304 );
nor ( n9684 , n9682 , n9683 );
xnor ( n9685 , n9684 , n5314 );
or ( n9686 , n9681 , n9685 );
and ( n9687 , n5246 , n5390 );
and ( n9688 , n5317 , n5387 );
nor ( n9689 , n9687 , n9688 );
xnor ( n9690 , n9689 , n5382 );
and ( n9691 , n5265 , n5414 );
and ( n9692 , n5233 , n5412 );
nor ( n9693 , n9691 , n9692 );
xnor ( n9694 , n9693 , n5420 );
and ( n9695 , n9690 , n9694 );
and ( n9696 , n5529 , n7865 );
and ( n9697 , n5274 , n7863 );
nor ( n9698 , n9696 , n9697 );
xnor ( n9699 , n9698 , n5429 );
and ( n9700 , n9694 , n9699 );
and ( n9701 , n9690 , n9699 );
or ( n9702 , n9695 , n9700 , n9701 );
and ( n9703 , n9686 , n9702 );
and ( n9704 , n7690 , n7722 );
and ( n9705 , n7660 , n7720 );
nor ( n9706 , n9704 , n9705 );
xnor ( n9707 , n9706 , n7728 );
and ( n9708 , n5340 , n5497 );
not ( n9709 , n9708 );
and ( n9710 , n9709 , n5505 );
and ( n9711 , n9707 , n9710 );
xor ( n9712 , n7284 , n7593 );
buf ( n9713 , n9712 );
buf ( n9714 , n9713 );
buf ( n9715 , n9714 );
and ( n9716 , n9710 , n9715 );
and ( n9717 , n9707 , n9715 );
or ( n9718 , n9711 , n9716 , n9717 );
and ( n9719 , n9702 , n9718 );
and ( n9720 , n9686 , n9718 );
or ( n9721 , n9703 , n9719 , n9720 );
xor ( n9722 , n9572 , n9582 );
xor ( n9723 , n9722 , n9584 );
and ( n9724 , n9721 , n9723 );
xor ( n9725 , n9631 , n9647 );
xor ( n9726 , n9725 , n9650 );
and ( n9727 , n9723 , n9726 );
and ( n9728 , n9721 , n9726 );
or ( n9729 , n9724 , n9727 , n9728 );
xor ( n9730 , n9531 , n9546 );
xor ( n9731 , n9730 , n9549 );
and ( n9732 , n9729 , n9731 );
xor ( n9733 , n9554 , n9567 );
xor ( n9734 , n9733 , n9587 );
and ( n9735 , n9731 , n9734 );
and ( n9736 , n9729 , n9734 );
or ( n9737 , n9732 , n9735 , n9736 );
and ( n9738 , n9676 , n9737 );
and ( n9739 , n9615 , n9737 );
or ( n9740 , n9677 , n9738 , n9739 );
and ( n9741 , n9613 , n9740 );
xor ( n9742 , n9512 , n9514 );
xor ( n9743 , n9742 , n9596 );
and ( n9744 , n9740 , n9743 );
and ( n9745 , n9613 , n9743 );
or ( n9746 , n9741 , n9744 , n9745 );
xor ( n9747 , n9510 , n9599 );
xor ( n9748 , n9747 , n9602 );
and ( n9749 , n9746 , n9748 );
xor ( n9750 , n9552 , n9590 );
xor ( n9751 , n9750 , n9593 );
xor ( n9752 , n9619 , n9623 );
xor ( n9753 , n9752 , n9628 );
xor ( n9754 , n9635 , n9639 );
xor ( n9755 , n9754 , n9644 );
and ( n9756 , n9753 , n9755 );
xnor ( n9757 , n9681 , n9685 );
and ( n9758 , n5254 , n5414 );
and ( n9759 , n5265 , n5412 );
nor ( n9760 , n9758 , n9759 );
xnor ( n9761 , n9760 , n5420 );
and ( n9762 , n5274 , n5468 );
and ( n9763 , n5285 , n5438 );
nor ( n9764 , n9762 , n9763 );
xnor ( n9765 , n9764 , n5405 );
and ( n9766 , n9761 , n9765 );
and ( n9767 , n7639 , n7722 );
and ( n9768 , n7690 , n7720 );
nor ( n9769 , n9767 , n9768 );
xnor ( n9770 , n9769 , n7728 );
and ( n9771 , n9765 , n9770 );
and ( n9772 , n9761 , n9770 );
or ( n9773 , n9766 , n9771 , n9772 );
and ( n9774 , n9757 , n9773 );
and ( n9775 , n7660 , n5306 );
and ( n9776 , n5536 , n5304 );
nor ( n9777 , n9775 , n9776 );
xnor ( n9778 , n9777 , n5314 );
and ( n9779 , n9778 , n9708 );
xor ( n9780 , n7287 , n7591 );
buf ( n9781 , n9780 );
buf ( n9782 , n9781 );
buf ( n9783 , n9782 );
and ( n9784 , n9708 , n9783 );
and ( n9785 , n9778 , n9783 );
or ( n9786 , n9779 , n9784 , n9785 );
and ( n9787 , n9773 , n9786 );
and ( n9788 , n9757 , n9786 );
or ( n9789 , n9774 , n9787 , n9788 );
and ( n9790 , n9755 , n9789 );
and ( n9791 , n9753 , n9789 );
or ( n9792 , n9756 , n9790 , n9791 );
xor ( n9793 , n9658 , n9660 );
xor ( n9794 , n9793 , n9670 );
and ( n9795 , n9792 , n9794 );
xor ( n9796 , n9721 , n9723 );
xor ( n9797 , n9796 , n9726 );
and ( n9798 , n9794 , n9797 );
and ( n9799 , n9792 , n9797 );
or ( n9800 , n9795 , n9798 , n9799 );
xor ( n9801 , n9653 , n9655 );
xor ( n9802 , n9801 , n9673 );
and ( n9803 , n9800 , n9802 );
xor ( n9804 , n9729 , n9731 );
xor ( n9805 , n9804 , n9734 );
and ( n9806 , n9802 , n9805 );
and ( n9807 , n9800 , n9805 );
or ( n9808 , n9803 , n9806 , n9807 );
and ( n9809 , n9751 , n9808 );
xor ( n9810 , n9615 , n9676 );
xor ( n9811 , n9810 , n9737 );
and ( n9812 , n9808 , n9811 );
and ( n9813 , n9751 , n9811 );
or ( n9814 , n9809 , n9812 , n9813 );
xor ( n9815 , n9613 , n9740 );
xor ( n9816 , n9815 , n9743 );
and ( n9817 , n9814 , n9816 );
xor ( n9818 , n9751 , n9808 );
xor ( n9819 , n9818 , n9811 );
xor ( n9820 , n9800 , n9802 );
xor ( n9821 , n9820 , n9805 );
xor ( n9822 , n9541 , n9665 );
xor ( n9823 , n9822 , n9667 );
xor ( n9824 , n9686 , n9702 );
xor ( n9825 , n9824 , n9718 );
and ( n9826 , n9823 , n9825 );
and ( n9827 , n5355 , n7865 );
and ( n9828 , n5368 , n7863 );
nor ( n9829 , n9827 , n9828 );
xnor ( n9830 , n9829 , n5429 );
and ( n9831 , n5536 , n5487 );
and ( n9832 , n5545 , n5485 );
nor ( n9833 , n9831 , n9832 );
xnor ( n9834 , n9833 , n5478 );
and ( n9835 , n9830 , n9834 );
and ( n9836 , n5368 , n7865 );
and ( n9837 , n5529 , n7863 );
nor ( n9838 , n9836 , n9837 );
xnor ( n9839 , n9838 , n5429 );
and ( n9840 , n9835 , n9839 );
and ( n9841 , n5545 , n5487 );
and ( n9842 , n5355 , n5485 );
nor ( n9843 , n9841 , n9842 );
xnor ( n9844 , n9843 , n5478 );
and ( n9845 , n9839 , n9844 );
and ( n9846 , n9835 , n9844 );
or ( n9847 , n9840 , n9845 , n9846 );
and ( n9848 , n5285 , n5468 );
and ( n9849 , n5254 , n5438 );
nor ( n9850 , n9848 , n9849 );
xnor ( n9851 , n9850 , n5405 );
and ( n9852 , n9847 , n9851 );
and ( n9853 , n5340 , n5499 );
and ( n9854 , n7639 , n5497 );
nor ( n9855 , n9853 , n9854 );
xnor ( n9856 , n9855 , n5505 );
and ( n9857 , n9851 , n9856 );
and ( n9858 , n9847 , n9856 );
or ( n9859 , n9852 , n9857 , n9858 );
and ( n9860 , n9825 , n9859 );
and ( n9861 , n9823 , n9859 );
or ( n9862 , n9826 , n9860 , n9861 );
xor ( n9863 , n9792 , n9794 );
xor ( n9864 , n9863 , n9797 );
and ( n9865 , n9862 , n9864 );
xor ( n9866 , n9690 , n9694 );
xor ( n9867 , n9866 , n9699 );
xor ( n9868 , n9707 , n9710 );
xor ( n9869 , n9868 , n9715 );
and ( n9870 , n9867 , n9869 );
xor ( n9871 , n9761 , n9765 );
xor ( n9872 , n9871 , n9770 );
and ( n9873 , n5285 , n5414 );
and ( n9874 , n5254 , n5412 );
nor ( n9875 , n9873 , n9874 );
xnor ( n9876 , n9875 , n5420 );
and ( n9877 , n5340 , n7722 );
and ( n9878 , n7639 , n7720 );
nor ( n9879 , n9877 , n9878 );
xnor ( n9880 , n9879 , n7728 );
and ( n9881 , n9876 , n9880 );
and ( n9882 , n5340 , n7720 );
not ( n9883 , n9882 );
and ( n9884 , n9883 , n7728 );
and ( n9885 , n9880 , n9884 );
and ( n9886 , n9876 , n9884 );
or ( n9887 , n9881 , n9885 , n9886 );
and ( n9888 , n9872 , n9887 );
xor ( n9889 , n9778 , n9708 );
xor ( n9890 , n9889 , n9783 );
and ( n9891 , n9887 , n9890 );
and ( n9892 , n9872 , n9890 );
or ( n9893 , n9888 , n9891 , n9892 );
and ( n9894 , n9869 , n9893 );
and ( n9895 , n9867 , n9893 );
or ( n9896 , n9870 , n9894 , n9895 );
xor ( n9897 , n9753 , n9755 );
xor ( n9898 , n9897 , n9789 );
and ( n9899 , n9896 , n9898 );
xor ( n9900 , n9757 , n9773 );
xor ( n9901 , n9900 , n9786 );
xor ( n9902 , n9847 , n9851 );
xor ( n9903 , n9902 , n9856 );
and ( n9904 , n9901 , n9903 );
xor ( n9905 , n9835 , n9839 );
xor ( n9906 , n9905 , n9844 );
xor ( n9907 , n7538 , n7589 );
buf ( n9908 , n9907 );
buf ( n9909 , n9908 );
buf ( n9910 , n9909 );
xor ( n9911 , n9830 , n9834 );
and ( n9912 , n9910 , n9911 );
and ( n9913 , n5368 , n5468 );
and ( n9914 , n5529 , n5438 );
nor ( n9915 , n9913 , n9914 );
xnor ( n9916 , n9915 , n5405 );
and ( n9917 , n7639 , n5306 );
and ( n9918 , n7690 , n5304 );
nor ( n9919 , n9917 , n9918 );
xnor ( n9920 , n9919 , n5314 );
and ( n9921 , n9916 , n9920 );
and ( n9922 , n9920 , n9882 );
and ( n9923 , n9916 , n9882 );
or ( n9924 , n9921 , n9922 , n9923 );
and ( n9925 , n9911 , n9924 );
and ( n9926 , n9910 , n9924 );
or ( n9927 , n9912 , n9925 , n9926 );
and ( n9928 , n9906 , n9927 );
xor ( n9929 , n9872 , n9887 );
xor ( n9930 , n9929 , n9890 );
and ( n9931 , n9927 , n9930 );
and ( n9932 , n9906 , n9930 );
or ( n9933 , n9928 , n9931 , n9932 );
and ( n9934 , n9903 , n9933 );
and ( n9935 , n9901 , n9933 );
or ( n9936 , n9904 , n9934 , n9935 );
and ( n9937 , n9898 , n9936 );
and ( n9938 , n9896 , n9936 );
or ( n9939 , n9899 , n9937 , n9938 );
and ( n9940 , n9864 , n9939 );
and ( n9941 , n9862 , n9939 );
or ( n9942 , n9865 , n9940 , n9941 );
and ( n9943 , n9821 , n9942 );
xor ( n9944 , n9823 , n9825 );
xor ( n9945 , n9944 , n9859 );
xor ( n9946 , n9867 , n9869 );
xor ( n9947 , n9946 , n9893 );
and ( n9948 , n5355 , n5468 );
and ( n9949 , n5368 , n5438 );
nor ( n9950 , n9948 , n9949 );
xnor ( n9951 , n9950 , n5405 );
and ( n9952 , n5340 , n5304 );
not ( n9953 , n9952 );
and ( n9954 , n9953 , n5314 );
and ( n9955 , n9951 , n9954 );
and ( n9956 , n5545 , n7865 );
and ( n9957 , n5355 , n7863 );
nor ( n9958 , n9956 , n9957 );
xnor ( n9959 , n9958 , n5429 );
and ( n9960 , n9955 , n9959 );
and ( n9961 , n7660 , n5487 );
and ( n9962 , n5536 , n5485 );
nor ( n9963 , n9961 , n9962 );
xnor ( n9964 , n9963 , n5478 );
and ( n9965 , n9959 , n9964 );
and ( n9966 , n9955 , n9964 );
or ( n9967 , n9960 , n9965 , n9966 );
and ( n9968 , n5529 , n5468 );
and ( n9969 , n5274 , n5438 );
nor ( n9970 , n9968 , n9969 );
xnor ( n9971 , n9970 , n5405 );
and ( n9972 , n9967 , n9971 );
and ( n9973 , n7690 , n5306 );
and ( n9974 , n7660 , n5304 );
nor ( n9975 , n9973 , n9974 );
xnor ( n9976 , n9975 , n5314 );
and ( n9977 , n9971 , n9976 );
and ( n9978 , n9967 , n9976 );
or ( n9979 , n9972 , n9977 , n9978 );
and ( n9980 , n5233 , n5390 );
and ( n9981 , n5246 , n5387 );
nor ( n9982 , n9980 , n9981 );
xnor ( n9983 , n9982 , n5382 );
or ( n9984 , n9979 , n9983 );
and ( n9985 , n9947 , n9984 );
xor ( n9986 , n9901 , n9903 );
xor ( n9987 , n9986 , n9933 );
and ( n9988 , n9984 , n9987 );
and ( n9989 , n9947 , n9987 );
or ( n9990 , n9985 , n9988 , n9989 );
and ( n9991 , n9945 , n9990 );
xor ( n9992 , n9896 , n9898 );
xor ( n9993 , n9992 , n9936 );
and ( n9994 , n9990 , n9993 );
and ( n9995 , n9945 , n9993 );
or ( n9996 , n9991 , n9994 , n9995 );
xor ( n9997 , n9862 , n9864 );
xor ( n9998 , n9997 , n9939 );
or ( n9999 , n9996 , n9998 );
and ( n10000 , n9942 , n9999 );
and ( n10001 , n9821 , n9999 );
or ( n10002 , n9943 , n10000 , n10001 );
or ( n10003 , n9819 , n10002 );
and ( n10004 , n9816 , n10003 );
and ( n10005 , n9814 , n10003 );
or ( n10006 , n9817 , n10004 , n10005 );
and ( n10007 , n9748 , n10006 );
and ( n10008 , n9746 , n10006 );
or ( n10009 , n9749 , n10007 , n10008 );
or ( n10010 , n9611 , n10009 );
and ( n10011 , n9608 , n10010 );
and ( n10012 , n9433 , n10010 );
or ( n10013 , n9609 , n10011 , n10012 );
and ( n10014 , n9430 , n10013 );
and ( n10015 , n9428 , n10013 );
or ( n10016 , n9431 , n10014 , n10015 );
and ( n10017 , n9334 , n10016 );
xor ( n10018 , n9334 , n10016 );
xor ( n10019 , n9428 , n9430 );
xor ( n10020 , n10019 , n10013 );
not ( n10021 , n10020 );
xor ( n10022 , n9433 , n9608 );
xor ( n10023 , n10022 , n10010 );
not ( n10024 , n10023 );
xnor ( n10025 , n9611 , n10009 );
xor ( n10026 , n9746 , n9748 );
xor ( n10027 , n10026 , n10006 );
not ( n10028 , n10027 );
xor ( n10029 , n9814 , n9816 );
xor ( n10030 , n10029 , n10003 );
xnor ( n10031 , n9819 , n10002 );
xor ( n10032 , n9821 , n9942 );
xor ( n10033 , n10032 , n9999 );
not ( n10034 , n10033 );
xnor ( n10035 , n9996 , n9998 );
xor ( n10036 , n9945 , n9990 );
xor ( n10037 , n10036 , n9993 );
xor ( n10038 , n9876 , n9880 );
xor ( n10039 , n10038 , n9884 );
and ( n10040 , n5254 , n5390 );
and ( n10041 , n5265 , n5387 );
nor ( n10042 , n10040 , n10041 );
xnor ( n10043 , n10042 , n5382 );
xor ( n10044 , n9916 , n9920 );
xor ( n10045 , n10044 , n9882 );
or ( n10046 , n10043 , n10045 );
and ( n10047 , n10039 , n10046 );
and ( n10048 , n5274 , n5414 );
and ( n10049 , n5285 , n5412 );
nor ( n10050 , n10048 , n10049 );
xnor ( n10051 , n10050 , n5420 );
xor ( n10052 , n7541 , n7587 );
buf ( n10053 , n10052 );
buf ( n10054 , n10053 );
buf ( n10055 , n10054 );
and ( n10056 , n10051 , n10055 );
and ( n10057 , n5285 , n5390 );
and ( n10058 , n5254 , n5387 );
nor ( n10059 , n10057 , n10058 );
xnor ( n10060 , n10059 , n5382 );
and ( n10061 , n5529 , n5414 );
and ( n10062 , n5274 , n5412 );
nor ( n10063 , n10061 , n10062 );
xnor ( n10064 , n10063 , n5420 );
and ( n10065 , n10060 , n10064 );
and ( n10066 , n5340 , n5306 );
and ( n10067 , n7639 , n5304 );
nor ( n10068 , n10066 , n10067 );
xnor ( n10069 , n10068 , n5314 );
and ( n10070 , n10064 , n10069 );
and ( n10071 , n10060 , n10069 );
or ( n10072 , n10065 , n10070 , n10071 );
and ( n10073 , n10055 , n10072 );
and ( n10074 , n10051 , n10072 );
or ( n10075 , n10056 , n10073 , n10074 );
and ( n10076 , n10046 , n10075 );
and ( n10077 , n10039 , n10075 );
or ( n10078 , n10047 , n10076 , n10077 );
xor ( n10079 , n9906 , n9927 );
xor ( n10080 , n10079 , n9930 );
and ( n10081 , n10078 , n10080 );
xnor ( n10082 , n9979 , n9983 );
and ( n10083 , n10080 , n10082 );
and ( n10084 , n10078 , n10082 );
or ( n10085 , n10081 , n10083 , n10084 );
xor ( n10086 , n9947 , n9984 );
xor ( n10087 , n10086 , n9987 );
and ( n10088 , n10085 , n10087 );
and ( n10089 , n5265 , n5390 );
and ( n10090 , n5233 , n5387 );
nor ( n10091 , n10089 , n10090 );
xnor ( n10092 , n10091 , n5382 );
xor ( n10093 , n9967 , n9971 );
xor ( n10094 , n10093 , n9976 );
or ( n10095 , n10092 , n10094 );
xor ( n10096 , n9910 , n9911 );
xor ( n10097 , n10096 , n9924 );
xor ( n10098 , n9955 , n9959 );
xor ( n10099 , n10098 , n9964 );
xnor ( n10100 , n10043 , n10045 );
and ( n10101 , n10099 , n10100 );
xor ( n10102 , n9951 , n9954 );
and ( n10103 , n5536 , n7865 );
and ( n10104 , n5545 , n7863 );
nor ( n10105 , n10103 , n10104 );
xnor ( n10106 , n10105 , n5429 );
and ( n10107 , n10102 , n10106 );
and ( n10108 , n7690 , n5487 );
and ( n10109 , n7660 , n5485 );
nor ( n10110 , n10108 , n10109 );
xnor ( n10111 , n10110 , n5478 );
and ( n10112 , n10106 , n10111 );
and ( n10113 , n10102 , n10111 );
or ( n10114 , n10107 , n10112 , n10113 );
and ( n10115 , n10100 , n10114 );
and ( n10116 , n10099 , n10114 );
or ( n10117 , n10101 , n10115 , n10116 );
and ( n10118 , n10097 , n10117 );
xor ( n10119 , n10039 , n10046 );
xor ( n10120 , n10119 , n10075 );
and ( n10121 , n10117 , n10120 );
and ( n10122 , n10097 , n10120 );
or ( n10123 , n10118 , n10121 , n10122 );
and ( n10124 , n10095 , n10123 );
xnor ( n10125 , n10092 , n10094 );
xor ( n10126 , n7542 , n7586 );
buf ( n10127 , n10126 );
buf ( n10128 , n10127 );
buf ( n10129 , n10128 );
and ( n10130 , n5545 , n5468 );
and ( n10131 , n5355 , n5438 );
nor ( n10132 , n10130 , n10131 );
xnor ( n10133 , n10132 , n5405 );
and ( n10134 , n7639 , n5487 );
and ( n10135 , n7690 , n5485 );
nor ( n10136 , n10134 , n10135 );
xnor ( n10137 , n10136 , n5478 );
and ( n10138 , n10133 , n10137 );
and ( n10139 , n10137 , n9952 );
and ( n10140 , n10133 , n9952 );
or ( n10141 , n10138 , n10139 , n10140 );
and ( n10142 , n10129 , n10141 );
and ( n10143 , n5274 , n5390 );
and ( n10144 , n5285 , n5387 );
nor ( n10145 , n10143 , n10144 );
xnor ( n10146 , n10145 , n5382 );
and ( n10147 , n5368 , n5414 );
and ( n10148 , n5529 , n5412 );
nor ( n10149 , n10147 , n10148 );
xnor ( n10150 , n10149 , n5420 );
and ( n10151 , n10146 , n10150 );
and ( n10152 , n7660 , n7865 );
and ( n10153 , n5536 , n7863 );
nor ( n10154 , n10152 , n10153 );
xnor ( n10155 , n10154 , n5429 );
and ( n10156 , n10150 , n10155 );
and ( n10157 , n10146 , n10155 );
or ( n10158 , n10151 , n10156 , n10157 );
and ( n10159 , n10141 , n10158 );
and ( n10160 , n10129 , n10158 );
or ( n10161 , n10142 , n10159 , n10160 );
xor ( n10162 , n10051 , n10055 );
xor ( n10163 , n10162 , n10072 );
and ( n10164 , n10161 , n10163 );
xor ( n10165 , n10060 , n10064 );
xor ( n10166 , n10165 , n10069 );
xor ( n10167 , n10102 , n10106 );
xor ( n10168 , n10167 , n10111 );
and ( n10169 , n10166 , n10168 );
xor ( n10170 , n7543 , n7585 );
buf ( n10171 , n10170 );
buf ( n10172 , n10171 );
buf ( n10173 , n10172 );
xor ( n10174 , n10133 , n10137 );
xor ( n10175 , n10174 , n9952 );
and ( n10176 , n10173 , n10175 );
and ( n10177 , n5536 , n5468 );
and ( n10178 , n5545 , n5438 );
nor ( n10179 , n10177 , n10178 );
xnor ( n10180 , n10179 , n5405 );
and ( n10181 , n7690 , n7865 );
and ( n10182 , n7660 , n7863 );
nor ( n10183 , n10181 , n10182 );
xnor ( n10184 , n10183 , n5429 );
and ( n10185 , n10180 , n10184 );
and ( n10186 , n5340 , n5487 );
and ( n10187 , n7639 , n5485 );
nor ( n10188 , n10186 , n10187 );
xnor ( n10189 , n10188 , n5478 );
and ( n10190 , n10184 , n10189 );
and ( n10191 , n10180 , n10189 );
or ( n10192 , n10185 , n10190 , n10191 );
and ( n10193 , n10175 , n10192 );
and ( n10194 , n10173 , n10192 );
or ( n10195 , n10176 , n10193 , n10194 );
and ( n10196 , n10168 , n10195 );
and ( n10197 , n10166 , n10195 );
or ( n10198 , n10169 , n10196 , n10197 );
and ( n10199 , n10163 , n10198 );
and ( n10200 , n10161 , n10198 );
or ( n10201 , n10164 , n10199 , n10200 );
and ( n10202 , n10125 , n10201 );
xor ( n10203 , n10097 , n10117 );
xor ( n10204 , n10203 , n10120 );
and ( n10205 , n10201 , n10204 );
and ( n10206 , n10125 , n10204 );
or ( n10207 , n10202 , n10205 , n10206 );
and ( n10208 , n10123 , n10207 );
and ( n10209 , n10095 , n10207 );
or ( n10210 , n10124 , n10208 , n10209 );
and ( n10211 , n10087 , n10210 );
and ( n10212 , n10085 , n10210 );
or ( n10213 , n10088 , n10211 , n10212 );
and ( n10214 , n10037 , n10213 );
xor ( n10215 , n10037 , n10213 );
xor ( n10216 , n10085 , n10087 );
xor ( n10217 , n10216 , n10210 );
xor ( n10218 , n10078 , n10080 );
xor ( n10219 , n10218 , n10082 );
xor ( n10220 , n10095 , n10123 );
xor ( n10221 , n10220 , n10207 );
and ( n10222 , n10219 , n10221 );
xor ( n10223 , n10219 , n10221 );
xor ( n10224 , n10099 , n10100 );
xor ( n10225 , n10224 , n10114 );
xor ( n10226 , n10129 , n10141 );
xor ( n10227 , n10226 , n10158 );
and ( n10228 , n5355 , n5414 );
and ( n10229 , n5368 , n5412 );
nor ( n10230 , n10228 , n10229 );
xnor ( n10231 , n10230 , n5420 );
and ( n10232 , n5340 , n5485 );
not ( n10233 , n10232 );
and ( n10234 , n10233 , n5478 );
and ( n10235 , n10231 , n10234 );
xor ( n10236 , n10146 , n10150 );
xor ( n10237 , n10236 , n10155 );
and ( n10238 , n10235 , n10237 );
and ( n10239 , n5529 , n5390 );
and ( n10240 , n5274 , n5387 );
nor ( n10241 , n10239 , n10240 );
xnor ( n10242 , n10241 , n5382 );
xor ( n10243 , n7544 , n7584 );
buf ( n10244 , n10243 );
buf ( n10245 , n10244 );
buf ( n10246 , n10245 );
and ( n10247 , n10242 , n10246 );
xor ( n10248 , n10180 , n10184 );
xor ( n10249 , n10248 , n10189 );
and ( n10250 , n10246 , n10249 );
and ( n10251 , n10242 , n10249 );
or ( n10252 , n10247 , n10250 , n10251 );
and ( n10253 , n10237 , n10252 );
and ( n10254 , n10235 , n10252 );
or ( n10255 , n10238 , n10253 , n10254 );
and ( n10256 , n10227 , n10255 );
xor ( n10257 , n10166 , n10168 );
xor ( n10258 , n10257 , n10195 );
and ( n10259 , n10255 , n10258 );
and ( n10260 , n10227 , n10258 );
or ( n10261 , n10256 , n10259 , n10260 );
and ( n10262 , n10225 , n10261 );
xor ( n10263 , n10161 , n10163 );
xor ( n10264 , n10263 , n10198 );
and ( n10265 , n10261 , n10264 );
and ( n10266 , n10225 , n10264 );
or ( n10267 , n10262 , n10265 , n10266 );
xor ( n10268 , n10125 , n10201 );
xor ( n10269 , n10268 , n10204 );
and ( n10270 , n10267 , n10269 );
xor ( n10271 , n10267 , n10269 );
xor ( n10272 , n10225 , n10261 );
xor ( n10273 , n10272 , n10264 );
xor ( n10274 , n10231 , n10234 );
and ( n10275 , n5545 , n5414 );
and ( n10276 , n5355 , n5412 );
nor ( n10277 , n10275 , n10276 );
xnor ( n10278 , n10277 , n5420 );
and ( n10279 , n7660 , n5468 );
and ( n10280 , n5536 , n5438 );
nor ( n10281 , n10279 , n10280 );
xnor ( n10282 , n10281 , n5405 );
or ( n10283 , n10278 , n10282 );
and ( n10284 , n10274 , n10283 );
and ( n10285 , n5368 , n5390 );
and ( n10286 , n5529 , n5387 );
nor ( n10287 , n10285 , n10286 );
xnor ( n10288 , n10287 , n5382 );
and ( n10289 , n7639 , n7865 );
and ( n10290 , n7690 , n7863 );
nor ( n10291 , n10289 , n10290 );
xnor ( n10292 , n10291 , n5429 );
and ( n10293 , n10288 , n10292 );
and ( n10294 , n10292 , n10232 );
and ( n10295 , n10288 , n10232 );
or ( n10296 , n10293 , n10294 , n10295 );
and ( n10297 , n10283 , n10296 );
and ( n10298 , n10274 , n10296 );
or ( n10299 , n10284 , n10297 , n10298 );
xor ( n10300 , n10173 , n10175 );
xor ( n10301 , n10300 , n10192 );
and ( n10302 , n10299 , n10301 );
xor ( n10303 , n7547 , n7582 );
buf ( n10304 , n10303 );
buf ( n10305 , n10304 );
buf ( n10306 , n10305 );
xnor ( n10307 , n10278 , n10282 );
and ( n10308 , n10306 , n10307 );
and ( n10309 , n5536 , n5414 );
and ( n10310 , n5545 , n5412 );
nor ( n10311 , n10309 , n10310 );
xnor ( n10312 , n10311 , n5420 );
and ( n10313 , n7690 , n5468 );
and ( n10314 , n7660 , n5438 );
nor ( n10315 , n10313 , n10314 );
xnor ( n10316 , n10315 , n5405 );
and ( n10317 , n10312 , n10316 );
and ( n10318 , n5340 , n7865 );
and ( n10319 , n7639 , n7863 );
nor ( n10320 , n10318 , n10319 );
xnor ( n10321 , n10320 , n5429 );
and ( n10322 , n10316 , n10321 );
and ( n10323 , n10312 , n10321 );
or ( n10324 , n10317 , n10322 , n10323 );
and ( n10325 , n10307 , n10324 );
and ( n10326 , n10306 , n10324 );
or ( n10327 , n10308 , n10325 , n10326 );
xor ( n10328 , n10242 , n10246 );
xor ( n10329 , n10328 , n10249 );
and ( n10330 , n10327 , n10329 );
xor ( n10331 , n10274 , n10283 );
xor ( n10332 , n10331 , n10296 );
and ( n10333 , n10329 , n10332 );
and ( n10334 , n10327 , n10332 );
or ( n10335 , n10330 , n10333 , n10334 );
and ( n10336 , n10301 , n10335 );
and ( n10337 , n10299 , n10335 );
or ( n10338 , n10302 , n10336 , n10337 );
xor ( n10339 , n10227 , n10255 );
xor ( n10340 , n10339 , n10258 );
and ( n10341 , n10338 , n10340 );
xor ( n10342 , n10235 , n10237 );
xor ( n10343 , n10342 , n10252 );
xor ( n10344 , n10299 , n10301 );
xor ( n10345 , n10344 , n10335 );
and ( n10346 , n10343 , n10345 );
and ( n10347 , n5355 , n5390 );
and ( n10348 , n5368 , n5387 );
nor ( n10349 , n10347 , n10348 );
xnor ( n10350 , n10349 , n5382 );
and ( n10351 , n5340 , n7863 );
not ( n10352 , n10351 );
and ( n10353 , n10352 , n5429 );
and ( n10354 , n10350 , n10353 );
xor ( n10355 , n7548 , n7581 );
buf ( n10356 , n10355 );
buf ( n10357 , n10356 );
buf ( n10358 , n10357 );
and ( n10359 , n10353 , n10358 );
and ( n10360 , n10350 , n10358 );
or ( n10361 , n10354 , n10359 , n10360 );
xor ( n10362 , n10288 , n10292 );
xor ( n10363 , n10362 , n10232 );
and ( n10364 , n10361 , n10363 );
xor ( n10365 , n10312 , n10316 );
xor ( n10366 , n10365 , n10321 );
and ( n10367 , n5545 , n5390 );
and ( n10368 , n5355 , n5387 );
nor ( n10369 , n10367 , n10368 );
xnor ( n10370 , n10369 , n5382 );
and ( n10371 , n7660 , n5414 );
and ( n10372 , n5536 , n5412 );
nor ( n10373 , n10371 , n10372 );
xnor ( n10374 , n10373 , n5420 );
and ( n10375 , n10370 , n10374 );
and ( n10376 , n7639 , n5468 );
and ( n10377 , n7690 , n5438 );
nor ( n10378 , n10376 , n10377 );
xnor ( n10379 , n10378 , n5405 );
and ( n10380 , n10374 , n10379 );
and ( n10381 , n10370 , n10379 );
or ( n10382 , n10375 , n10380 , n10381 );
and ( n10383 , n10366 , n10382 );
xor ( n10384 , n10350 , n10353 );
xor ( n10385 , n10384 , n10358 );
and ( n10386 , n10382 , n10385 );
and ( n10387 , n10366 , n10385 );
or ( n10388 , n10383 , n10386 , n10387 );
and ( n10389 , n10363 , n10388 );
and ( n10390 , n10361 , n10388 );
or ( n10391 , n10364 , n10389 , n10390 );
xor ( n10392 , n10327 , n10329 );
xor ( n10393 , n10392 , n10332 );
and ( n10394 , n10391 , n10393 );
xor ( n10395 , n10306 , n10307 );
xor ( n10396 , n10395 , n10324 );
xor ( n10397 , n10361 , n10363 );
xor ( n10398 , n10397 , n10388 );
and ( n10399 , n10396 , n10398 );
xor ( n10400 , n7549 , n7580 );
buf ( n10401 , n10400 );
buf ( n10402 , n10401 );
buf ( n10403 , n10402 );
and ( n10404 , n10351 , n10403 );
and ( n10405 , n5536 , n5390 );
and ( n10406 , n5545 , n5387 );
nor ( n10407 , n10405 , n10406 );
xnor ( n10408 , n10407 , n5382 );
and ( n10409 , n7690 , n5414 );
and ( n10410 , n7660 , n5412 );
nor ( n10411 , n10409 , n10410 );
xnor ( n10412 , n10411 , n5420 );
and ( n10413 , n10408 , n10412 );
and ( n10414 , n5340 , n5468 );
and ( n10415 , n7639 , n5438 );
nor ( n10416 , n10414 , n10415 );
xnor ( n10417 , n10416 , n5405 );
and ( n10418 , n10412 , n10417 );
and ( n10419 , n10408 , n10417 );
or ( n10420 , n10413 , n10418 , n10419 );
and ( n10421 , n10403 , n10420 );
and ( n10422 , n10351 , n10420 );
or ( n10423 , n10404 , n10421 , n10422 );
xor ( n10424 , n10366 , n10382 );
xor ( n10425 , n10424 , n10385 );
and ( n10426 , n10423 , n10425 );
xor ( n10427 , n10370 , n10374 );
xor ( n10428 , n10427 , n10379 );
and ( n10429 , n5340 , n5438 );
not ( n10430 , n10429 );
and ( n10431 , n10430 , n5405 );
xor ( n10432 , n7576 , n7578 );
buf ( n10433 , n10432 );
buf ( n10434 , n10433 );
buf ( n10435 , n10434 );
and ( n10436 , n10431 , n10435 );
and ( n10437 , n7660 , n5390 );
and ( n10438 , n5536 , n5387 );
nor ( n10439 , n10437 , n10438 );
xnor ( n10440 , n10439 , n5382 );
and ( n10441 , n7639 , n5414 );
and ( n10442 , n7690 , n5412 );
nor ( n10443 , n10441 , n10442 );
xnor ( n10444 , n10443 , n5420 );
and ( n10445 , n10440 , n10444 );
and ( n10446 , n10444 , n10429 );
and ( n10447 , n10440 , n10429 );
or ( n10448 , n10445 , n10446 , n10447 );
and ( n10449 , n10435 , n10448 );
and ( n10450 , n10431 , n10448 );
or ( n10451 , n10436 , n10449 , n10450 );
and ( n10452 , n10428 , n10451 );
xor ( n10453 , n10351 , n10403 );
xor ( n10454 , n10453 , n10420 );
and ( n10455 , n10451 , n10454 );
and ( n10456 , n10428 , n10454 );
or ( n10457 , n10452 , n10455 , n10456 );
and ( n10458 , n10425 , n10457 );
and ( n10459 , n10423 , n10457 );
or ( n10460 , n10426 , n10458 , n10459 );
and ( n10461 , n10398 , n10460 );
and ( n10462 , n10396 , n10460 );
or ( n10463 , n10399 , n10461 , n10462 );
and ( n10464 , n10393 , n10463 );
and ( n10465 , n10391 , n10463 );
or ( n10466 , n10394 , n10464 , n10465 );
and ( n10467 , n10345 , n10466 );
and ( n10468 , n10343 , n10466 );
or ( n10469 , n10346 , n10467 , n10468 );
and ( n10470 , n10340 , n10469 );
and ( n10471 , n10338 , n10469 );
or ( n10472 , n10341 , n10470 , n10471 );
and ( n10473 , n10273 , n10472 );
xor ( n10474 , n10273 , n10472 );
xor ( n10475 , n10338 , n10340 );
xor ( n10476 , n10475 , n10469 );
not ( n10477 , n10476 );
xor ( n10478 , n10343 , n10345 );
xor ( n10479 , n10478 , n10466 );
not ( n10480 , n10479 );
xor ( n10481 , n10391 , n10393 );
xor ( n10482 , n10481 , n10463 );
not ( n10483 , n10482 );
xor ( n10484 , n10396 , n10398 );
xor ( n10485 , n10484 , n10460 );
not ( n10486 , n10485 );
xor ( n10487 , n10423 , n10425 );
xor ( n10488 , n10487 , n10457 );
xor ( n10489 , n10408 , n10412 );
xor ( n10490 , n10489 , n10417 );
not ( n10491 , n7578 );
buf ( n10492 , n10491 );
buf ( n10493 , n10492 );
buf ( n10494 , n10493 );
and ( n10495 , n7690 , n5390 );
and ( n10496 , n7660 , n5387 );
nor ( n10497 , n10495 , n10496 );
xnor ( n10498 , n10497 , n5382 );
and ( n10499 , n5340 , n5414 );
and ( n10500 , n7639 , n5412 );
nor ( n10501 , n10499 , n10500 );
xnor ( n10502 , n10501 , n5420 );
and ( n10503 , n10498 , n10502 );
and ( n10504 , n5340 , n5412 );
not ( n10505 , n10504 );
and ( n10506 , n10505 , n5420 );
and ( n10507 , n10502 , n10506 );
and ( n10508 , n10498 , n10506 );
or ( n10509 , n10503 , n10507 , n10508 );
and ( n10510 , n10494 , n10509 );
xor ( n10511 , n10440 , n10444 );
xor ( n10512 , n10511 , n10429 );
and ( n10513 , n10509 , n10512 );
and ( n10514 , n10494 , n10512 );
or ( n10515 , n10510 , n10513 , n10514 );
and ( n10516 , n10490 , n10515 );
xor ( n10517 , n10431 , n10435 );
xor ( n10518 , n10517 , n10448 );
and ( n10519 , n10515 , n10518 );
and ( n10520 , n10490 , n10518 );
or ( n10521 , n10516 , n10519 , n10520 );
xor ( n10522 , n10428 , n10451 );
xor ( n10523 , n10522 , n10454 );
and ( n10524 , n10521 , n10523 );
xor ( n10525 , n10521 , n10523 );
xor ( n10526 , n10490 , n10515 );
xor ( n10527 , n10526 , n10518 );
xnor ( n10528 , n7568 , n7570 );
buf ( n10529 , n10528 );
buf ( n10530 , n10529 );
buf ( n10531 , n10530 );
and ( n10532 , n7639 , n5390 );
and ( n10533 , n7690 , n5387 );
nor ( n10534 , n10532 , n10533 );
xnor ( n10535 , n10534 , n5382 );
and ( n10536 , n10504 , n10535 );
and ( n10537 , n10531 , n10536 );
xor ( n10538 , n10498 , n10502 );
xor ( n10539 , n10538 , n10506 );
and ( n10540 , n10536 , n10539 );
and ( n10541 , n10531 , n10539 );
or ( n10542 , n10537 , n10540 , n10541 );
xor ( n10543 , n10494 , n10509 );
xor ( n10544 , n10543 , n10512 );
and ( n10545 , n10542 , n10544 );
xor ( n10546 , n10542 , n10544 );
xnor ( n10547 , n7566 , n7567 );
buf ( n10548 , n10547 );
buf ( n10549 , n10548 );
buf ( n10550 , n10549 );
xor ( n10551 , n10504 , n10535 );
and ( n10552 , n10550 , n10551 );
and ( n10553 , n5340 , n5390 );
and ( n10554 , n7639 , n5387 );
nor ( n10555 , n10553 , n10554 );
xnor ( n10556 , n10555 , n5382 );
buf ( n10557 , n5340 );
not ( n10558 , n10557 );
and ( n10559 , n10558 , n5382 );
and ( n10560 , n10556 , n10559 );
and ( n10561 , n10551 , n10560 );
and ( n10562 , n10550 , n10560 );
or ( n10563 , n10552 , n10561 , n10562 );
xor ( n10564 , n10531 , n10536 );
xor ( n10565 , n10564 , n10539 );
and ( n10566 , n10563 , n10565 );
xor ( n10567 , n10563 , n10565 );
xor ( n10568 , n10550 , n10551 );
xor ( n10569 , n10568 , n10560 );
xor ( n10570 , n10556 , n10559 );
buf ( n10571 , n6314 );
buf ( n10572 , n10571 );
buf ( n10573 , n10572 );
buf ( n10574 , n10573 );
and ( n10575 , n10557 , n10574 );
and ( n10576 , n10570 , n10575 );
and ( n10577 , n10569 , n10576 );
and ( n10578 , n10567 , n10577 );
or ( n10579 , n10566 , n10578 );
and ( n10580 , n10546 , n10579 );
or ( n10581 , n10545 , n10580 );
and ( n10582 , n10527 , n10581 );
and ( n10583 , n10525 , n10582 );
or ( n10584 , n10524 , n10583 );
and ( n10585 , n10488 , n10584 );
and ( n10586 , n10486 , n10585 );
or ( n10587 , n10485 , n10586 );
and ( n10588 , n10483 , n10587 );
or ( n10589 , n10482 , n10588 );
and ( n10590 , n10480 , n10589 );
or ( n10591 , n10479 , n10590 );
and ( n10592 , n10477 , n10591 );
or ( n10593 , n10476 , n10592 );
and ( n10594 , n10474 , n10593 );
or ( n10595 , n10473 , n10594 );
and ( n10596 , n10271 , n10595 );
or ( n10597 , n10270 , n10596 );
and ( n10598 , n10223 , n10597 );
or ( n10599 , n10222 , n10598 );
and ( n10600 , n10217 , n10599 );
and ( n10601 , n10215 , n10600 );
or ( n10602 , n10214 , n10601 );
and ( n10603 , n10035 , n10602 );
and ( n10604 , n10034 , n10603 );
or ( n10605 , n10033 , n10604 );
and ( n10606 , n10031 , n10605 );
and ( n10607 , n10030 , n10606 );
and ( n10608 , n10028 , n10607 );
or ( n10609 , n10027 , n10608 );
and ( n10610 , n10025 , n10609 );
and ( n10611 , n10024 , n10610 );
or ( n10612 , n10023 , n10611 );
and ( n10613 , n10021 , n10612 );
or ( n10614 , n10020 , n10613 );
and ( n10615 , n10018 , n10614 );
or ( n10616 , n10017 , n10615 );
and ( n10617 , n9332 , n10616 );
and ( n10618 , n9331 , n10617 );
or ( n10619 , n9330 , n10618 );
and ( n10620 , n9328 , n10619 );
or ( n10621 , n9327 , n10620 );
and ( n10622 , n9325 , n10621 );
and ( n10623 , n9324 , n10622 );
or ( n10624 , n9323 , n10623 );
and ( n10625 , n8860 , n10624 );
or ( n10626 , n8859 , n10625 );
and ( n10627 , n8502 , n10626 );
xor ( n10628 , n8500 , n10627 );
buf ( n10629 , n10628 );
buf ( n10630 , n10629 );
buf ( n10631 , n10630 );
and ( n10632 , n5230 , n10631 );
and ( n10633 , n5229 , n10631 );
or ( n10634 , n5231 , n10632 , n10633 );
and ( n10635 , n5228 , n10634 );
xor ( n10636 , n4992 , n4993 );
and ( n10637 , n10634 , n10636 );
and ( n10638 , n5228 , n10636 );
or ( n10639 , n10635 , n10637 , n10638 );
and ( n10640 , n5224 , n10639 );
and ( n10641 , n5215 , n10639 );
or ( n10642 , n5225 , n10640 , n10641 );
xor ( n10643 , n4928 , n4929 );
xor ( n10644 , n10643 , n4931 );
xor ( n10645 , n4941 , n4942 );
xor ( n10646 , n10645 , n4944 );
and ( n10647 , n10644 , n10646 );
xor ( n10648 , n4948 , n4949 );
xor ( n10649 , n10648 , n4951 );
and ( n10650 , n10646 , n10649 );
and ( n10651 , n10644 , n10649 );
or ( n10652 , n10647 , n10650 , n10651 );
and ( n10653 , n10642 , n10652 );
xor ( n10654 , n4874 , n4875 );
xor ( n10655 , n10654 , n4878 );
and ( n10656 , n10652 , n10655 );
and ( n10657 , n10642 , n10655 );
or ( n10658 , n10653 , n10656 , n10657 );
and ( n10659 , n5207 , n10658 );
and ( n10660 , n5139 , n10658 );
or ( n10661 , n5208 , n10659 , n10660 );
xor ( n10662 , n4882 , n4895 );
xor ( n10663 , n10662 , n4905 );
xor ( n10664 , n4920 , n4925 );
xor ( n10665 , n10664 , n4934 );
and ( n10666 , n10663 , n10665 );
xor ( n10667 , n4947 , n4954 );
xor ( n10668 , n10667 , n4974 );
and ( n10669 , n10665 , n10668 );
and ( n10670 , n10663 , n10668 );
or ( n10671 , n10666 , n10669 , n10670 );
xor ( n10672 , n4795 , n4797 );
xor ( n10673 , n10672 , n4800 );
and ( n10674 , n10671 , n10673 );
xor ( n10675 , n4805 , n4807 );
xor ( n10676 , n10675 , n4810 );
and ( n10677 , n10673 , n10676 );
and ( n10678 , n10671 , n10676 );
or ( n10679 , n10674 , n10677 , n10678 );
and ( n10680 , n10661 , n10679 );
xor ( n10681 , n4843 , n4853 );
xor ( n10682 , n10681 , n4864 );
xor ( n10683 , n4881 , n4908 );
xor ( n10684 , n10683 , n4937 );
and ( n10685 , n10682 , n10684 );
xor ( n10686 , n4977 , n5007 );
xor ( n10687 , n10686 , n5010 );
and ( n10688 , n10684 , n10687 );
and ( n10689 , n10682 , n10687 );
or ( n10690 , n10685 , n10688 , n10689 );
and ( n10691 , n10679 , n10690 );
and ( n10692 , n10661 , n10690 );
or ( n10693 , n10680 , n10691 , n10692 );
xor ( n10694 , n4785 , n4787 );
xor ( n10695 , n10694 , n4790 );
xor ( n10696 , n4803 , n4813 );
xor ( n10697 , n10696 , n4867 );
and ( n10698 , n10695 , n10697 );
xor ( n10699 , n4940 , n5013 );
xor ( n10700 , n10699 , n5016 );
and ( n10701 , n10697 , n10700 );
and ( n10702 , n10695 , n10700 );
or ( n10703 , n10698 , n10701 , n10702 );
and ( n10704 , n10693 , n10703 );
xor ( n10705 , n4774 , n4776 );
xor ( n10706 , n10705 , n4779 );
and ( n10707 , n10703 , n10706 );
and ( n10708 , n10693 , n10706 );
or ( n10709 , n10704 , n10707 , n10708 );
and ( n10710 , n5069 , n10709 );
and ( n10711 , n5035 , n10709 );
or ( n10712 , n5070 , n10710 , n10711 );
xor ( n10713 , n4631 , n4649 );
xor ( n10714 , n10713 , n4652 );
and ( n10715 , n10712 , n10714 );
xor ( n10716 , n4770 , n5025 );
xor ( n10717 , n10716 , n5028 );
and ( n10718 , n10714 , n10717 );
and ( n10719 , n10712 , n10717 );
or ( n10720 , n10715 , n10718 , n10719 );
and ( n10721 , n5032 , n10720 );
and ( n10722 , n5031 , n10720 );
or ( n10723 , n5033 , n10721 , n10722 );
and ( n10724 , n4658 , n10723 );
xor ( n10725 , n4438 , n4440 );
xor ( n10726 , n10725 , n4446 );
and ( n10727 , n10723 , n10726 );
and ( n10728 , n4658 , n10726 );
or ( n10729 , n10724 , n10727 , n10728 );
xor ( n10730 , n4436 , n4449 );
xor ( n10731 , n10730 , n4452 );
and ( n10732 , n10729 , n10731 );
xor ( n10733 , n10729 , n10731 );
xor ( n10734 , n4658 , n10723 );
xor ( n10735 , n10734 , n10726 );
xor ( n10736 , n4461 , n4514 );
xor ( n10737 , n10736 , n4655 );
xor ( n10738 , n5031 , n5032 );
xor ( n10739 , n10738 , n10720 );
and ( n10740 , n10737 , n10739 );
xor ( n10741 , n4762 , n4764 );
xor ( n10742 , n10741 , n4767 );
xor ( n10743 , n4772 , n4782 );
xor ( n10744 , n10743 , n5022 );
and ( n10745 , n10742 , n10744 );
xor ( n10746 , n4793 , n4870 );
xor ( n10747 , n10746 , n5019 );
xor ( n10748 , n4999 , n5001 );
xor ( n10749 , n10748 , n5004 );
xor ( n10750 , n4956 , n4963 );
xor ( n10751 , n10750 , n4971 );
xor ( n10752 , n4987 , n4994 );
xor ( n10753 , n10752 , n4996 );
and ( n10754 , n10751 , n10753 );
xor ( n10755 , n5081 , n5103 );
xor ( n10756 , n10755 , n5115 );
and ( n10757 , n10753 , n10756 );
and ( n10758 , n10751 , n10756 );
or ( n10759 , n10754 , n10757 , n10758 );
and ( n10760 , n10749 , n10759 );
xor ( n10761 , n5128 , n5130 );
xor ( n10762 , n10761 , n5133 );
xor ( n10763 , n5141 , n5143 );
xor ( n10764 , n10763 , n5146 );
and ( n10765 , n10762 , n10764 );
and ( n10766 , n4579 , n1530 );
and ( n10767 , n3246 , n2948 );
and ( n10768 , n10766 , n10767 );
and ( n10769 , n2764 , n3929 );
and ( n10770 , n10767 , n10769 );
and ( n10771 , n10766 , n10769 );
or ( n10772 , n10768 , n10770 , n10771 );
and ( n10773 , n4385 , n1711 );
and ( n10774 , n3339 , n2577 );
and ( n10775 , n10773 , n10774 );
and ( n10776 , n2937 , n3627 );
and ( n10777 , n10774 , n10776 );
and ( n10778 , n10773 , n10776 );
or ( n10779 , n10775 , n10777 , n10778 );
and ( n10780 , n10772 , n10779 );
and ( n10781 , n1995 , n2718 );
and ( n10782 , n2723 , n1990 );
and ( n10783 , n10781 , n10782 );
and ( n10784 , n4138 , n1860 );
and ( n10785 , n10783 , n10784 );
and ( n10786 , n2477 , n5077 );
and ( n10787 , n10784 , n10786 );
and ( n10788 , n10783 , n10786 );
or ( n10789 , n10785 , n10787 , n10788 );
and ( n10790 , n10779 , n10789 );
and ( n10791 , n10772 , n10789 );
or ( n10792 , n10780 , n10790 , n10791 );
and ( n10793 , n10764 , n10792 );
and ( n10794 , n10762 , n10792 );
or ( n10795 , n10765 , n10793 , n10794 );
and ( n10796 , n10759 , n10795 );
and ( n10797 , n10749 , n10795 );
or ( n10798 , n10760 , n10796 , n10797 );
xor ( n10799 , n4965 , n4966 );
xor ( n10800 , n10799 , n4968 );
xor ( n10801 , n5107 , n5110 );
xor ( n10802 , n10801 , n5112 );
and ( n10803 , n10800 , n10802 );
xor ( n10804 , n5122 , n5123 );
xor ( n10805 , n10804 , n5125 );
xor ( n10806 , n5095 , n5098 );
xor ( n10807 , n10806 , n5100 );
and ( n10808 , n10805 , n10807 );
xor ( n10809 , n5160 , n5167 );
and ( n10810 , n10807 , n10809 );
and ( n10811 , n10805 , n10809 );
or ( n10812 , n10808 , n10810 , n10811 );
and ( n10813 , n10803 , n10812 );
and ( n10814 , n1724 , n3288 );
and ( n10815 , n3293 , n1719 );
and ( n10816 , n10814 , n10815 );
and ( n10817 , n4721 , n1465 );
and ( n10818 , n10816 , n10817 );
and ( n10819 , n3833 , n2040 );
and ( n10820 , n10817 , n10819 );
and ( n10821 , n10816 , n10819 );
or ( n10822 , n10818 , n10820 , n10821 );
and ( n10823 , n2048 , n2586 );
and ( n10824 , n2591 , n2059 );
and ( n10825 , n10823 , n10824 );
and ( n10826 , n5177 , n1360 );
and ( n10827 , n10825 , n10826 );
and ( n10828 , n2634 , n4522 );
and ( n10829 , n10826 , n10828 );
and ( n10830 , n10825 , n10828 );
or ( n10831 , n10827 , n10829 , n10830 );
and ( n10832 , n10822 , n10831 );
and ( n10833 , n1778 , n3146 );
and ( n10834 , n3151 , n1789 );
and ( n10835 , n10833 , n10834 );
and ( n10836 , n2255 , n2492 );
and ( n10837 , n2497 , n2250 );
and ( n10838 , n10836 , n10837 );
and ( n10839 , n10835 , n10838 );
and ( n10840 , n3645 , n2407 );
and ( n10841 , n10838 , n10840 );
and ( n10842 , n10835 , n10840 );
or ( n10843 , n10839 , n10841 , n10842 );
and ( n10844 , n10831 , n10843 );
and ( n10845 , n10822 , n10843 );
or ( n10846 , n10832 , n10844 , n10845 );
and ( n10847 , n10812 , n10846 );
and ( n10848 , n10803 , n10846 );
or ( n10849 , n10813 , n10847 , n10848 );
and ( n10850 , n1694 , n3449 );
and ( n10851 , n3454 , n1689 );
and ( n10852 , n10850 , n10851 );
and ( n10853 , n1911 , n2923 );
and ( n10854 , n2928 , n1906 );
and ( n10855 , n10853 , n10854 );
and ( n10856 , n10852 , n10855 );
and ( n10857 , n3169 , n3301 );
and ( n10858 , n10855 , n10857 );
and ( n10859 , n10852 , n10857 );
or ( n10860 , n10856 , n10858 , n10859 );
buf ( n10861 , n7637 );
buf ( n10862 , n10861 );
not ( n10863 , n10862 );
and ( n10864 , n1279 , n10862 );
nor ( n10865 , n10863 , n10864 );
and ( n10866 , n4739 , n1348 );
and ( n10867 , n10865 , n10866 );
buf ( n10868 , n7637 );
buf ( n10869 , n10868 );
and ( n10870 , n1291 , n10869 );
not ( n10871 , n10869 );
nor ( n10872 , n10870 , n10871 );
and ( n10873 , n1353 , n4734 );
and ( n10874 , n10872 , n10873 );
and ( n10875 , n10867 , n10874 );
and ( n10876 , n10860 , n10875 );
xor ( n10877 , n5154 , n5155 );
xor ( n10878 , n10877 , n5157 );
xor ( n10879 , n5161 , n5162 );
xor ( n10880 , n10879 , n5164 );
and ( n10881 , n10878 , n10880 );
and ( n10882 , n10875 , n10881 );
and ( n10883 , n10860 , n10881 );
or ( n10884 , n10876 , n10882 , n10883 );
buf ( n10885 , n5380 );
buf ( n10886 , n10885 );
and ( n10887 , n10886 , n1287 );
xnor ( n10888 , n5219 , n5220 );
and ( n10889 , n10887 , n10888 );
xor ( n10890 , n5089 , n5094 );
and ( n10891 , n10888 , n10890 );
and ( n10892 , n10887 , n10890 );
or ( n10893 , n10889 , n10891 , n10892 );
xor ( n10894 , n5105 , n5106 );
xor ( n10895 , n5120 , n5121 );
and ( n10896 , n10894 , n10895 );
xor ( n10897 , n5108 , n5109 );
and ( n10898 , n10895 , n10897 );
and ( n10899 , n10894 , n10897 );
or ( n10900 , n10896 , n10898 , n10899 );
and ( n10901 , n10893 , n10900 );
xor ( n10902 , n5096 , n5097 );
xor ( n10903 , n5226 , n5227 );
and ( n10904 , n10902 , n10903 );
and ( n10905 , n10886 , n1360 );
and ( n10906 , n3246 , n3301 );
and ( n10907 , n10905 , n10906 );
and ( n10908 , n3169 , n3627 );
and ( n10909 , n10906 , n10908 );
and ( n10910 , n10905 , n10908 );
or ( n10911 , n10907 , n10909 , n10910 );
and ( n10912 , n10903 , n10911 );
and ( n10913 , n10902 , n10911 );
or ( n10914 , n10904 , n10912 , n10913 );
and ( n10915 , n10900 , n10914 );
and ( n10916 , n10893 , n10914 );
or ( n10917 , n10901 , n10915 , n10916 );
and ( n10918 , n10884 , n10917 );
buf ( n10919 , n2309 );
xor ( n10920 , n8502 , n10626 );
buf ( n10921 , n10920 );
buf ( n10922 , n10921 );
buf ( n10923 , n10922 );
and ( n10924 , n10919 , n10923 );
and ( n10925 , n1275 , n5086 );
and ( n10926 , n1317 , n4982 );
or ( n10927 , n10925 , n10926 );
and ( n10928 , n10924 , n10927 );
and ( n10929 , n5091 , n1293 );
and ( n10930 , n4989 , n1312 );
and ( n10931 , n10929 , n10930 );
buf ( n10932 , n5385 );
buf ( n10933 , n10932 );
and ( n10934 , n10933 , n1287 );
and ( n10935 , n10930 , n10934 );
and ( n10936 , n10929 , n10934 );
or ( n10937 , n10931 , n10935 , n10936 );
and ( n10938 , n10927 , n10937 );
and ( n10939 , n10924 , n10937 );
or ( n10940 , n10928 , n10938 , n10939 );
xor ( n10941 , n5178 , n5179 );
xor ( n10942 , n10941 , n5182 );
and ( n10943 , n10940 , n10942 );
xor ( n10944 , n5187 , n5188 );
xor ( n10945 , n10944 , n5190 );
and ( n10946 , n10942 , n10945 );
and ( n10947 , n10940 , n10945 );
or ( n10948 , n10943 , n10946 , n10947 );
and ( n10949 , n10917 , n10948 );
and ( n10950 , n10884 , n10948 );
or ( n10951 , n10918 , n10949 , n10950 );
and ( n10952 , n10849 , n10951 );
xor ( n10953 , n5195 , n5196 );
xor ( n10954 , n10953 , n5198 );
xor ( n10955 , n5209 , n5210 );
xor ( n10956 , n10955 , n5212 );
and ( n10957 , n10954 , n10956 );
xor ( n10958 , n5216 , n5217 );
xor ( n10959 , n10958 , n5221 );
and ( n10960 , n10956 , n10959 );
and ( n10961 , n10954 , n10959 );
or ( n10962 , n10957 , n10960 , n10961 );
xor ( n10963 , n5151 , n5152 );
xor ( n10964 , n10963 , n5168 );
and ( n10965 , n10962 , n10964 );
xor ( n10966 , n5185 , n5193 );
xor ( n10967 , n10966 , n5201 );
and ( n10968 , n10964 , n10967 );
and ( n10969 , n10962 , n10967 );
or ( n10970 , n10965 , n10968 , n10969 );
and ( n10971 , n10951 , n10970 );
and ( n10972 , n10849 , n10970 );
or ( n10973 , n10952 , n10971 , n10972 );
and ( n10974 , n10798 , n10973 );
xor ( n10975 , n5052 , n5054 );
xor ( n10976 , n10975 , n5057 );
xor ( n10977 , n5072 , n5118 );
xor ( n10978 , n10977 , n5136 );
and ( n10979 , n10976 , n10978 );
xor ( n10980 , n5149 , n5171 );
xor ( n10981 , n10980 , n5204 );
and ( n10982 , n10978 , n10981 );
and ( n10983 , n10976 , n10981 );
or ( n10984 , n10979 , n10982 , n10983 );
and ( n10985 , n10973 , n10984 );
and ( n10986 , n10798 , n10984 );
or ( n10987 , n10974 , n10985 , n10986 );
xor ( n10988 , n5047 , n5049 );
xor ( n10989 , n10988 , n5060 );
xor ( n10990 , n5139 , n5207 );
xor ( n10991 , n10990 , n10658 );
and ( n10992 , n10989 , n10991 );
xor ( n10993 , n10671 , n10673 );
xor ( n10994 , n10993 , n10676 );
and ( n10995 , n10991 , n10994 );
and ( n10996 , n10989 , n10994 );
or ( n10997 , n10992 , n10995 , n10996 );
and ( n10998 , n10987 , n10997 );
xor ( n10999 , n5042 , n5044 );
xor ( n11000 , n10999 , n5063 );
and ( n11001 , n10997 , n11000 );
and ( n11002 , n10987 , n11000 );
or ( n11003 , n10998 , n11001 , n11002 );
and ( n11004 , n10747 , n11003 );
xor ( n11005 , n5037 , n5039 );
xor ( n11006 , n11005 , n5066 );
and ( n11007 , n11003 , n11006 );
and ( n11008 , n10747 , n11006 );
or ( n11009 , n11004 , n11007 , n11008 );
and ( n11010 , n10744 , n11009 );
and ( n11011 , n10742 , n11009 );
or ( n11012 , n10745 , n11010 , n11011 );
xor ( n11013 , n10712 , n10714 );
xor ( n11014 , n11013 , n10717 );
and ( n11015 , n11012 , n11014 );
xor ( n11016 , n5035 , n5069 );
xor ( n11017 , n11016 , n10709 );
xor ( n11018 , n10693 , n10703 );
xor ( n11019 , n11018 , n10706 );
xor ( n11020 , n10661 , n10679 );
xor ( n11021 , n11020 , n10690 );
xor ( n11022 , n10695 , n10697 );
xor ( n11023 , n11022 , n10700 );
and ( n11024 , n11021 , n11023 );
xor ( n11025 , n10682 , n10684 );
xor ( n11026 , n11025 , n10687 );
xor ( n11027 , n10642 , n10652 );
xor ( n11028 , n11027 , n10655 );
xor ( n11029 , n10663 , n10665 );
xor ( n11030 , n11029 , n10668 );
and ( n11031 , n11028 , n11030 );
xor ( n11032 , n5215 , n5224 );
xor ( n11033 , n11032 , n10639 );
xor ( n11034 , n10644 , n10646 );
xor ( n11035 , n11034 , n10649 );
and ( n11036 , n11033 , n11035 );
xor ( n11037 , n5228 , n10634 );
xor ( n11038 , n11037 , n10636 );
xor ( n11039 , n10772 , n10779 );
xor ( n11040 , n11039 , n10789 );
and ( n11041 , n11038 , n11040 );
xor ( n11042 , n10800 , n10802 );
and ( n11043 , n11040 , n11042 );
and ( n11044 , n11038 , n11042 );
or ( n11045 , n11041 , n11043 , n11044 );
and ( n11046 , n11035 , n11045 );
and ( n11047 , n11033 , n11045 );
or ( n11048 , n11036 , n11046 , n11047 );
and ( n11049 , n11030 , n11048 );
and ( n11050 , n11028 , n11048 );
or ( n11051 , n11031 , n11049 , n11050 );
and ( n11052 , n11026 , n11051 );
and ( n11053 , n1317 , n5086 );
and ( n11054 , n5091 , n1312 );
and ( n11055 , n11053 , n11054 );
and ( n11056 , n1911 , n3146 );
and ( n11057 , n3151 , n1906 );
and ( n11058 , n11056 , n11057 );
and ( n11059 , n11055 , n11058 );
and ( n11060 , n2764 , n4522 );
and ( n11061 , n11058 , n11060 );
and ( n11062 , n11055 , n11060 );
or ( n11063 , n11059 , n11061 , n11062 );
and ( n11064 , n2255 , n2586 );
and ( n11065 , n2591 , n2250 );
and ( n11066 , n11064 , n11065 );
and ( n11067 , n3339 , n2948 );
and ( n11068 , n11066 , n11067 );
and ( n11069 , n2634 , n5077 );
and ( n11070 , n11067 , n11069 );
and ( n11071 , n11066 , n11069 );
or ( n11072 , n11068 , n11070 , n11071 );
and ( n11073 , n11063 , n11072 );
and ( n11074 , n2309 , n2492 );
and ( n11075 , n2497 , n2304 );
and ( n11076 , n11074 , n11075 );
and ( n11077 , n4138 , n2040 );
and ( n11078 , n11076 , n11077 );
and ( n11079 , n3833 , n2407 );
and ( n11080 , n11077 , n11079 );
and ( n11081 , n11076 , n11079 );
or ( n11082 , n11078 , n11080 , n11081 );
and ( n11083 , n11072 , n11082 );
and ( n11084 , n11063 , n11082 );
or ( n11085 , n11073 , n11083 , n11084 );
xor ( n11086 , n10766 , n10767 );
xor ( n11087 , n11086 , n10769 );
xor ( n11088 , n10816 , n10817 );
xor ( n11089 , n11088 , n10819 );
and ( n11090 , n11087 , n11089 );
xor ( n11091 , n10825 , n10826 );
xor ( n11092 , n11091 , n10828 );
and ( n11093 , n11089 , n11092 );
and ( n11094 , n11087 , n11092 );
or ( n11095 , n11090 , n11093 , n11094 );
and ( n11096 , n11085 , n11095 );
xor ( n11097 , n10773 , n10774 );
xor ( n11098 , n11097 , n10776 );
xor ( n11099 , n10783 , n10784 );
xor ( n11100 , n11099 , n10786 );
and ( n11101 , n11098 , n11100 );
xor ( n11102 , n10835 , n10838 );
xor ( n11103 , n11102 , n10840 );
and ( n11104 , n11100 , n11103 );
and ( n11105 , n11098 , n11103 );
or ( n11106 , n11101 , n11104 , n11105 );
and ( n11107 , n11095 , n11106 );
and ( n11108 , n11085 , n11106 );
or ( n11109 , n11096 , n11107 , n11108 );
buf ( n11110 , n5338 );
buf ( n11111 , n11110 );
and ( n11112 , n1291 , n11111 );
not ( n11113 , n11111 );
nor ( n11114 , n11112 , n11113 );
buf ( n11115 , n5338 );
buf ( n11116 , n11115 );
not ( n11117 , n11116 );
and ( n11118 , n1279 , n11116 );
nor ( n11119 , n11117 , n11118 );
and ( n11120 , n11114 , n11119 );
and ( n11121 , n1724 , n3449 );
and ( n11122 , n3454 , n1719 );
and ( n11123 , n11121 , n11122 );
and ( n11124 , n11120 , n11123 );
and ( n11125 , n4579 , n1711 );
and ( n11126 , n11123 , n11125 );
and ( n11127 , n11120 , n11125 );
or ( n11128 , n11124 , n11126 , n11127 );
and ( n11129 , n1353 , n4982 );
and ( n11130 , n4989 , n1348 );
and ( n11131 , n11129 , n11130 );
and ( n11132 , n3645 , n2577 );
and ( n11133 , n11131 , n11132 );
and ( n11134 , n2937 , n3929 );
and ( n11135 , n11132 , n11134 );
and ( n11136 , n11131 , n11134 );
or ( n11137 , n11133 , n11135 , n11136 );
and ( n11138 , n11128 , n11137 );
xor ( n11139 , n5229 , n5230 );
xor ( n11140 , n11139 , n10631 );
xor ( n11141 , n10852 , n10855 );
xor ( n11142 , n11141 , n10857 );
and ( n11143 , n11140 , n11142 );
xor ( n11144 , n10867 , n10874 );
and ( n11145 , n11142 , n11144 );
and ( n11146 , n11140 , n11144 );
or ( n11147 , n11143 , n11145 , n11146 );
and ( n11148 , n11138 , n11147 );
xor ( n11149 , n10878 , n10880 );
and ( n11150 , n1778 , n3288 );
and ( n11151 , n3293 , n1789 );
and ( n11152 , n11150 , n11151 );
and ( n11153 , n4385 , n1860 );
and ( n11154 , n11152 , n11153 );
buf ( n11155 , n2284 );
buf ( n11156 , n11155 );
and ( n11157 , n2477 , n11156 );
and ( n11158 , n11153 , n11157 );
and ( n11159 , n11152 , n11157 );
or ( n11160 , n11154 , n11158 , n11159 );
and ( n11161 , n11149 , n11160 );
and ( n11162 , n1275 , n10869 );
and ( n11163 , n10862 , n1293 );
and ( n11164 , n11162 , n11163 );
and ( n11165 , n5177 , n1465 );
and ( n11166 , n11164 , n11165 );
and ( n11167 , n4721 , n1530 );
and ( n11168 , n11165 , n11167 );
and ( n11169 , n11164 , n11167 );
or ( n11170 , n11166 , n11168 , n11169 );
and ( n11171 , n11160 , n11170 );
and ( n11172 , n11149 , n11170 );
or ( n11173 , n11161 , n11171 , n11172 );
and ( n11174 , n11147 , n11173 );
and ( n11175 , n11138 , n11173 );
or ( n11176 , n11148 , n11174 , n11175 );
and ( n11177 , n11109 , n11176 );
and ( n11178 , n1995 , n2923 );
and ( n11179 , n2928 , n1990 );
and ( n11180 , n11178 , n11179 );
buf ( n11181 , n2286 );
and ( n11182 , n11180 , n11181 );
and ( n11183 , n3728 , n1689 );
and ( n11184 , n2723 , n2059 );
and ( n11185 , n11183 , n11184 );
and ( n11186 , n1694 , n3739 );
and ( n11187 , n2048 , n2718 );
and ( n11188 , n11186 , n11187 );
and ( n11189 , n11185 , n11188 );
and ( n11190 , n11182 , n11189 );
xor ( n11191 , n10865 , n10866 );
xor ( n11192 , n10872 , n10873 );
and ( n11193 , n11191 , n11192 );
and ( n11194 , n11189 , n11193 );
and ( n11195 , n11182 , n11193 );
or ( n11196 , n11190 , n11194 , n11195 );
xnor ( n11197 , n10925 , n10926 );
xor ( n11198 , n10850 , n10851 );
and ( n11199 , n11197 , n11198 );
xor ( n11200 , n10814 , n10815 );
and ( n11201 , n11198 , n11200 );
and ( n11202 , n11197 , n11200 );
or ( n11203 , n11199 , n11201 , n11202 );
xor ( n11204 , n10833 , n10834 );
xor ( n11205 , n10853 , n10854 );
and ( n11206 , n11204 , n11205 );
xor ( n11207 , n10781 , n10782 );
and ( n11208 , n11205 , n11207 );
and ( n11209 , n11204 , n11207 );
or ( n11210 , n11206 , n11208 , n11209 );
and ( n11211 , n11203 , n11210 );
xor ( n11212 , n10823 , n10824 );
xor ( n11213 , n10836 , n10837 );
and ( n11214 , n11212 , n11213 );
xor ( n11215 , n10929 , n10930 );
xor ( n11216 , n11215 , n10934 );
and ( n11217 , n11213 , n11216 );
and ( n11218 , n11212 , n11216 );
or ( n11219 , n11214 , n11217 , n11218 );
and ( n11220 , n11210 , n11219 );
and ( n11221 , n11203 , n11219 );
or ( n11222 , n11211 , n11220 , n11221 );
and ( n11223 , n11196 , n11222 );
xor ( n11224 , n10887 , n10888 );
xor ( n11225 , n11224 , n10890 );
xor ( n11226 , n10894 , n10895 );
xor ( n11227 , n11226 , n10897 );
and ( n11228 , n11225 , n11227 );
xor ( n11229 , n10902 , n10903 );
xor ( n11230 , n11229 , n10911 );
and ( n11231 , n11227 , n11230 );
and ( n11232 , n11225 , n11230 );
or ( n11233 , n11228 , n11231 , n11232 );
and ( n11234 , n11222 , n11233 );
and ( n11235 , n11196 , n11233 );
or ( n11236 , n11223 , n11234 , n11235 );
and ( n11237 , n11176 , n11236 );
and ( n11238 , n11109 , n11236 );
or ( n11239 , n11177 , n11237 , n11238 );
xor ( n11240 , n10805 , n10807 );
xor ( n11241 , n11240 , n10809 );
xor ( n11242 , n10822 , n10831 );
xor ( n11243 , n11242 , n10843 );
and ( n11244 , n11241 , n11243 );
xor ( n11245 , n10860 , n10875 );
xor ( n11246 , n11245 , n10881 );
and ( n11247 , n11243 , n11246 );
and ( n11248 , n11241 , n11246 );
or ( n11249 , n11244 , n11247 , n11248 );
xor ( n11250 , n10893 , n10900 );
xor ( n11251 , n11250 , n10914 );
xor ( n11252 , n10940 , n10942 );
xor ( n11253 , n11252 , n10945 );
and ( n11254 , n11251 , n11253 );
xor ( n11255 , n10954 , n10956 );
xor ( n11256 , n11255 , n10959 );
and ( n11257 , n11253 , n11256 );
and ( n11258 , n11251 , n11256 );
or ( n11259 , n11254 , n11257 , n11258 );
and ( n11260 , n11249 , n11259 );
xor ( n11261 , n10751 , n10753 );
xor ( n11262 , n11261 , n10756 );
and ( n11263 , n11259 , n11262 );
and ( n11264 , n11249 , n11262 );
or ( n11265 , n11260 , n11263 , n11264 );
and ( n11266 , n11239 , n11265 );
xor ( n11267 , n10762 , n10764 );
xor ( n11268 , n11267 , n10792 );
xor ( n11269 , n10803 , n10812 );
xor ( n11270 , n11269 , n10846 );
and ( n11271 , n11268 , n11270 );
xor ( n11272 , n10884 , n10917 );
xor ( n11273 , n11272 , n10948 );
and ( n11274 , n11270 , n11273 );
and ( n11275 , n11268 , n11273 );
or ( n11276 , n11271 , n11274 , n11275 );
and ( n11277 , n11265 , n11276 );
and ( n11278 , n11239 , n11276 );
or ( n11279 , n11266 , n11277 , n11278 );
and ( n11280 , n11051 , n11279 );
and ( n11281 , n11026 , n11279 );
or ( n11282 , n11052 , n11280 , n11281 );
and ( n11283 , n11023 , n11282 );
and ( n11284 , n11021 , n11282 );
or ( n11285 , n11024 , n11283 , n11284 );
and ( n11286 , n11019 , n11285 );
xor ( n11287 , n10747 , n11003 );
xor ( n11288 , n11287 , n11006 );
and ( n11289 , n11285 , n11288 );
and ( n11290 , n11019 , n11288 );
or ( n11291 , n11286 , n11289 , n11290 );
and ( n11292 , n11017 , n11291 );
xor ( n11293 , n10742 , n10744 );
xor ( n11294 , n11293 , n11009 );
and ( n11295 , n11291 , n11294 );
and ( n11296 , n11017 , n11294 );
or ( n11297 , n11292 , n11295 , n11296 );
and ( n11298 , n11014 , n11297 );
and ( n11299 , n11012 , n11297 );
or ( n11300 , n11015 , n11298 , n11299 );
and ( n11301 , n10739 , n11300 );
and ( n11302 , n10737 , n11300 );
or ( n11303 , n10740 , n11301 , n11302 );
and ( n11304 , n10735 , n11303 );
xor ( n11305 , n10735 , n11303 );
xor ( n11306 , n10737 , n10739 );
xor ( n11307 , n11306 , n11300 );
xor ( n11308 , n11012 , n11014 );
xor ( n11309 , n11308 , n11297 );
xor ( n11310 , n11017 , n11291 );
xor ( n11311 , n11310 , n11294 );
xor ( n11312 , n10749 , n10759 );
xor ( n11313 , n11312 , n10795 );
xor ( n11314 , n10849 , n10951 );
xor ( n11315 , n11314 , n10970 );
and ( n11316 , n11313 , n11315 );
xor ( n11317 , n10976 , n10978 );
xor ( n11318 , n11317 , n10981 );
and ( n11319 , n11315 , n11318 );
and ( n11320 , n11313 , n11318 );
or ( n11321 , n11316 , n11319 , n11320 );
xor ( n11322 , n10798 , n10973 );
xor ( n11323 , n11322 , n10984 );
and ( n11324 , n11321 , n11323 );
xor ( n11325 , n10989 , n10991 );
xor ( n11326 , n11325 , n10994 );
and ( n11327 , n11323 , n11326 );
and ( n11328 , n11321 , n11326 );
or ( n11329 , n11324 , n11327 , n11328 );
xor ( n11330 , n10987 , n10997 );
xor ( n11331 , n11330 , n11000 );
and ( n11332 , n11329 , n11331 );
xor ( n11333 , n10962 , n10964 );
xor ( n11334 , n11333 , n10967 );
and ( n11335 , n1995 , n3146 );
and ( n11336 , n3151 , n1990 );
and ( n11337 , n11335 , n11336 );
and ( n11338 , n4721 , n1711 );
and ( n11339 , n11337 , n11338 );
and ( n11340 , n3246 , n3627 );
and ( n11341 , n11338 , n11340 );
and ( n11342 , n11337 , n11340 );
or ( n11343 , n11339 , n11341 , n11342 );
and ( n11344 , n5177 , n1530 );
and ( n11345 , n3339 , n3301 );
and ( n11346 , n11344 , n11345 );
and ( n11347 , n2937 , n4522 );
and ( n11348 , n11345 , n11347 );
and ( n11349 , n11344 , n11347 );
or ( n11350 , n11346 , n11348 , n11349 );
and ( n11351 , n11343 , n11350 );
and ( n11352 , n2048 , n2923 );
and ( n11353 , n2928 , n2059 );
and ( n11354 , n11352 , n11353 );
and ( n11355 , n3645 , n2948 );
and ( n11356 , n11354 , n11355 );
and ( n11357 , n3169 , n3929 );
and ( n11358 , n11355 , n11357 );
and ( n11359 , n11354 , n11357 );
or ( n11360 , n11356 , n11358 , n11359 );
and ( n11361 , n11350 , n11360 );
and ( n11362 , n11343 , n11360 );
or ( n11363 , n11351 , n11361 , n11362 );
xor ( n11364 , n10919 , n10923 );
and ( n11365 , n1724 , n3739 );
and ( n11366 , n3728 , n1719 );
and ( n11367 , n11365 , n11366 );
and ( n11368 , n2255 , n2718 );
and ( n11369 , n2723 , n2250 );
and ( n11370 , n11368 , n11369 );
and ( n11371 , n11367 , n11370 );
and ( n11372 , n2764 , n5077 );
and ( n11373 , n11370 , n11372 );
and ( n11374 , n11367 , n11372 );
or ( n11375 , n11371 , n11373 , n11374 );
and ( n11376 , n11364 , n11375 );
xor ( n11377 , n8860 , n10624 );
buf ( n11378 , n11377 );
buf ( n11379 , n11378 );
buf ( n11380 , n11379 );
buf ( n11381 , n11380 );
and ( n11382 , n11375 , n11381 );
and ( n11383 , n11364 , n11381 );
or ( n11384 , n11376 , n11382 , n11383 );
and ( n11385 , n11363 , n11384 );
and ( n11386 , n1275 , n11111 );
and ( n11387 , n11116 , n1293 );
and ( n11388 , n11386 , n11387 );
not ( n11389 , n11380 );
and ( n11390 , n11388 , n11389 );
and ( n11391 , n4385 , n2040 );
and ( n11392 , n11389 , n11391 );
and ( n11393 , n11388 , n11391 );
or ( n11394 , n11390 , n11392 , n11393 );
xor ( n11395 , n11120 , n11123 );
xor ( n11396 , n11395 , n11125 );
and ( n11397 , n11394 , n11396 );
xor ( n11398 , n11066 , n11067 );
xor ( n11399 , n11398 , n11069 );
and ( n11400 , n11396 , n11399 );
and ( n11401 , n11394 , n11399 );
or ( n11402 , n11397 , n11400 , n11401 );
and ( n11403 , n11384 , n11402 );
and ( n11404 , n11363 , n11402 );
or ( n11405 , n11385 , n11403 , n11404 );
xor ( n11406 , n10924 , n10927 );
xor ( n11407 , n11406 , n10937 );
xor ( n11408 , n11063 , n11072 );
xor ( n11409 , n11408 , n11082 );
and ( n11410 , n11407 , n11409 );
xor ( n11411 , n11087 , n11089 );
xor ( n11412 , n11411 , n11092 );
and ( n11413 , n11409 , n11412 );
and ( n11414 , n11407 , n11412 );
or ( n11415 , n11410 , n11413 , n11414 );
and ( n11416 , n11405 , n11415 );
xor ( n11417 , n11098 , n11100 );
xor ( n11418 , n11417 , n11103 );
xor ( n11419 , n11128 , n11137 );
and ( n11420 , n11418 , n11419 );
xor ( n11421 , n11152 , n11153 );
xor ( n11422 , n11421 , n11157 );
xor ( n11423 , n11055 , n11058 );
xor ( n11424 , n11423 , n11060 );
and ( n11425 , n11422 , n11424 );
xor ( n11426 , n10905 , n10906 );
xor ( n11427 , n11426 , n10908 );
and ( n11428 , n11424 , n11427 );
and ( n11429 , n11422 , n11427 );
or ( n11430 , n11425 , n11428 , n11429 );
and ( n11431 , n11419 , n11430 );
and ( n11432 , n11418 , n11430 );
or ( n11433 , n11420 , n11431 , n11432 );
and ( n11434 , n11415 , n11433 );
and ( n11435 , n11405 , n11433 );
or ( n11436 , n11416 , n11434 , n11435 );
and ( n11437 , n11334 , n11436 );
xor ( n11438 , n11164 , n11165 );
xor ( n11439 , n11438 , n11167 );
xor ( n11440 , n11076 , n11077 );
xor ( n11441 , n11440 , n11079 );
and ( n11442 , n11439 , n11441 );
xor ( n11443 , n11131 , n11132 );
xor ( n11444 , n11443 , n11134 );
and ( n11445 , n11441 , n11444 );
and ( n11446 , n11439 , n11444 );
or ( n11447 , n11442 , n11445 , n11446 );
and ( n11448 , n10886 , n1465 );
and ( n11449 , n4579 , n1860 );
and ( n11450 , n11448 , n11449 );
and ( n11451 , n2634 , n11156 );
and ( n11452 , n11449 , n11451 );
and ( n11453 , n11448 , n11451 );
or ( n11454 , n11450 , n11452 , n11453 );
xor ( n11455 , n11180 , n11181 );
and ( n11456 , n11454 , n11455 );
and ( n11457 , n11447 , n11456 );
xor ( n11458 , n11185 , n11188 );
xor ( n11459 , n11191 , n11192 );
and ( n11460 , n11458 , n11459 );
and ( n11461 , n1694 , n3903 );
and ( n11462 , n3892 , n1689 );
and ( n11463 , n11461 , n11462 );
and ( n11464 , n1778 , n3449 );
and ( n11465 , n3454 , n1789 );
and ( n11466 , n11464 , n11465 );
and ( n11467 , n11463 , n11466 );
and ( n11468 , n4138 , n2407 );
and ( n11469 , n11466 , n11468 );
and ( n11470 , n11463 , n11468 );
or ( n11471 , n11467 , n11469 , n11470 );
and ( n11472 , n11459 , n11471 );
and ( n11473 , n11458 , n11471 );
or ( n11474 , n11460 , n11472 , n11473 );
and ( n11475 , n11456 , n11474 );
and ( n11476 , n11447 , n11474 );
or ( n11477 , n11457 , n11475 , n11476 );
and ( n11478 , n1317 , n10869 );
and ( n11479 , n10862 , n1312 );
and ( n11480 , n11478 , n11479 );
and ( n11481 , n1353 , n5086 );
and ( n11482 , n5091 , n1348 );
and ( n11483 , n11481 , n11482 );
and ( n11484 , n11480 , n11483 );
and ( n11485 , n10933 , n1360 );
and ( n11486 , n11483 , n11485 );
and ( n11487 , n11480 , n11485 );
or ( n11488 , n11484 , n11486 , n11487 );
xor ( n11489 , n11183 , n11184 );
xor ( n11490 , n11186 , n11187 );
and ( n11491 , n11489 , n11490 );
and ( n11492 , n11488 , n11491 );
and ( n11493 , n3833 , n2577 );
xor ( n11494 , n11344 , n11345 );
xor ( n11495 , n11494 , n11347 );
and ( n11496 , n11493 , n11495 );
xor ( n11497 , n11114 , n11119 );
and ( n11498 , n11495 , n11497 );
and ( n11499 , n11493 , n11497 );
or ( n11500 , n11496 , n11498 , n11499 );
and ( n11501 , n11491 , n11500 );
and ( n11502 , n11488 , n11500 );
or ( n11503 , n11492 , n11501 , n11502 );
xor ( n11504 , n11162 , n11163 );
xor ( n11505 , n11053 , n11054 );
and ( n11506 , n11504 , n11505 );
xor ( n11507 , n11129 , n11130 );
and ( n11508 , n11505 , n11507 );
and ( n11509 , n11504 , n11507 );
or ( n11510 , n11506 , n11508 , n11509 );
xor ( n11511 , n11121 , n11122 );
xor ( n11512 , n11150 , n11151 );
and ( n11513 , n11511 , n11512 );
xor ( n11514 , n11056 , n11057 );
and ( n11515 , n11512 , n11514 );
and ( n11516 , n11511 , n11514 );
or ( n11517 , n11513 , n11515 , n11516 );
and ( n11518 , n11510 , n11517 );
xor ( n11519 , n11178 , n11179 );
xor ( n11520 , n11064 , n11065 );
and ( n11521 , n11519 , n11520 );
xor ( n11522 , n11074 , n11075 );
and ( n11523 , n11520 , n11522 );
and ( n11524 , n11519 , n11522 );
or ( n11525 , n11521 , n11523 , n11524 );
and ( n11526 , n11517 , n11525 );
and ( n11527 , n11510 , n11525 );
or ( n11528 , n11518 , n11526 , n11527 );
and ( n11529 , n11503 , n11528 );
xor ( n11530 , n11197 , n11198 );
xor ( n11531 , n11530 , n11200 );
xor ( n11532 , n11204 , n11205 );
xor ( n11533 , n11532 , n11207 );
and ( n11534 , n11531 , n11533 );
xor ( n11535 , n11212 , n11213 );
xor ( n11536 , n11535 , n11216 );
and ( n11537 , n11533 , n11536 );
and ( n11538 , n11531 , n11536 );
or ( n11539 , n11534 , n11537 , n11538 );
and ( n11540 , n11528 , n11539 );
and ( n11541 , n11503 , n11539 );
or ( n11542 , n11529 , n11540 , n11541 );
and ( n11543 , n11477 , n11542 );
xor ( n11544 , n11140 , n11142 );
xor ( n11545 , n11544 , n11144 );
xor ( n11546 , n11149 , n11160 );
xor ( n11547 , n11546 , n11170 );
and ( n11548 , n11545 , n11547 );
xor ( n11549 , n11182 , n11189 );
xor ( n11550 , n11549 , n11193 );
and ( n11551 , n11547 , n11550 );
and ( n11552 , n11545 , n11550 );
or ( n11553 , n11548 , n11551 , n11552 );
and ( n11554 , n11542 , n11553 );
and ( n11555 , n11477 , n11553 );
or ( n11556 , n11543 , n11554 , n11555 );
and ( n11557 , n11436 , n11556 );
and ( n11558 , n11334 , n11556 );
or ( n11559 , n11437 , n11557 , n11558 );
xor ( n11560 , n11038 , n11040 );
xor ( n11561 , n11560 , n11042 );
xor ( n11562 , n11085 , n11095 );
xor ( n11563 , n11562 , n11106 );
and ( n11564 , n11561 , n11563 );
xor ( n11565 , n11138 , n11147 );
xor ( n11566 , n11565 , n11173 );
and ( n11567 , n11563 , n11566 );
and ( n11568 , n11561 , n11566 );
or ( n11569 , n11564 , n11567 , n11568 );
xor ( n11570 , n11196 , n11222 );
xor ( n11571 , n11570 , n11233 );
xor ( n11572 , n11241 , n11243 );
xor ( n11573 , n11572 , n11246 );
and ( n11574 , n11571 , n11573 );
xor ( n11575 , n11251 , n11253 );
xor ( n11576 , n11575 , n11256 );
and ( n11577 , n11573 , n11576 );
and ( n11578 , n11571 , n11576 );
or ( n11579 , n11574 , n11577 , n11578 );
and ( n11580 , n11569 , n11579 );
xor ( n11581 , n11033 , n11035 );
xor ( n11582 , n11581 , n11045 );
and ( n11583 , n11579 , n11582 );
and ( n11584 , n11569 , n11582 );
or ( n11585 , n11580 , n11583 , n11584 );
and ( n11586 , n11559 , n11585 );
xor ( n11587 , n11109 , n11176 );
xor ( n11588 , n11587 , n11236 );
xor ( n11589 , n11249 , n11259 );
xor ( n11590 , n11589 , n11262 );
and ( n11591 , n11588 , n11590 );
xor ( n11592 , n11268 , n11270 );
xor ( n11593 , n11592 , n11273 );
and ( n11594 , n11590 , n11593 );
and ( n11595 , n11588 , n11593 );
or ( n11596 , n11591 , n11594 , n11595 );
and ( n11597 , n11585 , n11596 );
and ( n11598 , n11559 , n11596 );
or ( n11599 , n11586 , n11597 , n11598 );
xor ( n11600 , n11028 , n11030 );
xor ( n11601 , n11600 , n11048 );
xor ( n11602 , n11239 , n11265 );
xor ( n11603 , n11602 , n11276 );
and ( n11604 , n11601 , n11603 );
xor ( n11605 , n11313 , n11315 );
xor ( n11606 , n11605 , n11318 );
and ( n11607 , n11603 , n11606 );
and ( n11608 , n11601 , n11606 );
or ( n11609 , n11604 , n11607 , n11608 );
and ( n11610 , n11599 , n11609 );
xor ( n11611 , n11026 , n11051 );
xor ( n11612 , n11611 , n11279 );
and ( n11613 , n11609 , n11612 );
and ( n11614 , n11599 , n11612 );
or ( n11615 , n11610 , n11613 , n11614 );
and ( n11616 , n11331 , n11615 );
and ( n11617 , n11329 , n11615 );
or ( n11618 , n11332 , n11616 , n11617 );
xor ( n11619 , n11019 , n11285 );
xor ( n11620 , n11619 , n11288 );
and ( n11621 , n11618 , n11620 );
xor ( n11622 , n11021 , n11023 );
xor ( n11623 , n11622 , n11282 );
xor ( n11624 , n11321 , n11323 );
xor ( n11625 , n11624 , n11326 );
xor ( n11626 , n11203 , n11210 );
xor ( n11627 , n11626 , n11219 );
xor ( n11628 , n11225 , n11227 );
xor ( n11629 , n11628 , n11230 );
and ( n11630 , n11627 , n11629 );
xor ( n11631 , n11363 , n11384 );
xor ( n11632 , n11631 , n11402 );
and ( n11633 , n11629 , n11632 );
and ( n11634 , n11627 , n11632 );
or ( n11635 , n11630 , n11633 , n11634 );
xor ( n11636 , n11343 , n11350 );
xor ( n11637 , n11636 , n11360 );
xor ( n11638 , n11364 , n11375 );
xor ( n11639 , n11638 , n11381 );
and ( n11640 , n11637 , n11639 );
xor ( n11641 , n11422 , n11424 );
xor ( n11642 , n11641 , n11427 );
and ( n11643 , n11639 , n11642 );
and ( n11644 , n11637 , n11642 );
or ( n11645 , n11640 , n11643 , n11644 );
xor ( n11646 , n11439 , n11441 );
xor ( n11647 , n11646 , n11444 );
xor ( n11648 , n11394 , n11396 );
xor ( n11649 , n11648 , n11399 );
and ( n11650 , n11647 , n11649 );
xor ( n11651 , n11454 , n11455 );
and ( n11652 , n11649 , n11651 );
and ( n11653 , n11647 , n11651 );
or ( n11654 , n11650 , n11652 , n11653 );
and ( n11655 , n11645 , n11654 );
and ( n11656 , n10886 , n1530 );
and ( n11657 , n3645 , n3301 );
and ( n11658 , n11656 , n11657 );
and ( n11659 , n3169 , n4522 );
and ( n11660 , n11657 , n11659 );
and ( n11661 , n11656 , n11659 );
or ( n11662 , n11658 , n11660 , n11661 );
and ( n11663 , n1353 , n10869 );
and ( n11664 , n10862 , n1348 );
and ( n11665 , n11663 , n11664 );
and ( n11666 , n2048 , n3146 );
and ( n11667 , n3151 , n2059 );
and ( n11668 , n11666 , n11667 );
and ( n11669 , n11665 , n11668 );
and ( n11670 , n2937 , n5077 );
and ( n11671 , n11668 , n11670 );
and ( n11672 , n11665 , n11670 );
or ( n11673 , n11669 , n11671 , n11672 );
and ( n11674 , n11662 , n11673 );
and ( n11675 , n2255 , n2923 );
and ( n11676 , n2928 , n2250 );
and ( n11677 , n11675 , n11676 );
and ( n11678 , n5177 , n1711 );
and ( n11679 , n11677 , n11678 );
and ( n11680 , n3246 , n3929 );
and ( n11681 , n11678 , n11680 );
and ( n11682 , n11677 , n11680 );
or ( n11683 , n11679 , n11681 , n11682 );
and ( n11684 , n11673 , n11683 );
and ( n11685 , n11662 , n11683 );
or ( n11686 , n11674 , n11684 , n11685 );
and ( n11687 , n2497 , n2586 );
and ( n11688 , n2591 , n2492 );
and ( n11689 , n11687 , n11688 );
and ( n11690 , n10933 , n1465 );
and ( n11691 , n11689 , n11690 );
and ( n11692 , n4385 , n2407 );
and ( n11693 , n11690 , n11692 );
and ( n11694 , n11689 , n11692 );
or ( n11695 , n11691 , n11693 , n11694 );
and ( n11696 , n1995 , n3288 );
and ( n11697 , n3293 , n1990 );
and ( n11698 , n11696 , n11697 );
and ( n11699 , n4138 , n2577 );
and ( n11700 , n11698 , n11699 );
and ( n11701 , n3339 , n3627 );
and ( n11702 , n11699 , n11701 );
and ( n11703 , n11698 , n11701 );
or ( n11704 , n11700 , n11702 , n11703 );
and ( n11705 , n11695 , n11704 );
buf ( n11706 , n2497 );
xor ( n11707 , n9324 , n10622 );
buf ( n11708 , n11707 );
buf ( n11709 , n11708 );
buf ( n11710 , n11709 );
and ( n11711 , n11706 , n11710 );
and ( n11712 , n11704 , n11711 );
and ( n11713 , n11695 , n11711 );
or ( n11714 , n11705 , n11712 , n11713 );
and ( n11715 , n11686 , n11714 );
xor ( n11716 , n11367 , n11370 );
xor ( n11717 , n11716 , n11372 );
xor ( n11718 , n11463 , n11466 );
xor ( n11719 , n11718 , n11468 );
and ( n11720 , n11717 , n11719 );
xor ( n11721 , n11354 , n11355 );
xor ( n11722 , n11721 , n11357 );
and ( n11723 , n11719 , n11722 );
and ( n11724 , n11717 , n11722 );
or ( n11725 , n11720 , n11723 , n11724 );
and ( n11726 , n11714 , n11725 );
and ( n11727 , n11686 , n11725 );
or ( n11728 , n11715 , n11726 , n11727 );
and ( n11729 , n11654 , n11728 );
and ( n11730 , n11645 , n11728 );
or ( n11731 , n11655 , n11729 , n11730 );
and ( n11732 , n11635 , n11731 );
and ( n11733 , n1911 , n3288 );
and ( n11734 , n2309 , n2586 );
or ( n11735 , n11733 , n11734 );
and ( n11736 , n3293 , n1906 );
and ( n11737 , n2591 , n2304 );
and ( n11738 , n11736 , n11737 );
and ( n11739 , n4721 , n1860 );
and ( n11740 , n11737 , n11739 );
and ( n11741 , n11736 , n11739 );
or ( n11742 , n11738 , n11740 , n11741 );
and ( n11743 , n11735 , n11742 );
xor ( n11744 , n11337 , n11338 );
xor ( n11745 , n11744 , n11340 );
and ( n11746 , n11742 , n11745 );
and ( n11747 , n11735 , n11745 );
or ( n11748 , n11743 , n11746 , n11747 );
xor ( n11749 , n11480 , n11483 );
xor ( n11750 , n11749 , n11485 );
xor ( n11751 , n11388 , n11389 );
xor ( n11752 , n11751 , n11391 );
and ( n11753 , n11750 , n11752 );
xor ( n11754 , n11489 , n11490 );
and ( n11755 , n11752 , n11754 );
and ( n11756 , n11750 , n11754 );
or ( n11757 , n11753 , n11755 , n11756 );
and ( n11758 , n11748 , n11757 );
and ( n11759 , n1724 , n3903 );
and ( n11760 , n3892 , n1719 );
and ( n11761 , n11759 , n11760 );
and ( n11762 , n3833 , n2948 );
and ( n11763 , n11761 , n11762 );
and ( n11764 , n2764 , n11156 );
and ( n11765 , n11762 , n11764 );
and ( n11766 , n11761 , n11764 );
or ( n11767 , n11763 , n11765 , n11766 );
and ( n11768 , n4150 , n1689 );
and ( n11769 , n3454 , n1906 );
and ( n11770 , n11768 , n11769 );
and ( n11771 , n1694 , n4161 );
and ( n11772 , n1911 , n3449 );
and ( n11773 , n11771 , n11772 );
and ( n11774 , n11770 , n11773 );
and ( n11775 , n11767 , n11774 );
buf ( n11776 , n2475 );
buf ( n11777 , n11776 );
and ( n11778 , n2634 , n11777 );
buf ( n11779 , n2477 );
and ( n11780 , n11778 , n11779 );
xor ( n11781 , n11656 , n11657 );
xor ( n11782 , n11781 , n11659 );
and ( n11783 , n11779 , n11782 );
and ( n11784 , n11778 , n11782 );
or ( n11785 , n11780 , n11783 , n11784 );
and ( n11786 , n11774 , n11785 );
and ( n11787 , n11767 , n11785 );
or ( n11788 , n11775 , n11786 , n11787 );
and ( n11789 , n11757 , n11788 );
and ( n11790 , n11748 , n11788 );
or ( n11791 , n11758 , n11789 , n11790 );
xnor ( n11792 , n11733 , n11734 );
xor ( n11793 , n11706 , n11710 );
and ( n11794 , n11792 , n11793 );
xor ( n11795 , n11386 , n11387 );
and ( n11796 , n11793 , n11795 );
and ( n11797 , n11792 , n11795 );
or ( n11798 , n11794 , n11796 , n11797 );
xor ( n11799 , n11478 , n11479 );
xor ( n11800 , n11481 , n11482 );
and ( n11801 , n11799 , n11800 );
xor ( n11802 , n11461 , n11462 );
and ( n11803 , n11800 , n11802 );
and ( n11804 , n11799 , n11802 );
or ( n11805 , n11801 , n11803 , n11804 );
and ( n11806 , n11798 , n11805 );
xor ( n11807 , n11365 , n11366 );
xor ( n11808 , n11464 , n11465 );
and ( n11809 , n11807 , n11808 );
xor ( n11810 , n11335 , n11336 );
and ( n11811 , n11808 , n11810 );
and ( n11812 , n11807 , n11810 );
or ( n11813 , n11809 , n11811 , n11812 );
and ( n11814 , n11805 , n11813 );
and ( n11815 , n11798 , n11813 );
or ( n11816 , n11806 , n11814 , n11815 );
xor ( n11817 , n11352 , n11353 );
xor ( n11818 , n11368 , n11369 );
and ( n11819 , n11817 , n11818 );
and ( n11820 , n4721 , n2040 );
and ( n11821 , n3833 , n3301 );
and ( n11822 , n11820 , n11821 );
and ( n11823 , n2937 , n11156 );
and ( n11824 , n11821 , n11823 );
and ( n11825 , n11820 , n11823 );
or ( n11826 , n11822 , n11824 , n11825 );
and ( n11827 , n11818 , n11826 );
and ( n11828 , n11817 , n11826 );
or ( n11829 , n11819 , n11827 , n11828 );
and ( n11830 , n1317 , n11111 );
and ( n11831 , n2309 , n2718 );
or ( n11832 , n11830 , n11831 );
and ( n11833 , n1778 , n3739 );
xor ( n11834 , n9325 , n10621 );
buf ( n11835 , n11834 );
buf ( n11836 , n11835 );
buf ( n11837 , n11836 );
and ( n11838 , n11833 , n11837 );
and ( n11839 , n11832 , n11838 );
and ( n11840 , n11116 , n1312 );
and ( n11841 , n3728 , n1789 );
and ( n11842 , n11840 , n11841 );
and ( n11843 , n2723 , n2304 );
and ( n11844 , n11841 , n11843 );
and ( n11845 , n11840 , n11843 );
or ( n11846 , n11842 , n11844 , n11845 );
and ( n11847 , n11838 , n11846 );
and ( n11848 , n11832 , n11846 );
or ( n11849 , n11839 , n11847 , n11848 );
and ( n11850 , n11829 , n11849 );
xor ( n11851 , n11493 , n11495 );
xor ( n11852 , n11851 , n11497 );
and ( n11853 , n11849 , n11852 );
and ( n11854 , n11829 , n11852 );
or ( n11855 , n11850 , n11853 , n11854 );
and ( n11856 , n11816 , n11855 );
xor ( n11857 , n11504 , n11505 );
xor ( n11858 , n11857 , n11507 );
xor ( n11859 , n11511 , n11512 );
xor ( n11860 , n11859 , n11514 );
and ( n11861 , n11858 , n11860 );
xor ( n11862 , n11519 , n11520 );
xor ( n11863 , n11862 , n11522 );
and ( n11864 , n11860 , n11863 );
and ( n11865 , n11858 , n11863 );
or ( n11866 , n11861 , n11864 , n11865 );
and ( n11867 , n11855 , n11866 );
and ( n11868 , n11816 , n11866 );
or ( n11869 , n11856 , n11867 , n11868 );
and ( n11870 , n11791 , n11869 );
xor ( n11871 , n11458 , n11459 );
xor ( n11872 , n11871 , n11471 );
xor ( n11873 , n11488 , n11491 );
xor ( n11874 , n11873 , n11500 );
and ( n11875 , n11872 , n11874 );
xor ( n11876 , n11510 , n11517 );
xor ( n11877 , n11876 , n11525 );
and ( n11878 , n11874 , n11877 );
and ( n11879 , n11872 , n11877 );
or ( n11880 , n11875 , n11878 , n11879 );
and ( n11881 , n11869 , n11880 );
and ( n11882 , n11791 , n11880 );
or ( n11883 , n11870 , n11881 , n11882 );
and ( n11884 , n11731 , n11883 );
and ( n11885 , n11635 , n11883 );
or ( n11886 , n11732 , n11884 , n11885 );
xor ( n11887 , n11407 , n11409 );
xor ( n11888 , n11887 , n11412 );
xor ( n11889 , n11418 , n11419 );
xor ( n11890 , n11889 , n11430 );
and ( n11891 , n11888 , n11890 );
xor ( n11892 , n11447 , n11456 );
xor ( n11893 , n11892 , n11474 );
and ( n11894 , n11890 , n11893 );
and ( n11895 , n11888 , n11893 );
or ( n11896 , n11891 , n11894 , n11895 );
xor ( n11897 , n11405 , n11415 );
xor ( n11898 , n11897 , n11433 );
and ( n11899 , n11896 , n11898 );
xor ( n11900 , n11477 , n11542 );
xor ( n11901 , n11900 , n11553 );
and ( n11902 , n11898 , n11901 );
and ( n11903 , n11896 , n11901 );
or ( n11904 , n11899 , n11902 , n11903 );
and ( n11905 , n11886 , n11904 );
xor ( n11906 , n11334 , n11436 );
xor ( n11907 , n11906 , n11556 );
and ( n11908 , n11904 , n11907 );
and ( n11909 , n11886 , n11907 );
or ( n11910 , n11905 , n11908 , n11909 );
xor ( n11911 , n11559 , n11585 );
xor ( n11912 , n11911 , n11596 );
and ( n11913 , n11910 , n11912 );
xor ( n11914 , n11601 , n11603 );
xor ( n11915 , n11914 , n11606 );
and ( n11916 , n11912 , n11915 );
and ( n11917 , n11910 , n11915 );
or ( n11918 , n11913 , n11916 , n11917 );
and ( n11919 , n11625 , n11918 );
xor ( n11920 , n11599 , n11609 );
xor ( n11921 , n11920 , n11612 );
and ( n11922 , n11918 , n11921 );
and ( n11923 , n11625 , n11921 );
or ( n11924 , n11919 , n11922 , n11923 );
and ( n11925 , n11623 , n11924 );
xor ( n11926 , n11329 , n11331 );
xor ( n11927 , n11926 , n11615 );
and ( n11928 , n11924 , n11927 );
and ( n11929 , n11623 , n11927 );
or ( n11930 , n11925 , n11928 , n11929 );
and ( n11931 , n11620 , n11930 );
and ( n11932 , n11618 , n11930 );
or ( n11933 , n11621 , n11931 , n11932 );
and ( n11934 , n11311 , n11933 );
xor ( n11935 , n11311 , n11933 );
xor ( n11936 , n11618 , n11620 );
xor ( n11937 , n11936 , n11930 );
xor ( n11938 , n11623 , n11924 );
xor ( n11939 , n11938 , n11927 );
xor ( n11940 , n11625 , n11918 );
xor ( n11941 , n11940 , n11921 );
xor ( n11942 , n11569 , n11579 );
xor ( n11943 , n11942 , n11582 );
xor ( n11944 , n11588 , n11590 );
xor ( n11945 , n11944 , n11593 );
and ( n11946 , n11943 , n11945 );
xor ( n11947 , n11561 , n11563 );
xor ( n11948 , n11947 , n11566 );
xor ( n11949 , n11571 , n11573 );
xor ( n11950 , n11949 , n11576 );
and ( n11951 , n11948 , n11950 );
xor ( n11952 , n11503 , n11528 );
xor ( n11953 , n11952 , n11539 );
xor ( n11954 , n11545 , n11547 );
xor ( n11955 , n11954 , n11550 );
and ( n11956 , n11953 , n11955 );
xor ( n11957 , n11531 , n11533 );
xor ( n11958 , n11957 , n11536 );
and ( n11959 , n1353 , n11111 );
and ( n11960 , n11116 , n1348 );
and ( n11961 , n11959 , n11960 );
and ( n11962 , n1995 , n3449 );
and ( n11963 , n3454 , n1990 );
and ( n11964 , n11962 , n11963 );
and ( n11965 , n11961 , n11964 );
and ( n11966 , n5177 , n1860 );
and ( n11967 , n11964 , n11966 );
and ( n11968 , n11961 , n11966 );
or ( n11969 , n11965 , n11967 , n11968 );
and ( n11970 , n1911 , n3739 );
and ( n11971 , n3728 , n1906 );
and ( n11972 , n11970 , n11971 );
and ( n11973 , n3169 , n5077 );
and ( n11974 , n11972 , n11973 );
and ( n11975 , n2764 , n11777 );
and ( n11976 , n11973 , n11975 );
and ( n11977 , n11972 , n11975 );
or ( n11978 , n11974 , n11976 , n11977 );
and ( n11979 , n11969 , n11978 );
and ( n11980 , n10933 , n1530 );
and ( n11981 , n4385 , n2577 );
and ( n11982 , n11980 , n11981 );
and ( n11983 , n4138 , n2948 );
and ( n11984 , n11981 , n11983 );
and ( n11985 , n11980 , n11983 );
or ( n11986 , n11982 , n11984 , n11985 );
and ( n11987 , n11978 , n11986 );
and ( n11988 , n11969 , n11986 );
or ( n11989 , n11979 , n11987 , n11988 );
xor ( n11990 , n11448 , n11449 );
xor ( n11991 , n11990 , n11451 );
and ( n11992 , n11989 , n11991 );
and ( n11993 , n11958 , n11992 );
xor ( n11994 , n11665 , n11668 );
xor ( n11995 , n11994 , n11670 );
xor ( n11996 , n11761 , n11762 );
xor ( n11997 , n11996 , n11764 );
and ( n11998 , n11995 , n11997 );
xor ( n11999 , n11698 , n11699 );
xor ( n12000 , n11999 , n11701 );
and ( n12001 , n11997 , n12000 );
and ( n12002 , n11995 , n12000 );
or ( n12003 , n11998 , n12001 , n12002 );
xor ( n12004 , n11717 , n11719 );
xor ( n12005 , n12004 , n11722 );
and ( n12006 , n12003 , n12005 );
and ( n12007 , n11992 , n12006 );
and ( n12008 , n11958 , n12006 );
or ( n12009 , n11993 , n12007 , n12008 );
and ( n12010 , n11955 , n12009 );
and ( n12011 , n11953 , n12009 );
or ( n12012 , n11956 , n12010 , n12011 );
and ( n12013 , n11950 , n12012 );
and ( n12014 , n11948 , n12012 );
or ( n12015 , n11951 , n12013 , n12014 );
and ( n12016 , n11945 , n12015 );
and ( n12017 , n11943 , n12015 );
or ( n12018 , n11946 , n12016 , n12017 );
xor ( n12019 , n11910 , n11912 );
xor ( n12020 , n12019 , n11915 );
and ( n12021 , n12018 , n12020 );
xor ( n12022 , n11662 , n11673 );
xor ( n12023 , n12022 , n11683 );
xor ( n12024 , n11695 , n11704 );
xor ( n12025 , n12024 , n11711 );
and ( n12026 , n12023 , n12025 );
and ( n12027 , n1694 , n4362 );
and ( n12028 , n4367 , n1689 );
and ( n12029 , n12027 , n12028 );
and ( n12030 , n1778 , n3903 );
and ( n12031 , n3892 , n1789 );
and ( n12032 , n12030 , n12031 );
and ( n12033 , n12029 , n12032 );
and ( n12034 , n3645 , n3627 );
and ( n12035 , n12032 , n12034 );
and ( n12036 , n12029 , n12034 );
or ( n12037 , n12033 , n12035 , n12036 );
and ( n12038 , n2255 , n3146 );
and ( n12039 , n3151 , n2250 );
and ( n12040 , n12038 , n12039 );
and ( n12041 , n4579 , n2407 );
and ( n12042 , n12040 , n12041 );
and ( n12043 , n3246 , n4522 );
and ( n12044 , n12041 , n12043 );
and ( n12045 , n12040 , n12043 );
or ( n12046 , n12042 , n12044 , n12045 );
and ( n12047 , n12037 , n12046 );
and ( n12048 , n2309 , n2923 );
and ( n12049 , n2928 , n2304 );
and ( n12050 , n12048 , n12049 );
and ( n12051 , n2497 , n2718 );
and ( n12052 , n2723 , n2492 );
and ( n12053 , n12051 , n12052 );
and ( n12054 , n12050 , n12053 );
and ( n12055 , n10886 , n1711 );
and ( n12056 , n12053 , n12055 );
and ( n12057 , n12050 , n12055 );
or ( n12058 , n12054 , n12056 , n12057 );
and ( n12059 , n12046 , n12058 );
and ( n12060 , n12037 , n12058 );
or ( n12061 , n12047 , n12059 , n12060 );
and ( n12062 , n12025 , n12061 );
and ( n12063 , n12023 , n12061 );
or ( n12064 , n12026 , n12062 , n12063 );
xor ( n12065 , n11768 , n11769 );
xor ( n12066 , n11771 , n11772 );
and ( n12067 , n12065 , n12066 );
and ( n12068 , n4579 , n2040 );
and ( n12069 , n12067 , n12068 );
xor ( n12070 , n11736 , n11737 );
xor ( n12071 , n12070 , n11739 );
xor ( n12072 , n11689 , n11690 );
xor ( n12073 , n12072 , n11692 );
and ( n12074 , n12071 , n12073 );
xor ( n12075 , n11770 , n11773 );
and ( n12076 , n12073 , n12075 );
and ( n12077 , n12071 , n12075 );
or ( n12078 , n12074 , n12076 , n12077 );
and ( n12079 , n12069 , n12078 );
and ( n12080 , n3339 , n3929 );
xnor ( n12081 , n11830 , n11831 );
and ( n12082 , n12080 , n12081 );
xor ( n12083 , n11833 , n11837 );
and ( n12084 , n12081 , n12083 );
and ( n12085 , n12080 , n12083 );
or ( n12086 , n12082 , n12084 , n12085 );
xor ( n12087 , n11663 , n11664 );
xor ( n12088 , n11759 , n11760 );
and ( n12089 , n12087 , n12088 );
xor ( n12090 , n11696 , n11697 );
and ( n12091 , n12088 , n12090 );
and ( n12092 , n12087 , n12090 );
or ( n12093 , n12089 , n12091 , n12092 );
and ( n12094 , n12086 , n12093 );
xor ( n12095 , n11666 , n11667 );
xor ( n12096 , n11675 , n11676 );
and ( n12097 , n12095 , n12096 );
xor ( n12098 , n11687 , n11688 );
and ( n12099 , n12096 , n12098 );
and ( n12100 , n12095 , n12098 );
or ( n12101 , n12097 , n12099 , n12100 );
and ( n12102 , n12093 , n12101 );
and ( n12103 , n12086 , n12101 );
or ( n12104 , n12094 , n12102 , n12103 );
and ( n12105 , n12078 , n12104 );
and ( n12106 , n12069 , n12104 );
or ( n12107 , n12079 , n12105 , n12106 );
and ( n12108 , n12064 , n12107 );
and ( n12109 , n1724 , n4161 );
and ( n12110 , n2048 , n3288 );
or ( n12111 , n12109 , n12110 );
buf ( n12112 , n2591 );
buf ( n12113 , n2634 );
and ( n12114 , n12112 , n12113 );
and ( n12115 , n12111 , n12114 );
and ( n12116 , n4150 , n1719 );
and ( n12117 , n3293 , n2059 );
and ( n12118 , n12116 , n12117 );
xor ( n12119 , n9328 , n10619 );
buf ( n12120 , n12119 );
buf ( n12121 , n12120 );
buf ( n12122 , n12121 );
and ( n12123 , n12117 , n12122 );
and ( n12124 , n12116 , n12122 );
or ( n12125 , n12118 , n12123 , n12124 );
and ( n12126 , n12114 , n12125 );
and ( n12127 , n12111 , n12125 );
or ( n12128 , n12115 , n12126 , n12127 );
xor ( n12129 , n11778 , n11779 );
xor ( n12130 , n12129 , n11782 );
and ( n12131 , n12128 , n12130 );
xor ( n12132 , n11792 , n11793 );
xor ( n12133 , n12132 , n11795 );
and ( n12134 , n12130 , n12133 );
and ( n12135 , n12128 , n12133 );
or ( n12136 , n12131 , n12134 , n12135 );
xor ( n12137 , n11799 , n11800 );
xor ( n12138 , n12137 , n11802 );
xor ( n12139 , n11807 , n11808 );
xor ( n12140 , n12139 , n11810 );
and ( n12141 , n12138 , n12140 );
xor ( n12142 , n11817 , n11818 );
xor ( n12143 , n12142 , n11826 );
and ( n12144 , n12140 , n12143 );
and ( n12145 , n12138 , n12143 );
or ( n12146 , n12141 , n12144 , n12145 );
and ( n12147 , n12136 , n12146 );
xor ( n12148 , n11735 , n11742 );
xor ( n12149 , n12148 , n11745 );
and ( n12150 , n12146 , n12149 );
and ( n12151 , n12136 , n12149 );
or ( n12152 , n12147 , n12150 , n12151 );
and ( n12153 , n12107 , n12152 );
and ( n12154 , n12064 , n12152 );
or ( n12155 , n12108 , n12153 , n12154 );
xor ( n12156 , n11750 , n11752 );
xor ( n12157 , n12156 , n11754 );
xor ( n12158 , n11767 , n11774 );
xor ( n12159 , n12158 , n11785 );
and ( n12160 , n12157 , n12159 );
xor ( n12161 , n11798 , n11805 );
xor ( n12162 , n12161 , n11813 );
and ( n12163 , n12159 , n12162 );
and ( n12164 , n12157 , n12162 );
or ( n12165 , n12160 , n12163 , n12164 );
xor ( n12166 , n11637 , n11639 );
xor ( n12167 , n12166 , n11642 );
and ( n12168 , n12165 , n12167 );
xor ( n12169 , n11647 , n11649 );
xor ( n12170 , n12169 , n11651 );
and ( n12171 , n12167 , n12170 );
and ( n12172 , n12165 , n12170 );
or ( n12173 , n12168 , n12171 , n12172 );
and ( n12174 , n12155 , n12173 );
xor ( n12175 , n11686 , n11714 );
xor ( n12176 , n12175 , n11725 );
xor ( n12177 , n11748 , n11757 );
xor ( n12178 , n12177 , n11788 );
and ( n12179 , n12176 , n12178 );
xor ( n12180 , n11816 , n11855 );
xor ( n12181 , n12180 , n11866 );
and ( n12182 , n12178 , n12181 );
and ( n12183 , n12176 , n12181 );
or ( n12184 , n12179 , n12182 , n12183 );
and ( n12185 , n12173 , n12184 );
and ( n12186 , n12155 , n12184 );
or ( n12187 , n12174 , n12185 , n12186 );
xor ( n12188 , n11627 , n11629 );
xor ( n12189 , n12188 , n11632 );
xor ( n12190 , n11645 , n11654 );
xor ( n12191 , n12190 , n11728 );
and ( n12192 , n12189 , n12191 );
xor ( n12193 , n11791 , n11869 );
xor ( n12194 , n12193 , n11880 );
and ( n12195 , n12191 , n12194 );
and ( n12196 , n12189 , n12194 );
or ( n12197 , n12192 , n12195 , n12196 );
and ( n12198 , n12187 , n12197 );
xor ( n12199 , n11635 , n11731 );
xor ( n12200 , n12199 , n11883 );
and ( n12201 , n12197 , n12200 );
and ( n12202 , n12187 , n12200 );
or ( n12203 , n12198 , n12201 , n12202 );
xor ( n12204 , n11886 , n11904 );
xor ( n12205 , n12204 , n11907 );
and ( n12206 , n12203 , n12205 );
xor ( n12207 , n11896 , n11898 );
xor ( n12208 , n12207 , n11901 );
xor ( n12209 , n11888 , n11890 );
xor ( n12210 , n12209 , n11893 );
xor ( n12211 , n11872 , n11874 );
xor ( n12212 , n12211 , n11877 );
xor ( n12213 , n11829 , n11849 );
xor ( n12214 , n12213 , n11852 );
xor ( n12215 , n11858 , n11860 );
xor ( n12216 , n12215 , n11863 );
and ( n12217 , n12214 , n12216 );
xor ( n12218 , n11989 , n11991 );
and ( n12219 , n12216 , n12218 );
and ( n12220 , n12214 , n12218 );
or ( n12221 , n12217 , n12219 , n12220 );
and ( n12222 , n12212 , n12221 );
xor ( n12223 , n12003 , n12005 );
xor ( n12224 , n11677 , n11678 );
xor ( n12225 , n12224 , n11680 );
xor ( n12226 , n12067 , n12068 );
and ( n12227 , n12225 , n12226 );
and ( n12228 , n12223 , n12227 );
xor ( n12229 , n11832 , n11838 );
xor ( n12230 , n12229 , n11846 );
xor ( n12231 , n11969 , n11978 );
xor ( n12232 , n12231 , n11986 );
and ( n12233 , n12230 , n12232 );
xor ( n12234 , n12037 , n12046 );
xor ( n12235 , n12234 , n12058 );
and ( n12236 , n12232 , n12235 );
and ( n12237 , n12230 , n12235 );
or ( n12238 , n12233 , n12236 , n12237 );
and ( n12239 , n12227 , n12238 );
and ( n12240 , n12223 , n12238 );
or ( n12241 , n12228 , n12239 , n12240 );
and ( n12242 , n12221 , n12241 );
and ( n12243 , n12212 , n12241 );
or ( n12244 , n12222 , n12242 , n12243 );
and ( n12245 , n12210 , n12244 );
xor ( n12246 , n11995 , n11997 );
xor ( n12247 , n12246 , n12000 );
and ( n12248 , n1995 , n3739 );
and ( n12249 , n3728 , n1990 );
and ( n12250 , n12248 , n12249 );
and ( n12251 , n2591 , n2718 );
and ( n12252 , n2723 , n2586 );
and ( n12253 , n12251 , n12252 );
and ( n12254 , n12250 , n12253 );
and ( n12255 , n3246 , n5077 );
and ( n12256 , n12253 , n12255 );
and ( n12257 , n12250 , n12255 );
or ( n12258 , n12254 , n12256 , n12257 );
and ( n12259 , n1778 , n4161 );
and ( n12260 , n4150 , n1789 );
and ( n12261 , n12259 , n12260 );
and ( n12262 , n2497 , n2923 );
and ( n12263 , n2928 , n2492 );
and ( n12264 , n12262 , n12263 );
and ( n12265 , n12261 , n12264 );
and ( n12266 , n4579 , n2577 );
and ( n12267 , n12264 , n12266 );
and ( n12268 , n12261 , n12266 );
or ( n12269 , n12265 , n12267 , n12268 );
and ( n12270 , n12258 , n12269 );
and ( n12271 , n1694 , n4734 );
and ( n12272 , n4739 , n1689 );
and ( n12273 , n12271 , n12272 );
and ( n12274 , n5177 , n2040 );
and ( n12275 , n12273 , n12274 );
and ( n12276 , n3339 , n4522 );
and ( n12277 , n12274 , n12276 );
and ( n12278 , n12273 , n12276 );
or ( n12279 , n12275 , n12277 , n12278 );
and ( n12280 , n12269 , n12279 );
and ( n12281 , n12258 , n12279 );
or ( n12282 , n12270 , n12280 , n12281 );
and ( n12283 , n12247 , n12282 );
and ( n12284 , n1911 , n3903 );
and ( n12285 , n3892 , n1906 );
and ( n12286 , n12284 , n12285 );
and ( n12287 , n3833 , n3627 );
and ( n12288 , n12286 , n12287 );
buf ( n12289 , n2632 );
buf ( n12290 , n12289 );
and ( n12291 , n2764 , n12290 );
and ( n12292 , n12287 , n12291 );
and ( n12293 , n12286 , n12291 );
or ( n12294 , n12288 , n12292 , n12293 );
xor ( n12295 , n11961 , n11964 );
xor ( n12296 , n12295 , n11966 );
and ( n12297 , n12294 , n12296 );
xor ( n12298 , n12029 , n12032 );
xor ( n12299 , n12298 , n12034 );
and ( n12300 , n12296 , n12299 );
and ( n12301 , n12294 , n12299 );
or ( n12302 , n12297 , n12300 , n12301 );
and ( n12303 , n12282 , n12302 );
and ( n12304 , n12247 , n12302 );
or ( n12305 , n12283 , n12303 , n12304 );
xor ( n12306 , n11980 , n11981 );
xor ( n12307 , n12306 , n11983 );
xor ( n12308 , n11820 , n11821 );
xor ( n12309 , n12308 , n11823 );
and ( n12310 , n12307 , n12309 );
xor ( n12311 , n12050 , n12053 );
xor ( n12312 , n12311 , n12055 );
and ( n12313 , n12309 , n12312 );
and ( n12314 , n12307 , n12312 );
or ( n12315 , n12310 , n12313 , n12314 );
xor ( n12316 , n11840 , n11841 );
xor ( n12317 , n12316 , n11843 );
xor ( n12318 , n11972 , n11973 );
xor ( n12319 , n12318 , n11975 );
and ( n12320 , n12317 , n12319 );
xor ( n12321 , n12040 , n12041 );
xor ( n12322 , n12321 , n12043 );
and ( n12323 , n12319 , n12322 );
and ( n12324 , n12317 , n12322 );
or ( n12325 , n12320 , n12323 , n12324 );
and ( n12326 , n12315 , n12325 );
xor ( n12327 , n12065 , n12066 );
and ( n12328 , n2309 , n3146 );
and ( n12329 , n3151 , n2304 );
and ( n12330 , n12328 , n12329 );
and ( n12331 , n10933 , n1711 );
and ( n12332 , n12330 , n12331 );
and ( n12333 , n4721 , n2407 );
and ( n12334 , n12331 , n12333 );
and ( n12335 , n12330 , n12333 );
or ( n12336 , n12332 , n12334 , n12335 );
and ( n12337 , n12327 , n12336 );
and ( n12338 , n2255 , n3288 );
and ( n12339 , n3293 , n2250 );
and ( n12340 , n12338 , n12339 );
and ( n12341 , n10886 , n1860 );
and ( n12342 , n12340 , n12341 );
and ( n12343 , n2937 , n11777 );
and ( n12344 , n12341 , n12343 );
and ( n12345 , n12340 , n12343 );
or ( n12346 , n12342 , n12344 , n12345 );
and ( n12347 , n12336 , n12346 );
and ( n12348 , n12327 , n12346 );
or ( n12349 , n12337 , n12347 , n12348 );
and ( n12350 , n12325 , n12349 );
and ( n12351 , n12315 , n12349 );
or ( n12352 , n12326 , n12350 , n12351 );
and ( n12353 , n12305 , n12352 );
and ( n12354 , n2048 , n3449 );
and ( n12355 , n3454 , n2059 );
and ( n12356 , n12354 , n12355 );
and ( n12357 , n4138 , n3301 );
and ( n12358 , n12356 , n12357 );
and ( n12359 , n3645 , n3929 );
and ( n12360 , n12357 , n12359 );
and ( n12361 , n12356 , n12359 );
or ( n12362 , n12358 , n12360 , n12361 );
and ( n12363 , n3169 , n11156 );
xnor ( n12364 , n12109 , n12110 );
and ( n12365 , n12363 , n12364 );
xor ( n12366 , n12112 , n12113 );
and ( n12367 , n12364 , n12366 );
and ( n12368 , n12363 , n12366 );
or ( n12369 , n12365 , n12367 , n12368 );
and ( n12370 , n12362 , n12369 );
xor ( n12371 , n11959 , n11960 );
xor ( n12372 , n12027 , n12028 );
and ( n12373 , n12371 , n12372 );
xor ( n12374 , n12030 , n12031 );
and ( n12375 , n12372 , n12374 );
and ( n12376 , n12371 , n12374 );
or ( n12377 , n12373 , n12375 , n12376 );
and ( n12378 , n12369 , n12377 );
and ( n12379 , n12362 , n12377 );
or ( n12380 , n12370 , n12378 , n12379 );
xor ( n12381 , n11970 , n11971 );
xor ( n12382 , n11962 , n11963 );
and ( n12383 , n12381 , n12382 );
xor ( n12384 , n12038 , n12039 );
and ( n12385 , n12382 , n12384 );
and ( n12386 , n12381 , n12384 );
or ( n12387 , n12383 , n12385 , n12386 );
xor ( n12388 , n12048 , n12049 );
xor ( n12389 , n12051 , n12052 );
and ( n12390 , n12388 , n12389 );
and ( n12391 , n1724 , n4362 );
and ( n12392 , n4367 , n1719 );
and ( n12393 , n12391 , n12392 );
and ( n12394 , n12389 , n12393 );
and ( n12395 , n12388 , n12393 );
or ( n12396 , n12390 , n12394 , n12395 );
and ( n12397 , n12387 , n12396 );
xor ( n12398 , n12080 , n12081 );
xor ( n12399 , n12398 , n12083 );
and ( n12400 , n12396 , n12399 );
and ( n12401 , n12387 , n12399 );
or ( n12402 , n12397 , n12400 , n12401 );
and ( n12403 , n12380 , n12402 );
xor ( n12404 , n12087 , n12088 );
xor ( n12405 , n12404 , n12090 );
xor ( n12406 , n12095 , n12096 );
xor ( n12407 , n12406 , n12098 );
and ( n12408 , n12405 , n12407 );
xor ( n12409 , n12111 , n12114 );
xor ( n12410 , n12409 , n12125 );
and ( n12411 , n12407 , n12410 );
and ( n12412 , n12405 , n12410 );
or ( n12413 , n12408 , n12411 , n12412 );
and ( n12414 , n12402 , n12413 );
and ( n12415 , n12380 , n12413 );
or ( n12416 , n12403 , n12414 , n12415 );
and ( n12417 , n12352 , n12416 );
and ( n12418 , n12305 , n12416 );
or ( n12419 , n12353 , n12417 , n12418 );
xor ( n12420 , n12071 , n12073 );
xor ( n12421 , n12420 , n12075 );
xor ( n12422 , n12086 , n12093 );
xor ( n12423 , n12422 , n12101 );
and ( n12424 , n12421 , n12423 );
xor ( n12425 , n12128 , n12130 );
xor ( n12426 , n12425 , n12133 );
and ( n12427 , n12423 , n12426 );
and ( n12428 , n12421 , n12426 );
or ( n12429 , n12424 , n12427 , n12428 );
xor ( n12430 , n12023 , n12025 );
xor ( n12431 , n12430 , n12061 );
and ( n12432 , n12429 , n12431 );
xor ( n12433 , n12069 , n12078 );
xor ( n12434 , n12433 , n12104 );
and ( n12435 , n12431 , n12434 );
and ( n12436 , n12429 , n12434 );
or ( n12437 , n12432 , n12435 , n12436 );
and ( n12438 , n12419 , n12437 );
xor ( n12439 , n11958 , n11992 );
xor ( n12440 , n12439 , n12006 );
and ( n12441 , n12437 , n12440 );
and ( n12442 , n12419 , n12440 );
or ( n12443 , n12438 , n12441 , n12442 );
and ( n12444 , n12244 , n12443 );
and ( n12445 , n12210 , n12443 );
or ( n12446 , n12245 , n12444 , n12445 );
and ( n12447 , n12208 , n12446 );
xor ( n12448 , n12064 , n12107 );
xor ( n12449 , n12448 , n12152 );
xor ( n12450 , n12165 , n12167 );
xor ( n12451 , n12450 , n12170 );
and ( n12452 , n12449 , n12451 );
xor ( n12453 , n12176 , n12178 );
xor ( n12454 , n12453 , n12181 );
and ( n12455 , n12451 , n12454 );
and ( n12456 , n12449 , n12454 );
or ( n12457 , n12452 , n12455 , n12456 );
xor ( n12458 , n11953 , n11955 );
xor ( n12459 , n12458 , n12009 );
and ( n12460 , n12457 , n12459 );
xor ( n12461 , n12155 , n12173 );
xor ( n12462 , n12461 , n12184 );
and ( n12463 , n12459 , n12462 );
and ( n12464 , n12457 , n12462 );
or ( n12465 , n12460 , n12463 , n12464 );
and ( n12466 , n12446 , n12465 );
and ( n12467 , n12208 , n12465 );
or ( n12468 , n12447 , n12466 , n12467 );
and ( n12469 , n12205 , n12468 );
and ( n12470 , n12203 , n12468 );
or ( n12471 , n12206 , n12469 , n12470 );
and ( n12472 , n12020 , n12471 );
and ( n12473 , n12018 , n12471 );
or ( n12474 , n12021 , n12472 , n12473 );
and ( n12475 , n11941 , n12474 );
xor ( n12476 , n11941 , n12474 );
xor ( n12477 , n11943 , n11945 );
xor ( n12478 , n12477 , n12015 );
xor ( n12479 , n11948 , n11950 );
xor ( n12480 , n12479 , n12012 );
xor ( n12481 , n12187 , n12197 );
xor ( n12482 , n12481 , n12200 );
and ( n12483 , n12480 , n12482 );
xor ( n12484 , n12189 , n12191 );
xor ( n12485 , n12484 , n12194 );
xor ( n12486 , n12136 , n12146 );
xor ( n12487 , n12486 , n12149 );
xor ( n12488 , n12157 , n12159 );
xor ( n12489 , n12488 , n12162 );
and ( n12490 , n12487 , n12489 );
xor ( n12491 , n12138 , n12140 );
xor ( n12492 , n12491 , n12143 );
xor ( n12493 , n12225 , n12226 );
and ( n12494 , n12492 , n12493 );
xor ( n12495 , n12258 , n12269 );
xor ( n12496 , n12495 , n12279 );
xor ( n12497 , n12294 , n12296 );
xor ( n12498 , n12497 , n12299 );
and ( n12499 , n12496 , n12498 );
xor ( n12500 , n12307 , n12309 );
xor ( n12501 , n12500 , n12312 );
and ( n12502 , n12498 , n12501 );
and ( n12503 , n12496 , n12501 );
or ( n12504 , n12499 , n12502 , n12503 );
and ( n12505 , n12493 , n12504 );
and ( n12506 , n12492 , n12504 );
or ( n12507 , n12494 , n12505 , n12506 );
and ( n12508 , n12489 , n12507 );
and ( n12509 , n12487 , n12507 );
or ( n12510 , n12490 , n12508 , n12509 );
and ( n12511 , n1911 , n4161 );
and ( n12512 , n4150 , n1906 );
and ( n12513 , n12511 , n12512 );
and ( n12514 , n4385 , n3301 );
and ( n12515 , n12513 , n12514 );
and ( n12516 , n3246 , n11156 );
and ( n12517 , n12514 , n12516 );
and ( n12518 , n12513 , n12516 );
or ( n12519 , n12515 , n12517 , n12518 );
and ( n12520 , n1694 , n4982 );
and ( n12521 , n4989 , n1689 );
and ( n12522 , n12520 , n12521 );
and ( n12523 , n4721 , n2577 );
and ( n12524 , n12522 , n12523 );
and ( n12525 , n3169 , n11777 );
and ( n12526 , n12523 , n12525 );
and ( n12527 , n12522 , n12525 );
or ( n12528 , n12524 , n12526 , n12527 );
and ( n12529 , n12519 , n12528 );
and ( n12530 , n2591 , n2923 );
and ( n12531 , n2928 , n2586 );
and ( n12532 , n12530 , n12531 );
and ( n12533 , n5177 , n2407 );
and ( n12534 , n12532 , n12533 );
and ( n12535 , n4138 , n3627 );
and ( n12536 , n12533 , n12535 );
and ( n12537 , n12532 , n12535 );
or ( n12538 , n12534 , n12536 , n12537 );
and ( n12539 , n12528 , n12538 );
and ( n12540 , n12519 , n12538 );
or ( n12541 , n12529 , n12539 , n12540 );
and ( n12542 , n1724 , n4734 );
and ( n12543 , n4739 , n1719 );
and ( n12544 , n12542 , n12543 );
and ( n12545 , n2048 , n3739 );
and ( n12546 , n3728 , n2059 );
and ( n12547 , n12545 , n12546 );
and ( n12548 , n12544 , n12547 );
and ( n12549 , n10933 , n1860 );
and ( n12550 , n12547 , n12549 );
and ( n12551 , n12544 , n12549 );
or ( n12552 , n12548 , n12550 , n12551 );
and ( n12553 , n2497 , n3146 );
and ( n12554 , n3151 , n2492 );
and ( n12555 , n12553 , n12554 );
and ( n12556 , n3833 , n3929 );
and ( n12557 , n12555 , n12556 );
and ( n12558 , n2937 , n12290 );
and ( n12559 , n12556 , n12558 );
and ( n12560 , n12555 , n12558 );
or ( n12561 , n12557 , n12559 , n12560 );
and ( n12562 , n12552 , n12561 );
and ( n12563 , n4385 , n2948 );
and ( n12564 , n12561 , n12563 );
and ( n12565 , n12552 , n12563 );
or ( n12566 , n12562 , n12564 , n12565 );
and ( n12567 , n12541 , n12566 );
and ( n12568 , n2309 , n3288 );
and ( n12569 , n3293 , n2304 );
and ( n12570 , n12568 , n12569 );
and ( n12571 , n4579 , n2948 );
and ( n12572 , n12570 , n12571 );
and ( n12573 , n3339 , n5077 );
and ( n12574 , n12571 , n12573 );
and ( n12575 , n12570 , n12573 );
or ( n12576 , n12572 , n12574 , n12575 );
xor ( n12577 , n12356 , n12357 );
xor ( n12578 , n12577 , n12359 );
and ( n12579 , n12576 , n12578 );
xor ( n12580 , n12261 , n12264 );
xor ( n12581 , n12580 , n12266 );
and ( n12582 , n12578 , n12581 );
and ( n12583 , n12576 , n12581 );
or ( n12584 , n12579 , n12582 , n12583 );
and ( n12585 , n12566 , n12584 );
and ( n12586 , n12541 , n12584 );
or ( n12587 , n12567 , n12585 , n12586 );
xor ( n12588 , n12330 , n12331 );
xor ( n12589 , n12588 , n12333 );
xor ( n12590 , n12250 , n12253 );
xor ( n12591 , n12590 , n12255 );
and ( n12592 , n12589 , n12591 );
xor ( n12593 , n12340 , n12341 );
xor ( n12594 , n12593 , n12343 );
and ( n12595 , n12591 , n12594 );
and ( n12596 , n12589 , n12594 );
or ( n12597 , n12592 , n12595 , n12596 );
xor ( n12598 , n12116 , n12117 );
xor ( n12599 , n12598 , n12122 );
xor ( n12600 , n12286 , n12287 );
xor ( n12601 , n12600 , n12291 );
and ( n12602 , n12599 , n12601 );
xor ( n12603 , n12273 , n12274 );
xor ( n12604 , n12603 , n12276 );
and ( n12605 , n12601 , n12604 );
and ( n12606 , n12599 , n12604 );
or ( n12607 , n12602 , n12605 , n12606 );
and ( n12608 , n12597 , n12607 );
and ( n12609 , n1995 , n3903 );
and ( n12610 , n3892 , n1990 );
and ( n12611 , n12609 , n12610 );
and ( n12612 , n10886 , n2040 );
and ( n12613 , n12611 , n12612 );
and ( n12614 , n3645 , n4522 );
and ( n12615 , n12612 , n12614 );
and ( n12616 , n12611 , n12614 );
or ( n12617 , n12613 , n12615 , n12616 );
xor ( n12618 , n9331 , n10617 );
buf ( n12619 , n12618 );
buf ( n12620 , n12619 );
buf ( n12621 , n12620 );
xor ( n12622 , n12271 , n12272 );
and ( n12623 , n12621 , n12622 );
xor ( n12624 , n12391 , n12392 );
and ( n12625 , n12622 , n12624 );
and ( n12626 , n12621 , n12624 );
or ( n12627 , n12623 , n12625 , n12626 );
and ( n12628 , n12617 , n12627 );
xor ( n12629 , n12259 , n12260 );
xor ( n12630 , n12284 , n12285 );
and ( n12631 , n12629 , n12630 );
xor ( n12632 , n12248 , n12249 );
and ( n12633 , n12630 , n12632 );
and ( n12634 , n12629 , n12632 );
or ( n12635 , n12631 , n12633 , n12634 );
and ( n12636 , n12627 , n12635 );
and ( n12637 , n12617 , n12635 );
or ( n12638 , n12628 , n12636 , n12637 );
and ( n12639 , n12607 , n12638 );
and ( n12640 , n12597 , n12638 );
or ( n12641 , n12608 , n12639 , n12640 );
and ( n12642 , n12587 , n12641 );
xor ( n12643 , n12354 , n12355 );
xor ( n12644 , n12338 , n12339 );
and ( n12645 , n12643 , n12644 );
xor ( n12646 , n12328 , n12329 );
and ( n12647 , n12644 , n12646 );
and ( n12648 , n12643 , n12646 );
or ( n12649 , n12645 , n12647 , n12648 );
xor ( n12650 , n12262 , n12263 );
xor ( n12651 , n12251 , n12252 );
and ( n12652 , n12650 , n12651 );
buf ( n12653 , n2723 );
buf ( n12654 , n2764 );
or ( n12655 , n12653 , n12654 );
and ( n12656 , n12651 , n12655 );
and ( n12657 , n12650 , n12655 );
or ( n12658 , n12652 , n12656 , n12657 );
and ( n12659 , n12649 , n12658 );
and ( n12660 , n1778 , n4362 );
and ( n12661 , n4367 , n1789 );
and ( n12662 , n12660 , n12661 );
and ( n12663 , n2255 , n3449 );
and ( n12664 , n3454 , n2250 );
and ( n12665 , n12663 , n12664 );
and ( n12666 , n12662 , n12665 );
xor ( n12667 , n9332 , n10616 );
buf ( n12668 , n12667 );
buf ( n12669 , n12668 );
buf ( n12670 , n12669 );
and ( n12671 , n4385 , n3627 );
and ( n12672 , n12670 , n12671 );
and ( n12673 , n3833 , n4522 );
and ( n12674 , n12671 , n12673 );
and ( n12675 , n12670 , n12673 );
or ( n12676 , n12672 , n12674 , n12675 );
and ( n12677 , n12665 , n12676 );
and ( n12678 , n12662 , n12676 );
or ( n12679 , n12666 , n12677 , n12678 );
and ( n12680 , n12658 , n12679 );
and ( n12681 , n12649 , n12679 );
or ( n12682 , n12659 , n12680 , n12681 );
xor ( n12683 , n12363 , n12364 );
xor ( n12684 , n12683 , n12366 );
xor ( n12685 , n12371 , n12372 );
xor ( n12686 , n12685 , n12374 );
and ( n12687 , n12684 , n12686 );
xor ( n12688 , n12381 , n12382 );
xor ( n12689 , n12688 , n12384 );
and ( n12690 , n12686 , n12689 );
and ( n12691 , n12684 , n12689 );
or ( n12692 , n12687 , n12690 , n12691 );
and ( n12693 , n12682 , n12692 );
xor ( n12694 , n12317 , n12319 );
xor ( n12695 , n12694 , n12322 );
and ( n12696 , n12692 , n12695 );
and ( n12697 , n12682 , n12695 );
or ( n12698 , n12693 , n12696 , n12697 );
and ( n12699 , n12641 , n12698 );
and ( n12700 , n12587 , n12698 );
or ( n12701 , n12642 , n12699 , n12700 );
xor ( n12702 , n12327 , n12336 );
xor ( n12703 , n12702 , n12346 );
xor ( n12704 , n12362 , n12369 );
xor ( n12705 , n12704 , n12377 );
and ( n12706 , n12703 , n12705 );
xor ( n12707 , n12387 , n12396 );
xor ( n12708 , n12707 , n12399 );
and ( n12709 , n12705 , n12708 );
and ( n12710 , n12703 , n12708 );
or ( n12711 , n12706 , n12709 , n12710 );
xor ( n12712 , n12230 , n12232 );
xor ( n12713 , n12712 , n12235 );
and ( n12714 , n12711 , n12713 );
xor ( n12715 , n12247 , n12282 );
xor ( n12716 , n12715 , n12302 );
and ( n12717 , n12713 , n12716 );
and ( n12718 , n12711 , n12716 );
or ( n12719 , n12714 , n12717 , n12718 );
and ( n12720 , n12701 , n12719 );
xor ( n12721 , n12315 , n12325 );
xor ( n12722 , n12721 , n12349 );
xor ( n12723 , n12380 , n12402 );
xor ( n12724 , n12723 , n12413 );
and ( n12725 , n12722 , n12724 );
xor ( n12726 , n12421 , n12423 );
xor ( n12727 , n12726 , n12426 );
and ( n12728 , n12724 , n12727 );
and ( n12729 , n12722 , n12727 );
or ( n12730 , n12725 , n12728 , n12729 );
and ( n12731 , n12719 , n12730 );
and ( n12732 , n12701 , n12730 );
or ( n12733 , n12720 , n12731 , n12732 );
and ( n12734 , n12510 , n12733 );
xor ( n12735 , n12214 , n12216 );
xor ( n12736 , n12735 , n12218 );
xor ( n12737 , n12223 , n12227 );
xor ( n12738 , n12737 , n12238 );
and ( n12739 , n12736 , n12738 );
xor ( n12740 , n12305 , n12352 );
xor ( n12741 , n12740 , n12416 );
and ( n12742 , n12738 , n12741 );
and ( n12743 , n12736 , n12741 );
or ( n12744 , n12739 , n12742 , n12743 );
and ( n12745 , n12733 , n12744 );
and ( n12746 , n12510 , n12744 );
or ( n12747 , n12734 , n12745 , n12746 );
and ( n12748 , n12485 , n12747 );
xor ( n12749 , n12212 , n12221 );
xor ( n12750 , n12749 , n12241 );
xor ( n12751 , n12419 , n12437 );
xor ( n12752 , n12751 , n12440 );
and ( n12753 , n12750 , n12752 );
xor ( n12754 , n12449 , n12451 );
xor ( n12755 , n12754 , n12454 );
and ( n12756 , n12752 , n12755 );
and ( n12757 , n12750 , n12755 );
or ( n12758 , n12753 , n12756 , n12757 );
and ( n12759 , n12747 , n12758 );
and ( n12760 , n12485 , n12758 );
or ( n12761 , n12748 , n12759 , n12760 );
and ( n12762 , n12482 , n12761 );
and ( n12763 , n12480 , n12761 );
or ( n12764 , n12483 , n12762 , n12763 );
and ( n12765 , n12478 , n12764 );
xor ( n12766 , n12203 , n12205 );
xor ( n12767 , n12766 , n12468 );
and ( n12768 , n12764 , n12767 );
and ( n12769 , n12478 , n12767 );
or ( n12770 , n12765 , n12768 , n12769 );
xor ( n12771 , n12018 , n12020 );
xor ( n12772 , n12771 , n12471 );
and ( n12773 , n12770 , n12772 );
xor ( n12774 , n12770 , n12772 );
xor ( n12775 , n12208 , n12446 );
xor ( n12776 , n12775 , n12465 );
xor ( n12777 , n12210 , n12244 );
xor ( n12778 , n12777 , n12443 );
xor ( n12779 , n12457 , n12459 );
xor ( n12780 , n12779 , n12462 );
and ( n12781 , n12778 , n12780 );
xor ( n12782 , n12429 , n12431 );
xor ( n12783 , n12782 , n12434 );
xor ( n12784 , n12405 , n12407 );
xor ( n12785 , n12784 , n12410 );
and ( n12786 , n1778 , n4734 );
and ( n12787 , n4739 , n1789 );
and ( n12788 , n12786 , n12787 );
and ( n12789 , n10933 , n2040 );
and ( n12790 , n12788 , n12789 );
and ( n12791 , n4721 , n2948 );
and ( n12792 , n12789 , n12791 );
and ( n12793 , n12788 , n12791 );
or ( n12794 , n12790 , n12792 , n12793 );
and ( n12795 , n2591 , n3146 );
and ( n12796 , n3151 , n2586 );
and ( n12797 , n12795 , n12796 );
and ( n12798 , n4579 , n3301 );
and ( n12799 , n12797 , n12798 );
and ( n12800 , n3645 , n5077 );
and ( n12801 , n12798 , n12800 );
and ( n12802 , n12797 , n12800 );
or ( n12803 , n12799 , n12801 , n12802 );
and ( n12804 , n12794 , n12803 );
xor ( n12805 , n12522 , n12523 );
xor ( n12806 , n12805 , n12525 );
and ( n12807 , n12803 , n12806 );
and ( n12808 , n12794 , n12806 );
or ( n12809 , n12804 , n12807 , n12808 );
xor ( n12810 , n12611 , n12612 );
xor ( n12811 , n12810 , n12614 );
xor ( n12812 , n12555 , n12556 );
xor ( n12813 , n12812 , n12558 );
and ( n12814 , n12811 , n12813 );
xor ( n12815 , n12532 , n12533 );
xor ( n12816 , n12815 , n12535 );
and ( n12817 , n12813 , n12816 );
and ( n12818 , n12811 , n12816 );
or ( n12819 , n12814 , n12817 , n12818 );
and ( n12820 , n12809 , n12819 );
xor ( n12821 , n12552 , n12561 );
xor ( n12822 , n12821 , n12563 );
and ( n12823 , n12819 , n12822 );
and ( n12824 , n12809 , n12822 );
or ( n12825 , n12820 , n12823 , n12824 );
and ( n12826 , n12785 , n12825 );
xor ( n12827 , n12513 , n12514 );
xor ( n12828 , n12827 , n12516 );
xor ( n12829 , n12570 , n12571 );
xor ( n12830 , n12829 , n12573 );
and ( n12831 , n12828 , n12830 );
xor ( n12832 , n12544 , n12547 );
xor ( n12833 , n12832 , n12549 );
and ( n12834 , n12830 , n12833 );
and ( n12835 , n12828 , n12833 );
or ( n12836 , n12831 , n12834 , n12835 );
xor ( n12837 , n12519 , n12528 );
xor ( n12838 , n12837 , n12538 );
and ( n12839 , n12836 , n12838 );
and ( n12840 , n12825 , n12839 );
and ( n12841 , n12785 , n12839 );
or ( n12842 , n12826 , n12840 , n12841 );
xor ( n12843 , n12388 , n12389 );
xor ( n12844 , n12843 , n12393 );
xor ( n12845 , n12576 , n12578 );
xor ( n12846 , n12845 , n12581 );
and ( n12847 , n12844 , n12846 );
xor ( n12848 , n12589 , n12591 );
xor ( n12849 , n12848 , n12594 );
and ( n12850 , n12846 , n12849 );
and ( n12851 , n12844 , n12849 );
or ( n12852 , n12847 , n12850 , n12851 );
and ( n12853 , n2048 , n3903 );
and ( n12854 , n3892 , n2059 );
and ( n12855 , n12853 , n12854 );
and ( n12856 , n3339 , n11156 );
and ( n12857 , n12855 , n12856 );
and ( n12858 , n3246 , n11777 );
and ( n12859 , n12856 , n12858 );
and ( n12860 , n12855 , n12858 );
or ( n12861 , n12857 , n12859 , n12860 );
and ( n12862 , n2309 , n3449 );
and ( n12863 , n3454 , n2304 );
and ( n12864 , n12862 , n12863 );
and ( n12865 , n5177 , n2577 );
and ( n12866 , n12864 , n12865 );
and ( n12867 , n3169 , n12290 );
and ( n12868 , n12865 , n12867 );
and ( n12869 , n12864 , n12867 );
or ( n12870 , n12866 , n12868 , n12869 );
and ( n12871 , n12861 , n12870 );
and ( n12872 , n5091 , n1689 );
and ( n12873 , n3293 , n2492 );
and ( n12874 , n12872 , n12873 );
and ( n12875 , n2928 , n2718 );
and ( n12876 , n12873 , n12875 );
and ( n12877 , n12872 , n12875 );
or ( n12878 , n12874 , n12876 , n12877 );
and ( n12879 , n1694 , n5086 );
and ( n12880 , n2497 , n3288 );
and ( n12881 , n12879 , n12880 );
and ( n12882 , n2723 , n2923 );
and ( n12883 , n12880 , n12882 );
and ( n12884 , n12879 , n12882 );
or ( n12885 , n12881 , n12883 , n12884 );
and ( n12886 , n12878 , n12885 );
and ( n12887 , n12870 , n12886 );
and ( n12888 , n12861 , n12886 );
or ( n12889 , n12871 , n12887 , n12888 );
and ( n12890 , n1724 , n4982 );
and ( n12891 , n4989 , n1719 );
and ( n12892 , n12890 , n12891 );
and ( n12893 , n10886 , n2407 );
and ( n12894 , n12892 , n12893 );
and ( n12895 , n4138 , n3929 );
and ( n12896 , n12893 , n12895 );
and ( n12897 , n12892 , n12895 );
or ( n12898 , n12894 , n12896 , n12897 );
buf ( n12899 , n2762 );
buf ( n12900 , n12899 );
and ( n12901 , n2937 , n12900 );
xnor ( n12902 , n12653 , n12654 );
and ( n12903 , n12901 , n12902 );
xor ( n12904 , n12520 , n12521 );
and ( n12905 , n12902 , n12904 );
and ( n12906 , n12901 , n12904 );
or ( n12907 , n12903 , n12905 , n12906 );
and ( n12908 , n12898 , n12907 );
xor ( n12909 , n12542 , n12543 );
xor ( n12910 , n12660 , n12661 );
and ( n12911 , n12909 , n12910 );
xor ( n12912 , n12511 , n12512 );
and ( n12913 , n12910 , n12912 );
and ( n12914 , n12909 , n12912 );
or ( n12915 , n12911 , n12913 , n12914 );
and ( n12916 , n12907 , n12915 );
and ( n12917 , n12898 , n12915 );
or ( n12918 , n12908 , n12916 , n12917 );
and ( n12919 , n12889 , n12918 );
xor ( n12920 , n12609 , n12610 );
xor ( n12921 , n12545 , n12546 );
and ( n12922 , n12920 , n12921 );
xor ( n12923 , n12663 , n12664 );
and ( n12924 , n12921 , n12923 );
and ( n12925 , n12920 , n12923 );
or ( n12926 , n12922 , n12924 , n12925 );
xor ( n12927 , n12568 , n12569 );
xor ( n12928 , n12553 , n12554 );
and ( n12929 , n12927 , n12928 );
xor ( n12930 , n12530 , n12531 );
and ( n12931 , n12928 , n12930 );
and ( n12932 , n12927 , n12930 );
or ( n12933 , n12929 , n12931 , n12932 );
and ( n12934 , n12926 , n12933 );
and ( n12935 , n10933 , n2407 );
and ( n12936 , n5177 , n2948 );
and ( n12937 , n12935 , n12936 );
and ( n12938 , n3339 , n11777 );
and ( n12939 , n12936 , n12938 );
and ( n12940 , n12935 , n12938 );
or ( n12941 , n12937 , n12939 , n12940 );
and ( n12942 , n1995 , n4161 );
and ( n12943 , n2255 , n3739 );
or ( n12944 , n12942 , n12943 );
and ( n12945 , n12941 , n12944 );
and ( n12946 , n1911 , n4362 );
and ( n12947 , n4367 , n1906 );
and ( n12948 , n12946 , n12947 );
and ( n12949 , n12944 , n12948 );
and ( n12950 , n12941 , n12948 );
or ( n12951 , n12945 , n12949 , n12950 );
and ( n12952 , n12933 , n12951 );
and ( n12953 , n12926 , n12951 );
or ( n12954 , n12934 , n12952 , n12953 );
and ( n12955 , n12918 , n12954 );
and ( n12956 , n12889 , n12954 );
or ( n12957 , n12919 , n12955 , n12956 );
and ( n12958 , n12852 , n12957 );
and ( n12959 , n4150 , n1990 );
and ( n12960 , n3728 , n2250 );
and ( n12961 , n12959 , n12960 );
xor ( n12962 , n10018 , n10614 );
buf ( n12963 , n12962 );
buf ( n12964 , n12963 );
buf ( n12965 , n12964 );
and ( n12966 , n12960 , n12965 );
and ( n12967 , n12959 , n12965 );
or ( n12968 , n12961 , n12966 , n12967 );
and ( n12969 , n4385 , n3929 );
and ( n12970 , n3645 , n11156 );
and ( n12971 , n12969 , n12970 );
and ( n12972 , n3246 , n12290 );
and ( n12973 , n12970 , n12972 );
and ( n12974 , n12969 , n12972 );
or ( n12975 , n12971 , n12973 , n12974 );
and ( n12976 , n12968 , n12975 );
xor ( n12977 , n12670 , n12671 );
xor ( n12978 , n12977 , n12673 );
and ( n12979 , n12975 , n12978 );
and ( n12980 , n12968 , n12978 );
or ( n12981 , n12976 , n12979 , n12980 );
xor ( n12982 , n12621 , n12622 );
xor ( n12983 , n12982 , n12624 );
and ( n12984 , n12981 , n12983 );
xor ( n12985 , n12629 , n12630 );
xor ( n12986 , n12985 , n12632 );
and ( n12987 , n12983 , n12986 );
and ( n12988 , n12981 , n12986 );
or ( n12989 , n12984 , n12987 , n12988 );
xor ( n12990 , n12643 , n12644 );
xor ( n12991 , n12990 , n12646 );
xor ( n12992 , n12650 , n12651 );
xor ( n12993 , n12992 , n12655 );
and ( n12994 , n12991 , n12993 );
xor ( n12995 , n12662 , n12665 );
xor ( n12996 , n12995 , n12676 );
and ( n12997 , n12993 , n12996 );
and ( n12998 , n12991 , n12996 );
or ( n12999 , n12994 , n12997 , n12998 );
and ( n13000 , n12989 , n12999 );
xor ( n13001 , n12599 , n12601 );
xor ( n13002 , n13001 , n12604 );
and ( n13003 , n12999 , n13002 );
and ( n13004 , n12989 , n13002 );
or ( n13005 , n13000 , n13003 , n13004 );
and ( n13006 , n12957 , n13005 );
and ( n13007 , n12852 , n13005 );
or ( n13008 , n12958 , n13006 , n13007 );
and ( n13009 , n12842 , n13008 );
xor ( n13010 , n12617 , n12627 );
xor ( n13011 , n13010 , n12635 );
xor ( n13012 , n12649 , n12658 );
xor ( n13013 , n13012 , n12679 );
and ( n13014 , n13011 , n13013 );
xor ( n13015 , n12684 , n12686 );
xor ( n13016 , n13015 , n12689 );
and ( n13017 , n13013 , n13016 );
and ( n13018 , n13011 , n13016 );
or ( n13019 , n13014 , n13017 , n13018 );
xor ( n13020 , n12496 , n12498 );
xor ( n13021 , n13020 , n12501 );
and ( n13022 , n13019 , n13021 );
xor ( n13023 , n12541 , n12566 );
xor ( n13024 , n13023 , n12584 );
and ( n13025 , n13021 , n13024 );
and ( n13026 , n13019 , n13024 );
or ( n13027 , n13022 , n13025 , n13026 );
and ( n13028 , n13008 , n13027 );
and ( n13029 , n12842 , n13027 );
or ( n13030 , n13009 , n13028 , n13029 );
and ( n13031 , n12783 , n13030 );
xor ( n13032 , n12597 , n12607 );
xor ( n13033 , n13032 , n12638 );
xor ( n13034 , n12682 , n12692 );
xor ( n13035 , n13034 , n12695 );
and ( n13036 , n13033 , n13035 );
xor ( n13037 , n12703 , n12705 );
xor ( n13038 , n13037 , n12708 );
and ( n13039 , n13035 , n13038 );
and ( n13040 , n13033 , n13038 );
or ( n13041 , n13036 , n13039 , n13040 );
xor ( n13042 , n12492 , n12493 );
xor ( n13043 , n13042 , n12504 );
and ( n13044 , n13041 , n13043 );
xor ( n13045 , n12587 , n12641 );
xor ( n13046 , n13045 , n12698 );
and ( n13047 , n13043 , n13046 );
and ( n13048 , n13041 , n13046 );
or ( n13049 , n13044 , n13047 , n13048 );
and ( n13050 , n13030 , n13049 );
and ( n13051 , n12783 , n13049 );
or ( n13052 , n13031 , n13050 , n13051 );
xor ( n13053 , n12487 , n12489 );
xor ( n13054 , n13053 , n12507 );
xor ( n13055 , n12701 , n12719 );
xor ( n13056 , n13055 , n12730 );
and ( n13057 , n13054 , n13056 );
xor ( n13058 , n12736 , n12738 );
xor ( n13059 , n13058 , n12741 );
and ( n13060 , n13056 , n13059 );
and ( n13061 , n13054 , n13059 );
or ( n13062 , n13057 , n13060 , n13061 );
and ( n13063 , n13052 , n13062 );
xor ( n13064 , n12510 , n12733 );
xor ( n13065 , n13064 , n12744 );
and ( n13066 , n13062 , n13065 );
and ( n13067 , n13052 , n13065 );
or ( n13068 , n13063 , n13066 , n13067 );
and ( n13069 , n12780 , n13068 );
and ( n13070 , n12778 , n13068 );
or ( n13071 , n12781 , n13069 , n13070 );
and ( n13072 , n12776 , n13071 );
xor ( n13073 , n12480 , n12482 );
xor ( n13074 , n13073 , n12761 );
and ( n13075 , n13071 , n13074 );
and ( n13076 , n12776 , n13074 );
or ( n13077 , n13072 , n13075 , n13076 );
xor ( n13078 , n12478 , n12764 );
xor ( n13079 , n13078 , n12767 );
and ( n13080 , n13077 , n13079 );
xor ( n13081 , n13077 , n13079 );
xor ( n13082 , n12485 , n12747 );
xor ( n13083 , n13082 , n12758 );
xor ( n13084 , n12750 , n12752 );
xor ( n13085 , n13084 , n12755 );
xor ( n13086 , n12711 , n12713 );
xor ( n13087 , n13086 , n12716 );
xor ( n13088 , n12722 , n12724 );
xor ( n13089 , n13088 , n12727 );
and ( n13090 , n13087 , n13089 );
xor ( n13091 , n12809 , n12819 );
xor ( n13092 , n13091 , n12822 );
xor ( n13093 , n12836 , n12838 );
and ( n13094 , n13092 , n13093 );
xor ( n13095 , n12788 , n12789 );
xor ( n13096 , n13095 , n12791 );
xor ( n13097 , n12864 , n12865 );
xor ( n13098 , n13097 , n12867 );
and ( n13099 , n13096 , n13098 );
xor ( n13100 , n12797 , n12798 );
xor ( n13101 , n13100 , n12800 );
and ( n13102 , n13098 , n13101 );
and ( n13103 , n13096 , n13101 );
or ( n13104 , n13099 , n13102 , n13103 );
not ( n13105 , n13104 );
xor ( n13106 , n12861 , n12870 );
xor ( n13107 , n13106 , n12886 );
and ( n13108 , n13105 , n13107 );
and ( n13109 , n13093 , n13108 );
and ( n13110 , n13092 , n13108 );
or ( n13111 , n13094 , n13109 , n13110 );
buf ( n13112 , n13104 );
xor ( n13113 , n12794 , n12803 );
xor ( n13114 , n13113 , n12806 );
xor ( n13115 , n12828 , n12830 );
xor ( n13116 , n13115 , n12833 );
and ( n13117 , n13114 , n13116 );
xor ( n13118 , n12811 , n12813 );
xor ( n13119 , n13118 , n12816 );
and ( n13120 , n13116 , n13119 );
and ( n13121 , n13114 , n13119 );
or ( n13122 , n13117 , n13120 , n13121 );
and ( n13123 , n13112 , n13122 );
and ( n13124 , n5091 , n1719 );
and ( n13125 , n4989 , n1789 );
and ( n13126 , n13124 , n13125 );
and ( n13127 , n3454 , n2492 );
and ( n13128 , n13125 , n13127 );
and ( n13129 , n13124 , n13127 );
or ( n13130 , n13126 , n13128 , n13129 );
and ( n13131 , n1724 , n5086 );
and ( n13132 , n1778 , n4982 );
and ( n13133 , n13131 , n13132 );
and ( n13134 , n2497 , n3449 );
and ( n13135 , n13132 , n13134 );
and ( n13136 , n13131 , n13134 );
or ( n13137 , n13133 , n13135 , n13136 );
and ( n13138 , n13130 , n13137 );
xor ( n13139 , n12892 , n12893 );
xor ( n13140 , n13139 , n12895 );
and ( n13141 , n13138 , n13140 );
and ( n13142 , n2309 , n3739 );
and ( n13143 , n3728 , n2304 );
and ( n13144 , n13142 , n13143 );
and ( n13145 , n4721 , n3301 );
and ( n13146 , n13144 , n13145 );
and ( n13147 , n4138 , n4522 );
and ( n13148 , n13145 , n13147 );
and ( n13149 , n13144 , n13147 );
or ( n13150 , n13146 , n13148 , n13149 );
and ( n13151 , n1694 , n10869 );
and ( n13152 , n10862 , n1689 );
and ( n13153 , n13151 , n13152 );
and ( n13154 , n10886 , n2577 );
and ( n13155 , n13153 , n13154 );
and ( n13156 , n4579 , n3627 );
and ( n13157 , n13154 , n13156 );
and ( n13158 , n13153 , n13156 );
or ( n13159 , n13155 , n13157 , n13158 );
and ( n13160 , n13150 , n13159 );
and ( n13161 , n13141 , n13160 );
xor ( n13162 , n12855 , n12856 );
xor ( n13163 , n13162 , n12858 );
xor ( n13164 , n12878 , n12885 );
and ( n13165 , n13163 , n13164 );
and ( n13166 , n1995 , n4362 );
and ( n13167 , n4367 , n1990 );
and ( n13168 , n13166 , n13167 );
and ( n13169 , n2048 , n4161 );
and ( n13170 , n4150 , n2059 );
and ( n13171 , n13169 , n13170 );
and ( n13172 , n13168 , n13171 );
and ( n13173 , n3833 , n5077 );
and ( n13174 , n13171 , n13173 );
and ( n13175 , n13168 , n13173 );
or ( n13176 , n13172 , n13174 , n13175 );
and ( n13177 , n13164 , n13176 );
and ( n13178 , n13163 , n13176 );
or ( n13179 , n13165 , n13177 , n13178 );
and ( n13180 , n13160 , n13179 );
and ( n13181 , n13141 , n13179 );
or ( n13182 , n13161 , n13180 , n13181 );
and ( n13183 , n13122 , n13182 );
and ( n13184 , n13112 , n13182 );
or ( n13185 , n13123 , n13183 , n13184 );
and ( n13186 , n13111 , n13185 );
and ( n13187 , n2255 , n3903 );
and ( n13188 , n3892 , n2250 );
and ( n13189 , n13187 , n13188 );
and ( n13190 , n2591 , n3288 );
and ( n13191 , n3293 , n2586 );
and ( n13192 , n13190 , n13191 );
and ( n13193 , n13189 , n13192 );
and ( n13194 , n3169 , n12900 );
and ( n13195 , n13192 , n13194 );
and ( n13196 , n13189 , n13194 );
or ( n13197 , n13193 , n13195 , n13196 );
xor ( n13198 , n12872 , n12873 );
xor ( n13199 , n13198 , n12875 );
xor ( n13200 , n12879 , n12880 );
xor ( n13201 , n13200 , n12882 );
and ( n13202 , n13199 , n13201 );
and ( n13203 , n13197 , n13202 );
xnor ( n13204 , n12942 , n12943 );
xor ( n13205 , n12890 , n12891 );
and ( n13206 , n13204 , n13205 );
xor ( n13207 , n12786 , n12787 );
and ( n13208 , n13205 , n13207 );
and ( n13209 , n13204 , n13207 );
or ( n13210 , n13206 , n13208 , n13209 );
and ( n13211 , n13202 , n13210 );
and ( n13212 , n13197 , n13210 );
or ( n13213 , n13203 , n13211 , n13212 );
xor ( n13214 , n12946 , n12947 );
xor ( n13215 , n12853 , n12854 );
and ( n13216 , n13214 , n13215 );
xor ( n13217 , n12862 , n12863 );
and ( n13218 , n13215 , n13217 );
and ( n13219 , n13214 , n13217 );
or ( n13220 , n13216 , n13218 , n13219 );
xor ( n13221 , n12795 , n12796 );
and ( n13222 , n1911 , n4734 );
and ( n13223 , n2723 , n3146 );
or ( n13224 , n13222 , n13223 );
and ( n13225 , n13221 , n13224 );
xor ( n13226 , n12959 , n12960 );
xor ( n13227 , n13226 , n12965 );
and ( n13228 , n13224 , n13227 );
and ( n13229 , n13221 , n13227 );
or ( n13230 , n13225 , n13228 , n13229 );
and ( n13231 , n13220 , n13230 );
xor ( n13232 , n12901 , n12902 );
xor ( n13233 , n13232 , n12904 );
and ( n13234 , n13230 , n13233 );
and ( n13235 , n13220 , n13233 );
or ( n13236 , n13231 , n13234 , n13235 );
and ( n13237 , n13213 , n13236 );
xor ( n13238 , n12909 , n12910 );
xor ( n13239 , n13238 , n12912 );
xor ( n13240 , n12920 , n12921 );
xor ( n13241 , n13240 , n12923 );
and ( n13242 , n13239 , n13241 );
xor ( n13243 , n12927 , n12928 );
xor ( n13244 , n13243 , n12930 );
and ( n13245 , n13241 , n13244 );
and ( n13246 , n13239 , n13244 );
or ( n13247 , n13242 , n13245 , n13246 );
and ( n13248 , n13236 , n13247 );
and ( n13249 , n13213 , n13247 );
or ( n13250 , n13237 , n13248 , n13249 );
xor ( n13251 , n12898 , n12907 );
xor ( n13252 , n13251 , n12915 );
xor ( n13253 , n12926 , n12933 );
xor ( n13254 , n13253 , n12951 );
and ( n13255 , n13252 , n13254 );
xor ( n13256 , n12981 , n12983 );
xor ( n13257 , n13256 , n12986 );
and ( n13258 , n13254 , n13257 );
and ( n13259 , n13252 , n13257 );
or ( n13260 , n13255 , n13258 , n13259 );
and ( n13261 , n13250 , n13260 );
xor ( n13262 , n12844 , n12846 );
xor ( n13263 , n13262 , n12849 );
and ( n13264 , n13260 , n13263 );
and ( n13265 , n13250 , n13263 );
or ( n13266 , n13261 , n13264 , n13265 );
and ( n13267 , n13185 , n13266 );
and ( n13268 , n13111 , n13266 );
or ( n13269 , n13186 , n13267 , n13268 );
and ( n13270 , n13089 , n13269 );
and ( n13271 , n13087 , n13269 );
or ( n13272 , n13090 , n13270 , n13271 );
xor ( n13273 , n12889 , n12918 );
xor ( n13274 , n13273 , n12954 );
xor ( n13275 , n12989 , n12999 );
xor ( n13276 , n13275 , n13002 );
and ( n13277 , n13274 , n13276 );
xor ( n13278 , n13011 , n13013 );
xor ( n13279 , n13278 , n13016 );
and ( n13280 , n13276 , n13279 );
and ( n13281 , n13274 , n13279 );
or ( n13282 , n13277 , n13280 , n13281 );
xor ( n13283 , n12785 , n12825 );
xor ( n13284 , n13283 , n12839 );
and ( n13285 , n13282 , n13284 );
xor ( n13286 , n12852 , n12957 );
xor ( n13287 , n13286 , n13005 );
and ( n13288 , n13284 , n13287 );
and ( n13289 , n13282 , n13287 );
or ( n13290 , n13285 , n13288 , n13289 );
xor ( n13291 , n12842 , n13008 );
xor ( n13292 , n13291 , n13027 );
and ( n13293 , n13290 , n13292 );
xor ( n13294 , n13041 , n13043 );
xor ( n13295 , n13294 , n13046 );
and ( n13296 , n13292 , n13295 );
and ( n13297 , n13290 , n13295 );
or ( n13298 , n13293 , n13296 , n13297 );
and ( n13299 , n13272 , n13298 );
xor ( n13300 , n12783 , n13030 );
xor ( n13301 , n13300 , n13049 );
and ( n13302 , n13298 , n13301 );
and ( n13303 , n13272 , n13301 );
or ( n13304 , n13299 , n13302 , n13303 );
and ( n13305 , n13085 , n13304 );
xor ( n13306 , n13052 , n13062 );
xor ( n13307 , n13306 , n13065 );
and ( n13308 , n13304 , n13307 );
and ( n13309 , n13085 , n13307 );
or ( n13310 , n13305 , n13308 , n13309 );
and ( n13311 , n13083 , n13310 );
xor ( n13312 , n12778 , n12780 );
xor ( n13313 , n13312 , n13068 );
and ( n13314 , n13310 , n13313 );
and ( n13315 , n13083 , n13313 );
or ( n13316 , n13311 , n13314 , n13315 );
xor ( n13317 , n12776 , n13071 );
xor ( n13318 , n13317 , n13074 );
and ( n13319 , n13316 , n13318 );
xor ( n13320 , n13316 , n13318 );
xor ( n13321 , n13083 , n13310 );
xor ( n13322 , n13321 , n13313 );
xor ( n13323 , n13054 , n13056 );
xor ( n13324 , n13323 , n13059 );
xor ( n13325 , n13019 , n13021 );
xor ( n13326 , n13325 , n13024 );
xor ( n13327 , n13033 , n13035 );
xor ( n13328 , n13327 , n13038 );
and ( n13329 , n13326 , n13328 );
xor ( n13330 , n12991 , n12993 );
xor ( n13331 , n13330 , n12996 );
xor ( n13332 , n13105 , n13107 );
and ( n13333 , n13331 , n13332 );
xor ( n13334 , n12941 , n12944 );
xor ( n13335 , n13334 , n12948 );
xor ( n13336 , n12968 , n12975 );
xor ( n13337 , n13336 , n12978 );
and ( n13338 , n13335 , n13337 );
xor ( n13339 , n13096 , n13098 );
xor ( n13340 , n13339 , n13101 );
and ( n13341 , n13337 , n13340 );
and ( n13342 , n13335 , n13340 );
or ( n13343 , n13338 , n13341 , n13342 );
and ( n13344 , n13332 , n13343 );
and ( n13345 , n13331 , n13343 );
or ( n13346 , n13333 , n13344 , n13345 );
xor ( n13347 , n13138 , n13140 );
xor ( n13348 , n13150 , n13159 );
and ( n13349 , n13347 , n13348 );
and ( n13350 , n2591 , n3449 );
and ( n13351 , n3454 , n2586 );
and ( n13352 , n13350 , n13351 );
and ( n13353 , n4721 , n3627 );
and ( n13354 , n13352 , n13353 );
and ( n13355 , n3645 , n11777 );
and ( n13356 , n13353 , n13355 );
and ( n13357 , n13352 , n13355 );
or ( n13358 , n13354 , n13356 , n13357 );
and ( n13359 , n4579 , n3929 );
and ( n13360 , n4385 , n4522 );
and ( n13361 , n13359 , n13360 );
and ( n13362 , n4138 , n5077 );
and ( n13363 , n13360 , n13362 );
and ( n13364 , n13359 , n13362 );
or ( n13365 , n13361 , n13363 , n13364 );
and ( n13366 , n13358 , n13365 );
and ( n13367 , n4150 , n2250 );
and ( n13368 , n3728 , n2492 );
and ( n13369 , n13367 , n13368 );
and ( n13370 , n3151 , n2923 );
and ( n13371 , n13368 , n13370 );
and ( n13372 , n13367 , n13370 );
or ( n13373 , n13369 , n13371 , n13372 );
and ( n13374 , n2255 , n4161 );
and ( n13375 , n2497 , n3739 );
and ( n13376 , n13374 , n13375 );
and ( n13377 , n2928 , n3146 );
and ( n13378 , n13375 , n13377 );
and ( n13379 , n13374 , n13377 );
or ( n13380 , n13376 , n13378 , n13379 );
and ( n13381 , n13373 , n13380 );
and ( n13382 , n13365 , n13381 );
and ( n13383 , n13358 , n13381 );
or ( n13384 , n13366 , n13382 , n13383 );
and ( n13385 , n13348 , n13384 );
and ( n13386 , n13347 , n13384 );
or ( n13387 , n13349 , n13385 , n13386 );
and ( n13388 , n1778 , n5086 );
and ( n13389 , n5091 , n1789 );
and ( n13390 , n13388 , n13389 );
and ( n13391 , n3833 , n11156 );
and ( n13392 , n13390 , n13391 );
and ( n13393 , n3339 , n12290 );
and ( n13394 , n13391 , n13393 );
and ( n13395 , n13390 , n13393 );
or ( n13396 , n13392 , n13394 , n13395 );
and ( n13397 , n1694 , n11111 );
and ( n13398 , n11116 , n1689 );
and ( n13399 , n13397 , n13398 );
and ( n13400 , n1911 , n4982 );
and ( n13401 , n4989 , n1906 );
and ( n13402 , n13400 , n13401 );
and ( n13403 , n13399 , n13402 );
and ( n13404 , n5177 , n3301 );
and ( n13405 , n13402 , n13404 );
and ( n13406 , n13399 , n13404 );
or ( n13407 , n13403 , n13405 , n13406 );
and ( n13408 , n13396 , n13407 );
buf ( n13409 , n2928 );
xor ( n13410 , n10021 , n10612 );
buf ( n13411 , n13410 );
buf ( n13412 , n13411 );
buf ( n13413 , n13412 );
and ( n13414 , n13409 , n13413 );
buf ( n13415 , n2937 );
and ( n13416 , n13413 , n13415 );
and ( n13417 , n13409 , n13415 );
or ( n13418 , n13414 , n13416 , n13417 );
and ( n13419 , n13407 , n13418 );
and ( n13420 , n13396 , n13418 );
or ( n13421 , n13408 , n13419 , n13420 );
xor ( n13422 , n13189 , n13192 );
xor ( n13423 , n13422 , n13194 );
xor ( n13424 , n12935 , n12936 );
xor ( n13425 , n13424 , n12938 );
and ( n13426 , n13423 , n13425 );
and ( n13427 , n13421 , n13426 );
xor ( n13428 , n13144 , n13145 );
xor ( n13429 , n13428 , n13147 );
xor ( n13430 , n13153 , n13154 );
xor ( n13431 , n13430 , n13156 );
and ( n13432 , n13429 , n13431 );
and ( n13433 , n13426 , n13432 );
and ( n13434 , n13421 , n13432 );
or ( n13435 , n13427 , n13433 , n13434 );
and ( n13436 , n13387 , n13435 );
xor ( n13437 , n12969 , n12970 );
xor ( n13438 , n13437 , n12972 );
xor ( n13439 , n13168 , n13171 );
xor ( n13440 , n13439 , n13173 );
and ( n13441 , n13438 , n13440 );
xor ( n13442 , n13130 , n13137 );
and ( n13443 , n13440 , n13442 );
and ( n13444 , n13438 , n13442 );
or ( n13445 , n13441 , n13443 , n13444 );
xor ( n13446 , n13199 , n13201 );
and ( n13447 , n1724 , n10869 );
and ( n13448 , n10862 , n1719 );
and ( n13449 , n13447 , n13448 );
and ( n13450 , n10933 , n2577 );
and ( n13451 , n13449 , n13450 );
and ( n13452 , n10886 , n2948 );
and ( n13453 , n13450 , n13452 );
and ( n13454 , n13449 , n13452 );
or ( n13455 , n13451 , n13453 , n13454 );
and ( n13456 , n13446 , n13455 );
and ( n13457 , n2309 , n3903 );
and ( n13458 , n3892 , n2304 );
and ( n13459 , n13457 , n13458 );
and ( n13460 , n2723 , n3288 );
and ( n13461 , n3293 , n2718 );
and ( n13462 , n13460 , n13461 );
and ( n13463 , n13459 , n13462 );
buf ( n13464 , n2935 );
buf ( n13465 , n13464 );
and ( n13466 , n3169 , n13465 );
and ( n13467 , n13462 , n13466 );
and ( n13468 , n13459 , n13466 );
or ( n13469 , n13463 , n13467 , n13468 );
and ( n13470 , n13455 , n13469 );
and ( n13471 , n13446 , n13469 );
or ( n13472 , n13456 , n13470 , n13471 );
and ( n13473 , n13445 , n13472 );
xor ( n13474 , n13124 , n13125 );
xor ( n13475 , n13474 , n13127 );
xor ( n13476 , n13131 , n13132 );
xor ( n13477 , n13476 , n13134 );
and ( n13478 , n13475 , n13477 );
and ( n13479 , n4739 , n1906 );
and ( n13480 , n3151 , n2718 );
and ( n13481 , n13479 , n13480 );
xor ( n13482 , n13359 , n13360 );
xor ( n13483 , n13482 , n13362 );
and ( n13484 , n13480 , n13483 );
and ( n13485 , n13479 , n13483 );
or ( n13486 , n13481 , n13484 , n13485 );
and ( n13487 , n13478 , n13486 );
xnor ( n13488 , n13222 , n13223 );
xor ( n13489 , n13151 , n13152 );
and ( n13490 , n13488 , n13489 );
xor ( n13491 , n13166 , n13167 );
and ( n13492 , n13489 , n13491 );
and ( n13493 , n13488 , n13491 );
or ( n13494 , n13490 , n13492 , n13493 );
and ( n13495 , n13486 , n13494 );
and ( n13496 , n13478 , n13494 );
or ( n13497 , n13487 , n13495 , n13496 );
and ( n13498 , n13472 , n13497 );
and ( n13499 , n13445 , n13497 );
or ( n13500 , n13473 , n13498 , n13499 );
and ( n13501 , n13435 , n13500 );
and ( n13502 , n13387 , n13500 );
or ( n13503 , n13436 , n13501 , n13502 );
and ( n13504 , n13346 , n13503 );
xor ( n13505 , n13169 , n13170 );
xor ( n13506 , n13187 , n13188 );
and ( n13507 , n13505 , n13506 );
xor ( n13508 , n13142 , n13143 );
and ( n13509 , n13506 , n13508 );
and ( n13510 , n13505 , n13508 );
or ( n13511 , n13507 , n13509 , n13510 );
xor ( n13512 , n13190 , n13191 );
and ( n13513 , n1995 , n4734 );
and ( n13514 , n4739 , n1990 );
and ( n13515 , n13513 , n13514 );
and ( n13516 , n13512 , n13515 );
and ( n13517 , n2048 , n4362 );
and ( n13518 , n4367 , n2059 );
and ( n13519 , n13517 , n13518 );
and ( n13520 , n13515 , n13519 );
and ( n13521 , n13512 , n13519 );
or ( n13522 , n13516 , n13520 , n13521 );
and ( n13523 , n13511 , n13522 );
xor ( n13524 , n13204 , n13205 );
xor ( n13525 , n13524 , n13207 );
and ( n13526 , n13522 , n13525 );
and ( n13527 , n13511 , n13525 );
or ( n13528 , n13523 , n13526 , n13527 );
xor ( n13529 , n13163 , n13164 );
xor ( n13530 , n13529 , n13176 );
and ( n13531 , n13528 , n13530 );
xor ( n13532 , n13197 , n13202 );
xor ( n13533 , n13532 , n13210 );
and ( n13534 , n13530 , n13533 );
and ( n13535 , n13528 , n13533 );
or ( n13536 , n13531 , n13534 , n13535 );
xor ( n13537 , n13114 , n13116 );
xor ( n13538 , n13537 , n13119 );
and ( n13539 , n13536 , n13538 );
xor ( n13540 , n13141 , n13160 );
xor ( n13541 , n13540 , n13179 );
and ( n13542 , n13538 , n13541 );
and ( n13543 , n13536 , n13541 );
or ( n13544 , n13539 , n13542 , n13543 );
and ( n13545 , n13503 , n13544 );
and ( n13546 , n13346 , n13544 );
or ( n13547 , n13504 , n13545 , n13546 );
and ( n13548 , n13328 , n13547 );
and ( n13549 , n13326 , n13547 );
or ( n13550 , n13329 , n13548 , n13549 );
xor ( n13551 , n13092 , n13093 );
xor ( n13552 , n13551 , n13108 );
xor ( n13553 , n13112 , n13122 );
xor ( n13554 , n13553 , n13182 );
and ( n13555 , n13552 , n13554 );
xor ( n13556 , n13250 , n13260 );
xor ( n13557 , n13556 , n13263 );
and ( n13558 , n13554 , n13557 );
and ( n13559 , n13552 , n13557 );
or ( n13560 , n13555 , n13558 , n13559 );
xor ( n13561 , n13111 , n13185 );
xor ( n13562 , n13561 , n13266 );
and ( n13563 , n13560 , n13562 );
xor ( n13564 , n13282 , n13284 );
xor ( n13565 , n13564 , n13287 );
and ( n13566 , n13562 , n13565 );
and ( n13567 , n13560 , n13565 );
or ( n13568 , n13563 , n13566 , n13567 );
and ( n13569 , n13550 , n13568 );
xor ( n13570 , n13087 , n13089 );
xor ( n13571 , n13570 , n13269 );
and ( n13572 , n13568 , n13571 );
and ( n13573 , n13550 , n13571 );
or ( n13574 , n13569 , n13572 , n13573 );
and ( n13575 , n13324 , n13574 );
xor ( n13576 , n13272 , n13298 );
xor ( n13577 , n13576 , n13301 );
and ( n13578 , n13574 , n13577 );
and ( n13579 , n13324 , n13577 );
or ( n13580 , n13575 , n13578 , n13579 );
xor ( n13581 , n13085 , n13304 );
xor ( n13582 , n13581 , n13307 );
and ( n13583 , n13580 , n13582 );
xor ( n13584 , n13580 , n13582 );
xor ( n13585 , n13290 , n13292 );
xor ( n13586 , n13585 , n13295 );
xor ( n13587 , n13274 , n13276 );
xor ( n13588 , n13587 , n13279 );
xor ( n13589 , n13213 , n13236 );
xor ( n13590 , n13589 , n13247 );
xor ( n13591 , n13252 , n13254 );
xor ( n13592 , n13591 , n13257 );
and ( n13593 , n13590 , n13592 );
xor ( n13594 , n13220 , n13230 );
xor ( n13595 , n13594 , n13233 );
xor ( n13596 , n13239 , n13241 );
xor ( n13597 , n13596 , n13244 );
and ( n13598 , n13595 , n13597 );
xor ( n13599 , n13214 , n13215 );
xor ( n13600 , n13599 , n13217 );
xor ( n13601 , n13221 , n13224 );
xor ( n13602 , n13601 , n13227 );
and ( n13603 , n13600 , n13602 );
xor ( n13604 , n13358 , n13365 );
xor ( n13605 , n13604 , n13381 );
and ( n13606 , n13602 , n13605 );
and ( n13607 , n13600 , n13605 );
or ( n13608 , n13603 , n13606 , n13607 );
and ( n13609 , n13597 , n13608 );
and ( n13610 , n13595 , n13608 );
or ( n13611 , n13598 , n13609 , n13610 );
and ( n13612 , n13592 , n13611 );
and ( n13613 , n13590 , n13611 );
or ( n13614 , n13593 , n13612 , n13613 );
and ( n13615 , n13588 , n13614 );
xor ( n13616 , n13396 , n13407 );
xor ( n13617 , n13616 , n13418 );
xor ( n13618 , n13423 , n13425 );
and ( n13619 , n13617 , n13618 );
xor ( n13620 , n13429 , n13431 );
and ( n13621 , n13618 , n13620 );
and ( n13622 , n13617 , n13620 );
or ( n13623 , n13619 , n13621 , n13622 );
and ( n13624 , n2255 , n4362 );
and ( n13625 , n4367 , n2250 );
and ( n13626 , n13624 , n13625 );
and ( n13627 , n4138 , n11156 );
and ( n13628 , n13626 , n13627 );
and ( n13629 , n3339 , n12900 );
and ( n13630 , n13627 , n13629 );
and ( n13631 , n13626 , n13629 );
or ( n13632 , n13628 , n13630 , n13631 );
and ( n13633 , n10933 , n2948 );
and ( n13634 , n4579 , n4522 );
and ( n13635 , n13633 , n13634 );
and ( n13636 , n3645 , n12290 );
and ( n13637 , n13634 , n13636 );
and ( n13638 , n13633 , n13636 );
or ( n13639 , n13635 , n13637 , n13638 );
and ( n13640 , n13632 , n13639 );
and ( n13641 , n3246 , n12900 );
and ( n13642 , n13639 , n13641 );
and ( n13643 , n13632 , n13641 );
or ( n13644 , n13640 , n13642 , n13643 );
and ( n13645 , n2309 , n4161 );
and ( n13646 , n4150 , n2304 );
and ( n13647 , n13645 , n13646 );
and ( n13648 , n2591 , n3739 );
and ( n13649 , n3728 , n2586 );
and ( n13650 , n13648 , n13649 );
and ( n13651 , n13647 , n13650 );
and ( n13652 , n3833 , n11777 );
and ( n13653 , n13650 , n13652 );
and ( n13654 , n13647 , n13652 );
or ( n13655 , n13651 , n13653 , n13654 );
and ( n13656 , n1778 , n10869 );
and ( n13657 , n10862 , n1789 );
and ( n13658 , n13656 , n13657 );
and ( n13659 , n2497 , n3903 );
and ( n13660 , n3892 , n2492 );
and ( n13661 , n13659 , n13660 );
and ( n13662 , n13658 , n13661 );
and ( n13663 , n3246 , n13465 );
and ( n13664 , n13661 , n13663 );
and ( n13665 , n13658 , n13663 );
or ( n13666 , n13662 , n13664 , n13665 );
and ( n13667 , n13655 , n13666 );
xor ( n13668 , n13409 , n13413 );
xor ( n13669 , n13668 , n13415 );
and ( n13670 , n13666 , n13669 );
and ( n13671 , n13655 , n13669 );
or ( n13672 , n13667 , n13670 , n13671 );
and ( n13673 , n13644 , n13672 );
xor ( n13674 , n13459 , n13462 );
xor ( n13675 , n13674 , n13466 );
xor ( n13676 , n13352 , n13353 );
xor ( n13677 , n13676 , n13355 );
and ( n13678 , n13675 , n13677 );
xor ( n13679 , n13390 , n13391 );
xor ( n13680 , n13679 , n13393 );
and ( n13681 , n13677 , n13680 );
and ( n13682 , n13675 , n13680 );
or ( n13683 , n13678 , n13681 , n13682 );
and ( n13684 , n13672 , n13683 );
and ( n13685 , n13644 , n13683 );
or ( n13686 , n13673 , n13684 , n13685 );
and ( n13687 , n13623 , n13686 );
xor ( n13688 , n10024 , n10610 );
buf ( n13689 , n13688 );
buf ( n13690 , n13689 );
buf ( n13691 , n13690 );
and ( n13692 , n10886 , n3301 );
and ( n13693 , n13691 , n13692 );
and ( n13694 , n4721 , n3929 );
and ( n13695 , n13692 , n13694 );
and ( n13696 , n13691 , n13694 );
or ( n13697 , n13693 , n13695 , n13696 );
xor ( n13698 , n13449 , n13450 );
xor ( n13699 , n13698 , n13452 );
and ( n13700 , n13697 , n13699 );
xor ( n13701 , n13399 , n13402 );
xor ( n13702 , n13701 , n13404 );
and ( n13703 , n13699 , n13702 );
and ( n13704 , n13697 , n13702 );
or ( n13705 , n13700 , n13703 , n13704 );
xor ( n13706 , n13373 , n13380 );
xor ( n13707 , n13475 , n13477 );
and ( n13708 , n13706 , n13707 );
and ( n13709 , n1724 , n11111 );
and ( n13710 , n11116 , n1719 );
and ( n13711 , n13709 , n13710 );
and ( n13712 , n5177 , n3627 );
and ( n13713 , n13711 , n13712 );
and ( n13714 , n4385 , n5077 );
and ( n13715 , n13712 , n13714 );
and ( n13716 , n13711 , n13714 );
or ( n13717 , n13713 , n13715 , n13716 );
and ( n13718 , n13707 , n13717 );
and ( n13719 , n13706 , n13717 );
or ( n13720 , n13708 , n13718 , n13719 );
and ( n13721 , n13705 , n13720 );
and ( n13722 , n5091 , n1906 );
and ( n13723 , n4989 , n1990 );
and ( n13724 , n13722 , n13723 );
and ( n13725 , n3454 , n2718 );
and ( n13726 , n13723 , n13725 );
and ( n13727 , n13722 , n13725 );
or ( n13728 , n13724 , n13726 , n13727 );
and ( n13729 , n1911 , n5086 );
and ( n13730 , n1995 , n4982 );
and ( n13731 , n13729 , n13730 );
and ( n13732 , n2723 , n3449 );
and ( n13733 , n13730 , n13732 );
and ( n13734 , n13729 , n13732 );
or ( n13735 , n13731 , n13733 , n13734 );
and ( n13736 , n13728 , n13735 );
xor ( n13737 , n13367 , n13368 );
xor ( n13738 , n13737 , n13370 );
xor ( n13739 , n13374 , n13375 );
xor ( n13740 , n13739 , n13377 );
and ( n13741 , n13738 , n13740 );
and ( n13742 , n13736 , n13741 );
xor ( n13743 , n13397 , n13398 );
xor ( n13744 , n13447 , n13448 );
and ( n13745 , n13743 , n13744 );
xor ( n13746 , n13388 , n13389 );
and ( n13747 , n13744 , n13746 );
and ( n13748 , n13743 , n13746 );
or ( n13749 , n13745 , n13747 , n13748 );
and ( n13750 , n13741 , n13749 );
and ( n13751 , n13736 , n13749 );
or ( n13752 , n13742 , n13750 , n13751 );
and ( n13753 , n13720 , n13752 );
and ( n13754 , n13705 , n13752 );
or ( n13755 , n13721 , n13753 , n13754 );
and ( n13756 , n13686 , n13755 );
and ( n13757 , n13623 , n13755 );
or ( n13758 , n13687 , n13756 , n13757 );
xor ( n13759 , n13400 , n13401 );
xor ( n13760 , n13513 , n13514 );
and ( n13761 , n13759 , n13760 );
xor ( n13762 , n13517 , n13518 );
and ( n13763 , n13760 , n13762 );
and ( n13764 , n13759 , n13762 );
or ( n13765 , n13761 , n13763 , n13764 );
xor ( n13766 , n13457 , n13458 );
xor ( n13767 , n13350 , n13351 );
and ( n13768 , n13766 , n13767 );
xor ( n13769 , n13460 , n13461 );
and ( n13770 , n13767 , n13769 );
and ( n13771 , n13766 , n13769 );
or ( n13772 , n13768 , n13770 , n13771 );
and ( n13773 , n13765 , n13772 );
and ( n13774 , n2048 , n4734 );
and ( n13775 , n2928 , n3288 );
or ( n13776 , n13774 , n13775 );
and ( n13777 , n4739 , n2059 );
and ( n13778 , n3293 , n2923 );
and ( n13779 , n13777 , n13778 );
xor ( n13780 , n10025 , n10609 );
buf ( n13781 , n13780 );
buf ( n13782 , n13781 );
buf ( n13783 , n13782 );
and ( n13784 , n13778 , n13783 );
and ( n13785 , n13777 , n13783 );
or ( n13786 , n13779 , n13784 , n13785 );
and ( n13787 , n13776 , n13786 );
xor ( n13788 , n13691 , n13692 );
xor ( n13789 , n13788 , n13694 );
and ( n13790 , n13786 , n13789 );
and ( n13791 , n13776 , n13789 );
or ( n13792 , n13787 , n13790 , n13791 );
and ( n13793 , n13772 , n13792 );
and ( n13794 , n13765 , n13792 );
or ( n13795 , n13773 , n13793 , n13794 );
xor ( n13796 , n13479 , n13480 );
xor ( n13797 , n13796 , n13483 );
xor ( n13798 , n13488 , n13489 );
xor ( n13799 , n13798 , n13491 );
and ( n13800 , n13797 , n13799 );
xor ( n13801 , n13505 , n13506 );
xor ( n13802 , n13801 , n13508 );
and ( n13803 , n13799 , n13802 );
and ( n13804 , n13797 , n13802 );
or ( n13805 , n13800 , n13803 , n13804 );
and ( n13806 , n13795 , n13805 );
xor ( n13807 , n13438 , n13440 );
xor ( n13808 , n13807 , n13442 );
and ( n13809 , n13805 , n13808 );
and ( n13810 , n13795 , n13808 );
or ( n13811 , n13806 , n13809 , n13810 );
xor ( n13812 , n13446 , n13455 );
xor ( n13813 , n13812 , n13469 );
xor ( n13814 , n13478 , n13486 );
xor ( n13815 , n13814 , n13494 );
and ( n13816 , n13813 , n13815 );
xor ( n13817 , n13511 , n13522 );
xor ( n13818 , n13817 , n13525 );
and ( n13819 , n13815 , n13818 );
and ( n13820 , n13813 , n13818 );
or ( n13821 , n13816 , n13819 , n13820 );
and ( n13822 , n13811 , n13821 );
xor ( n13823 , n13335 , n13337 );
xor ( n13824 , n13823 , n13340 );
and ( n13825 , n13821 , n13824 );
and ( n13826 , n13811 , n13824 );
or ( n13827 , n13822 , n13825 , n13826 );
and ( n13828 , n13758 , n13827 );
xor ( n13829 , n13347 , n13348 );
xor ( n13830 , n13829 , n13384 );
xor ( n13831 , n13421 , n13426 );
xor ( n13832 , n13831 , n13432 );
and ( n13833 , n13830 , n13832 );
xor ( n13834 , n13445 , n13472 );
xor ( n13835 , n13834 , n13497 );
and ( n13836 , n13832 , n13835 );
and ( n13837 , n13830 , n13835 );
or ( n13838 , n13833 , n13836 , n13837 );
and ( n13839 , n13827 , n13838 );
and ( n13840 , n13758 , n13838 );
or ( n13841 , n13828 , n13839 , n13840 );
and ( n13842 , n13614 , n13841 );
and ( n13843 , n13588 , n13841 );
or ( n13844 , n13615 , n13842 , n13843 );
xor ( n13845 , n13331 , n13332 );
xor ( n13846 , n13845 , n13343 );
xor ( n13847 , n13387 , n13435 );
xor ( n13848 , n13847 , n13500 );
and ( n13849 , n13846 , n13848 );
xor ( n13850 , n13536 , n13538 );
xor ( n13851 , n13850 , n13541 );
and ( n13852 , n13848 , n13851 );
and ( n13853 , n13846 , n13851 );
or ( n13854 , n13849 , n13852 , n13853 );
xor ( n13855 , n13346 , n13503 );
xor ( n13856 , n13855 , n13544 );
and ( n13857 , n13854 , n13856 );
xor ( n13858 , n13552 , n13554 );
xor ( n13859 , n13858 , n13557 );
and ( n13860 , n13856 , n13859 );
and ( n13861 , n13854 , n13859 );
or ( n13862 , n13857 , n13860 , n13861 );
and ( n13863 , n13844 , n13862 );
xor ( n13864 , n13326 , n13328 );
xor ( n13865 , n13864 , n13547 );
and ( n13866 , n13862 , n13865 );
and ( n13867 , n13844 , n13865 );
or ( n13868 , n13863 , n13866 , n13867 );
and ( n13869 , n13586 , n13868 );
xor ( n13870 , n13550 , n13568 );
xor ( n13871 , n13870 , n13571 );
and ( n13872 , n13868 , n13871 );
and ( n13873 , n13586 , n13871 );
or ( n13874 , n13869 , n13872 , n13873 );
xor ( n13875 , n13324 , n13574 );
xor ( n13876 , n13875 , n13577 );
and ( n13877 , n13874 , n13876 );
xor ( n13878 , n13874 , n13876 );
xor ( n13879 , n13560 , n13562 );
xor ( n13880 , n13879 , n13565 );
xor ( n13881 , n13528 , n13530 );
xor ( n13882 , n13881 , n13533 );
and ( n13883 , n2591 , n3903 );
and ( n13884 , n3892 , n2586 );
and ( n13885 , n13883 , n13884 );
and ( n13886 , n10886 , n3627 );
and ( n13887 , n13885 , n13886 );
buf ( n13888 , n3167 );
buf ( n13889 , n13888 );
and ( n13890 , n3246 , n13889 );
and ( n13891 , n13886 , n13890 );
and ( n13892 , n13885 , n13890 );
or ( n13893 , n13887 , n13891 , n13892 );
and ( n13894 , n1911 , n10869 );
and ( n13895 , n10862 , n1906 );
and ( n13896 , n13894 , n13895 );
and ( n13897 , n1995 , n5086 );
and ( n13898 , n5091 , n1990 );
and ( n13899 , n13897 , n13898 );
and ( n13900 , n13896 , n13899 );
and ( n13901 , n4138 , n11777 );
and ( n13902 , n13899 , n13901 );
and ( n13903 , n13896 , n13901 );
or ( n13904 , n13900 , n13902 , n13903 );
and ( n13905 , n13893 , n13904 );
and ( n13906 , n2048 , n4982 );
and ( n13907 , n4989 , n2059 );
and ( n13908 , n13906 , n13907 );
and ( n13909 , n4579 , n5077 );
and ( n13910 , n13908 , n13909 );
and ( n13911 , n3645 , n12900 );
and ( n13912 , n13909 , n13911 );
and ( n13913 , n13908 , n13911 );
or ( n13914 , n13910 , n13912 , n13913 );
and ( n13915 , n13904 , n13914 );
and ( n13916 , n13893 , n13914 );
or ( n13917 , n13905 , n13915 , n13916 );
and ( n13918 , n3151 , n3288 );
and ( n13919 , n3293 , n3146 );
and ( n13920 , n13918 , n13919 );
and ( n13921 , n5177 , n3929 );
and ( n13922 , n13920 , n13921 );
and ( n13923 , n4385 , n11156 );
and ( n13924 , n13921 , n13923 );
and ( n13925 , n13920 , n13923 );
or ( n13926 , n13922 , n13924 , n13925 );
and ( n13927 , n2255 , n4734 );
and ( n13928 , n4739 , n2250 );
and ( n13929 , n13927 , n13928 );
and ( n13930 , n2928 , n3449 );
and ( n13931 , n3454 , n2923 );
and ( n13932 , n13930 , n13931 );
and ( n13933 , n13929 , n13932 );
and ( n13934 , n3339 , n13465 );
and ( n13935 , n13932 , n13934 );
and ( n13936 , n13929 , n13934 );
or ( n13937 , n13933 , n13935 , n13936 );
and ( n13938 , n13926 , n13937 );
and ( n13939 , n1778 , n11111 );
and ( n13940 , n11116 , n1789 );
and ( n13941 , n13939 , n13940 );
and ( n13942 , n2497 , n4161 );
and ( n13943 , n4150 , n2492 );
and ( n13944 , n13942 , n13943 );
and ( n13945 , n13941 , n13944 );
and ( n13946 , n3833 , n12290 );
and ( n13947 , n13944 , n13946 );
and ( n13948 , n13941 , n13946 );
or ( n13949 , n13945 , n13947 , n13948 );
and ( n13950 , n13937 , n13949 );
and ( n13951 , n13926 , n13949 );
or ( n13952 , n13938 , n13950 , n13951 );
and ( n13953 , n13917 , n13952 );
xor ( n13954 , n13512 , n13515 );
xor ( n13955 , n13954 , n13519 );
xor ( n13956 , n13632 , n13639 );
xor ( n13957 , n13956 , n13641 );
and ( n13958 , n13955 , n13957 );
xor ( n13959 , n13655 , n13666 );
xor ( n13960 , n13959 , n13669 );
and ( n13961 , n13957 , n13960 );
and ( n13962 , n13955 , n13960 );
or ( n13963 , n13958 , n13961 , n13962 );
and ( n13964 , n13953 , n13963 );
xor ( n13965 , n13675 , n13677 );
xor ( n13966 , n13965 , n13680 );
xor ( n13967 , n13626 , n13627 );
xor ( n13968 , n13967 , n13629 );
xor ( n13969 , n13633 , n13634 );
xor ( n13970 , n13969 , n13636 );
and ( n13971 , n13968 , n13970 );
xor ( n13972 , n13711 , n13712 );
xor ( n13973 , n13972 , n13714 );
and ( n13974 , n13970 , n13973 );
and ( n13975 , n13968 , n13973 );
or ( n13976 , n13971 , n13974 , n13975 );
and ( n13977 , n13966 , n13976 );
xor ( n13978 , n13647 , n13650 );
xor ( n13979 , n13978 , n13652 );
xor ( n13980 , n13658 , n13661 );
xor ( n13981 , n13980 , n13663 );
or ( n13982 , n13979 , n13981 );
and ( n13983 , n13976 , n13982 );
and ( n13984 , n13966 , n13982 );
or ( n13985 , n13977 , n13983 , n13984 );
and ( n13986 , n13963 , n13985 );
and ( n13987 , n13953 , n13985 );
or ( n13988 , n13964 , n13986 , n13987 );
and ( n13989 , n13882 , n13988 );
xor ( n13990 , n13728 , n13735 );
xor ( n13991 , n13738 , n13740 );
and ( n13992 , n13990 , n13991 );
and ( n13993 , n2309 , n4362 );
and ( n13994 , n4367 , n2304 );
and ( n13995 , n13993 , n13994 );
buf ( n13996 , n3151 );
and ( n13997 , n13995 , n13996 );
and ( n13998 , n4721 , n4522 );
and ( n13999 , n13996 , n13998 );
and ( n14000 , n13995 , n13998 );
or ( n14001 , n13997 , n13999 , n14000 );
and ( n14002 , n13991 , n14001 );
and ( n14003 , n13990 , n14001 );
or ( n14004 , n13992 , n14002 , n14003 );
buf ( n14005 , n3169 );
xnor ( n14006 , n13774 , n13775 );
and ( n14007 , n14005 , n14006 );
xor ( n14008 , n13709 , n13710 );
and ( n14009 , n14006 , n14008 );
and ( n14010 , n14005 , n14008 );
or ( n14011 , n14007 , n14009 , n14010 );
xor ( n14012 , n13656 , n13657 );
xor ( n14013 , n13624 , n13625 );
and ( n14014 , n14012 , n14013 );
xor ( n14015 , n13645 , n13646 );
and ( n14016 , n14013 , n14015 );
and ( n14017 , n14012 , n14015 );
or ( n14018 , n14014 , n14016 , n14017 );
and ( n14019 , n14011 , n14018 );
xor ( n14020 , n13659 , n13660 );
xor ( n14021 , n13648 , n13649 );
and ( n14022 , n14020 , n14021 );
xor ( n14023 , n13777 , n13778 );
xor ( n14024 , n14023 , n13783 );
and ( n14025 , n14021 , n14024 );
and ( n14026 , n14020 , n14024 );
or ( n14027 , n14022 , n14025 , n14026 );
and ( n14028 , n14018 , n14027 );
and ( n14029 , n14011 , n14027 );
or ( n14030 , n14019 , n14028 , n14029 );
and ( n14031 , n14004 , n14030 );
xor ( n14032 , n13743 , n13744 );
xor ( n14033 , n14032 , n13746 );
xor ( n14034 , n13759 , n13760 );
xor ( n14035 , n14034 , n13762 );
and ( n14036 , n14033 , n14035 );
xor ( n14037 , n13766 , n13767 );
xor ( n14038 , n14037 , n13769 );
and ( n14039 , n14035 , n14038 );
and ( n14040 , n14033 , n14038 );
or ( n14041 , n14036 , n14039 , n14040 );
and ( n14042 , n14030 , n14041 );
and ( n14043 , n14004 , n14041 );
or ( n14044 , n14031 , n14042 , n14043 );
xor ( n14045 , n13697 , n13699 );
xor ( n14046 , n14045 , n13702 );
xor ( n14047 , n13706 , n13707 );
xor ( n14048 , n14047 , n13717 );
and ( n14049 , n14046 , n14048 );
xor ( n14050 , n13736 , n13741 );
xor ( n14051 , n14050 , n13749 );
and ( n14052 , n14048 , n14051 );
and ( n14053 , n14046 , n14051 );
or ( n14054 , n14049 , n14052 , n14053 );
and ( n14055 , n14044 , n14054 );
xor ( n14056 , n13600 , n13602 );
xor ( n14057 , n14056 , n13605 );
and ( n14058 , n14054 , n14057 );
and ( n14059 , n14044 , n14057 );
or ( n14060 , n14055 , n14058 , n14059 );
and ( n14061 , n13988 , n14060 );
and ( n14062 , n13882 , n14060 );
or ( n14063 , n13989 , n14061 , n14062 );
xor ( n14064 , n13617 , n13618 );
xor ( n14065 , n14064 , n13620 );
xor ( n14066 , n13644 , n13672 );
xor ( n14067 , n14066 , n13683 );
and ( n14068 , n14065 , n14067 );
xor ( n14069 , n13705 , n13720 );
xor ( n14070 , n14069 , n13752 );
and ( n14071 , n14067 , n14070 );
and ( n14072 , n14065 , n14070 );
or ( n14073 , n14068 , n14071 , n14072 );
xor ( n14074 , n13595 , n13597 );
xor ( n14075 , n14074 , n13608 );
and ( n14076 , n14073 , n14075 );
xor ( n14077 , n13623 , n13686 );
xor ( n14078 , n14077 , n13755 );
and ( n14079 , n14075 , n14078 );
and ( n14080 , n14073 , n14078 );
or ( n14081 , n14076 , n14079 , n14080 );
and ( n14082 , n14063 , n14081 );
xor ( n14083 , n13590 , n13592 );
xor ( n14084 , n14083 , n13611 );
and ( n14085 , n14081 , n14084 );
and ( n14086 , n14063 , n14084 );
or ( n14087 , n14082 , n14085 , n14086 );
xor ( n14088 , n13588 , n13614 );
xor ( n14089 , n14088 , n13841 );
and ( n14090 , n14087 , n14089 );
xor ( n14091 , n13854 , n13856 );
xor ( n14092 , n14091 , n13859 );
and ( n14093 , n14089 , n14092 );
and ( n14094 , n14087 , n14092 );
or ( n14095 , n14090 , n14093 , n14094 );
and ( n14096 , n13880 , n14095 );
xor ( n14097 , n13844 , n13862 );
xor ( n14098 , n14097 , n13865 );
and ( n14099 , n14095 , n14098 );
and ( n14100 , n13880 , n14098 );
or ( n14101 , n14096 , n14099 , n14100 );
xor ( n14102 , n13586 , n13868 );
xor ( n14103 , n14102 , n13871 );
and ( n14104 , n14101 , n14103 );
xor ( n14105 , n14101 , n14103 );
xor ( n14106 , n13880 , n14095 );
xor ( n14107 , n14106 , n14098 );
xor ( n14108 , n13758 , n13827 );
xor ( n14109 , n14108 , n13838 );
xor ( n14110 , n13846 , n13848 );
xor ( n14111 , n14110 , n13851 );
and ( n14112 , n14109 , n14111 );
xor ( n14113 , n13811 , n13821 );
xor ( n14114 , n14113 , n13824 );
xor ( n14115 , n13830 , n13832 );
xor ( n14116 , n14115 , n13835 );
and ( n14117 , n14114 , n14116 );
xor ( n14118 , n13795 , n13805 );
xor ( n14119 , n14118 , n13808 );
xor ( n14120 , n13813 , n13815 );
xor ( n14121 , n14120 , n13818 );
and ( n14122 , n14119 , n14121 );
xor ( n14123 , n13765 , n13772 );
xor ( n14124 , n14123 , n13792 );
xor ( n14125 , n13797 , n13799 );
xor ( n14126 , n14125 , n13802 );
and ( n14127 , n14124 , n14126 );
xor ( n14128 , n13917 , n13952 );
and ( n14129 , n14126 , n14128 );
and ( n14130 , n14124 , n14128 );
or ( n14131 , n14127 , n14129 , n14130 );
and ( n14132 , n14121 , n14131 );
and ( n14133 , n14119 , n14131 );
or ( n14134 , n14122 , n14132 , n14133 );
and ( n14135 , n14116 , n14134 );
and ( n14136 , n14114 , n14134 );
or ( n14137 , n14117 , n14135 , n14136 );
and ( n14138 , n14111 , n14137 );
and ( n14139 , n14109 , n14137 );
or ( n14140 , n14112 , n14138 , n14139 );
xor ( n14141 , n14087 , n14089 );
xor ( n14142 , n14141 , n14092 );
and ( n14143 , n14140 , n14142 );
and ( n14144 , n2255 , n4982 );
and ( n14145 , n4989 , n2250 );
and ( n14146 , n14144 , n14145 );
and ( n14147 , n4721 , n5077 );
and ( n14148 , n14146 , n14147 );
and ( n14149 , n3339 , n13889 );
and ( n14150 , n14147 , n14149 );
and ( n14151 , n14146 , n14149 );
or ( n14152 , n14148 , n14150 , n14151 );
and ( n14153 , n2723 , n3739 );
and ( n14154 , n3728 , n2718 );
and ( n14155 , n14153 , n14154 );
and ( n14156 , n14152 , n14155 );
and ( n14157 , n10933 , n3301 );
and ( n14158 , n14155 , n14157 );
and ( n14159 , n14152 , n14157 );
or ( n14160 , n14156 , n14158 , n14159 );
and ( n14161 , n2928 , n3739 );
and ( n14162 , n3728 , n2923 );
and ( n14163 , n14161 , n14162 );
and ( n14164 , n10933 , n3627 );
and ( n14165 , n14163 , n14164 );
and ( n14166 , n4385 , n11777 );
and ( n14167 , n14164 , n14166 );
and ( n14168 , n14163 , n14166 );
or ( n14169 , n14165 , n14167 , n14168 );
and ( n14170 , n2048 , n5086 );
and ( n14171 , n5091 , n2059 );
and ( n14172 , n14170 , n14171 );
and ( n14173 , n3151 , n3449 );
and ( n14174 , n3454 , n3146 );
and ( n14175 , n14173 , n14174 );
and ( n14176 , n14172 , n14175 );
and ( n14177 , n4138 , n12290 );
and ( n14178 , n14175 , n14177 );
and ( n14179 , n14172 , n14177 );
or ( n14180 , n14176 , n14178 , n14179 );
and ( n14181 , n14169 , n14180 );
and ( n14182 , n2497 , n4362 );
and ( n14183 , n4367 , n2492 );
and ( n14184 , n14182 , n14183 );
and ( n14185 , n2591 , n4161 );
and ( n14186 , n4150 , n2586 );
and ( n14187 , n14185 , n14186 );
and ( n14188 , n14184 , n14187 );
and ( n14189 , n3645 , n13465 );
and ( n14190 , n14187 , n14189 );
and ( n14191 , n14184 , n14189 );
or ( n14192 , n14188 , n14190 , n14191 );
and ( n14193 , n14180 , n14192 );
and ( n14194 , n14169 , n14192 );
or ( n14195 , n14181 , n14193 , n14194 );
and ( n14196 , n14160 , n14195 );
xor ( n14197 , n13722 , n13723 );
xor ( n14198 , n14197 , n13725 );
xor ( n14199 , n13729 , n13730 );
xor ( n14200 , n14199 , n13732 );
and ( n14201 , n14198 , n14200 );
and ( n14202 , n14195 , n14201 );
and ( n14203 , n14160 , n14201 );
or ( n14204 , n14196 , n14202 , n14203 );
xor ( n14205 , n13929 , n13932 );
xor ( n14206 , n14205 , n13934 );
xor ( n14207 , n13896 , n13899 );
xor ( n14208 , n14207 , n13901 );
and ( n14209 , n14206 , n14208 );
xor ( n14210 , n13995 , n13996 );
xor ( n14211 , n14210 , n13998 );
and ( n14212 , n14208 , n14211 );
and ( n14213 , n14206 , n14211 );
or ( n14214 , n14209 , n14212 , n14213 );
xor ( n14215 , n13926 , n13937 );
xor ( n14216 , n14215 , n13949 );
and ( n14217 , n14214 , n14216 );
and ( n14218 , n14204 , n14217 );
xor ( n14219 , n13776 , n13786 );
xor ( n14220 , n14219 , n13789 );
xor ( n14221 , n13893 , n13904 );
xor ( n14222 , n14221 , n13914 );
and ( n14223 , n14220 , n14222 );
xor ( n14224 , n13968 , n13970 );
xor ( n14225 , n14224 , n13973 );
and ( n14226 , n14222 , n14225 );
and ( n14227 , n14220 , n14225 );
or ( n14228 , n14223 , n14226 , n14227 );
and ( n14229 , n14217 , n14228 );
and ( n14230 , n14204 , n14228 );
or ( n14231 , n14218 , n14229 , n14230 );
xnor ( n14232 , n13979 , n13981 );
xor ( n14233 , n13920 , n13921 );
xor ( n14234 , n14233 , n13923 );
xor ( n14235 , n13885 , n13886 );
xor ( n14236 , n14235 , n13890 );
and ( n14237 , n14234 , n14236 );
xor ( n14238 , n14198 , n14200 );
and ( n14239 , n14236 , n14238 );
and ( n14240 , n14234 , n14238 );
or ( n14241 , n14237 , n14239 , n14240 );
and ( n14242 , n14232 , n14241 );
and ( n14243 , n1995 , n10869 );
and ( n14244 , n10862 , n1990 );
and ( n14245 , n14243 , n14244 );
and ( n14246 , n2309 , n4734 );
and ( n14247 , n4739 , n2304 );
and ( n14248 , n14246 , n14247 );
and ( n14249 , n14245 , n14248 );
and ( n14250 , n4579 , n11156 );
and ( n14251 , n14248 , n14250 );
and ( n14252 , n14245 , n14250 );
or ( n14253 , n14249 , n14251 , n14252 );
and ( n14254 , n2723 , n3903 );
and ( n14255 , n3892 , n2718 );
and ( n14256 , n14254 , n14255 );
and ( n14257 , n10886 , n3929 );
and ( n14258 , n14256 , n14257 );
and ( n14259 , n3833 , n12900 );
and ( n14260 , n14257 , n14259 );
and ( n14261 , n14256 , n14259 );
or ( n14262 , n14258 , n14260 , n14261 );
and ( n14263 , n14253 , n14262 );
xor ( n14264 , n10028 , n10607 );
buf ( n14265 , n14264 );
buf ( n14266 , n14265 );
buf ( n14267 , n14266 );
and ( n14268 , n5177 , n4522 );
and ( n14269 , n14267 , n14268 );
xor ( n14270 , n13939 , n13940 );
and ( n14271 , n14268 , n14270 );
and ( n14272 , n14267 , n14270 );
or ( n14273 , n14269 , n14271 , n14272 );
and ( n14274 , n14262 , n14273 );
and ( n14275 , n14253 , n14273 );
or ( n14276 , n14263 , n14274 , n14275 );
and ( n14277 , n14241 , n14276 );
and ( n14278 , n14232 , n14276 );
or ( n14279 , n14242 , n14277 , n14278 );
xor ( n14280 , n13894 , n13895 );
xor ( n14281 , n13897 , n13898 );
and ( n14282 , n14280 , n14281 );
xor ( n14283 , n13906 , n13907 );
and ( n14284 , n14281 , n14283 );
and ( n14285 , n14280 , n14283 );
or ( n14286 , n14282 , n14284 , n14285 );
xor ( n14287 , n13927 , n13928 );
xor ( n14288 , n13993 , n13994 );
and ( n14289 , n14287 , n14288 );
xor ( n14290 , n13942 , n13943 );
and ( n14291 , n14288 , n14290 );
and ( n14292 , n14287 , n14290 );
or ( n14293 , n14289 , n14291 , n14292 );
and ( n14294 , n14286 , n14293 );
xor ( n14295 , n13883 , n13884 );
xor ( n14296 , n14153 , n14154 );
and ( n14297 , n14295 , n14296 );
xor ( n14298 , n13930 , n13931 );
and ( n14299 , n14296 , n14298 );
and ( n14300 , n14295 , n14298 );
or ( n14301 , n14297 , n14299 , n14300 );
and ( n14302 , n14293 , n14301 );
and ( n14303 , n14286 , n14301 );
or ( n14304 , n14294 , n14302 , n14303 );
xor ( n14305 , n14005 , n14006 );
xor ( n14306 , n14305 , n14008 );
xor ( n14307 , n14012 , n14013 );
xor ( n14308 , n14307 , n14015 );
and ( n14309 , n14306 , n14308 );
xor ( n14310 , n14020 , n14021 );
xor ( n14311 , n14310 , n14024 );
and ( n14312 , n14308 , n14311 );
and ( n14313 , n14306 , n14311 );
or ( n14314 , n14309 , n14312 , n14313 );
and ( n14315 , n14304 , n14314 );
xor ( n14316 , n13990 , n13991 );
xor ( n14317 , n14316 , n14001 );
and ( n14318 , n14314 , n14317 );
and ( n14319 , n14304 , n14317 );
or ( n14320 , n14315 , n14318 , n14319 );
and ( n14321 , n14279 , n14320 );
xor ( n14322 , n13955 , n13957 );
xor ( n14323 , n14322 , n13960 );
and ( n14324 , n14320 , n14323 );
and ( n14325 , n14279 , n14323 );
or ( n14326 , n14321 , n14324 , n14325 );
and ( n14327 , n14231 , n14326 );
xor ( n14328 , n13966 , n13976 );
xor ( n14329 , n14328 , n13982 );
xor ( n14330 , n14004 , n14030 );
xor ( n14331 , n14330 , n14041 );
and ( n14332 , n14329 , n14331 );
xor ( n14333 , n14046 , n14048 );
xor ( n14334 , n14333 , n14051 );
and ( n14335 , n14331 , n14334 );
and ( n14336 , n14329 , n14334 );
or ( n14337 , n14332 , n14335 , n14336 );
and ( n14338 , n14326 , n14337 );
and ( n14339 , n14231 , n14337 );
or ( n14340 , n14327 , n14338 , n14339 );
xor ( n14341 , n13953 , n13963 );
xor ( n14342 , n14341 , n13985 );
xor ( n14343 , n14044 , n14054 );
xor ( n14344 , n14343 , n14057 );
and ( n14345 , n14342 , n14344 );
xor ( n14346 , n14065 , n14067 );
xor ( n14347 , n14346 , n14070 );
and ( n14348 , n14344 , n14347 );
and ( n14349 , n14342 , n14347 );
or ( n14350 , n14345 , n14348 , n14349 );
and ( n14351 , n14340 , n14350 );
xor ( n14352 , n13882 , n13988 );
xor ( n14353 , n14352 , n14060 );
and ( n14354 , n14350 , n14353 );
and ( n14355 , n14340 , n14353 );
or ( n14356 , n14351 , n14354 , n14355 );
xor ( n14357 , n14063 , n14081 );
xor ( n14358 , n14357 , n14084 );
and ( n14359 , n14356 , n14358 );
xor ( n14360 , n14073 , n14075 );
xor ( n14361 , n14360 , n14078 );
xor ( n14362 , n13941 , n13944 );
xor ( n14363 , n14362 , n13946 );
xor ( n14364 , n13908 , n13909 );
xor ( n14365 , n14364 , n13911 );
and ( n14366 , n14363 , n14365 );
xor ( n14367 , n14152 , n14155 );
xor ( n14368 , n14367 , n14157 );
and ( n14369 , n14365 , n14368 );
and ( n14370 , n14363 , n14368 );
or ( n14371 , n14366 , n14369 , n14370 );
and ( n14372 , n11116 , n1990 );
and ( n14373 , n10862 , n2059 );
and ( n14374 , n14372 , n14373 );
and ( n14375 , n4989 , n2304 );
and ( n14376 , n14373 , n14375 );
and ( n14377 , n14372 , n14375 );
or ( n14378 , n14374 , n14376 , n14377 );
and ( n14379 , n1995 , n11111 );
and ( n14380 , n2048 , n10869 );
and ( n14381 , n14379 , n14380 );
and ( n14382 , n2309 , n4982 );
and ( n14383 , n14380 , n14382 );
and ( n14384 , n14379 , n14382 );
or ( n14385 , n14381 , n14383 , n14384 );
and ( n14386 , n14378 , n14385 );
xor ( n14387 , n14245 , n14248 );
xor ( n14388 , n14387 , n14250 );
and ( n14389 , n14386 , n14388 );
xor ( n14390 , n14163 , n14164 );
xor ( n14391 , n14390 , n14166 );
and ( n14392 , n14388 , n14391 );
and ( n14393 , n14386 , n14391 );
or ( n14394 , n14389 , n14392 , n14393 );
xor ( n14395 , n14172 , n14175 );
xor ( n14396 , n14395 , n14177 );
xor ( n14397 , n14256 , n14257 );
xor ( n14398 , n14397 , n14259 );
and ( n14399 , n14396 , n14398 );
xor ( n14400 , n14146 , n14147 );
xor ( n14401 , n14400 , n14149 );
and ( n14402 , n14398 , n14401 );
and ( n14403 , n14396 , n14401 );
or ( n14404 , n14399 , n14402 , n14403 );
and ( n14405 , n14394 , n14404 );
xor ( n14406 , n14169 , n14180 );
xor ( n14407 , n14406 , n14192 );
and ( n14408 , n14404 , n14407 );
and ( n14409 , n14394 , n14407 );
or ( n14410 , n14405 , n14408 , n14409 );
and ( n14411 , n14371 , n14410 );
xor ( n14412 , n14160 , n14195 );
xor ( n14413 , n14412 , n14201 );
and ( n14414 , n14410 , n14413 );
and ( n14415 , n14371 , n14413 );
or ( n14416 , n14411 , n14414 , n14415 );
xor ( n14417 , n14011 , n14018 );
xor ( n14418 , n14417 , n14027 );
xor ( n14419 , n14033 , n14035 );
xor ( n14420 , n14419 , n14038 );
and ( n14421 , n14418 , n14420 );
xor ( n14422 , n14214 , n14216 );
and ( n14423 , n14420 , n14422 );
and ( n14424 , n14418 , n14422 );
or ( n14425 , n14421 , n14423 , n14424 );
and ( n14426 , n14416 , n14425 );
xor ( n14427 , n14206 , n14208 );
xor ( n14428 , n14427 , n14211 );
and ( n14429 , n2591 , n4362 );
and ( n14430 , n4367 , n2586 );
and ( n14431 , n14429 , n14430 );
buf ( n14432 , n3293 );
and ( n14433 , n14431 , n14432 );
and ( n14434 , n4579 , n11777 );
and ( n14435 , n14432 , n14434 );
and ( n14436 , n14431 , n14434 );
or ( n14437 , n14433 , n14435 , n14436 );
and ( n14438 , n2928 , n3903 );
and ( n14439 , n3892 , n2923 );
and ( n14440 , n14438 , n14439 );
and ( n14441 , n10886 , n4522 );
and ( n14442 , n14440 , n14441 );
and ( n14443 , n4138 , n12900 );
and ( n14444 , n14441 , n14443 );
and ( n14445 , n14440 , n14443 );
or ( n14446 , n14442 , n14444 , n14445 );
and ( n14447 , n14437 , n14446 );
and ( n14448 , n2497 , n4734 );
and ( n14449 , n4739 , n2492 );
and ( n14450 , n14448 , n14449 );
and ( n14451 , n4385 , n12290 );
and ( n14452 , n14450 , n14451 );
buf ( n14453 , n3244 );
buf ( n14454 , n14453 );
and ( n14455 , n3339 , n14454 );
and ( n14456 , n14451 , n14455 );
and ( n14457 , n14450 , n14455 );
or ( n14458 , n14452 , n14456 , n14457 );
and ( n14459 , n14446 , n14458 );
and ( n14460 , n14437 , n14458 );
or ( n14461 , n14447 , n14459 , n14460 );
and ( n14462 , n14428 , n14461 );
and ( n14463 , n2723 , n4161 );
and ( n14464 , n4150 , n2718 );
and ( n14465 , n14463 , n14464 );
and ( n14466 , n3151 , n3739 );
and ( n14467 , n3728 , n3146 );
and ( n14468 , n14466 , n14467 );
and ( n14469 , n14465 , n14468 );
and ( n14470 , n3645 , n13889 );
and ( n14471 , n14468 , n14470 );
and ( n14472 , n14465 , n14470 );
or ( n14473 , n14469 , n14471 , n14472 );
and ( n14474 , n10933 , n3929 );
and ( n14475 , n4721 , n11156 );
and ( n14476 , n14474 , n14475 );
and ( n14477 , n3833 , n13465 );
and ( n14478 , n14475 , n14477 );
and ( n14479 , n14474 , n14477 );
or ( n14480 , n14476 , n14478 , n14479 );
or ( n14481 , n14473 , n14480 );
and ( n14482 , n14461 , n14481 );
and ( n14483 , n14428 , n14481 );
or ( n14484 , n14462 , n14482 , n14483 );
xor ( n14485 , n13918 , n13919 );
and ( n14486 , n1911 , n11111 );
and ( n14487 , n11116 , n1906 );
and ( n14488 , n14486 , n14487 );
and ( n14489 , n14485 , n14488 );
xor ( n14490 , n14184 , n14187 );
xor ( n14491 , n14490 , n14189 );
and ( n14492 , n14488 , n14491 );
and ( n14493 , n14485 , n14491 );
or ( n14494 , n14489 , n14492 , n14493 );
and ( n14495 , n2255 , n5086 );
and ( n14496 , n5091 , n2250 );
and ( n14497 , n14495 , n14496 );
and ( n14498 , n3293 , n3449 );
and ( n14499 , n3454 , n3288 );
and ( n14500 , n14498 , n14499 );
and ( n14501 , n14497 , n14500 );
and ( n14502 , n5177 , n5077 );
and ( n14503 , n14500 , n14502 );
and ( n14504 , n14497 , n14502 );
or ( n14505 , n14501 , n14503 , n14504 );
xor ( n14506 , n10030 , n10606 );
buf ( n14507 , n14506 );
buf ( n14508 , n14507 );
buf ( n14509 , n14508 );
buf ( n14510 , n3246 );
and ( n14511 , n14509 , n14510 );
xor ( n14512 , n14486 , n14487 );
and ( n14513 , n14510 , n14512 );
and ( n14514 , n14509 , n14512 );
or ( n14515 , n14511 , n14513 , n14514 );
and ( n14516 , n14505 , n14515 );
xor ( n14517 , n14243 , n14244 );
xor ( n14518 , n14170 , n14171 );
and ( n14519 , n14517 , n14518 );
xor ( n14520 , n14144 , n14145 );
and ( n14521 , n14518 , n14520 );
and ( n14522 , n14517 , n14520 );
or ( n14523 , n14519 , n14521 , n14522 );
and ( n14524 , n14515 , n14523 );
and ( n14525 , n14505 , n14523 );
or ( n14526 , n14516 , n14524 , n14525 );
and ( n14527 , n14494 , n14526 );
xor ( n14528 , n14246 , n14247 );
xor ( n14529 , n14182 , n14183 );
and ( n14530 , n14528 , n14529 );
xor ( n14531 , n14185 , n14186 );
and ( n14532 , n14529 , n14531 );
and ( n14533 , n14528 , n14531 );
or ( n14534 , n14530 , n14532 , n14533 );
xor ( n14535 , n14254 , n14255 );
xor ( n14536 , n14161 , n14162 );
and ( n14537 , n14535 , n14536 );
xor ( n14538 , n14173 , n14174 );
and ( n14539 , n14536 , n14538 );
and ( n14540 , n14535 , n14538 );
or ( n14541 , n14537 , n14539 , n14540 );
and ( n14542 , n14534 , n14541 );
xor ( n14543 , n14267 , n14268 );
xor ( n14544 , n14543 , n14270 );
and ( n14545 , n14541 , n14544 );
and ( n14546 , n14534 , n14544 );
or ( n14547 , n14542 , n14545 , n14546 );
and ( n14548 , n14526 , n14547 );
and ( n14549 , n14494 , n14547 );
or ( n14550 , n14527 , n14548 , n14549 );
and ( n14551 , n14484 , n14550 );
xor ( n14552 , n14280 , n14281 );
xor ( n14553 , n14552 , n14283 );
xor ( n14554 , n14287 , n14288 );
xor ( n14555 , n14554 , n14290 );
and ( n14556 , n14553 , n14555 );
xor ( n14557 , n14295 , n14296 );
xor ( n14558 , n14557 , n14298 );
and ( n14559 , n14555 , n14558 );
and ( n14560 , n14553 , n14558 );
or ( n14561 , n14556 , n14559 , n14560 );
xor ( n14562 , n14234 , n14236 );
xor ( n14563 , n14562 , n14238 );
and ( n14564 , n14561 , n14563 );
xor ( n14565 , n14253 , n14262 );
xor ( n14566 , n14565 , n14273 );
and ( n14567 , n14563 , n14566 );
and ( n14568 , n14561 , n14566 );
or ( n14569 , n14564 , n14567 , n14568 );
and ( n14570 , n14550 , n14569 );
and ( n14571 , n14484 , n14569 );
or ( n14572 , n14551 , n14570 , n14571 );
and ( n14573 , n14425 , n14572 );
and ( n14574 , n14416 , n14572 );
or ( n14575 , n14426 , n14573 , n14574 );
xor ( n14576 , n14220 , n14222 );
xor ( n14577 , n14576 , n14225 );
xor ( n14578 , n14232 , n14241 );
xor ( n14579 , n14578 , n14276 );
and ( n14580 , n14577 , n14579 );
xor ( n14581 , n14304 , n14314 );
xor ( n14582 , n14581 , n14317 );
and ( n14583 , n14579 , n14582 );
and ( n14584 , n14577 , n14582 );
or ( n14585 , n14580 , n14583 , n14584 );
xor ( n14586 , n14124 , n14126 );
xor ( n14587 , n14586 , n14128 );
and ( n14588 , n14585 , n14587 );
xor ( n14589 , n14204 , n14217 );
xor ( n14590 , n14589 , n14228 );
and ( n14591 , n14587 , n14590 );
and ( n14592 , n14585 , n14590 );
or ( n14593 , n14588 , n14591 , n14592 );
and ( n14594 , n14575 , n14593 );
xor ( n14595 , n14119 , n14121 );
xor ( n14596 , n14595 , n14131 );
and ( n14597 , n14593 , n14596 );
and ( n14598 , n14575 , n14596 );
or ( n14599 , n14594 , n14597 , n14598 );
and ( n14600 , n14361 , n14599 );
xor ( n14601 , n14114 , n14116 );
xor ( n14602 , n14601 , n14134 );
and ( n14603 , n14599 , n14602 );
and ( n14604 , n14361 , n14602 );
or ( n14605 , n14600 , n14603 , n14604 );
and ( n14606 , n14358 , n14605 );
and ( n14607 , n14356 , n14605 );
or ( n14608 , n14359 , n14606 , n14607 );
and ( n14609 , n14142 , n14608 );
and ( n14610 , n14140 , n14608 );
or ( n14611 , n14143 , n14609 , n14610 );
and ( n14612 , n14107 , n14611 );
xor ( n14613 , n14107 , n14611 );
xor ( n14614 , n14109 , n14111 );
xor ( n14615 , n14614 , n14137 );
xor ( n14616 , n14340 , n14350 );
xor ( n14617 , n14616 , n14353 );
xor ( n14618 , n14231 , n14326 );
xor ( n14619 , n14618 , n14337 );
xor ( n14620 , n14342 , n14344 );
xor ( n14621 , n14620 , n14347 );
and ( n14622 , n14619 , n14621 );
xor ( n14623 , n14279 , n14320 );
xor ( n14624 , n14623 , n14323 );
xor ( n14625 , n14329 , n14331 );
xor ( n14626 , n14625 , n14334 );
and ( n14627 , n14624 , n14626 );
xor ( n14628 , n14371 , n14410 );
xor ( n14629 , n14628 , n14413 );
xor ( n14630 , n14286 , n14293 );
xor ( n14631 , n14630 , n14301 );
xor ( n14632 , n14306 , n14308 );
xor ( n14633 , n14632 , n14311 );
and ( n14634 , n14631 , n14633 );
xor ( n14635 , n14363 , n14365 );
xor ( n14636 , n14635 , n14368 );
and ( n14637 , n14633 , n14636 );
and ( n14638 , n14631 , n14636 );
or ( n14639 , n14634 , n14637 , n14638 );
and ( n14640 , n14629 , n14639 );
xor ( n14641 , n14394 , n14404 );
xor ( n14642 , n14641 , n14407 );
xor ( n14643 , n14386 , n14388 );
xor ( n14644 , n14643 , n14391 );
xor ( n14645 , n14396 , n14398 );
xor ( n14646 , n14645 , n14401 );
and ( n14647 , n14644 , n14646 );
and ( n14648 , n14642 , n14647 );
xor ( n14649 , n14437 , n14446 );
xor ( n14650 , n14649 , n14458 );
xnor ( n14651 , n14473 , n14480 );
and ( n14652 , n14650 , n14651 );
xor ( n14653 , n14372 , n14373 );
xor ( n14654 , n14653 , n14375 );
xor ( n14655 , n14379 , n14380 );
xor ( n14656 , n14655 , n14382 );
and ( n14657 , n14654 , n14656 );
xor ( n14658 , n14465 , n14468 );
xor ( n14659 , n14658 , n14470 );
and ( n14660 , n14657 , n14659 );
xor ( n14661 , n14431 , n14432 );
xor ( n14662 , n14661 , n14434 );
and ( n14663 , n14659 , n14662 );
and ( n14664 , n14657 , n14662 );
or ( n14665 , n14660 , n14663 , n14664 );
and ( n14666 , n14651 , n14665 );
and ( n14667 , n14650 , n14665 );
or ( n14668 , n14652 , n14666 , n14667 );
and ( n14669 , n14647 , n14668 );
and ( n14670 , n14642 , n14668 );
or ( n14671 , n14648 , n14669 , n14670 );
and ( n14672 , n14639 , n14671 );
and ( n14673 , n14629 , n14671 );
or ( n14674 , n14640 , n14672 , n14673 );
and ( n14675 , n14626 , n14674 );
and ( n14676 , n14624 , n14674 );
or ( n14677 , n14627 , n14675 , n14676 );
and ( n14678 , n14621 , n14677 );
and ( n14679 , n14619 , n14677 );
or ( n14680 , n14622 , n14678 , n14679 );
and ( n14681 , n14617 , n14680 );
xor ( n14682 , n14361 , n14599 );
xor ( n14683 , n14682 , n14602 );
and ( n14684 , n14680 , n14683 );
and ( n14685 , n14617 , n14683 );
or ( n14686 , n14681 , n14684 , n14685 );
and ( n14687 , n14615 , n14686 );
xor ( n14688 , n14356 , n14358 );
xor ( n14689 , n14688 , n14605 );
and ( n14690 , n14686 , n14689 );
and ( n14691 , n14615 , n14689 );
or ( n14692 , n14687 , n14690 , n14691 );
xor ( n14693 , n14140 , n14142 );
xor ( n14694 , n14693 , n14608 );
and ( n14695 , n14692 , n14694 );
xor ( n14696 , n14692 , n14694 );
xor ( n14697 , n14615 , n14686 );
xor ( n14698 , n14697 , n14689 );
xor ( n14699 , n10031 , n10605 );
buf ( n14700 , n14699 );
buf ( n14701 , n14700 );
buf ( n14702 , n14701 );
and ( n14703 , n4721 , n11777 );
or ( n14704 , n14702 , n14703 );
xor ( n14705 , n14497 , n14500 );
xor ( n14706 , n14705 , n14502 );
and ( n14707 , n14704 , n14706 );
xor ( n14708 , n14450 , n14451 );
xor ( n14709 , n14708 , n14455 );
and ( n14710 , n14706 , n14709 );
and ( n14711 , n14704 , n14709 );
or ( n14712 , n14707 , n14710 , n14711 );
and ( n14713 , n2309 , n5086 );
and ( n14714 , n5091 , n2304 );
and ( n14715 , n14713 , n14714 );
and ( n14716 , n3151 , n3903 );
and ( n14717 , n3892 , n3146 );
and ( n14718 , n14716 , n14717 );
and ( n14719 , n14715 , n14718 );
and ( n14720 , n3645 , n14454 );
and ( n14721 , n14718 , n14720 );
and ( n14722 , n14715 , n14720 );
or ( n14723 , n14719 , n14721 , n14722 );
and ( n14724 , n2048 , n11111 );
and ( n14725 , n11116 , n2059 );
and ( n14726 , n14724 , n14725 );
and ( n14727 , n3293 , n3739 );
and ( n14728 , n3728 , n3288 );
and ( n14729 , n14727 , n14728 );
and ( n14730 , n14726 , n14729 );
and ( n14731 , n4138 , n13465 );
and ( n14732 , n14729 , n14731 );
and ( n14733 , n14726 , n14731 );
or ( n14734 , n14730 , n14732 , n14733 );
or ( n14735 , n14723 , n14734 );
and ( n14736 , n14712 , n14735 );
xor ( n14737 , n14474 , n14475 );
xor ( n14738 , n14737 , n14477 );
xor ( n14739 , n14440 , n14441 );
xor ( n14740 , n14739 , n14443 );
and ( n14741 , n14738 , n14740 );
and ( n14742 , n14735 , n14741 );
and ( n14743 , n14712 , n14741 );
or ( n14744 , n14736 , n14742 , n14743 );
xor ( n14745 , n14378 , n14385 );
and ( n14746 , n2591 , n4734 );
and ( n14747 , n4739 , n2586 );
and ( n14748 , n14746 , n14747 );
and ( n14749 , n5177 , n11156 );
and ( n14750 , n14748 , n14749 );
and ( n14751 , n4579 , n12290 );
and ( n14752 , n14749 , n14751 );
and ( n14753 , n14748 , n14751 );
or ( n14754 , n14750 , n14752 , n14753 );
and ( n14755 , n14745 , n14754 );
and ( n14756 , n2255 , n10869 );
and ( n14757 , n10862 , n2250 );
and ( n14758 , n14756 , n14757 );
and ( n14759 , n10886 , n5077 );
and ( n14760 , n14758 , n14759 );
and ( n14761 , n3833 , n13889 );
and ( n14762 , n14759 , n14761 );
and ( n14763 , n14758 , n14761 );
or ( n14764 , n14760 , n14762 , n14763 );
and ( n14765 , n14754 , n14764 );
and ( n14766 , n14745 , n14764 );
or ( n14767 , n14755 , n14765 , n14766 );
and ( n14768 , n10933 , n4522 );
and ( n14769 , n4385 , n12900 );
and ( n14770 , n14768 , n14769 );
xor ( n14771 , n14495 , n14496 );
and ( n14772 , n14769 , n14771 );
and ( n14773 , n14768 , n14771 );
or ( n14774 , n14770 , n14772 , n14773 );
xor ( n14775 , n14448 , n14449 );
xor ( n14776 , n14429 , n14430 );
and ( n14777 , n14775 , n14776 );
xor ( n14778 , n14463 , n14464 );
and ( n14779 , n14776 , n14778 );
and ( n14780 , n14775 , n14778 );
or ( n14781 , n14777 , n14779 , n14780 );
and ( n14782 , n14774 , n14781 );
xor ( n14783 , n14438 , n14439 );
xor ( n14784 , n14466 , n14467 );
and ( n14785 , n14783 , n14784 );
xor ( n14786 , n14498 , n14499 );
and ( n14787 , n14784 , n14786 );
and ( n14788 , n14783 , n14786 );
or ( n14789 , n14785 , n14787 , n14788 );
and ( n14790 , n14781 , n14789 );
and ( n14791 , n14774 , n14789 );
or ( n14792 , n14782 , n14790 , n14791 );
and ( n14793 , n14767 , n14792 );
and ( n14794 , n2723 , n4362 );
and ( n14795 , n2928 , n4161 );
or ( n14796 , n14794 , n14795 );
and ( n14797 , n2497 , n4982 );
and ( n14798 , n4989 , n2492 );
and ( n14799 , n14797 , n14798 );
and ( n14800 , n14796 , n14799 );
and ( n14801 , n4367 , n2718 );
and ( n14802 , n4150 , n2923 );
and ( n14803 , n14801 , n14802 );
buf ( n14804 , n3454 );
and ( n14805 , n14802 , n14804 );
and ( n14806 , n14801 , n14804 );
or ( n14807 , n14803 , n14805 , n14806 );
and ( n14808 , n14799 , n14807 );
and ( n14809 , n14796 , n14807 );
or ( n14810 , n14800 , n14808 , n14809 );
xor ( n14811 , n14509 , n14510 );
xor ( n14812 , n14811 , n14512 );
and ( n14813 , n14810 , n14812 );
xor ( n14814 , n14517 , n14518 );
xor ( n14815 , n14814 , n14520 );
and ( n14816 , n14812 , n14815 );
and ( n14817 , n14810 , n14815 );
or ( n14818 , n14813 , n14816 , n14817 );
and ( n14819 , n14792 , n14818 );
and ( n14820 , n14767 , n14818 );
or ( n14821 , n14793 , n14819 , n14820 );
and ( n14822 , n14744 , n14821 );
xor ( n14823 , n14485 , n14488 );
xor ( n14824 , n14823 , n14491 );
xor ( n14825 , n14505 , n14515 );
xor ( n14826 , n14825 , n14523 );
and ( n14827 , n14824 , n14826 );
xor ( n14828 , n14534 , n14541 );
xor ( n14829 , n14828 , n14544 );
and ( n14830 , n14826 , n14829 );
and ( n14831 , n14824 , n14829 );
or ( n14832 , n14827 , n14830 , n14831 );
and ( n14833 , n14821 , n14832 );
and ( n14834 , n14744 , n14832 );
or ( n14835 , n14822 , n14833 , n14834 );
xor ( n14836 , n14428 , n14461 );
xor ( n14837 , n14836 , n14481 );
xor ( n14838 , n14494 , n14526 );
xor ( n14839 , n14838 , n14547 );
and ( n14840 , n14837 , n14839 );
xor ( n14841 , n14561 , n14563 );
xor ( n14842 , n14841 , n14566 );
and ( n14843 , n14839 , n14842 );
and ( n14844 , n14837 , n14842 );
or ( n14845 , n14840 , n14843 , n14844 );
and ( n14846 , n14835 , n14845 );
xor ( n14847 , n14418 , n14420 );
xor ( n14848 , n14847 , n14422 );
and ( n14849 , n14845 , n14848 );
and ( n14850 , n14835 , n14848 );
or ( n14851 , n14846 , n14849 , n14850 );
xor ( n14852 , n14416 , n14425 );
xor ( n14853 , n14852 , n14572 );
and ( n14854 , n14851 , n14853 );
xor ( n14855 , n14585 , n14587 );
xor ( n14856 , n14855 , n14590 );
and ( n14857 , n14853 , n14856 );
and ( n14858 , n14851 , n14856 );
or ( n14859 , n14854 , n14857 , n14858 );
xor ( n14860 , n14575 , n14593 );
xor ( n14861 , n14860 , n14596 );
and ( n14862 , n14859 , n14861 );
xor ( n14863 , n14484 , n14550 );
xor ( n14864 , n14863 , n14569 );
xor ( n14865 , n14577 , n14579 );
xor ( n14866 , n14865 , n14582 );
and ( n14867 , n14864 , n14866 );
xor ( n14868 , n14553 , n14555 );
xor ( n14869 , n14868 , n14558 );
xor ( n14870 , n14644 , n14646 );
and ( n14871 , n14869 , n14870 );
xor ( n14872 , n14528 , n14529 );
xor ( n14873 , n14872 , n14531 );
xor ( n14874 , n14535 , n14536 );
xor ( n14875 , n14874 , n14538 );
and ( n14876 , n14873 , n14875 );
xor ( n14877 , n14657 , n14659 );
xor ( n14878 , n14877 , n14662 );
and ( n14879 , n14875 , n14878 );
and ( n14880 , n14873 , n14878 );
or ( n14881 , n14876 , n14879 , n14880 );
and ( n14882 , n14870 , n14881 );
and ( n14883 , n14869 , n14881 );
or ( n14884 , n14871 , n14882 , n14883 );
xor ( n14885 , n14704 , n14706 );
xor ( n14886 , n14885 , n14709 );
xnor ( n14887 , n14723 , n14734 );
and ( n14888 , n14886 , n14887 );
xor ( n14889 , n14738 , n14740 );
and ( n14890 , n14887 , n14889 );
and ( n14891 , n14886 , n14889 );
or ( n14892 , n14888 , n14890 , n14891 );
and ( n14893 , n4721 , n12290 );
and ( n14894 , n4138 , n13889 );
and ( n14895 , n14893 , n14894 );
buf ( n14896 , n3337 );
buf ( n14897 , n14896 );
and ( n14898 , n3645 , n14897 );
and ( n14899 , n14894 , n14898 );
and ( n14900 , n14893 , n14898 );
or ( n14901 , n14895 , n14899 , n14900 );
and ( n14902 , n3293 , n3903 );
and ( n14903 , n3892 , n3288 );
and ( n14904 , n14902 , n14903 );
and ( n14905 , n4579 , n12900 );
and ( n14906 , n14904 , n14905 );
and ( n14907 , n3833 , n14454 );
and ( n14908 , n14905 , n14907 );
and ( n14909 , n14904 , n14907 );
or ( n14910 , n14906 , n14908 , n14909 );
and ( n14911 , n14901 , n14910 );
and ( n14912 , n2497 , n5086 );
and ( n14913 , n5091 , n2492 );
and ( n14914 , n14912 , n14913 );
and ( n14915 , n10886 , n11156 );
and ( n14916 , n14914 , n14915 );
and ( n14917 , n5177 , n11777 );
and ( n14918 , n14915 , n14917 );
and ( n14919 , n14914 , n14917 );
or ( n14920 , n14916 , n14918 , n14919 );
and ( n14921 , n14910 , n14920 );
and ( n14922 , n14901 , n14920 );
or ( n14923 , n14911 , n14921 , n14922 );
xnor ( n14924 , n14702 , n14703 );
and ( n14925 , n2309 , n10869 );
and ( n14926 , n10862 , n2304 );
and ( n14927 , n14925 , n14926 );
and ( n14928 , n3151 , n4161 );
and ( n14929 , n4150 , n3146 );
and ( n14930 , n14928 , n14929 );
and ( n14931 , n14927 , n14930 );
and ( n14932 , n4385 , n13465 );
and ( n14933 , n14930 , n14932 );
and ( n14934 , n14927 , n14932 );
or ( n14935 , n14931 , n14933 , n14934 );
and ( n14936 , n14924 , n14935 );
and ( n14937 , n2255 , n11111 );
and ( n14938 , n11116 , n2250 );
and ( n14939 , n14937 , n14938 );
and ( n14940 , n2723 , n4734 );
and ( n14941 , n4739 , n2718 );
and ( n14942 , n14940 , n14941 );
and ( n14943 , n14939 , n14942 );
buf ( n14944 , n3339 );
and ( n14945 , n14942 , n14944 );
and ( n14946 , n14939 , n14944 );
or ( n14947 , n14943 , n14945 , n14946 );
and ( n14948 , n14935 , n14947 );
and ( n14949 , n14924 , n14947 );
or ( n14950 , n14936 , n14948 , n14949 );
and ( n14951 , n14923 , n14950 );
and ( n14952 , n4989 , n2586 );
and ( n14953 , n4367 , n2923 );
and ( n14954 , n14952 , n14953 );
and ( n14955 , n3728 , n3449 );
and ( n14956 , n14953 , n14955 );
and ( n14957 , n14952 , n14955 );
or ( n14958 , n14954 , n14956 , n14957 );
and ( n14959 , n2591 , n4982 );
and ( n14960 , n2928 , n4362 );
and ( n14961 , n14959 , n14960 );
and ( n14962 , n3454 , n3739 );
and ( n14963 , n14960 , n14962 );
and ( n14964 , n14959 , n14962 );
or ( n14965 , n14961 , n14963 , n14964 );
and ( n14966 , n14958 , n14965 );
xor ( n14967 , n14748 , n14749 );
xor ( n14968 , n14967 , n14751 );
and ( n14969 , n14966 , n14968 );
xor ( n14970 , n14758 , n14759 );
xor ( n14971 , n14970 , n14761 );
and ( n14972 , n14968 , n14971 );
and ( n14973 , n14966 , n14971 );
or ( n14974 , n14969 , n14972 , n14973 );
and ( n14975 , n14950 , n14974 );
and ( n14976 , n14923 , n14974 );
or ( n14977 , n14951 , n14975 , n14976 );
and ( n14978 , n14892 , n14977 );
xor ( n14979 , n14715 , n14718 );
xor ( n14980 , n14979 , n14720 );
xor ( n14981 , n14726 , n14729 );
xor ( n14982 , n14981 , n14731 );
and ( n14983 , n14980 , n14982 );
xor ( n14984 , n14654 , n14656 );
and ( n14985 , n14982 , n14984 );
and ( n14986 , n14980 , n14984 );
or ( n14987 , n14983 , n14985 , n14986 );
xor ( n14988 , n10034 , n10603 );
buf ( n14989 , n14988 );
buf ( n14990 , n14989 );
buf ( n14991 , n14990 );
and ( n14992 , n10933 , n5077 );
and ( n14993 , n14991 , n14992 );
xnor ( n14994 , n14794 , n14795 );
and ( n14995 , n14992 , n14994 );
and ( n14996 , n14991 , n14994 );
or ( n14997 , n14993 , n14995 , n14996 );
xor ( n14998 , n14724 , n14725 );
xor ( n14999 , n14756 , n14757 );
and ( n15000 , n14998 , n14999 );
xor ( n15001 , n14713 , n14714 );
and ( n15002 , n14999 , n15001 );
and ( n15003 , n14998 , n15001 );
or ( n15004 , n15000 , n15002 , n15003 );
and ( n15005 , n14997 , n15004 );
xor ( n15006 , n14797 , n14798 );
xor ( n15007 , n14746 , n14747 );
and ( n15008 , n15006 , n15007 );
xor ( n15009 , n14716 , n14717 );
and ( n15010 , n15007 , n15009 );
and ( n15011 , n15006 , n15009 );
or ( n15012 , n15008 , n15010 , n15011 );
and ( n15013 , n15004 , n15012 );
and ( n15014 , n14997 , n15012 );
or ( n15015 , n15005 , n15013 , n15014 );
and ( n15016 , n14987 , n15015 );
xor ( n15017 , n14727 , n14728 );
xor ( n15018 , n10035 , n10602 );
buf ( n15019 , n15018 );
buf ( n15020 , n15019 );
buf ( n15021 , n15020 );
and ( n15022 , n4579 , n13465 );
or ( n15023 , n15021 , n15022 );
and ( n15024 , n15017 , n15023 );
xor ( n15025 , n14801 , n14802 );
xor ( n15026 , n15025 , n14804 );
and ( n15027 , n15023 , n15026 );
and ( n15028 , n15017 , n15026 );
or ( n15029 , n15024 , n15027 , n15028 );
xor ( n15030 , n14768 , n14769 );
xor ( n15031 , n15030 , n14771 );
and ( n15032 , n15029 , n15031 );
xor ( n15033 , n14775 , n14776 );
xor ( n15034 , n15033 , n14778 );
and ( n15035 , n15031 , n15034 );
and ( n15036 , n15029 , n15034 );
or ( n15037 , n15032 , n15035 , n15036 );
and ( n15038 , n15015 , n15037 );
and ( n15039 , n14987 , n15037 );
or ( n15040 , n15016 , n15038 , n15039 );
and ( n15041 , n14977 , n15040 );
and ( n15042 , n14892 , n15040 );
or ( n15043 , n14978 , n15041 , n15042 );
and ( n15044 , n14884 , n15043 );
xor ( n15045 , n14745 , n14754 );
xor ( n15046 , n15045 , n14764 );
xor ( n15047 , n14774 , n14781 );
xor ( n15048 , n15047 , n14789 );
and ( n15049 , n15046 , n15048 );
xor ( n15050 , n14810 , n14812 );
xor ( n15051 , n15050 , n14815 );
and ( n15052 , n15048 , n15051 );
and ( n15053 , n15046 , n15051 );
or ( n15054 , n15049 , n15052 , n15053 );
xor ( n15055 , n14650 , n14651 );
xor ( n15056 , n15055 , n14665 );
and ( n15057 , n15054 , n15056 );
xor ( n15058 , n14712 , n14735 );
xor ( n15059 , n15058 , n14741 );
and ( n15060 , n15056 , n15059 );
and ( n15061 , n15054 , n15059 );
or ( n15062 , n15057 , n15060 , n15061 );
and ( n15063 , n15043 , n15062 );
and ( n15064 , n14884 , n15062 );
or ( n15065 , n15044 , n15063 , n15064 );
and ( n15066 , n14866 , n15065 );
and ( n15067 , n14864 , n15065 );
or ( n15068 , n14867 , n15066 , n15067 );
xor ( n15069 , n14631 , n14633 );
xor ( n15070 , n15069 , n14636 );
xor ( n15071 , n14642 , n14647 );
xor ( n15072 , n15071 , n14668 );
and ( n15073 , n15070 , n15072 );
xor ( n15074 , n14744 , n14821 );
xor ( n15075 , n15074 , n14832 );
and ( n15076 , n15072 , n15075 );
and ( n15077 , n15070 , n15075 );
or ( n15078 , n15073 , n15076 , n15077 );
xor ( n15079 , n14629 , n14639 );
xor ( n15080 , n15079 , n14671 );
and ( n15081 , n15078 , n15080 );
xor ( n15082 , n14835 , n14845 );
xor ( n15083 , n15082 , n14848 );
and ( n15084 , n15080 , n15083 );
and ( n15085 , n15078 , n15083 );
or ( n15086 , n15081 , n15084 , n15085 );
and ( n15087 , n15068 , n15086 );
xor ( n15088 , n14624 , n14626 );
xor ( n15089 , n15088 , n14674 );
and ( n15090 , n15086 , n15089 );
and ( n15091 , n15068 , n15089 );
or ( n15092 , n15087 , n15090 , n15091 );
and ( n15093 , n14861 , n15092 );
and ( n15094 , n14859 , n15092 );
or ( n15095 , n14862 , n15093 , n15094 );
xor ( n15096 , n14617 , n14680 );
xor ( n15097 , n15096 , n14683 );
and ( n15098 , n15095 , n15097 );
xor ( n15099 , n14619 , n14621 );
xor ( n15100 , n15099 , n14677 );
xor ( n15101 , n14851 , n14853 );
xor ( n15102 , n15101 , n14856 );
xor ( n15103 , n14837 , n14839 );
xor ( n15104 , n15103 , n14842 );
xor ( n15105 , n14767 , n14792 );
xor ( n15106 , n15105 , n14818 );
xor ( n15107 , n14824 , n14826 );
xor ( n15108 , n15107 , n14829 );
and ( n15109 , n15106 , n15108 );
and ( n15110 , n2497 , n10869 );
and ( n15111 , n10862 , n2492 );
and ( n15112 , n15110 , n15111 );
and ( n15113 , n4721 , n12900 );
and ( n15114 , n15112 , n15113 );
and ( n15115 , n3833 , n14897 );
and ( n15116 , n15113 , n15115 );
and ( n15117 , n15112 , n15115 );
or ( n15118 , n15114 , n15116 , n15117 );
and ( n15119 , n2723 , n4982 );
and ( n15120 , n4989 , n2718 );
and ( n15121 , n15119 , n15120 );
and ( n15122 , n3293 , n4161 );
and ( n15123 , n4150 , n3288 );
and ( n15124 , n15122 , n15123 );
and ( n15125 , n15121 , n15124 );
and ( n15126 , n10886 , n11777 );
and ( n15127 , n15124 , n15126 );
and ( n15128 , n15121 , n15126 );
or ( n15129 , n15125 , n15127 , n15128 );
and ( n15130 , n15118 , n15129 );
xor ( n15131 , n14939 , n14942 );
xor ( n15132 , n15131 , n14944 );
and ( n15133 , n15129 , n15132 );
and ( n15134 , n15118 , n15132 );
or ( n15135 , n15130 , n15133 , n15134 );
xor ( n15136 , n14901 , n14910 );
xor ( n15137 , n15136 , n14920 );
and ( n15138 , n15135 , n15137 );
xor ( n15139 , n14924 , n14935 );
xor ( n15140 , n15139 , n14947 );
and ( n15141 , n15137 , n15140 );
and ( n15142 , n15135 , n15140 );
or ( n15143 , n15138 , n15141 , n15142 );
xor ( n15144 , n14783 , n14784 );
xor ( n15145 , n15144 , n14786 );
xor ( n15146 , n14796 , n14799 );
xor ( n15147 , n15146 , n14807 );
and ( n15148 , n15145 , n15147 );
xor ( n15149 , n14966 , n14968 );
xor ( n15150 , n15149 , n14971 );
and ( n15151 , n15147 , n15150 );
and ( n15152 , n15145 , n15150 );
or ( n15153 , n15148 , n15151 , n15152 );
and ( n15154 , n15143 , n15153 );
xor ( n15155 , n14952 , n14953 );
xor ( n15156 , n15155 , n14955 );
xor ( n15157 , n14959 , n14960 );
xor ( n15158 , n15157 , n14962 );
and ( n15159 , n15156 , n15158 );
xor ( n15160 , n14927 , n14930 );
xor ( n15161 , n15160 , n14932 );
and ( n15162 , n15159 , n15161 );
xor ( n15163 , n14893 , n14894 );
xor ( n15164 , n15163 , n14898 );
and ( n15165 , n15161 , n15164 );
and ( n15166 , n15159 , n15164 );
or ( n15167 , n15162 , n15165 , n15166 );
and ( n15168 , n2928 , n4734 );
and ( n15169 , n4739 , n2923 );
and ( n15170 , n15168 , n15169 );
and ( n15171 , n10933 , n11156 );
and ( n15172 , n15170 , n15171 );
and ( n15173 , n5177 , n12290 );
and ( n15174 , n15171 , n15173 );
and ( n15175 , n15170 , n15173 );
or ( n15176 , n15172 , n15174 , n15175 );
and ( n15177 , n2309 , n11111 );
and ( n15178 , n11116 , n2304 );
and ( n15179 , n15177 , n15178 );
and ( n15180 , n3151 , n4362 );
and ( n15181 , n4367 , n3146 );
and ( n15182 , n15180 , n15181 );
and ( n15183 , n15179 , n15182 );
and ( n15184 , n4385 , n13889 );
and ( n15185 , n15182 , n15184 );
and ( n15186 , n15179 , n15184 );
or ( n15187 , n15183 , n15185 , n15186 );
and ( n15188 , n15176 , n15187 );
and ( n15189 , n15167 , n15188 );
xor ( n15190 , n14958 , n14965 );
and ( n15191 , n2591 , n5086 );
and ( n15192 , n5091 , n2586 );
and ( n15193 , n15191 , n15192 );
and ( n15194 , n3454 , n3903 );
and ( n15195 , n3892 , n3449 );
and ( n15196 , n15194 , n15195 );
and ( n15197 , n15193 , n15196 );
and ( n15198 , n4138 , n14454 );
and ( n15199 , n15196 , n15198 );
and ( n15200 , n15193 , n15198 );
or ( n15201 , n15197 , n15199 , n15200 );
and ( n15202 , n15190 , n15201 );
buf ( n15203 , n3728 );
buf ( n15204 , n15203 );
xnor ( n15205 , n15021 , n15022 );
and ( n15206 , n15204 , n15205 );
xor ( n15207 , n14937 , n14938 );
and ( n15208 , n15205 , n15207 );
and ( n15209 , n15204 , n15207 );
or ( n15210 , n15206 , n15208 , n15209 );
and ( n15211 , n15201 , n15210 );
and ( n15212 , n15190 , n15210 );
or ( n15213 , n15202 , n15211 , n15212 );
and ( n15214 , n15188 , n15213 );
and ( n15215 , n15167 , n15213 );
or ( n15216 , n15189 , n15214 , n15215 );
and ( n15217 , n15153 , n15216 );
and ( n15218 , n15143 , n15216 );
or ( n15219 , n15154 , n15217 , n15218 );
and ( n15220 , n15108 , n15219 );
and ( n15221 , n15106 , n15219 );
or ( n15222 , n15109 , n15220 , n15221 );
and ( n15223 , n15104 , n15222 );
xor ( n15224 , n14925 , n14926 );
xor ( n15225 , n14912 , n14913 );
and ( n15226 , n15224 , n15225 );
xor ( n15227 , n14940 , n14941 );
and ( n15228 , n15225 , n15227 );
and ( n15229 , n15224 , n15227 );
or ( n15230 , n15226 , n15228 , n15229 );
xor ( n15231 , n14928 , n14929 );
xor ( n15232 , n14902 , n14903 );
and ( n15233 , n15231 , n15232 );
not ( n15234 , n15203 );
xor ( n15235 , n10215 , n10600 );
buf ( n15236 , n15235 );
buf ( n15237 , n15236 );
buf ( n15238 , n15237 );
and ( n15239 , n15234 , n15238 );
and ( n15240 , n15232 , n15239 );
and ( n15241 , n15231 , n15239 );
or ( n15242 , n15233 , n15240 , n15241 );
and ( n15243 , n15230 , n15242 );
xor ( n15244 , n14991 , n14992 );
xor ( n15245 , n15244 , n14994 );
and ( n15246 , n15242 , n15245 );
and ( n15247 , n15230 , n15245 );
or ( n15248 , n15243 , n15246 , n15247 );
xor ( n15249 , n14998 , n14999 );
xor ( n15250 , n15249 , n15001 );
xor ( n15251 , n15006 , n15007 );
xor ( n15252 , n15251 , n15009 );
and ( n15253 , n15250 , n15252 );
xor ( n15254 , n15017 , n15023 );
xor ( n15255 , n15254 , n15026 );
and ( n15256 , n15252 , n15255 );
and ( n15257 , n15250 , n15255 );
or ( n15258 , n15253 , n15256 , n15257 );
and ( n15259 , n15248 , n15258 );
xor ( n15260 , n14980 , n14982 );
xor ( n15261 , n15260 , n14984 );
and ( n15262 , n15258 , n15261 );
and ( n15263 , n15248 , n15261 );
or ( n15264 , n15259 , n15262 , n15263 );
xor ( n15265 , n14873 , n14875 );
xor ( n15266 , n15265 , n14878 );
and ( n15267 , n15264 , n15266 );
xor ( n15268 , n14886 , n14887 );
xor ( n15269 , n15268 , n14889 );
and ( n15270 , n15266 , n15269 );
and ( n15271 , n15264 , n15269 );
or ( n15272 , n15267 , n15270 , n15271 );
xor ( n15273 , n14923 , n14950 );
xor ( n15274 , n15273 , n14974 );
xor ( n15275 , n14987 , n15015 );
xor ( n15276 , n15275 , n15037 );
and ( n15277 , n15274 , n15276 );
xor ( n15278 , n15046 , n15048 );
xor ( n15279 , n15278 , n15051 );
and ( n15280 , n15276 , n15279 );
and ( n15281 , n15274 , n15279 );
or ( n15282 , n15277 , n15280 , n15281 );
and ( n15283 , n15272 , n15282 );
xor ( n15284 , n14869 , n14870 );
xor ( n15285 , n15284 , n14881 );
and ( n15286 , n15282 , n15285 );
and ( n15287 , n15272 , n15285 );
or ( n15288 , n15283 , n15286 , n15287 );
and ( n15289 , n15222 , n15288 );
and ( n15290 , n15104 , n15288 );
or ( n15291 , n15223 , n15289 , n15290 );
xor ( n15292 , n14864 , n14866 );
xor ( n15293 , n15292 , n15065 );
and ( n15294 , n15291 , n15293 );
xor ( n15295 , n15078 , n15080 );
xor ( n15296 , n15295 , n15083 );
and ( n15297 , n15293 , n15296 );
and ( n15298 , n15291 , n15296 );
or ( n15299 , n15294 , n15297 , n15298 );
and ( n15300 , n15102 , n15299 );
xor ( n15301 , n15068 , n15086 );
xor ( n15302 , n15301 , n15089 );
and ( n15303 , n15299 , n15302 );
and ( n15304 , n15102 , n15302 );
or ( n15305 , n15300 , n15303 , n15304 );
and ( n15306 , n15100 , n15305 );
xor ( n15307 , n14859 , n14861 );
xor ( n15308 , n15307 , n15092 );
and ( n15309 , n15305 , n15308 );
and ( n15310 , n15100 , n15308 );
or ( n15311 , n15306 , n15309 , n15310 );
and ( n15312 , n15097 , n15311 );
and ( n15313 , n15095 , n15311 );
or ( n15314 , n15098 , n15312 , n15313 );
and ( n15315 , n14698 , n15314 );
xor ( n15316 , n14698 , n15314 );
xor ( n15317 , n15095 , n15097 );
xor ( n15318 , n15317 , n15311 );
xor ( n15319 , n15100 , n15305 );
xor ( n15320 , n15319 , n15308 );
xor ( n15321 , n15102 , n15299 );
xor ( n15322 , n15321 , n15302 );
xor ( n15323 , n14884 , n15043 );
xor ( n15324 , n15323 , n15062 );
xor ( n15325 , n15070 , n15072 );
xor ( n15326 , n15325 , n15075 );
and ( n15327 , n15324 , n15326 );
xor ( n15328 , n14892 , n14977 );
xor ( n15329 , n15328 , n15040 );
xor ( n15330 , n15054 , n15056 );
xor ( n15331 , n15330 , n15059 );
and ( n15332 , n15329 , n15331 );
xor ( n15333 , n14997 , n15004 );
xor ( n15334 , n15333 , n15012 );
xor ( n15335 , n15029 , n15031 );
xor ( n15336 , n15335 , n15034 );
and ( n15337 , n15334 , n15336 );
xor ( n15338 , n15135 , n15137 );
xor ( n15339 , n15338 , n15140 );
and ( n15340 , n15336 , n15339 );
and ( n15341 , n15334 , n15339 );
or ( n15342 , n15337 , n15340 , n15341 );
and ( n15343 , n3454 , n4161 );
and ( n15344 , n4150 , n3449 );
and ( n15345 , n15343 , n15344 );
and ( n15346 , n3728 , n3903 );
and ( n15347 , n3892 , n3739 );
and ( n15348 , n15346 , n15347 );
and ( n15349 , n15345 , n15348 );
and ( n15350 , n10933 , n11777 );
and ( n15351 , n15348 , n15350 );
and ( n15352 , n15345 , n15350 );
or ( n15353 , n15349 , n15351 , n15352 );
and ( n15354 , n2591 , n10869 );
and ( n15355 , n10862 , n2586 );
and ( n15356 , n15354 , n15355 );
and ( n15357 , n10886 , n12290 );
and ( n15358 , n15356 , n15357 );
and ( n15359 , n4138 , n14897 );
and ( n15360 , n15357 , n15359 );
and ( n15361 , n15356 , n15359 );
or ( n15362 , n15358 , n15360 , n15361 );
and ( n15363 , n15353 , n15362 );
and ( n15364 , n2497 , n11111 );
and ( n15365 , n11116 , n2492 );
and ( n15366 , n15364 , n15365 );
and ( n15367 , n5177 , n12900 );
and ( n15368 , n15366 , n15367 );
and ( n15369 , n4721 , n13465 );
and ( n15370 , n15367 , n15369 );
and ( n15371 , n15366 , n15369 );
or ( n15372 , n15368 , n15370 , n15371 );
and ( n15373 , n15362 , n15372 );
and ( n15374 , n15353 , n15372 );
or ( n15375 , n15363 , n15373 , n15374 );
xor ( n15376 , n14904 , n14905 );
xor ( n15377 , n15376 , n14907 );
and ( n15378 , n15375 , n15377 );
xor ( n15379 , n14914 , n14915 );
xor ( n15380 , n15379 , n14917 );
and ( n15381 , n15377 , n15380 );
and ( n15382 , n15375 , n15380 );
or ( n15383 , n15378 , n15381 , n15382 );
xor ( n15384 , n15118 , n15129 );
xor ( n15385 , n15384 , n15132 );
xor ( n15386 , n15176 , n15187 );
and ( n15387 , n15385 , n15386 );
xor ( n15388 , n15112 , n15113 );
xor ( n15389 , n15388 , n15115 );
xor ( n15390 , n15121 , n15124 );
xor ( n15391 , n15390 , n15126 );
and ( n15392 , n15389 , n15391 );
xor ( n15393 , n15179 , n15182 );
xor ( n15394 , n15393 , n15184 );
and ( n15395 , n15391 , n15394 );
and ( n15396 , n15389 , n15394 );
or ( n15397 , n15392 , n15395 , n15396 );
and ( n15398 , n15386 , n15397 );
and ( n15399 , n15385 , n15397 );
or ( n15400 , n15387 , n15398 , n15399 );
and ( n15401 , n15383 , n15400 );
and ( n15402 , n2723 , n5086 );
and ( n15403 , n5091 , n2718 );
and ( n15404 , n15402 , n15403 );
and ( n15405 , n4579 , n13889 );
and ( n15406 , n15404 , n15405 );
buf ( n15407 , n3643 );
buf ( n15408 , n15407 );
and ( n15409 , n3833 , n15408 );
and ( n15410 , n15405 , n15409 );
and ( n15411 , n15404 , n15409 );
or ( n15412 , n15406 , n15410 , n15411 );
xor ( n15413 , n15170 , n15171 );
xor ( n15414 , n15413 , n15173 );
and ( n15415 , n15412 , n15414 );
xor ( n15416 , n15193 , n15196 );
xor ( n15417 , n15416 , n15198 );
and ( n15418 , n15414 , n15417 );
and ( n15419 , n15412 , n15417 );
or ( n15420 , n15415 , n15418 , n15419 );
xor ( n15421 , n15156 , n15158 );
and ( n15422 , n3151 , n4734 );
and ( n15423 , n4739 , n3146 );
and ( n15424 , n15422 , n15423 );
and ( n15425 , n3293 , n4362 );
and ( n15426 , n4367 , n3288 );
and ( n15427 , n15425 , n15426 );
and ( n15428 , n15424 , n15427 );
buf ( n15429 , n3645 );
and ( n15430 , n15427 , n15429 );
and ( n15431 , n15424 , n15429 );
or ( n15432 , n15428 , n15430 , n15431 );
and ( n15433 , n15421 , n15432 );
xor ( n15434 , n15234 , n15238 );
and ( n15435 , n2928 , n4982 );
and ( n15436 , n4989 , n2923 );
and ( n15437 , n15435 , n15436 );
and ( n15438 , n15434 , n15437 );
and ( n15439 , n4385 , n14454 );
and ( n15440 , n15437 , n15439 );
and ( n15441 , n15434 , n15439 );
or ( n15442 , n15438 , n15440 , n15441 );
and ( n15443 , n15432 , n15442 );
and ( n15444 , n15421 , n15442 );
or ( n15445 , n15433 , n15443 , n15444 );
and ( n15446 , n15420 , n15445 );
xor ( n15447 , n15177 , n15178 );
xor ( n15448 , n15110 , n15111 );
and ( n15449 , n15447 , n15448 );
xor ( n15450 , n15191 , n15192 );
and ( n15451 , n15448 , n15450 );
and ( n15452 , n15447 , n15450 );
or ( n15453 , n15449 , n15451 , n15452 );
xor ( n15454 , n15119 , n15120 );
xor ( n15455 , n15168 , n15169 );
and ( n15456 , n15454 , n15455 );
xor ( n15457 , n15180 , n15181 );
and ( n15458 , n15455 , n15457 );
and ( n15459 , n15454 , n15457 );
or ( n15460 , n15456 , n15458 , n15459 );
and ( n15461 , n15453 , n15460 );
xor ( n15462 , n15204 , n15205 );
xor ( n15463 , n15462 , n15207 );
and ( n15464 , n15460 , n15463 );
and ( n15465 , n15453 , n15463 );
or ( n15466 , n15461 , n15464 , n15465 );
and ( n15467 , n15445 , n15466 );
and ( n15468 , n15420 , n15466 );
or ( n15469 , n15446 , n15467 , n15468 );
and ( n15470 , n15400 , n15469 );
and ( n15471 , n15383 , n15469 );
or ( n15472 , n15401 , n15470 , n15471 );
and ( n15473 , n15342 , n15472 );
xor ( n15474 , n15190 , n15201 );
xor ( n15475 , n15474 , n15210 );
xor ( n15476 , n15230 , n15242 );
xor ( n15477 , n15476 , n15245 );
and ( n15478 , n15475 , n15477 );
xor ( n15479 , n15250 , n15252 );
xor ( n15480 , n15479 , n15255 );
and ( n15481 , n15477 , n15480 );
and ( n15482 , n15475 , n15480 );
or ( n15483 , n15478 , n15481 , n15482 );
xor ( n15484 , n15145 , n15147 );
xor ( n15485 , n15484 , n15150 );
and ( n15486 , n15483 , n15485 );
xor ( n15487 , n15167 , n15188 );
xor ( n15488 , n15487 , n15213 );
and ( n15489 , n15485 , n15488 );
and ( n15490 , n15483 , n15488 );
or ( n15491 , n15486 , n15489 , n15490 );
and ( n15492 , n15472 , n15491 );
and ( n15493 , n15342 , n15491 );
or ( n15494 , n15473 , n15492 , n15493 );
and ( n15495 , n15331 , n15494 );
and ( n15496 , n15329 , n15494 );
or ( n15497 , n15332 , n15495 , n15496 );
and ( n15498 , n15326 , n15497 );
and ( n15499 , n15324 , n15497 );
or ( n15500 , n15327 , n15498 , n15499 );
xor ( n15501 , n15291 , n15293 );
xor ( n15502 , n15501 , n15296 );
and ( n15503 , n15500 , n15502 );
xor ( n15504 , n15143 , n15153 );
xor ( n15505 , n15504 , n15216 );
xor ( n15506 , n15264 , n15266 );
xor ( n15507 , n15506 , n15269 );
and ( n15508 , n15505 , n15507 );
xor ( n15509 , n15274 , n15276 );
xor ( n15510 , n15509 , n15279 );
and ( n15511 , n15507 , n15510 );
and ( n15512 , n15505 , n15510 );
or ( n15513 , n15508 , n15511 , n15512 );
xor ( n15514 , n15106 , n15108 );
xor ( n15515 , n15514 , n15219 );
and ( n15516 , n15513 , n15515 );
xor ( n15517 , n15272 , n15282 );
xor ( n15518 , n15517 , n15285 );
and ( n15519 , n15515 , n15518 );
and ( n15520 , n15513 , n15518 );
or ( n15521 , n15516 , n15519 , n15520 );
xor ( n15522 , n15104 , n15222 );
xor ( n15523 , n15522 , n15288 );
and ( n15524 , n15521 , n15523 );
xor ( n15525 , n15248 , n15258 );
xor ( n15526 , n15525 , n15261 );
xor ( n15527 , n15159 , n15161 );
xor ( n15528 , n15527 , n15164 );
xor ( n15529 , n15375 , n15377 );
xor ( n15530 , n15529 , n15380 );
and ( n15531 , n15528 , n15530 );
and ( n15532 , n15526 , n15531 );
xor ( n15533 , n15389 , n15391 );
xor ( n15534 , n15533 , n15394 );
xor ( n15535 , n15412 , n15414 );
xor ( n15536 , n15535 , n15417 );
and ( n15537 , n15534 , n15536 );
xor ( n15538 , n15224 , n15225 );
xor ( n15539 , n15538 , n15227 );
xor ( n15540 , n15231 , n15232 );
xor ( n15541 , n15540 , n15239 );
and ( n15542 , n15539 , n15541 );
xor ( n15543 , n15353 , n15362 );
xor ( n15544 , n15543 , n15372 );
and ( n15545 , n15541 , n15544 );
and ( n15546 , n15539 , n15544 );
or ( n15547 , n15542 , n15545 , n15546 );
and ( n15548 , n15537 , n15547 );
and ( n15549 , n2591 , n11111 );
and ( n15550 , n11116 , n2586 );
and ( n15551 , n15549 , n15550 );
and ( n15552 , n10933 , n12290 );
and ( n15553 , n15551 , n15552 );
and ( n15554 , n10886 , n12900 );
and ( n15555 , n15552 , n15554 );
and ( n15556 , n15551 , n15554 );
or ( n15557 , n15553 , n15555 , n15556 );
and ( n15558 , n2928 , n5086 );
and ( n15559 , n5091 , n2923 );
and ( n15560 , n15558 , n15559 );
and ( n15561 , n4721 , n13889 );
and ( n15562 , n15560 , n15561 );
and ( n15563 , n4385 , n14897 );
and ( n15564 , n15561 , n15563 );
and ( n15565 , n15560 , n15563 );
or ( n15566 , n15562 , n15564 , n15565 );
and ( n15567 , n15557 , n15566 );
xor ( n15568 , n15366 , n15367 );
xor ( n15569 , n15568 , n15369 );
and ( n15570 , n15566 , n15569 );
and ( n15571 , n15557 , n15569 );
or ( n15572 , n15567 , n15570 , n15571 );
xor ( n15573 , n15424 , n15427 );
xor ( n15574 , n15573 , n15429 );
xor ( n15575 , n15345 , n15348 );
xor ( n15576 , n15575 , n15350 );
and ( n15577 , n15574 , n15576 );
xor ( n15578 , n15356 , n15357 );
xor ( n15579 , n15578 , n15359 );
and ( n15580 , n15576 , n15579 );
and ( n15581 , n15574 , n15579 );
or ( n15582 , n15577 , n15580 , n15581 );
and ( n15583 , n15572 , n15582 );
xor ( n15584 , n15122 , n15123 );
xor ( n15585 , n15194 , n15195 );
and ( n15586 , n15584 , n15585 );
xor ( n15587 , n15404 , n15405 );
xor ( n15588 , n15587 , n15409 );
and ( n15589 , n15585 , n15588 );
and ( n15590 , n15584 , n15588 );
or ( n15591 , n15586 , n15589 , n15590 );
and ( n15592 , n15582 , n15591 );
and ( n15593 , n15572 , n15591 );
or ( n15594 , n15583 , n15592 , n15593 );
and ( n15595 , n15547 , n15594 );
and ( n15596 , n15537 , n15594 );
or ( n15597 , n15548 , n15595 , n15596 );
and ( n15598 , n15531 , n15597 );
and ( n15599 , n15526 , n15597 );
or ( n15600 , n15532 , n15598 , n15599 );
xor ( n15601 , n15434 , n15437 );
xor ( n15602 , n15601 , n15439 );
and ( n15603 , n3151 , n4982 );
and ( n15604 , n4989 , n3146 );
and ( n15605 , n15603 , n15604 );
and ( n15606 , n3728 , n4161 );
and ( n15607 , n4150 , n3739 );
and ( n15608 , n15606 , n15607 );
and ( n15609 , n15605 , n15608 );
and ( n15610 , n5177 , n13465 );
and ( n15611 , n15608 , n15610 );
and ( n15612 , n15605 , n15610 );
or ( n15613 , n15609 , n15611 , n15612 );
and ( n15614 , n15602 , n15613 );
and ( n15615 , n3293 , n4734 );
and ( n15616 , n4739 , n3288 );
and ( n15617 , n15615 , n15616 );
and ( n15618 , n3454 , n4362 );
and ( n15619 , n4367 , n3449 );
and ( n15620 , n15618 , n15619 );
and ( n15621 , n15617 , n15620 );
and ( n15622 , n4138 , n15408 );
and ( n15623 , n15620 , n15622 );
and ( n15624 , n15617 , n15622 );
or ( n15625 , n15621 , n15623 , n15624 );
and ( n15626 , n15613 , n15625 );
and ( n15627 , n15602 , n15625 );
or ( n15628 , n15614 , n15626 , n15627 );
xor ( n15629 , n10217 , n10599 );
buf ( n15630 , n15629 );
buf ( n15631 , n15630 );
buf ( n15632 , n15631 );
xor ( n15633 , n15364 , n15365 );
and ( n15634 , n15632 , n15633 );
xor ( n15635 , n15354 , n15355 );
and ( n15636 , n15633 , n15635 );
and ( n15637 , n15632 , n15635 );
or ( n15638 , n15634 , n15636 , n15637 );
xor ( n15639 , n15402 , n15403 );
xor ( n15640 , n15435 , n15436 );
and ( n15641 , n15639 , n15640 );
xor ( n15642 , n15422 , n15423 );
and ( n15643 , n15640 , n15642 );
and ( n15644 , n15639 , n15642 );
or ( n15645 , n15641 , n15643 , n15644 );
and ( n15646 , n15638 , n15645 );
xor ( n15647 , n15425 , n15426 );
xor ( n15648 , n15343 , n15344 );
and ( n15649 , n15647 , n15648 );
xor ( n15650 , n15346 , n15347 );
and ( n15651 , n15648 , n15650 );
and ( n15652 , n15647 , n15650 );
or ( n15653 , n15649 , n15651 , n15652 );
and ( n15654 , n15645 , n15653 );
and ( n15655 , n15638 , n15653 );
or ( n15656 , n15646 , n15654 , n15655 );
and ( n15657 , n15628 , n15656 );
xor ( n15658 , n15421 , n15432 );
xor ( n15659 , n15658 , n15442 );
and ( n15660 , n15656 , n15659 );
and ( n15661 , n15628 , n15659 );
or ( n15662 , n15657 , n15660 , n15661 );
xor ( n15663 , n15385 , n15386 );
xor ( n15664 , n15663 , n15397 );
and ( n15665 , n15662 , n15664 );
xor ( n15666 , n15420 , n15445 );
xor ( n15667 , n15666 , n15466 );
and ( n15668 , n15664 , n15667 );
and ( n15669 , n15662 , n15667 );
or ( n15670 , n15665 , n15668 , n15669 );
xor ( n15671 , n15334 , n15336 );
xor ( n15672 , n15671 , n15339 );
and ( n15673 , n15670 , n15672 );
xor ( n15674 , n15383 , n15400 );
xor ( n15675 , n15674 , n15469 );
and ( n15676 , n15672 , n15675 );
and ( n15677 , n15670 , n15675 );
or ( n15678 , n15673 , n15676 , n15677 );
and ( n15679 , n15600 , n15678 );
xor ( n15680 , n15342 , n15472 );
xor ( n15681 , n15680 , n15491 );
and ( n15682 , n15678 , n15681 );
and ( n15683 , n15600 , n15681 );
or ( n15684 , n15679 , n15682 , n15683 );
xor ( n15685 , n15329 , n15331 );
xor ( n15686 , n15685 , n15494 );
and ( n15687 , n15684 , n15686 );
xor ( n15688 , n15513 , n15515 );
xor ( n15689 , n15688 , n15518 );
and ( n15690 , n15686 , n15689 );
and ( n15691 , n15684 , n15689 );
or ( n15692 , n15687 , n15690 , n15691 );
and ( n15693 , n15523 , n15692 );
and ( n15694 , n15521 , n15692 );
or ( n15695 , n15524 , n15693 , n15694 );
and ( n15696 , n15502 , n15695 );
and ( n15697 , n15500 , n15695 );
or ( n15698 , n15503 , n15696 , n15697 );
and ( n15699 , n15322 , n15698 );
xor ( n15700 , n15322 , n15698 );
xor ( n15701 , n15500 , n15502 );
xor ( n15702 , n15701 , n15695 );
xor ( n15703 , n15324 , n15326 );
xor ( n15704 , n15703 , n15497 );
xor ( n15705 , n15521 , n15523 );
xor ( n15706 , n15705 , n15692 );
and ( n15707 , n15704 , n15706 );
xor ( n15708 , n15505 , n15507 );
xor ( n15709 , n15708 , n15510 );
xor ( n15710 , n15483 , n15485 );
xor ( n15711 , n15710 , n15488 );
xor ( n15712 , n15475 , n15477 );
xor ( n15713 , n15712 , n15480 );
xor ( n15714 , n15528 , n15530 );
and ( n15715 , n15713 , n15714 );
xor ( n15716 , n15453 , n15460 );
xor ( n15717 , n15716 , n15463 );
xor ( n15718 , n15534 , n15536 );
and ( n15719 , n15717 , n15718 );
xor ( n15720 , n15551 , n15552 );
xor ( n15721 , n15720 , n15554 );
xor ( n15722 , n15605 , n15608 );
xor ( n15723 , n15722 , n15610 );
and ( n15724 , n15721 , n15723 );
xor ( n15725 , n15560 , n15561 );
xor ( n15726 , n15725 , n15563 );
and ( n15727 , n15723 , n15726 );
and ( n15728 , n15721 , n15726 );
or ( n15729 , n15724 , n15727 , n15728 );
xor ( n15730 , n15557 , n15566 );
xor ( n15731 , n15730 , n15569 );
and ( n15732 , n15729 , n15731 );
and ( n15733 , n15718 , n15732 );
and ( n15734 , n15717 , n15732 );
or ( n15735 , n15719 , n15733 , n15734 );
and ( n15736 , n15714 , n15735 );
and ( n15737 , n15713 , n15735 );
or ( n15738 , n15715 , n15736 , n15737 );
and ( n15739 , n15711 , n15738 );
and ( n15740 , n10886 , n13465 );
and ( n15741 , n5177 , n13889 );
and ( n15742 , n15740 , n15741 );
and ( n15743 , n4579 , n14897 );
and ( n15744 , n15741 , n15743 );
and ( n15745 , n15740 , n15743 );
or ( n15746 , n15742 , n15744 , n15745 );
and ( n15747 , n2928 , n10869 );
and ( n15748 , n10862 , n2923 );
and ( n15749 , n15747 , n15748 );
and ( n15750 , n3293 , n4982 );
and ( n15751 , n4989 , n3288 );
and ( n15752 , n15750 , n15751 );
and ( n15753 , n15749 , n15752 );
and ( n15754 , n4385 , n15408 );
and ( n15755 , n15752 , n15754 );
and ( n15756 , n15749 , n15754 );
or ( n15757 , n15753 , n15755 , n15756 );
and ( n15758 , n15746 , n15757 );
xor ( n15759 , n15617 , n15620 );
xor ( n15760 , n15759 , n15622 );
and ( n15761 , n15757 , n15760 );
and ( n15762 , n15746 , n15760 );
or ( n15763 , n15758 , n15761 , n15762 );
xor ( n15764 , n15574 , n15576 );
xor ( n15765 , n15764 , n15579 );
and ( n15766 , n15763 , n15765 );
xor ( n15767 , n15447 , n15448 );
xor ( n15768 , n15767 , n15450 );
xor ( n15769 , n15454 , n15455 );
xor ( n15770 , n15769 , n15457 );
and ( n15771 , n15768 , n15770 );
and ( n15772 , n3151 , n5086 );
buf ( n15773 , n15772 );
and ( n15774 , n3892 , n4161 );
and ( n15775 , n4150 , n3903 );
and ( n15776 , n15774 , n15775 );
and ( n15777 , n15773 , n15776 );
and ( n15778 , n10933 , n12900 );
and ( n15779 , n15776 , n15778 );
and ( n15780 , n15773 , n15778 );
or ( n15781 , n15777 , n15779 , n15780 );
and ( n15782 , n4579 , n14454 );
or ( n15783 , n15781 , n15782 );
and ( n15784 , n15770 , n15783 );
and ( n15785 , n15768 , n15783 );
or ( n15786 , n15771 , n15784 , n15785 );
and ( n15787 , n15766 , n15786 );
buf ( n15788 , n3892 );
buf ( n15789 , n3833 );
or ( n15790 , n15788 , n15789 );
and ( n15791 , n2723 , n10869 );
and ( n15792 , n10862 , n2718 );
and ( n15793 , n15791 , n15792 );
and ( n15794 , n15790 , n15793 );
and ( n15795 , n2723 , n11111 );
and ( n15796 , n11116 , n2718 );
and ( n15797 , n15795 , n15796 );
and ( n15798 , n4721 , n14454 );
and ( n15799 , n15797 , n15798 );
buf ( n15800 , n3831 );
buf ( n15801 , n15800 );
and ( n15802 , n4138 , n15801 );
and ( n15803 , n15798 , n15802 );
and ( n15804 , n15797 , n15802 );
or ( n15805 , n15799 , n15803 , n15804 );
and ( n15806 , n15793 , n15805 );
and ( n15807 , n15790 , n15805 );
or ( n15808 , n15794 , n15806 , n15807 );
xor ( n15809 , n10223 , n10597 );
buf ( n15810 , n15809 );
buf ( n15811 , n15810 );
buf ( n15812 , n15811 );
xor ( n15813 , n15740 , n15741 );
xor ( n15814 , n15813 , n15743 );
and ( n15815 , n15812 , n15814 );
xnor ( n15816 , n15788 , n15789 );
and ( n15817 , n15814 , n15816 );
and ( n15818 , n15812 , n15816 );
or ( n15819 , n15815 , n15817 , n15818 );
xor ( n15820 , n15549 , n15550 );
xor ( n15821 , n15791 , n15792 );
and ( n15822 , n15820 , n15821 );
xor ( n15823 , n15558 , n15559 );
and ( n15824 , n15821 , n15823 );
and ( n15825 , n15820 , n15823 );
or ( n15826 , n15822 , n15824 , n15825 );
and ( n15827 , n15819 , n15826 );
xor ( n15828 , n15603 , n15604 );
xor ( n15829 , n15615 , n15616 );
and ( n15830 , n15828 , n15829 );
xor ( n15831 , n15618 , n15619 );
and ( n15832 , n15829 , n15831 );
and ( n15833 , n15828 , n15831 );
or ( n15834 , n15830 , n15832 , n15833 );
and ( n15835 , n15826 , n15834 );
and ( n15836 , n15819 , n15834 );
or ( n15837 , n15827 , n15835 , n15836 );
and ( n15838 , n15808 , n15837 );
xor ( n15839 , n15606 , n15607 );
and ( n15840 , n10933 , n13465 );
and ( n15841 , n4721 , n14897 );
and ( n15842 , n15840 , n15841 );
and ( n15843 , n4385 , n15801 );
and ( n15844 , n15841 , n15843 );
and ( n15845 , n15840 , n15843 );
or ( n15846 , n15842 , n15844 , n15845 );
and ( n15847 , n15839 , n15846 );
and ( n15848 , n3454 , n4734 );
and ( n15849 , n4739 , n3449 );
and ( n15850 , n15848 , n15849 );
and ( n15851 , n15846 , n15850 );
and ( n15852 , n15839 , n15850 );
or ( n15853 , n15847 , n15851 , n15852 );
xor ( n15854 , n15632 , n15633 );
xor ( n15855 , n15854 , n15635 );
and ( n15856 , n15853 , n15855 );
xor ( n15857 , n15639 , n15640 );
xor ( n15858 , n15857 , n15642 );
and ( n15859 , n15855 , n15858 );
and ( n15860 , n15853 , n15858 );
or ( n15861 , n15856 , n15859 , n15860 );
and ( n15862 , n15837 , n15861 );
and ( n15863 , n15808 , n15861 );
or ( n15864 , n15838 , n15862 , n15863 );
and ( n15865 , n15786 , n15864 );
and ( n15866 , n15766 , n15864 );
or ( n15867 , n15787 , n15865 , n15866 );
xor ( n15868 , n15584 , n15585 );
xor ( n15869 , n15868 , n15588 );
xor ( n15870 , n15602 , n15613 );
xor ( n15871 , n15870 , n15625 );
and ( n15872 , n15869 , n15871 );
xor ( n15873 , n15638 , n15645 );
xor ( n15874 , n15873 , n15653 );
and ( n15875 , n15871 , n15874 );
and ( n15876 , n15869 , n15874 );
or ( n15877 , n15872 , n15875 , n15876 );
xor ( n15878 , n15539 , n15541 );
xor ( n15879 , n15878 , n15544 );
and ( n15880 , n15877 , n15879 );
xor ( n15881 , n15572 , n15582 );
xor ( n15882 , n15881 , n15591 );
and ( n15883 , n15879 , n15882 );
and ( n15884 , n15877 , n15882 );
or ( n15885 , n15880 , n15883 , n15884 );
and ( n15886 , n15867 , n15885 );
xor ( n15887 , n15537 , n15547 );
xor ( n15888 , n15887 , n15594 );
and ( n15889 , n15885 , n15888 );
and ( n15890 , n15867 , n15888 );
or ( n15891 , n15886 , n15889 , n15890 );
and ( n15892 , n15738 , n15891 );
and ( n15893 , n15711 , n15891 );
or ( n15894 , n15739 , n15892 , n15893 );
and ( n15895 , n15709 , n15894 );
xor ( n15896 , n15600 , n15678 );
xor ( n15897 , n15896 , n15681 );
and ( n15898 , n15894 , n15897 );
and ( n15899 , n15709 , n15897 );
or ( n15900 , n15895 , n15898 , n15899 );
xor ( n15901 , n15684 , n15686 );
xor ( n15902 , n15901 , n15689 );
and ( n15903 , n15900 , n15902 );
xor ( n15904 , n15526 , n15531 );
xor ( n15905 , n15904 , n15597 );
xor ( n15906 , n15670 , n15672 );
xor ( n15907 , n15906 , n15675 );
and ( n15908 , n15905 , n15907 );
xor ( n15909 , n15662 , n15664 );
xor ( n15910 , n15909 , n15667 );
xor ( n15911 , n15628 , n15656 );
xor ( n15912 , n15911 , n15659 );
xor ( n15913 , n15729 , n15731 );
xor ( n15914 , n15763 , n15765 );
and ( n15915 , n15913 , n15914 );
xor ( n15916 , n15647 , n15648 );
xor ( n15917 , n15916 , n15650 );
xor ( n15918 , n15746 , n15757 );
xor ( n15919 , n15918 , n15760 );
and ( n15920 , n15917 , n15919 );
xor ( n15921 , n15721 , n15723 );
xor ( n15922 , n15921 , n15726 );
and ( n15923 , n15919 , n15922 );
and ( n15924 , n15917 , n15922 );
or ( n15925 , n15920 , n15923 , n15924 );
and ( n15926 , n15914 , n15925 );
and ( n15927 , n15913 , n15925 );
or ( n15928 , n15915 , n15926 , n15927 );
and ( n15929 , n15912 , n15928 );
xnor ( n15930 , n15781 , n15782 );
and ( n15931 , n3728 , n4734 );
and ( n15932 , n4739 , n3739 );
and ( n15933 , n15931 , n15932 );
and ( n15934 , n3892 , n4362 );
and ( n15935 , n4367 , n3903 );
and ( n15936 , n15934 , n15935 );
and ( n15937 , n15933 , n15936 );
and ( n15938 , n10886 , n13889 );
and ( n15939 , n15936 , n15938 );
and ( n15940 , n15933 , n15938 );
or ( n15941 , n15937 , n15939 , n15940 );
and ( n15942 , n11116 , n2923 );
and ( n15943 , n5091 , n3288 );
and ( n15944 , n15942 , n15943 );
and ( n15945 , n4989 , n3449 );
and ( n15946 , n15943 , n15945 );
and ( n15947 , n15942 , n15945 );
or ( n15948 , n15944 , n15946 , n15947 );
and ( n15949 , n2928 , n11111 );
and ( n15950 , n3293 , n5086 );
and ( n15951 , n15949 , n15950 );
and ( n15952 , n3454 , n4982 );
and ( n15953 , n15950 , n15952 );
and ( n15954 , n15949 , n15952 );
or ( n15955 , n15951 , n15953 , n15954 );
and ( n15956 , n15948 , n15955 );
and ( n15957 , n15941 , n15956 );
and ( n15958 , n15930 , n15957 );
xor ( n15959 , n15773 , n15776 );
xor ( n15960 , n15959 , n15778 );
xor ( n15961 , n15749 , n15752 );
xor ( n15962 , n15961 , n15754 );
and ( n15963 , n15960 , n15962 );
and ( n15964 , n15957 , n15963 );
and ( n15965 , n15930 , n15963 );
or ( n15966 , n15958 , n15964 , n15965 );
and ( n15967 , n3728 , n4362 );
and ( n15968 , n4367 , n3739 );
and ( n15969 , n15967 , n15968 );
and ( n15970 , n5091 , n3146 );
xor ( n15971 , n10271 , n10595 );
buf ( n15972 , n15971 );
buf ( n15973 , n15972 );
buf ( n15974 , n15973 );
and ( n15975 , n15970 , n15974 );
and ( n15976 , n4579 , n15408 );
and ( n15977 , n15974 , n15976 );
and ( n15978 , n15970 , n15976 );
or ( n15979 , n15975 , n15977 , n15978 );
and ( n15980 , n15969 , n15979 );
xor ( n15981 , n15797 , n15798 );
xor ( n15982 , n15981 , n15802 );
and ( n15983 , n15979 , n15982 );
and ( n15984 , n15969 , n15982 );
or ( n15985 , n15980 , n15983 , n15984 );
xor ( n15986 , n15840 , n15841 );
xor ( n15987 , n15986 , n15843 );
not ( n15988 , n15772 );
and ( n15989 , n15987 , n15988 );
xor ( n15990 , n15795 , n15796 );
and ( n15991 , n15988 , n15990 );
and ( n15992 , n15987 , n15990 );
or ( n15993 , n15989 , n15991 , n15992 );
xor ( n15994 , n15747 , n15748 );
xor ( n15995 , n15750 , n15751 );
and ( n15996 , n15994 , n15995 );
xor ( n15997 , n15848 , n15849 );
and ( n15998 , n15995 , n15997 );
and ( n15999 , n15994 , n15997 );
or ( n16000 , n15996 , n15998 , n15999 );
and ( n16001 , n15993 , n16000 );
xor ( n16002 , n15967 , n15968 );
xor ( n16003 , n15774 , n15775 );
and ( n16004 , n16002 , n16003 );
and ( n16005 , n3151 , n10869 );
and ( n16006 , n10862 , n3146 );
and ( n16007 , n16005 , n16006 );
and ( n16008 , n16003 , n16007 );
and ( n16009 , n16002 , n16007 );
or ( n16010 , n16004 , n16008 , n16009 );
and ( n16011 , n16000 , n16010 );
and ( n16012 , n15993 , n16010 );
or ( n16013 , n16001 , n16011 , n16012 );
and ( n16014 , n15985 , n16013 );
xor ( n16015 , n15812 , n15814 );
xor ( n16016 , n16015 , n15816 );
xor ( n16017 , n15820 , n15821 );
xor ( n16018 , n16017 , n15823 );
and ( n16019 , n16016 , n16018 );
xor ( n16020 , n15828 , n15829 );
xor ( n16021 , n16020 , n15831 );
and ( n16022 , n16018 , n16021 );
and ( n16023 , n16016 , n16021 );
or ( n16024 , n16019 , n16022 , n16023 );
and ( n16025 , n16013 , n16024 );
and ( n16026 , n15985 , n16024 );
or ( n16027 , n16014 , n16025 , n16026 );
and ( n16028 , n15966 , n16027 );
xor ( n16029 , n15790 , n15793 );
xor ( n16030 , n16029 , n15805 );
xor ( n16031 , n15819 , n15826 );
xor ( n16032 , n16031 , n15834 );
and ( n16033 , n16030 , n16032 );
xor ( n16034 , n15853 , n15855 );
xor ( n16035 , n16034 , n15858 );
and ( n16036 , n16032 , n16035 );
and ( n16037 , n16030 , n16035 );
or ( n16038 , n16033 , n16036 , n16037 );
and ( n16039 , n16027 , n16038 );
and ( n16040 , n15966 , n16038 );
or ( n16041 , n16028 , n16039 , n16040 );
and ( n16042 , n15928 , n16041 );
and ( n16043 , n15912 , n16041 );
or ( n16044 , n15929 , n16042 , n16043 );
and ( n16045 , n15910 , n16044 );
xor ( n16046 , n15768 , n15770 );
xor ( n16047 , n16046 , n15783 );
xor ( n16048 , n15808 , n15837 );
xor ( n16049 , n16048 , n15861 );
and ( n16050 , n16047 , n16049 );
xor ( n16051 , n15869 , n15871 );
xor ( n16052 , n16051 , n15874 );
and ( n16053 , n16049 , n16052 );
and ( n16054 , n16047 , n16052 );
or ( n16055 , n16050 , n16053 , n16054 );
xor ( n16056 , n15717 , n15718 );
xor ( n16057 , n16056 , n15732 );
and ( n16058 , n16055 , n16057 );
xor ( n16059 , n15766 , n15786 );
xor ( n16060 , n16059 , n15864 );
and ( n16061 , n16057 , n16060 );
and ( n16062 , n16055 , n16060 );
or ( n16063 , n16058 , n16061 , n16062 );
and ( n16064 , n16044 , n16063 );
and ( n16065 , n15910 , n16063 );
or ( n16066 , n16045 , n16064 , n16065 );
and ( n16067 , n15907 , n16066 );
and ( n16068 , n15905 , n16066 );
or ( n16069 , n15908 , n16067 , n16068 );
xor ( n16070 , n15709 , n15894 );
xor ( n16071 , n16070 , n15897 );
and ( n16072 , n16069 , n16071 );
xor ( n16073 , n15711 , n15738 );
xor ( n16074 , n16073 , n15891 );
xor ( n16075 , n15713 , n15714 );
xor ( n16076 , n16075 , n15735 );
xor ( n16077 , n15867 , n15885 );
xor ( n16078 , n16077 , n15888 );
and ( n16079 , n16076 , n16078 );
xor ( n16080 , n15877 , n15879 );
xor ( n16081 , n16080 , n15882 );
xor ( n16082 , n15839 , n15846 );
xor ( n16083 , n16082 , n15850 );
xor ( n16084 , n15941 , n15956 );
and ( n16085 , n16083 , n16084 );
xor ( n16086 , n15960 , n15962 );
and ( n16087 , n16084 , n16086 );
and ( n16088 , n16083 , n16086 );
or ( n16089 , n16085 , n16087 , n16088 );
and ( n16090 , n3151 , n11111 );
and ( n16091 , n11116 , n3146 );
and ( n16092 , n16090 , n16091 );
and ( n16093 , n10886 , n14454 );
and ( n16094 , n16092 , n16093 );
and ( n16095 , n4721 , n15408 );
and ( n16096 , n16093 , n16095 );
and ( n16097 , n16092 , n16095 );
or ( n16098 , n16094 , n16096 , n16097 );
and ( n16099 , n3892 , n4734 );
and ( n16100 , n4739 , n3903 );
and ( n16101 , n16099 , n16100 );
and ( n16102 , n10933 , n13889 );
and ( n16103 , n16101 , n16102 );
and ( n16104 , n4579 , n15801 );
and ( n16105 , n16102 , n16104 );
and ( n16106 , n16101 , n16104 );
or ( n16107 , n16103 , n16105 , n16106 );
and ( n16108 , n16098 , n16107 );
and ( n16109 , n3293 , n10869 );
and ( n16110 , n10862 , n3288 );
and ( n16111 , n16109 , n16110 );
and ( n16112 , n3454 , n5086 );
and ( n16113 , n5091 , n3449 );
and ( n16114 , n16112 , n16113 );
and ( n16115 , n16111 , n16114 );
and ( n16116 , n5177 , n14897 );
and ( n16117 , n16114 , n16116 );
and ( n16118 , n16111 , n16116 );
or ( n16119 , n16115 , n16117 , n16118 );
and ( n16120 , n16107 , n16119 );
and ( n16121 , n16098 , n16119 );
or ( n16122 , n16108 , n16120 , n16121 );
buf ( n16123 , n4138 );
buf ( n16124 , n16123 );
xor ( n16125 , n15970 , n15974 );
xor ( n16126 , n16125 , n15976 );
and ( n16127 , n16124 , n16126 );
xor ( n16128 , n15933 , n15936 );
xor ( n16129 , n16128 , n15938 );
and ( n16130 , n16126 , n16129 );
and ( n16131 , n16124 , n16129 );
or ( n16132 , n16127 , n16130 , n16131 );
and ( n16133 , n16122 , n16132 );
xor ( n16134 , n15948 , n15955 );
buf ( n16135 , n4136 );
buf ( n16136 , n16135 );
and ( n16137 , n4385 , n16136 );
and ( n16138 , n4150 , n4362 );
and ( n16139 , n4367 , n4161 );
and ( n16140 , n16138 , n16139 );
and ( n16141 , n16137 , n16140 );
and ( n16142 , n16134 , n16141 );
xor ( n16143 , n15942 , n15943 );
xor ( n16144 , n16143 , n15945 );
xor ( n16145 , n15949 , n15950 );
xor ( n16146 , n16145 , n15952 );
and ( n16147 , n16144 , n16146 );
and ( n16148 , n16141 , n16147 );
and ( n16149 , n16134 , n16147 );
or ( n16150 , n16142 , n16148 , n16149 );
and ( n16151 , n16132 , n16150 );
and ( n16152 , n16122 , n16150 );
or ( n16153 , n16133 , n16151 , n16152 );
and ( n16154 , n16089 , n16153 );
xor ( n16155 , n16005 , n16006 );
xor ( n16156 , n15931 , n15932 );
and ( n16157 , n16155 , n16156 );
xor ( n16158 , n15934 , n15935 );
and ( n16159 , n16156 , n16158 );
and ( n16160 , n16155 , n16158 );
or ( n16161 , n16157 , n16159 , n16160 );
xor ( n16162 , n15987 , n15988 );
xor ( n16163 , n16162 , n15990 );
and ( n16164 , n16161 , n16163 );
xor ( n16165 , n15994 , n15995 );
xor ( n16166 , n16165 , n15997 );
and ( n16167 , n16163 , n16166 );
and ( n16168 , n16161 , n16166 );
or ( n16169 , n16164 , n16167 , n16168 );
xor ( n16170 , n15969 , n15979 );
xor ( n16171 , n16170 , n15982 );
and ( n16172 , n16169 , n16171 );
xor ( n16173 , n15993 , n16000 );
xor ( n16174 , n16173 , n16010 );
and ( n16175 , n16171 , n16174 );
and ( n16176 , n16169 , n16174 );
or ( n16177 , n16172 , n16175 , n16176 );
and ( n16178 , n16153 , n16177 );
and ( n16179 , n16089 , n16177 );
or ( n16180 , n16154 , n16178 , n16179 );
xor ( n16181 , n15917 , n15919 );
xor ( n16182 , n16181 , n15922 );
xor ( n16183 , n15930 , n15957 );
xor ( n16184 , n16183 , n15963 );
and ( n16185 , n16182 , n16184 );
xor ( n16186 , n15985 , n16013 );
xor ( n16187 , n16186 , n16024 );
and ( n16188 , n16184 , n16187 );
and ( n16189 , n16182 , n16187 );
or ( n16190 , n16185 , n16188 , n16189 );
and ( n16191 , n16180 , n16190 );
xor ( n16192 , n15913 , n15914 );
xor ( n16193 , n16192 , n15925 );
and ( n16194 , n16190 , n16193 );
and ( n16195 , n16180 , n16193 );
or ( n16196 , n16191 , n16194 , n16195 );
and ( n16197 , n16081 , n16196 );
xor ( n16198 , n15912 , n15928 );
xor ( n16199 , n16198 , n16041 );
and ( n16200 , n16196 , n16199 );
and ( n16201 , n16081 , n16199 );
or ( n16202 , n16197 , n16200 , n16201 );
and ( n16203 , n16078 , n16202 );
and ( n16204 , n16076 , n16202 );
or ( n16205 , n16079 , n16203 , n16204 );
and ( n16206 , n16074 , n16205 );
xor ( n16207 , n15905 , n15907 );
xor ( n16208 , n16207 , n16066 );
and ( n16209 , n16205 , n16208 );
and ( n16210 , n16074 , n16208 );
or ( n16211 , n16206 , n16209 , n16210 );
and ( n16212 , n16071 , n16211 );
and ( n16213 , n16069 , n16211 );
or ( n16214 , n16072 , n16212 , n16213 );
and ( n16215 , n15902 , n16214 );
and ( n16216 , n15900 , n16214 );
or ( n16217 , n15903 , n16215 , n16216 );
and ( n16218 , n15706 , n16217 );
and ( n16219 , n15704 , n16217 );
or ( n16220 , n15707 , n16218 , n16219 );
and ( n16221 , n15702 , n16220 );
xor ( n16222 , n15702 , n16220 );
xor ( n16223 , n15704 , n15706 );
xor ( n16224 , n16223 , n16217 );
xor ( n16225 , n15900 , n15902 );
xor ( n16226 , n16225 , n16214 );
xor ( n16227 , n16069 , n16071 );
xor ( n16228 , n16227 , n16211 );
xor ( n16229 , n15910 , n16044 );
xor ( n16230 , n16229 , n16063 );
xor ( n16231 , n16055 , n16057 );
xor ( n16232 , n16231 , n16060 );
xor ( n16233 , n15966 , n16027 );
xor ( n16234 , n16233 , n16038 );
xor ( n16235 , n16047 , n16049 );
xor ( n16236 , n16235 , n16052 );
and ( n16237 , n16234 , n16236 );
xor ( n16238 , n16030 , n16032 );
xor ( n16239 , n16238 , n16035 );
xor ( n16240 , n16016 , n16018 );
xor ( n16241 , n16240 , n16021 );
and ( n16242 , n4579 , n16136 );
and ( n16243 , n4150 , n4734 );
and ( n16244 , n4739 , n4161 );
and ( n16245 , n16243 , n16244 );
and ( n16246 , n16242 , n16245 );
xor ( n16247 , n10474 , n10593 );
buf ( n16248 , n16247 );
buf ( n16249 , n16248 );
buf ( n16250 , n16249 );
or ( n16251 , n16246 , n16250 );
and ( n16252 , n5177 , n14454 );
and ( n16253 , n16251 , n16252 );
and ( n16254 , n16241 , n16253 );
xor ( n16255 , n16002 , n16003 );
xor ( n16256 , n16255 , n16007 );
xor ( n16257 , n16098 , n16107 );
xor ( n16258 , n16257 , n16119 );
and ( n16259 , n16256 , n16258 );
xor ( n16260 , n16092 , n16093 );
xor ( n16261 , n16260 , n16095 );
xor ( n16262 , n16101 , n16102 );
xor ( n16263 , n16262 , n16104 );
and ( n16264 , n16261 , n16263 );
xor ( n16265 , n16111 , n16114 );
xor ( n16266 , n16265 , n16116 );
and ( n16267 , n16263 , n16266 );
and ( n16268 , n16261 , n16266 );
or ( n16269 , n16264 , n16267 , n16268 );
and ( n16270 , n16258 , n16269 );
and ( n16271 , n16256 , n16269 );
or ( n16272 , n16259 , n16270 , n16271 );
and ( n16273 , n16253 , n16272 );
and ( n16274 , n16241 , n16272 );
or ( n16275 , n16254 , n16273 , n16274 );
and ( n16276 , n16239 , n16275 );
and ( n16277 , n3728 , n4982 );
and ( n16278 , n4989 , n3739 );
and ( n16279 , n16277 , n16278 );
xor ( n16280 , n16137 , n16140 );
and ( n16281 , n16279 , n16280 );
buf ( n16282 , n16281 );
xor ( n16283 , n16144 , n16146 );
and ( n16284 , n3728 , n5086 );
and ( n16285 , n5091 , n3739 );
and ( n16286 , n16284 , n16285 );
and ( n16287 , n5177 , n15408 );
and ( n16288 , n16286 , n16287 );
and ( n16289 , n4721 , n15801 );
and ( n16290 , n16287 , n16289 );
and ( n16291 , n16286 , n16289 );
or ( n16292 , n16288 , n16290 , n16291 );
and ( n16293 , n16283 , n16292 );
and ( n16294 , n3293 , n11111 );
and ( n16295 , n11116 , n3288 );
and ( n16296 , n16294 , n16295 );
and ( n16297 , n3892 , n4982 );
and ( n16298 , n4989 , n3903 );
and ( n16299 , n16297 , n16298 );
and ( n16300 , n16296 , n16299 );
and ( n16301 , n10886 , n14897 );
and ( n16302 , n16299 , n16301 );
and ( n16303 , n16296 , n16301 );
or ( n16304 , n16300 , n16302 , n16303 );
and ( n16305 , n16292 , n16304 );
and ( n16306 , n16283 , n16304 );
or ( n16307 , n16293 , n16305 , n16306 );
and ( n16308 , n16282 , n16307 );
xor ( n16309 , n10477 , n10591 );
buf ( n16310 , n16309 );
buf ( n16311 , n16310 );
buf ( n16312 , n16311 );
and ( n16313 , n10933 , n14454 );
and ( n16314 , n16312 , n16313 );
xor ( n16315 , n16090 , n16091 );
and ( n16316 , n16313 , n16315 );
and ( n16317 , n16312 , n16315 );
or ( n16318 , n16314 , n16316 , n16317 );
xor ( n16319 , n16109 , n16110 );
xor ( n16320 , n16112 , n16113 );
and ( n16321 , n16319 , n16320 );
xor ( n16322 , n16277 , n16278 );
and ( n16323 , n16320 , n16322 );
and ( n16324 , n16319 , n16322 );
or ( n16325 , n16321 , n16323 , n16324 );
and ( n16326 , n16318 , n16325 );
xor ( n16327 , n16099 , n16100 );
xor ( n16328 , n16138 , n16139 );
and ( n16329 , n16327 , n16328 );
and ( n16330 , n3454 , n10869 );
and ( n16331 , n10862 , n3449 );
and ( n16332 , n16330 , n16331 );
and ( n16333 , n16328 , n16332 );
and ( n16334 , n16327 , n16332 );
or ( n16335 , n16329 , n16333 , n16334 );
and ( n16336 , n16325 , n16335 );
and ( n16337 , n16318 , n16335 );
or ( n16338 , n16326 , n16336 , n16337 );
and ( n16339 , n16307 , n16338 );
and ( n16340 , n16282 , n16338 );
or ( n16341 , n16308 , n16339 , n16340 );
xor ( n16342 , n16124 , n16126 );
xor ( n16343 , n16342 , n16129 );
xor ( n16344 , n16134 , n16141 );
xor ( n16345 , n16344 , n16147 );
and ( n16346 , n16343 , n16345 );
xor ( n16347 , n16161 , n16163 );
xor ( n16348 , n16347 , n16166 );
and ( n16349 , n16345 , n16348 );
and ( n16350 , n16343 , n16348 );
or ( n16351 , n16346 , n16349 , n16350 );
and ( n16352 , n16341 , n16351 );
xor ( n16353 , n16083 , n16084 );
xor ( n16354 , n16353 , n16086 );
and ( n16355 , n16351 , n16354 );
and ( n16356 , n16341 , n16354 );
or ( n16357 , n16352 , n16355 , n16356 );
and ( n16358 , n16275 , n16357 );
and ( n16359 , n16239 , n16357 );
or ( n16360 , n16276 , n16358 , n16359 );
and ( n16361 , n16236 , n16360 );
and ( n16362 , n16234 , n16360 );
or ( n16363 , n16237 , n16361 , n16362 );
and ( n16364 , n16232 , n16363 );
xor ( n16365 , n16081 , n16196 );
xor ( n16366 , n16365 , n16199 );
and ( n16367 , n16363 , n16366 );
and ( n16368 , n16232 , n16366 );
or ( n16369 , n16364 , n16367 , n16368 );
and ( n16370 , n16230 , n16369 );
xor ( n16371 , n16076 , n16078 );
xor ( n16372 , n16371 , n16202 );
and ( n16373 , n16369 , n16372 );
and ( n16374 , n16230 , n16372 );
or ( n16375 , n16370 , n16373 , n16374 );
xor ( n16376 , n16074 , n16205 );
xor ( n16377 , n16376 , n16208 );
and ( n16378 , n16375 , n16377 );
xor ( n16379 , n16375 , n16377 );
xor ( n16380 , n16230 , n16369 );
xor ( n16381 , n16380 , n16372 );
xor ( n16382 , n16180 , n16190 );
xor ( n16383 , n16382 , n16193 );
xor ( n16384 , n16089 , n16153 );
xor ( n16385 , n16384 , n16177 );
xor ( n16386 , n16182 , n16184 );
xor ( n16387 , n16386 , n16187 );
and ( n16388 , n16385 , n16387 );
xor ( n16389 , n16122 , n16132 );
xor ( n16390 , n16389 , n16150 );
xor ( n16391 , n16169 , n16171 );
xor ( n16392 , n16391 , n16174 );
and ( n16393 , n16390 , n16392 );
xor ( n16394 , n16251 , n16252 );
xor ( n16395 , n16155 , n16156 );
xor ( n16396 , n16395 , n16158 );
xor ( n16397 , n16261 , n16263 );
xor ( n16398 , n16397 , n16266 );
and ( n16399 , n16396 , n16398 );
xnor ( n16400 , n16246 , n16250 );
and ( n16401 , n16398 , n16400 );
and ( n16402 , n16396 , n16400 );
or ( n16403 , n16399 , n16401 , n16402 );
and ( n16404 , n16394 , n16403 );
xor ( n16405 , n16286 , n16287 );
xor ( n16406 , n16405 , n16289 );
xor ( n16407 , n16296 , n16299 );
xor ( n16408 , n16407 , n16301 );
and ( n16409 , n16406 , n16408 );
buf ( n16410 , n4385 );
buf ( n16411 , n16410 );
xor ( n16412 , n16242 , n16245 );
and ( n16413 , n16411 , n16412 );
and ( n16414 , n4721 , n16136 );
and ( n16415 , n4150 , n4982 );
and ( n16416 , n4989 , n4161 );
and ( n16417 , n16415 , n16416 );
and ( n16418 , n16414 , n16417 );
and ( n16419 , n16412 , n16418 );
and ( n16420 , n16411 , n16418 );
or ( n16421 , n16413 , n16419 , n16420 );
and ( n16422 , n16409 , n16421 );
buf ( n16423 , n4383 );
buf ( n16424 , n16423 );
and ( n16425 , n4579 , n16424 );
and ( n16426 , n4367 , n4734 );
and ( n16427 , n4739 , n4362 );
and ( n16428 , n16426 , n16427 );
and ( n16429 , n16425 , n16428 );
xor ( n16430 , n16294 , n16295 );
xor ( n16431 , n16330 , n16331 );
and ( n16432 , n16430 , n16431 );
xor ( n16433 , n16284 , n16285 );
and ( n16434 , n16431 , n16433 );
and ( n16435 , n16430 , n16433 );
or ( n16436 , n16432 , n16434 , n16435 );
and ( n16437 , n16429 , n16436 );
xor ( n16438 , n16297 , n16298 );
xor ( n16439 , n16243 , n16244 );
and ( n16440 , n16438 , n16439 );
buf ( n16441 , n16440 );
and ( n16442 , n16436 , n16441 );
and ( n16443 , n16429 , n16441 );
or ( n16444 , n16437 , n16442 , n16443 );
and ( n16445 , n16421 , n16444 );
and ( n16446 , n16409 , n16444 );
or ( n16447 , n16422 , n16445 , n16446 );
and ( n16448 , n16403 , n16447 );
and ( n16449 , n16394 , n16447 );
or ( n16450 , n16404 , n16448 , n16449 );
and ( n16451 , n16392 , n16450 );
and ( n16452 , n16390 , n16450 );
or ( n16453 , n16393 , n16451 , n16452 );
and ( n16454 , n16387 , n16453 );
and ( n16455 , n16385 , n16453 );
or ( n16456 , n16388 , n16454 , n16455 );
and ( n16457 , n16383 , n16456 );
xor ( n16458 , n16234 , n16236 );
xor ( n16459 , n16458 , n16360 );
and ( n16460 , n16456 , n16459 );
and ( n16461 , n16383 , n16459 );
or ( n16462 , n16457 , n16460 , n16461 );
xor ( n16463 , n16232 , n16363 );
xor ( n16464 , n16463 , n16366 );
and ( n16465 , n16462 , n16464 );
xor ( n16466 , n16312 , n16313 );
xor ( n16467 , n16466 , n16315 );
xor ( n16468 , n16319 , n16320 );
xor ( n16469 , n16468 , n16322 );
and ( n16470 , n16467 , n16469 );
xor ( n16471 , n16327 , n16328 );
xor ( n16472 , n16471 , n16332 );
and ( n16473 , n16469 , n16472 );
and ( n16474 , n16467 , n16472 );
or ( n16475 , n16470 , n16473 , n16474 );
buf ( n16476 , n16279 );
xor ( n16477 , n16476 , n16280 );
and ( n16478 , n16475 , n16477 );
xor ( n16479 , n16283 , n16292 );
xor ( n16480 , n16479 , n16304 );
and ( n16481 , n16477 , n16480 );
and ( n16482 , n16475 , n16480 );
or ( n16483 , n16478 , n16481 , n16482 );
xor ( n16484 , n16256 , n16258 );
xor ( n16485 , n16484 , n16269 );
and ( n16486 , n16483 , n16485 );
xor ( n16487 , n16282 , n16307 );
xor ( n16488 , n16487 , n16338 );
and ( n16489 , n16485 , n16488 );
and ( n16490 , n16483 , n16488 );
or ( n16491 , n16486 , n16489 , n16490 );
xor ( n16492 , n16241 , n16253 );
xor ( n16493 , n16492 , n16272 );
and ( n16494 , n16491 , n16493 );
xor ( n16495 , n16341 , n16351 );
xor ( n16496 , n16495 , n16354 );
and ( n16497 , n16493 , n16496 );
and ( n16498 , n16491 , n16496 );
or ( n16499 , n16494 , n16497 , n16498 );
xor ( n16500 , n16239 , n16275 );
xor ( n16501 , n16500 , n16357 );
and ( n16502 , n16499 , n16501 );
xor ( n16503 , n16343 , n16345 );
xor ( n16504 , n16503 , n16348 );
xor ( n16505 , n16318 , n16325 );
xor ( n16506 , n16505 , n16335 );
and ( n16507 , n3728 , n10869 );
and ( n16508 , n10862 , n3739 );
and ( n16509 , n16507 , n16508 );
and ( n16510 , n10886 , n15408 );
and ( n16511 , n16509 , n16510 );
and ( n16512 , n5177 , n15801 );
and ( n16513 , n16510 , n16512 );
and ( n16514 , n16509 , n16512 );
or ( n16515 , n16511 , n16513 , n16514 );
and ( n16516 , n4721 , n16424 );
and ( n16517 , n4367 , n4982 );
and ( n16518 , n4989 , n4362 );
and ( n16519 , n16517 , n16518 );
and ( n16520 , n16516 , n16519 );
and ( n16521 , n3454 , n11111 );
and ( n16522 , n11116 , n3449 );
and ( n16523 , n16521 , n16522 );
and ( n16524 , n16520 , n16523 );
and ( n16525 , n10933 , n14897 );
and ( n16526 , n16523 , n16525 );
and ( n16527 , n16520 , n16525 );
or ( n16528 , n16524 , n16526 , n16527 );
or ( n16529 , n16515 , n16528 );
and ( n16530 , n16506 , n16529 );
xor ( n16531 , n16406 , n16408 );
and ( n16532 , n5177 , n16136 );
and ( n16533 , n4150 , n5086 );
and ( n16534 , n5091 , n4161 );
and ( n16535 , n16533 , n16534 );
and ( n16536 , n16532 , n16535 );
xor ( n16537 , n10480 , n10589 );
buf ( n16538 , n16537 );
buf ( n16539 , n16538 );
buf ( n16540 , n16539 );
or ( n16541 , n16536 , n16540 );
and ( n16542 , n16531 , n16541 );
xor ( n16543 , n16414 , n16417 );
xor ( n16544 , n16425 , n16428 );
and ( n16545 , n16543 , n16544 );
xor ( n16546 , n16521 , n16522 );
xor ( n16547 , n16507 , n16508 );
and ( n16548 , n16546 , n16547 );
and ( n16549 , n3892 , n5086 );
and ( n16550 , n5091 , n3903 );
xor ( n16551 , n16549 , n16550 );
and ( n16552 , n16547 , n16551 );
and ( n16553 , n16546 , n16551 );
or ( n16554 , n16548 , n16552 , n16553 );
and ( n16555 , n16544 , n16554 );
and ( n16556 , n16543 , n16554 );
or ( n16557 , n16545 , n16555 , n16556 );
and ( n16558 , n16541 , n16557 );
and ( n16559 , n16531 , n16557 );
or ( n16560 , n16542 , n16558 , n16559 );
and ( n16561 , n16529 , n16560 );
and ( n16562 , n16506 , n16560 );
or ( n16563 , n16530 , n16561 , n16562 );
and ( n16564 , n16504 , n16563 );
xor ( n16565 , n16411 , n16412 );
xor ( n16566 , n16565 , n16418 );
xor ( n16567 , n16429 , n16436 );
xor ( n16568 , n16567 , n16441 );
and ( n16569 , n16566 , n16568 );
xor ( n16570 , n16467 , n16469 );
xor ( n16571 , n16570 , n16472 );
and ( n16572 , n16568 , n16571 );
and ( n16573 , n16566 , n16571 );
or ( n16574 , n16569 , n16572 , n16573 );
xor ( n16575 , n16396 , n16398 );
xor ( n16576 , n16575 , n16400 );
and ( n16577 , n16574 , n16576 );
xor ( n16578 , n16409 , n16421 );
xor ( n16579 , n16578 , n16444 );
and ( n16580 , n16576 , n16579 );
and ( n16581 , n16574 , n16579 );
or ( n16582 , n16577 , n16580 , n16581 );
and ( n16583 , n16563 , n16582 );
and ( n16584 , n16504 , n16582 );
or ( n16585 , n16564 , n16583 , n16584 );
xor ( n16586 , n16390 , n16392 );
xor ( n16587 , n16586 , n16450 );
and ( n16588 , n16585 , n16587 );
xor ( n16589 , n16491 , n16493 );
xor ( n16590 , n16589 , n16496 );
and ( n16591 , n16587 , n16590 );
and ( n16592 , n16585 , n16590 );
or ( n16593 , n16588 , n16591 , n16592 );
and ( n16594 , n16501 , n16593 );
and ( n16595 , n16499 , n16593 );
or ( n16596 , n16502 , n16594 , n16595 );
xor ( n16597 , n16383 , n16456 );
xor ( n16598 , n16597 , n16459 );
and ( n16599 , n16596 , n16598 );
xor ( n16600 , n16385 , n16387 );
xor ( n16601 , n16600 , n16453 );
xor ( n16602 , n16499 , n16501 );
xor ( n16603 , n16602 , n16593 );
and ( n16604 , n16601 , n16603 );
xor ( n16605 , n16394 , n16403 );
xor ( n16606 , n16605 , n16447 );
xor ( n16607 , n16483 , n16485 );
xor ( n16608 , n16607 , n16488 );
and ( n16609 , n16606 , n16608 );
xor ( n16610 , n16475 , n16477 );
xor ( n16611 , n16610 , n16480 );
xnor ( n16612 , n16515 , n16528 );
xnor ( n16613 , n16536 , n16540 );
and ( n16614 , n3728 , n11111 );
and ( n16615 , n11116 , n3739 );
and ( n16616 , n16614 , n16615 );
and ( n16617 , n10933 , n15408 );
and ( n16618 , n16616 , n16617 );
and ( n16619 , n10886 , n15801 );
and ( n16620 , n16617 , n16619 );
and ( n16621 , n16616 , n16619 );
or ( n16622 , n16618 , n16620 , n16621 );
and ( n16623 , n16613 , n16622 );
xor ( n16624 , n16509 , n16510 );
xor ( n16625 , n16624 , n16512 );
and ( n16626 , n16622 , n16625 );
and ( n16627 , n16613 , n16625 );
or ( n16628 , n16623 , n16626 , n16627 );
and ( n16629 , n16612 , n16628 );
and ( n16630 , n10886 , n16136 );
and ( n16631 , n4150 , n10869 );
and ( n16632 , n10862 , n4161 );
and ( n16633 , n16631 , n16632 );
and ( n16634 , n16630 , n16633 );
buf ( n16635 , n4577 );
buf ( n16636 , n16635 );
and ( n16637 , n4721 , n16636 );
and ( n16638 , n4739 , n4982 );
and ( n16639 , n4989 , n4734 );
and ( n16640 , n16638 , n16639 );
and ( n16641 , n16637 , n16640 );
or ( n16642 , n16634 , n16641 );
and ( n16643 , n16549 , n16550 );
and ( n16644 , n16642 , n16643 );
and ( n16645 , n16628 , n16644 );
and ( n16646 , n16612 , n16644 );
or ( n16647 , n16629 , n16645 , n16646 );
and ( n16648 , n16611 , n16647 );
xor ( n16649 , n16430 , n16431 );
xor ( n16650 , n16649 , n16433 );
xor ( n16651 , n16438 , n16439 );
buf ( n16652 , n16651 );
and ( n16653 , n16650 , n16652 );
xor ( n16654 , n16520 , n16523 );
xor ( n16655 , n16654 , n16525 );
and ( n16656 , n16652 , n16655 );
and ( n16657 , n16650 , n16655 );
or ( n16658 , n16653 , n16656 , n16657 );
and ( n16659 , n4367 , n5086 );
and ( n16660 , n5091 , n4362 );
and ( n16661 , n16659 , n16660 );
buf ( n16662 , n4739 );
and ( n16663 , n16661 , n16662 );
and ( n16664 , n5177 , n16424 );
buf ( n16665 , n4579 );
and ( n16666 , n16664 , n16665 );
and ( n16667 , n16663 , n16666 );
xor ( n16668 , n16415 , n16416 );
xor ( n16669 , n16426 , n16427 );
and ( n16670 , n16668 , n16669 );
xor ( n16671 , n16532 , n16535 );
and ( n16672 , n16669 , n16671 );
and ( n16673 , n16668 , n16671 );
or ( n16674 , n16670 , n16672 , n16673 );
and ( n16675 , n16667 , n16674 );
xor ( n16676 , n16516 , n16519 );
and ( n16677 , n3892 , n11111 );
and ( n16678 , n10933 , n16136 );
and ( n16679 , n16677 , n16678 );
and ( n16680 , n10886 , n16424 );
and ( n16681 , n16678 , n16680 );
and ( n16682 , n16677 , n16680 );
or ( n16683 , n16679 , n16681 , n16682 );
and ( n16684 , n3892 , n10869 );
and ( n16685 , n16683 , n16684 );
and ( n16686 , n16676 , n16685 );
and ( n16687 , n10862 , n3903 );
xor ( n16688 , n16614 , n16615 );
and ( n16689 , n16687 , n16688 );
xor ( n16690 , n16533 , n16534 );
and ( n16691 , n16688 , n16690 );
and ( n16692 , n16687 , n16690 );
or ( n16693 , n16689 , n16691 , n16692 );
and ( n16694 , n16685 , n16693 );
and ( n16695 , n16676 , n16693 );
or ( n16696 , n16686 , n16694 , n16695 );
and ( n16697 , n16674 , n16696 );
and ( n16698 , n16667 , n16696 );
or ( n16699 , n16675 , n16697 , n16698 );
and ( n16700 , n16658 , n16699 );
xor ( n16701 , n16531 , n16541 );
xor ( n16702 , n16701 , n16557 );
and ( n16703 , n16699 , n16702 );
and ( n16704 , n16658 , n16702 );
or ( n16705 , n16700 , n16703 , n16704 );
and ( n16706 , n16647 , n16705 );
and ( n16707 , n16611 , n16705 );
or ( n16708 , n16648 , n16706 , n16707 );
and ( n16709 , n16608 , n16708 );
and ( n16710 , n16606 , n16708 );
or ( n16711 , n16609 , n16709 , n16710 );
xor ( n16712 , n16585 , n16587 );
xor ( n16713 , n16712 , n16590 );
and ( n16714 , n16711 , n16713 );
xor ( n16715 , n16504 , n16563 );
xor ( n16716 , n16715 , n16582 );
xor ( n16717 , n16506 , n16529 );
xor ( n16718 , n16717 , n16560 );
xor ( n16719 , n16574 , n16576 );
xor ( n16720 , n16719 , n16579 );
and ( n16721 , n16718 , n16720 );
xor ( n16722 , n16566 , n16568 );
xor ( n16723 , n16722 , n16571 );
xor ( n16724 , n16543 , n16544 );
xor ( n16725 , n16724 , n16554 );
xor ( n16726 , n16642 , n16643 );
and ( n16727 , n16725 , n16726 );
xor ( n16728 , n16661 , n16662 );
xor ( n16729 , n16664 , n16665 );
and ( n16730 , n16728 , n16729 );
xor ( n16731 , n10483 , n10587 );
buf ( n16732 , n16731 );
buf ( n16733 , n16732 );
buf ( n16734 , n16733 );
and ( n16735 , n16730 , n16734 );
and ( n16736 , n16726 , n16735 );
and ( n16737 , n16725 , n16735 );
or ( n16738 , n16727 , n16736 , n16737 );
and ( n16739 , n16723 , n16738 );
xor ( n16740 , n16546 , n16547 );
xor ( n16741 , n16740 , n16551 );
xor ( n16742 , n16663 , n16666 );
and ( n16743 , n16741 , n16742 );
and ( n16744 , n5177 , n16636 );
and ( n16745 , n4739 , n5086 );
and ( n16746 , n5091 , n4734 );
and ( n16747 , n16745 , n16746 );
and ( n16748 , n16744 , n16747 );
xor ( n16749 , n10486 , n10585 );
buf ( n16750 , n16749 );
buf ( n16751 , n16750 );
buf ( n16752 , n16751 );
and ( n16753 , n16748 , n16752 );
and ( n16754 , n16742 , n16753 );
and ( n16755 , n16741 , n16753 );
or ( n16756 , n16743 , n16754 , n16755 );
xor ( n16757 , n16517 , n16518 );
xor ( n16758 , n16683 , n16684 );
and ( n16759 , n16757 , n16758 );
xor ( n16760 , n16630 , n16633 );
and ( n16761 , n16758 , n16760 );
and ( n16762 , n16757 , n16760 );
or ( n16763 , n16759 , n16761 , n16762 );
xor ( n16764 , n16637 , n16640 );
and ( n16765 , n11116 , n4161 );
and ( n16766 , n10862 , n4362 );
and ( n16767 , n16765 , n16766 );
and ( n16768 , n4150 , n11111 );
and ( n16769 , n4367 , n10869 );
and ( n16770 , n16768 , n16769 );
and ( n16771 , n16767 , n16770 );
and ( n16772 , n16764 , n16771 );
xor ( n16773 , n16631 , n16632 );
xor ( n16774 , n16659 , n16660 );
and ( n16775 , n16773 , n16774 );
xor ( n16776 , n16638 , n16639 );
and ( n16777 , n16774 , n16776 );
and ( n16778 , n16773 , n16776 );
or ( n16779 , n16775 , n16777 , n16778 );
and ( n16780 , n16771 , n16779 );
and ( n16781 , n16764 , n16779 );
or ( n16782 , n16772 , n16780 , n16781 );
and ( n16783 , n16763 , n16782 );
xor ( n16784 , n16668 , n16669 );
xor ( n16785 , n16784 , n16671 );
and ( n16786 , n16782 , n16785 );
and ( n16787 , n16763 , n16785 );
or ( n16788 , n16783 , n16786 , n16787 );
and ( n16789 , n16756 , n16788 );
xor ( n16790 , n16650 , n16652 );
xor ( n16791 , n16790 , n16655 );
and ( n16792 , n16788 , n16791 );
and ( n16793 , n16756 , n16791 );
or ( n16794 , n16789 , n16792 , n16793 );
and ( n16795 , n16738 , n16794 );
and ( n16796 , n16723 , n16794 );
or ( n16797 , n16739 , n16795 , n16796 );
and ( n16798 , n16720 , n16797 );
and ( n16799 , n16718 , n16797 );
or ( n16800 , n16721 , n16798 , n16799 );
and ( n16801 , n16716 , n16800 );
xor ( n16802 , n16606 , n16608 );
xor ( n16803 , n16802 , n16708 );
and ( n16804 , n16800 , n16803 );
and ( n16805 , n16716 , n16803 );
or ( n16806 , n16801 , n16804 , n16805 );
and ( n16807 , n16713 , n16806 );
and ( n16808 , n16711 , n16806 );
or ( n16809 , n16714 , n16807 , n16808 );
and ( n16810 , n16603 , n16809 );
and ( n16811 , n16601 , n16809 );
or ( n16812 , n16604 , n16810 , n16811 );
and ( n16813 , n16598 , n16812 );
and ( n16814 , n16596 , n16812 );
or ( n16815 , n16599 , n16813 , n16814 );
and ( n16816 , n16464 , n16815 );
and ( n16817 , n16462 , n16815 );
or ( n16818 , n16465 , n16816 , n16817 );
and ( n16819 , n16381 , n16818 );
xor ( n16820 , n16381 , n16818 );
xor ( n16821 , n16462 , n16464 );
xor ( n16822 , n16821 , n16815 );
xor ( n16823 , n16596 , n16598 );
xor ( n16824 , n16823 , n16812 );
xor ( n16825 , n16601 , n16603 );
xor ( n16826 , n16825 , n16809 );
xor ( n16827 , n16711 , n16713 );
xor ( n16828 , n16827 , n16806 );
xor ( n16829 , n16611 , n16647 );
xor ( n16830 , n16829 , n16705 );
xor ( n16831 , n16612 , n16628 );
xor ( n16832 , n16831 , n16644 );
xor ( n16833 , n16658 , n16699 );
xor ( n16834 , n16833 , n16702 );
and ( n16835 , n16832 , n16834 );
xor ( n16836 , n16730 , n16734 );
xor ( n16837 , n16616 , n16617 );
xor ( n16838 , n16837 , n16619 );
and ( n16839 , n16836 , n16838 );
xnor ( n16840 , n16634 , n16641 );
and ( n16841 , n16838 , n16840 );
and ( n16842 , n16836 , n16840 );
or ( n16843 , n16839 , n16841 , n16842 );
xor ( n16844 , n16613 , n16622 );
xor ( n16845 , n16844 , n16625 );
and ( n16846 , n16843 , n16845 );
and ( n16847 , n16834 , n16846 );
and ( n16848 , n16832 , n16846 );
or ( n16849 , n16835 , n16847 , n16848 );
and ( n16850 , n16830 , n16849 );
xor ( n16851 , n16718 , n16720 );
xor ( n16852 , n16851 , n16797 );
and ( n16853 , n16849 , n16852 );
and ( n16854 , n16830 , n16852 );
or ( n16855 , n16850 , n16853 , n16854 );
xor ( n16856 , n16716 , n16800 );
xor ( n16857 , n16856 , n16803 );
and ( n16858 , n16855 , n16857 );
xor ( n16859 , n16667 , n16674 );
xor ( n16860 , n16859 , n16696 );
xor ( n16861 , n16676 , n16685 );
xor ( n16862 , n16861 , n16693 );
xor ( n16863 , n16748 , n16752 );
and ( n16864 , n10886 , n16636 );
and ( n16865 , n4739 , n10869 );
and ( n16866 , n10862 , n4734 );
and ( n16867 , n16865 , n16866 );
and ( n16868 , n16864 , n16867 );
xor ( n16869 , n10488 , n10584 );
buf ( n16870 , n16869 );
buf ( n16871 , n16870 );
buf ( n16872 , n16871 );
and ( n16873 , n16868 , n16872 );
and ( n16874 , n16863 , n16873 );
and ( n16875 , n10933 , n15801 );
and ( n16876 , n16873 , n16875 );
and ( n16877 , n16863 , n16875 );
or ( n16878 , n16874 , n16876 , n16877 );
and ( n16879 , n16862 , n16878 );
xor ( n16880 , n16687 , n16688 );
xor ( n16881 , n16880 , n16690 );
xor ( n16882 , n16728 , n16729 );
and ( n16883 , n16881 , n16882 );
xor ( n16884 , n16765 , n16766 );
xor ( n16885 , n16768 , n16769 );
and ( n16886 , n16884 , n16885 );
and ( n16887 , n11116 , n3903 );
and ( n16888 , n16886 , n16887 );
and ( n16889 , n16882 , n16888 );
and ( n16890 , n16881 , n16888 );
or ( n16891 , n16883 , n16889 , n16890 );
and ( n16892 , n16878 , n16891 );
and ( n16893 , n16862 , n16891 );
or ( n16894 , n16879 , n16892 , n16893 );
and ( n16895 , n16860 , n16894 );
buf ( n16896 , n4721 );
buf ( n16897 , n16896 );
xor ( n16898 , n16767 , n16770 );
and ( n16899 , n16897 , n16898 );
xor ( n16900 , n16744 , n16747 );
and ( n16901 , n16898 , n16900 );
and ( n16902 , n16897 , n16900 );
or ( n16903 , n16899 , n16901 , n16902 );
and ( n16904 , n10933 , n16424 );
and ( n16905 , n4367 , n11111 );
and ( n16906 , n11116 , n4362 );
and ( n16907 , n16905 , n16906 );
and ( n16908 , n16904 , n16907 );
buf ( n16909 , n4719 );
buf ( n16910 , n16909 );
and ( n16911 , n5177 , n16910 );
and ( n16912 , n4989 , n5086 );
and ( n16913 , n5091 , n4982 );
and ( n16914 , n16912 , n16913 );
and ( n16915 , n16911 , n16914 );
and ( n16916 , n16908 , n16915 );
xor ( n16917 , n16773 , n16774 );
xor ( n16918 , n16917 , n16776 );
and ( n16919 , n16915 , n16918 );
and ( n16920 , n16908 , n16918 );
or ( n16921 , n16916 , n16919 , n16920 );
and ( n16922 , n16903 , n16921 );
xor ( n16923 , n16757 , n16758 );
xor ( n16924 , n16923 , n16760 );
and ( n16925 , n16921 , n16924 );
and ( n16926 , n16903 , n16924 );
or ( n16927 , n16922 , n16925 , n16926 );
xor ( n16928 , n16741 , n16742 );
xor ( n16929 , n16928 , n16753 );
and ( n16930 , n16927 , n16929 );
xor ( n16931 , n16763 , n16782 );
xor ( n16932 , n16931 , n16785 );
and ( n16933 , n16929 , n16932 );
and ( n16934 , n16927 , n16932 );
or ( n16935 , n16930 , n16933 , n16934 );
and ( n16936 , n16894 , n16935 );
and ( n16937 , n16860 , n16935 );
or ( n16938 , n16895 , n16936 , n16937 );
xor ( n16939 , n16723 , n16738 );
xor ( n16940 , n16939 , n16794 );
and ( n16941 , n16938 , n16940 );
xor ( n16942 , n16725 , n16726 );
xor ( n16943 , n16942 , n16735 );
xor ( n16944 , n16756 , n16788 );
xor ( n16945 , n16944 , n16791 );
and ( n16946 , n16943 , n16945 );
xor ( n16947 , n16843 , n16845 );
and ( n16948 , n16945 , n16947 );
and ( n16949 , n16943 , n16947 );
or ( n16950 , n16946 , n16948 , n16949 );
and ( n16951 , n16940 , n16950 );
and ( n16952 , n16938 , n16950 );
or ( n16953 , n16941 , n16951 , n16952 );
xor ( n16954 , n16830 , n16849 );
xor ( n16955 , n16954 , n16852 );
and ( n16956 , n16953 , n16955 );
xor ( n16957 , n16832 , n16834 );
xor ( n16958 , n16957 , n16846 );
xor ( n16959 , n16836 , n16838 );
xor ( n16960 , n16959 , n16840 );
xor ( n16961 , n16764 , n16771 );
xor ( n16962 , n16961 , n16779 );
xor ( n16963 , n16863 , n16873 );
xor ( n16964 , n16963 , n16875 );
and ( n16965 , n16962 , n16964 );
xor ( n16966 , n16886 , n16887 );
xor ( n16967 , n16677 , n16678 );
xor ( n16968 , n16967 , n16680 );
and ( n16969 , n16966 , n16968 );
and ( n16970 , n16964 , n16969 );
and ( n16971 , n16962 , n16969 );
or ( n16972 , n16965 , n16970 , n16971 );
and ( n16973 , n16960 , n16972 );
xor ( n16974 , n16868 , n16872 );
and ( n16975 , n10933 , n16636 );
and ( n16976 , n4739 , n11111 );
and ( n16977 , n11116 , n4734 );
and ( n16978 , n16976 , n16977 );
and ( n16979 , n16975 , n16978 );
xor ( n16980 , n10525 , n10582 );
buf ( n16981 , n16980 );
buf ( n16982 , n16981 );
buf ( n16983 , n16982 );
and ( n16984 , n16979 , n16983 );
and ( n16985 , n16974 , n16984 );
xor ( n16986 , n16745 , n16746 );
xor ( n16987 , n16904 , n16907 );
and ( n16988 , n16986 , n16987 );
buf ( n16989 , n16988 );
and ( n16990 , n16984 , n16989 );
and ( n16991 , n16974 , n16989 );
or ( n16992 , n16985 , n16990 , n16991 );
xor ( n16993 , n16864 , n16867 );
xor ( n16994 , n16911 , n16914 );
and ( n16995 , n16993 , n16994 );
xor ( n16996 , n16884 , n16885 );
and ( n16997 , n16994 , n16996 );
and ( n16998 , n16993 , n16996 );
or ( n16999 , n16995 , n16997 , n16998 );
xor ( n17000 , n16897 , n16898 );
xor ( n17001 , n17000 , n16900 );
and ( n17002 , n16999 , n17001 );
xor ( n17003 , n16908 , n16915 );
xor ( n17004 , n17003 , n16918 );
and ( n17005 , n17001 , n17004 );
and ( n17006 , n16999 , n17004 );
or ( n17007 , n17002 , n17005 , n17006 );
and ( n17008 , n16992 , n17007 );
xor ( n17009 , n16881 , n16882 );
xor ( n17010 , n17009 , n16888 );
and ( n17011 , n17007 , n17010 );
and ( n17012 , n16992 , n17010 );
or ( n17013 , n17008 , n17011 , n17012 );
and ( n17014 , n16972 , n17013 );
and ( n17015 , n16960 , n17013 );
or ( n17016 , n16973 , n17014 , n17015 );
xor ( n17017 , n16860 , n16894 );
xor ( n17018 , n17017 , n16935 );
and ( n17019 , n17016 , n17018 );
xor ( n17020 , n16862 , n16878 );
xor ( n17021 , n17020 , n16891 );
xor ( n17022 , n16927 , n16929 );
xor ( n17023 , n17022 , n16932 );
and ( n17024 , n17021 , n17023 );
xor ( n17025 , n16903 , n16921 );
xor ( n17026 , n17025 , n16924 );
xor ( n17027 , n16966 , n16968 );
xor ( n17028 , n16979 , n16983 );
and ( n17029 , n10933 , n16910 );
and ( n17030 , n4989 , n11111 );
and ( n17031 , n11116 , n4982 );
and ( n17032 , n17030 , n17031 );
and ( n17033 , n17029 , n17032 );
xor ( n17034 , n10527 , n10581 );
buf ( n17035 , n17034 );
buf ( n17036 , n17035 );
buf ( n17037 , n17036 );
or ( n17038 , n17033 , n17037 );
and ( n17039 , n17028 , n17038 );
and ( n17040 , n10886 , n16910 );
and ( n17041 , n4989 , n10869 );
and ( n17042 , n10862 , n4982 );
and ( n17043 , n17041 , n17042 );
and ( n17044 , n17040 , n17043 );
and ( n17045 , n17038 , n17044 );
and ( n17046 , n17028 , n17044 );
or ( n17047 , n17039 , n17045 , n17046 );
and ( n17048 , n17027 , n17047 );
xor ( n17049 , n16905 , n16906 );
xor ( n17050 , n16865 , n16866 );
and ( n17051 , n17049 , n17050 );
xor ( n17052 , n16912 , n16913 );
and ( n17053 , n17050 , n17052 );
and ( n17054 , n17049 , n17052 );
or ( n17055 , n17051 , n17053 , n17054 );
buf ( n17056 , n5177 );
buf ( n17057 , n17056 );
xor ( n17058 , n16975 , n16978 );
and ( n17059 , n17057 , n17058 );
xor ( n17060 , n17040 , n17043 );
and ( n17061 , n17058 , n17060 );
and ( n17062 , n17057 , n17060 );
or ( n17063 , n17059 , n17061 , n17062 );
and ( n17064 , n17055 , n17063 );
buf ( n17065 , n5175 );
buf ( n17066 , n17065 );
and ( n17067 , n10886 , n17066 );
and ( n17068 , n5091 , n10869 );
and ( n17069 , n10862 , n5086 );
and ( n17070 , n17068 , n17069 );
and ( n17071 , n17067 , n17070 );
xor ( n17072 , n16976 , n16977 );
xor ( n17073 , n17041 , n17042 );
and ( n17074 , n17072 , n17073 );
buf ( n17075 , n17074 );
and ( n17076 , n17071 , n17075 );
xor ( n17077 , n17049 , n17050 );
xor ( n17078 , n17077 , n17052 );
and ( n17079 , n17075 , n17078 );
and ( n17080 , n17071 , n17078 );
or ( n17081 , n17076 , n17079 , n17080 );
and ( n17082 , n17063 , n17081 );
and ( n17083 , n17055 , n17081 );
or ( n17084 , n17064 , n17082 , n17083 );
and ( n17085 , n17047 , n17084 );
and ( n17086 , n17027 , n17084 );
or ( n17087 , n17048 , n17085 , n17086 );
and ( n17088 , n17026 , n17087 );
xor ( n17089 , n16962 , n16964 );
xor ( n17090 , n17089 , n16969 );
and ( n17091 , n17087 , n17090 );
and ( n17092 , n17026 , n17090 );
or ( n17093 , n17088 , n17091 , n17092 );
and ( n17094 , n17023 , n17093 );
and ( n17095 , n17021 , n17093 );
or ( n17096 , n17024 , n17094 , n17095 );
and ( n17097 , n17018 , n17096 );
and ( n17098 , n17016 , n17096 );
or ( n17099 , n17019 , n17097 , n17098 );
and ( n17100 , n16958 , n17099 );
xor ( n17101 , n16938 , n16940 );
xor ( n17102 , n17101 , n16950 );
and ( n17103 , n17099 , n17102 );
and ( n17104 , n16958 , n17102 );
or ( n17105 , n17100 , n17103 , n17104 );
and ( n17106 , n16955 , n17105 );
and ( n17107 , n16953 , n17105 );
or ( n17108 , n16956 , n17106 , n17107 );
and ( n17109 , n16857 , n17108 );
and ( n17110 , n16855 , n17108 );
or ( n17111 , n16858 , n17109 , n17110 );
and ( n17112 , n16828 , n17111 );
xor ( n17113 , n16828 , n17111 );
xor ( n17114 , n16855 , n16857 );
xor ( n17115 , n17114 , n17108 );
xor ( n17116 , n16953 , n16955 );
xor ( n17117 , n17116 , n17105 );
xor ( n17118 , n16943 , n16945 );
xor ( n17119 , n17118 , n16947 );
xor ( n17120 , n16960 , n16972 );
xor ( n17121 , n17120 , n17013 );
xor ( n17122 , n16992 , n17007 );
xor ( n17123 , n17122 , n17010 );
xor ( n17124 , n16974 , n16984 );
xor ( n17125 , n17124 , n16989 );
xor ( n17126 , n16999 , n17001 );
xor ( n17127 , n17126 , n17004 );
and ( n17128 , n17125 , n17127 );
buf ( n17129 , n16986 );
xor ( n17130 , n17129 , n16987 );
xor ( n17131 , n16993 , n16994 );
xor ( n17132 , n17131 , n16996 );
and ( n17133 , n17130 , n17132 );
xor ( n17134 , n17028 , n17038 );
xor ( n17135 , n17134 , n17044 );
and ( n17136 , n17132 , n17135 );
and ( n17137 , n17130 , n17135 );
or ( n17138 , n17133 , n17136 , n17137 );
and ( n17139 , n17127 , n17138 );
and ( n17140 , n17125 , n17138 );
or ( n17141 , n17128 , n17139 , n17140 );
and ( n17142 , n17123 , n17141 );
xor ( n17143 , n17026 , n17087 );
xor ( n17144 , n17143 , n17090 );
and ( n17145 , n17141 , n17144 );
and ( n17146 , n17123 , n17144 );
or ( n17147 , n17142 , n17145 , n17146 );
and ( n17148 , n17121 , n17147 );
xor ( n17149 , n17021 , n17023 );
xor ( n17150 , n17149 , n17093 );
and ( n17151 , n17147 , n17150 );
and ( n17152 , n17121 , n17150 );
or ( n17153 , n17148 , n17151 , n17152 );
and ( n17154 , n17119 , n17153 );
xor ( n17155 , n17016 , n17018 );
xor ( n17156 , n17155 , n17096 );
and ( n17157 , n17153 , n17156 );
and ( n17158 , n17119 , n17156 );
or ( n17159 , n17154 , n17157 , n17158 );
xor ( n17160 , n16958 , n17099 );
xor ( n17161 , n17160 , n17102 );
and ( n17162 , n17159 , n17161 );
xor ( n17163 , n17159 , n17161 );
xor ( n17164 , n17119 , n17153 );
xor ( n17165 , n17164 , n17156 );
xor ( n17166 , n17121 , n17147 );
xor ( n17167 , n17166 , n17150 );
xor ( n17168 , n17027 , n17047 );
xor ( n17169 , n17168 , n17084 );
xnor ( n17170 , n17033 , n17037 );
and ( n17171 , n10933 , n17066 );
and ( n17172 , n5091 , n11111 );
buf ( n17173 , n17172 );
and ( n17174 , n17171 , n17173 );
xor ( n17175 , n10546 , n10579 );
buf ( n17176 , n17175 );
buf ( n17177 , n17176 );
buf ( n17178 , n17177 );
or ( n17179 , n17174 , n17178 );
and ( n17180 , n17170 , n17179 );
xor ( n17181 , n17029 , n17032 );
xor ( n17182 , n17067 , n17070 );
and ( n17183 , n17181 , n17182 );
xor ( n17184 , n17030 , n17031 );
xor ( n17185 , n17068 , n17069 );
and ( n17186 , n17184 , n17185 );
buf ( n17187 , n10886 );
buf ( n17188 , n17187 );
and ( n17189 , n17185 , n17188 );
and ( n17190 , n17184 , n17188 );
or ( n17191 , n17186 , n17189 , n17190 );
and ( n17192 , n17182 , n17191 );
and ( n17193 , n17181 , n17191 );
or ( n17194 , n17183 , n17192 , n17193 );
and ( n17195 , n17179 , n17194 );
and ( n17196 , n17170 , n17194 );
or ( n17197 , n17180 , n17195 , n17196 );
xor ( n17198 , n17055 , n17063 );
xor ( n17199 , n17198 , n17081 );
and ( n17200 , n17197 , n17199 );
xor ( n17201 , n17057 , n17058 );
xor ( n17202 , n17201 , n17060 );
xor ( n17203 , n17071 , n17075 );
xor ( n17204 , n17203 , n17078 );
and ( n17205 , n17202 , n17204 );
xor ( n17206 , n17072 , n17073 );
buf ( n17207 , n17206 );
xnor ( n17208 , n17174 , n17178 );
and ( n17209 , n17207 , n17208 );
buf ( n17210 , n5380 );
buf ( n17211 , n17210 );
and ( n17212 , n10933 , n17211 );
and ( n17213 , n10862 , n11111 );
buf ( n17214 , n17213 );
and ( n17215 , n17212 , n17214 );
xor ( n17216 , n10567 , n10577 );
buf ( n17217 , n17216 );
buf ( n17218 , n17217 );
buf ( n17219 , n17218 );
and ( n17220 , n17215 , n17219 );
and ( n17221 , n17208 , n17220 );
and ( n17222 , n17207 , n17220 );
or ( n17223 , n17209 , n17221 , n17222 );
and ( n17224 , n17204 , n17223 );
and ( n17225 , n17202 , n17223 );
or ( n17226 , n17205 , n17224 , n17225 );
and ( n17227 , n17199 , n17226 );
and ( n17228 , n17197 , n17226 );
or ( n17229 , n17200 , n17227 , n17228 );
and ( n17230 , n17169 , n17229 );
xor ( n17231 , n17125 , n17127 );
xor ( n17232 , n17231 , n17138 );
and ( n17233 , n17229 , n17232 );
and ( n17234 , n17169 , n17232 );
or ( n17235 , n17230 , n17233 , n17234 );
xor ( n17236 , n17123 , n17141 );
xor ( n17237 , n17236 , n17144 );
and ( n17238 , n17235 , n17237 );
xor ( n17239 , n17235 , n17237 );
xor ( n17240 , n17130 , n17132 );
xor ( n17241 , n17240 , n17135 );
xor ( n17242 , n17170 , n17179 );
xor ( n17243 , n17242 , n17194 );
xor ( n17244 , n17171 , n17173 );
and ( n17245 , n11116 , n5086 );
xor ( n17246 , n10569 , n10576 );
buf ( n17247 , n17246 );
buf ( n17248 , n17247 );
buf ( n17249 , n17248 );
and ( n17250 , n17245 , n17249 );
not ( n17251 , n17172 );
and ( n17252 , n17249 , n17251 );
and ( n17253 , n17245 , n17251 );
or ( n17254 , n17250 , n17252 , n17253 );
and ( n17255 , n17244 , n17254 );
xor ( n17256 , n17184 , n17185 );
xor ( n17257 , n17256 , n17188 );
and ( n17258 , n17254 , n17257 );
and ( n17259 , n17244 , n17257 );
or ( n17260 , n17255 , n17258 , n17259 );
xor ( n17261 , n17181 , n17182 );
xor ( n17262 , n17261 , n17191 );
and ( n17263 , n17260 , n17262 );
xor ( n17264 , n17215 , n17219 );
xor ( n17265 , n17212 , n17214 );
and ( n17266 , n11116 , n10869 );
xor ( n17267 , n10570 , n10575 );
buf ( n17268 , n17267 );
buf ( n17269 , n17268 );
buf ( n17270 , n17269 );
and ( n17271 , n17266 , n17270 );
not ( n17272 , n17213 );
and ( n17273 , n17270 , n17272 );
and ( n17274 , n17266 , n17272 );
or ( n17275 , n17271 , n17273 , n17274 );
and ( n17276 , n17265 , n17275 );
buf ( n17277 , n17276 );
and ( n17278 , n17264 , n17277 );
xor ( n17279 , n17244 , n17254 );
xor ( n17280 , n17279 , n17257 );
and ( n17281 , n17277 , n17280 );
and ( n17282 , n17264 , n17280 );
or ( n17283 , n17278 , n17281 , n17282 );
and ( n17284 , n17262 , n17283 );
and ( n17285 , n17260 , n17283 );
or ( n17286 , n17263 , n17284 , n17285 );
and ( n17287 , n17243 , n17286 );
xor ( n17288 , n17202 , n17204 );
xor ( n17289 , n17288 , n17223 );
and ( n17290 , n17286 , n17289 );
and ( n17291 , n17243 , n17289 );
or ( n17292 , n17287 , n17290 , n17291 );
and ( n17293 , n17241 , n17292 );
xor ( n17294 , n17197 , n17199 );
xor ( n17295 , n17294 , n17226 );
and ( n17296 , n17292 , n17295 );
and ( n17297 , n17241 , n17295 );
or ( n17298 , n17293 , n17296 , n17297 );
xor ( n17299 , n17169 , n17229 );
xor ( n17300 , n17299 , n17232 );
and ( n17301 , n17298 , n17300 );
xor ( n17302 , n17298 , n17300 );
xor ( n17303 , n17241 , n17292 );
xor ( n17304 , n17303 , n17295 );
xor ( n17305 , n17243 , n17286 );
xor ( n17306 , n17305 , n17289 );
xor ( n17307 , n17207 , n17208 );
xor ( n17308 , n17307 , n17220 );
xor ( n17309 , n17260 , n17262 );
xor ( n17310 , n17309 , n17283 );
and ( n17311 , n17308 , n17310 );
xor ( n17312 , n17308 , n17310 );
xor ( n17313 , n17245 , n17249 );
xor ( n17314 , n17313 , n17251 );
xor ( n17315 , n10557 , n10574 );
buf ( n17316 , n17315 );
buf ( n17317 , n17316 );
buf ( n17318 , n17317 );
buf ( n17319 , n17318 );
buf ( n17320 , n10933 );
buf ( n17321 , n17320 );
and ( n17322 , n17319 , n17321 );
not ( n17323 , n17318 );
buf ( n17324 , n17323 );
and ( n17325 , n17321 , n17324 );
or ( n17326 , n17322 , n17325 , C0 );
and ( n17327 , n17314 , n17326 );
buf ( n17328 , n17265 );
xor ( n17329 , n17328 , n17275 );
and ( n17330 , n17326 , n17329 );
and ( n17331 , n17314 , n17329 );
or ( n17332 , n17327 , n17330 , n17331 );
xor ( n17333 , n17264 , n17277 );
xor ( n17334 , n17333 , n17280 );
and ( n17335 , n17332 , n17334 );
xor ( n17336 , n17332 , n17334 );
xor ( n17337 , n17314 , n17326 );
xor ( n17338 , n17337 , n17329 );
xor ( n17339 , n17266 , n17270 );
xor ( n17340 , n17339 , n17272 );
xor ( n17341 , n17319 , n17321 );
xor ( n17342 , n17341 , n17324 );
and ( n17343 , n17340 , n17342 );
buf ( n17344 , n17343 );
and ( n17345 , n17338 , n17344 );
and ( n17346 , n17336 , n17345 );
or ( n17347 , n17335 , n17346 );
and ( n17348 , n17312 , n17347 );
or ( n17349 , n17311 , n17348 );
and ( n17350 , n17306 , n17349 );
and ( n17351 , n17304 , n17350 );
and ( n17352 , n17302 , n17351 );
or ( n17353 , n17301 , n17352 );
and ( n17354 , n17239 , n17353 );
or ( n17355 , n17238 , n17354 );
and ( n17356 , n17167 , n17355 );
and ( n17357 , n17165 , n17356 );
and ( n17358 , n17163 , n17357 );
or ( n17359 , n17162 , n17358 );
and ( n17360 , n17117 , n17359 );
and ( n17361 , n17115 , n17360 );
and ( n17362 , n17113 , n17361 );
or ( n17363 , n17112 , n17362 );
and ( n17364 , n16826 , n17363 );
and ( n17365 , n16824 , n17364 );
and ( n17366 , n16822 , n17365 );
and ( n17367 , n16820 , n17366 );
or ( n17368 , n16819 , n17367 );
and ( n17369 , n16379 , n17368 );
or ( n17370 , n16378 , n17369 );
and ( n17371 , n16228 , n17370 );
and ( n17372 , n16226 , n17371 );
and ( n17373 , n16224 , n17372 );
and ( n17374 , n16222 , n17373 );
or ( n17375 , n16221 , n17374 );
and ( n17376 , n15700 , n17375 );
or ( n17377 , n15699 , n17376 );
and ( n17378 , n15320 , n17377 );
and ( n17379 , n15318 , n17378 );
and ( n17380 , n15316 , n17379 );
or ( n17381 , n15315 , n17380 );
and ( n17382 , n14696 , n17381 );
or ( n17383 , n14695 , n17382 );
and ( n17384 , n14613 , n17383 );
or ( n17385 , n14612 , n17384 );
and ( n17386 , n14105 , n17385 );
or ( n17387 , n14104 , n17386 );
and ( n17388 , n13878 , n17387 );
or ( n17389 , n13877 , n17388 );
and ( n17390 , n13584 , n17389 );
or ( n17391 , n13583 , n17390 );
and ( n17392 , n13322 , n17391 );
and ( n17393 , n13320 , n17392 );
or ( n17394 , n13319 , n17393 );
and ( n17395 , n13081 , n17394 );
or ( n17396 , n13080 , n17395 );
and ( n17397 , n12774 , n17396 );
or ( n17398 , n12773 , n17397 );
and ( n17399 , n12476 , n17398 );
or ( n17400 , n12475 , n17399 );
and ( n17401 , n11939 , n17400 );
and ( n17402 , n11937 , n17401 );
and ( n17403 , n11935 , n17402 );
or ( n17404 , n11934 , n17403 );
and ( n17405 , n11309 , n17404 );
and ( n17406 , n11307 , n17405 );
and ( n17407 , n11305 , n17406 );
or ( n17408 , n11304 , n17407 );
and ( n17409 , n10733 , n17408 );
or ( n17410 , n10732 , n17409 );
and ( n17411 , n4459 , n17410 );
or ( n17412 , n4458 , n17411 );
and ( n17413 , n4123 , n17412 );
or ( n17414 , n4122 , n17413 );
and ( n17415 , n4011 , n17414 );
and ( n17416 , n4009 , n17415 );
or ( n17417 , n4008 , n17416 );
and ( n17418 , n3491 , n17417 );
or ( n17419 , n3490 , n17418 );
and ( n17420 , n3211 , n17419 );
or ( n17421 , n3210 , n17420 );
and ( n17422 , n2885 , n17421 );
or ( n17423 , n2884 , n17422 );
and ( n17424 , n2832 , n17423 );
and ( n17425 , n2830 , n17424 );
or ( n17426 , n2829 , n17425 );
and ( n17427 , n2441 , n17426 );
or ( n17428 , n2440 , n17427 );
and ( n17429 , n2244 , n17428 );
or ( n17430 , n2243 , n17429 );
and ( n17431 , n2187 , n17430 );
and ( n17432 , n2185 , n17431 );
or ( n17433 , n2184 , n17432 );
and ( n17434 , n1890 , n17433 );
or ( n17435 , n1889 , n17434 );
and ( n17436 , n1758 , n17435 );
or ( n17437 , n1757 , n17436 );
and ( n17438 , n1553 , n17437 );
or ( n17439 , n1552 , n17438 );
and ( n17440 , n1506 , n17439 );
or ( n17441 , n1505 , n17440 );
and ( n17442 , n1461 , n17441 );
or ( n17443 , n1460 , n17442 );
xor ( n17444 , n1400 , n17443 );
buf ( n17445 , n17444 );
xor ( n17446 , n1461 , n17441 );
buf ( n17447 , n17446 );
xor ( n17448 , n1506 , n17439 );
buf ( n17449 , n17448 );
xor ( n17450 , n1553 , n17437 );
buf ( n17451 , n17450 );
xor ( n17452 , n1758 , n17435 );
buf ( n17453 , n17452 );
xor ( n17454 , n1890 , n17433 );
buf ( n17455 , n17454 );
xor ( n17456 , n2185 , n17431 );
buf ( n17457 , n17456 );
xor ( n17458 , n2187 , n17430 );
buf ( n17459 , n17458 );
xor ( n17460 , n2244 , n17428 );
buf ( n17461 , n17460 );
xor ( n17462 , n2441 , n17426 );
buf ( n17463 , n17462 );
xor ( n17464 , n2830 , n17424 );
buf ( n17465 , n17464 );
xor ( n17466 , n2832 , n17423 );
buf ( n17467 , n17466 );
xor ( n17468 , n2885 , n17421 );
buf ( n17469 , n17468 );
xor ( n17470 , n3211 , n17419 );
buf ( n17471 , n17470 );
xor ( n17472 , n3491 , n17417 );
buf ( n17473 , n17472 );
xor ( n17474 , n4009 , n17415 );
buf ( n17475 , n17474 );
xor ( n17476 , n4011 , n17414 );
buf ( n17477 , n17476 );
xor ( n17478 , n4123 , n17412 );
buf ( n17479 , n17478 );
xor ( n17480 , n4459 , n17410 );
buf ( n17481 , n17480 );
xor ( n17482 , n10733 , n17408 );
buf ( n17483 , n17482 );
xor ( n17484 , n11305 , n17406 );
buf ( n17485 , n17484 );
xor ( n17486 , n11307 , n17405 );
buf ( n17487 , n17486 );
xor ( n17488 , n11309 , n17404 );
buf ( n17489 , n17488 );
xor ( n17490 , n11935 , n17402 );
buf ( n17491 , n17490 );
xor ( n17492 , n11937 , n17401 );
buf ( n17493 , n17492 );
xor ( n17494 , n11939 , n17400 );
buf ( n17495 , n17494 );
xor ( n17496 , n12476 , n17398 );
buf ( n17497 , n17496 );
xor ( n17498 , n12774 , n17396 );
buf ( n17499 , n17498 );
xor ( n17500 , n13081 , n17394 );
buf ( n17501 , n17500 );
xor ( n17502 , n13320 , n17392 );
buf ( n17503 , n17502 );
xor ( n17504 , n13322 , n17391 );
buf ( n17505 , n17504 );
xor ( n17506 , n13584 , n17389 );
buf ( n17507 , n17506 );
xor ( n17508 , n13878 , n17387 );
buf ( n17509 , n17508 );
xor ( n17510 , n14105 , n17385 );
buf ( n17511 , n17510 );
xor ( n17512 , n14613 , n17383 );
buf ( n17513 , n17512 );
xor ( n17514 , n14696 , n17381 );
buf ( n17515 , n17514 );
xor ( n17516 , n15316 , n17379 );
buf ( n17517 , n17516 );
xor ( n17518 , n15318 , n17378 );
buf ( n17519 , n17518 );
xor ( n17520 , n15320 , n17377 );
buf ( n17521 , n17520 );
xor ( n17522 , n15700 , n17375 );
buf ( n17523 , n17522 );
xor ( n17524 , n16222 , n17373 );
buf ( n17525 , n17524 );
xor ( n17526 , n16224 , n17372 );
buf ( n17527 , n17526 );
xor ( n17528 , n16226 , n17371 );
buf ( n17529 , n17528 );
xor ( n17530 , n16228 , n17370 );
buf ( n17531 , n17530 );
xor ( n17532 , n16379 , n17368 );
buf ( n17533 , n17532 );
xor ( n17534 , n16820 , n17366 );
buf ( n17535 , n17534 );
xor ( n17536 , n16822 , n17365 );
buf ( n17537 , n17536 );
xor ( n17538 , n16824 , n17364 );
buf ( n17539 , n17538 );
xor ( n17540 , n16826 , n17363 );
buf ( n17541 , n17540 );
xor ( n17542 , n17113 , n17361 );
buf ( n17543 , n17542 );
xor ( n17544 , n17115 , n17360 );
buf ( n17545 , n17544 );
xor ( n17546 , n17117 , n17359 );
buf ( n17547 , n17546 );
xor ( n17548 , n17163 , n17357 );
buf ( n17549 , n17548 );
xor ( n17550 , n17165 , n17356 );
buf ( n17551 , n17550 );
xor ( n17552 , n17167 , n17355 );
buf ( n17553 , n17552 );
xor ( n17554 , n17239 , n17353 );
buf ( n17555 , n17554 );
xor ( n17556 , n17302 , n17351 );
buf ( n17557 , n17556 );
xor ( n17558 , n17304 , n17350 );
buf ( n17559 , n17558 );
xor ( n17560 , n17306 , n17349 );
buf ( n17561 , n17560 );
xor ( n17562 , n17312 , n17347 );
buf ( n17563 , n17562 );
xor ( n17564 , n17336 , n17345 );
buf ( n17565 , n17564 );
xor ( n17566 , n17338 , n17344 );
buf ( n17567 , n17566 );
xor ( n17568 , n17340 , n17342 );
buf ( n17569 , n17568 );
buf ( n17570 , n17569 );
buf ( n17571 , n17318 );
buf ( n17572 , n17571 );
not ( n17573 , n7702 );
and ( n17574 , n5408 , n5342 );
and ( n17575 , n17573 , n17574 );
and ( n17576 , n5393 , n7633 );
not ( n17577 , n17576 );
xnor ( n17578 , n17577 , n5561 );
xor ( n17579 , n17575 , n17578 );
and ( n17580 , n5377 , n5342 );
not ( n17581 , n17580 );
xor ( n17582 , n17579 , n17581 );
xor ( n17583 , n17573 , n17574 );
and ( n17584 , n5393 , n7696 );
not ( n17585 , n17584 );
xnor ( n17586 , n17585 , n7702 );
and ( n17587 , n5437 , n5342 );
or ( n17588 , n17586 , n17587 );
and ( n17589 , n17583 , n17588 );
and ( n17590 , n5377 , n7633 );
and ( n17591 , n5393 , n5512 );
nor ( n17592 , n17590 , n17591 );
xnor ( n17593 , n17592 , n5561 );
and ( n17594 , n17588 , n17593 );
and ( n17595 , n17583 , n17593 );
or ( n17596 , n17589 , n17594 , n17595 );
and ( n17597 , n17582 , n17596 );
and ( n17598 , n17575 , n17578 );
and ( n17599 , n17578 , n17581 );
and ( n17600 , n17575 , n17581 );
or ( n17601 , n17598 , n17599 , n17600 );
buf ( n17602 , n17580 );
not ( n17603 , n5561 );
xor ( n17604 , n17602 , n17603 );
and ( n17605 , n5393 , n5342 );
xor ( n17606 , n17604 , n17605 );
xor ( n17607 , n17601 , n17606 );
xor ( n17608 , n17597 , n17607 );
xor ( n17609 , n17583 , n17588 );
xor ( n17610 , n17609 , n17593 );
xnor ( n17611 , n17586 , n17587 );
not ( n17612 , n5373 );
and ( n17613 , n5377 , n7696 );
and ( n17614 , n5393 , n7694 );
nor ( n17615 , n17613 , n17614 );
xnor ( n17616 , n17615 , n7702 );
and ( n17617 , n17612 , n17616 );
and ( n17618 , n5437 , n7633 );
and ( n17619 , n5408 , n5512 );
nor ( n17620 , n17618 , n17619 );
xnor ( n17621 , n17620 , n5561 );
and ( n17622 , n17616 , n17621 );
and ( n17623 , n17612 , n17621 );
or ( n17624 , n17617 , n17622 , n17623 );
and ( n17625 , n17611 , n17624 );
and ( n17626 , n5408 , n7633 );
and ( n17627 , n5377 , n5512 );
nor ( n17628 , n17626 , n17627 );
xnor ( n17629 , n17628 , n5561 );
and ( n17630 , n17624 , n17629 );
and ( n17631 , n17611 , n17629 );
or ( n17632 , n17625 , n17630 , n17631 );
and ( n17633 , n17610 , n17632 );
xor ( n17634 , n17582 , n17596 );
and ( n17635 , n17633 , n17634 );
xor ( n17636 , n17611 , n17624 );
xor ( n17637 , n17636 , n17629 );
and ( n17638 , n5393 , n5365 );
not ( n17639 , n17638 );
xnor ( n17640 , n17639 , n5373 );
not ( n17641 , n17640 );
and ( n17642 , n5408 , n7696 );
and ( n17643 , n5377 , n7694 );
nor ( n17644 , n17642 , n17643 );
xnor ( n17645 , n17644 , n7702 );
and ( n17646 , n17641 , n17645 );
and ( n17647 , n5437 , n5512 );
not ( n17648 , n17647 );
xnor ( n17649 , n17648 , n5561 );
and ( n17650 , n17645 , n17649 );
and ( n17651 , n17641 , n17649 );
or ( n17652 , n17646 , n17650 , n17651 );
buf ( n17653 , n17640 );
and ( n17654 , n17652 , n17653 );
xor ( n17655 , n17612 , n17616 );
xor ( n17656 , n17655 , n17621 );
and ( n17657 , n17653 , n17656 );
and ( n17658 , n17652 , n17656 );
or ( n17659 , n17654 , n17657 , n17658 );
and ( n17660 , n17637 , n17659 );
xor ( n17661 , n17610 , n17632 );
and ( n17662 , n17660 , n17661 );
xor ( n17663 , n17637 , n17659 );
xor ( n17664 , n17652 , n17653 );
xor ( n17665 , n17664 , n17656 );
and ( n17666 , n5377 , n5365 );
and ( n17667 , n5393 , n5363 );
nor ( n17668 , n17666 , n17667 );
xnor ( n17669 , n17668 , n5373 );
and ( n17670 , n5437 , n7696 );
and ( n17671 , n5408 , n7694 );
nor ( n17672 , n17670 , n17671 );
xnor ( n17673 , n17672 , n7702 );
and ( n17674 , n17669 , n17673 );
and ( n17675 , n17673 , n5561 );
and ( n17676 , n17669 , n5561 );
or ( n17677 , n17674 , n17675 , n17676 );
and ( n17678 , n5393 , n5542 );
not ( n17679 , n17678 );
xnor ( n17680 , n17679 , n5550 );
and ( n17681 , n5408 , n5365 );
and ( n17682 , n5377 , n5363 );
nor ( n17683 , n17681 , n17682 );
xnor ( n17684 , n17683 , n5373 );
or ( n17685 , n17680 , n17684 );
not ( n17686 , n5550 );
and ( n17687 , n17685 , n17686 );
xor ( n17688 , n17669 , n17673 );
xor ( n17689 , n17688 , n5561 );
and ( n17690 , n17686 , n17689 );
and ( n17691 , n17685 , n17689 );
or ( n17692 , n17687 , n17690 , n17691 );
and ( n17693 , n17677 , n17692 );
xor ( n17694 , n17641 , n17645 );
xor ( n17695 , n17694 , n17649 );
and ( n17696 , n17692 , n17695 );
and ( n17697 , n17677 , n17695 );
or ( n17698 , n17693 , n17696 , n17697 );
and ( n17699 , n17665 , n17698 );
and ( n17700 , n17663 , n17699 );
xor ( n17701 , n17665 , n17698 );
xor ( n17702 , n17677 , n17692 );
xor ( n17703 , n17702 , n17695 );
and ( n17704 , n5377 , n5542 );
and ( n17705 , n5393 , n5540 );
nor ( n17706 , n17704 , n17705 );
xnor ( n17707 , n17706 , n5550 );
and ( n17708 , n17707 , n7702 );
and ( n17709 , n7702 , n5561 );
and ( n17710 , n17707 , n5561 );
or ( n17711 , n17708 , n17709 , n17710 );
and ( n17712 , n5437 , n7694 );
not ( n17713 , n17712 );
xnor ( n17714 , n17713 , n7702 );
and ( n17715 , n17711 , n17714 );
and ( n17716 , n17714 , n5561 );
and ( n17717 , n17711 , n5561 );
or ( n17718 , n17715 , n17716 , n17717 );
xnor ( n17719 , n17680 , n17684 );
not ( n17720 , n5290 );
and ( n17721 , n5437 , n5365 );
and ( n17722 , n5408 , n5363 );
nor ( n17723 , n17721 , n17722 );
xnor ( n17724 , n17723 , n5373 );
and ( n17725 , n17720 , n17724 );
and ( n17726 , n7711 , n5342 );
and ( n17727 , n17724 , n17726 );
and ( n17728 , n17720 , n17726 );
or ( n17729 , n17725 , n17727 , n17728 );
and ( n17730 , n17719 , n17729 );
and ( n17731 , n5408 , n5542 );
and ( n17732 , n5377 , n5540 );
nor ( n17733 , n17731 , n17732 );
xnor ( n17734 , n17733 , n5550 );
and ( n17735 , n5437 , n5363 );
not ( n17736 , n17735 );
xnor ( n17737 , n17736 , n5373 );
and ( n17738 , n17734 , n17737 );
and ( n17739 , n17737 , n7702 );
and ( n17740 , n17734 , n7702 );
or ( n17741 , n17738 , n17739 , n17740 );
and ( n17742 , n5393 , n5282 );
not ( n17743 , n17742 );
xnor ( n17744 , n17743 , n5290 );
buf ( n17745 , n17744 );
and ( n17746 , n17741 , n17745 );
xor ( n17747 , n17720 , n17724 );
xor ( n17748 , n17747 , n17726 );
and ( n17749 , n17745 , n17748 );
and ( n17750 , n17741 , n17748 );
or ( n17751 , n17746 , n17749 , n17750 );
and ( n17752 , n17729 , n17751 );
and ( n17753 , n17719 , n17751 );
or ( n17754 , n17730 , n17752 , n17753 );
and ( n17755 , n17718 , n17754 );
xor ( n17756 , n17685 , n17686 );
xor ( n17757 , n17756 , n17689 );
and ( n17758 , n17754 , n17757 );
and ( n17759 , n17718 , n17757 );
or ( n17760 , n17755 , n17758 , n17759 );
and ( n17761 , n17703 , n17760 );
and ( n17762 , n17701 , n17761 );
xor ( n17763 , n17718 , n17754 );
xor ( n17764 , n17763 , n17757 );
not ( n17765 , n17744 );
and ( n17766 , n7711 , n7633 );
not ( n17767 , n17766 );
xnor ( n17768 , n17767 , n5561 );
and ( n17769 , n17765 , n17768 );
and ( n17770 , n5309 , n5342 );
and ( n17771 , n17768 , n17770 );
and ( n17772 , n17765 , n17770 );
or ( n17773 , n17769 , n17771 , n17772 );
xor ( n17774 , n17707 , n7702 );
xor ( n17775 , n17774 , n5561 );
and ( n17776 , n17773 , n17775 );
xor ( n17777 , n17741 , n17745 );
xor ( n17778 , n17777 , n17748 );
and ( n17779 , n17775 , n17778 );
and ( n17780 , n17773 , n17778 );
or ( n17781 , n17776 , n17779 , n17780 );
xor ( n17782 , n17711 , n17714 );
xor ( n17783 , n17782 , n5561 );
and ( n17784 , n17781 , n17783 );
xor ( n17785 , n17719 , n17729 );
xor ( n17786 , n17785 , n17751 );
and ( n17787 , n17783 , n17786 );
and ( n17788 , n17781 , n17786 );
or ( n17789 , n17784 , n17787 , n17788 );
and ( n17790 , n17764 , n17789 );
xor ( n17791 , n17703 , n17760 );
and ( n17792 , n17790 , n17791 );
xor ( n17793 , n17764 , n17789 );
xor ( n17794 , n17781 , n17783 );
xor ( n17795 , n17794 , n17786 );
and ( n17796 , n5437 , n5542 );
and ( n17797 , n5408 , n5540 );
nor ( n17798 , n17796 , n17797 );
xnor ( n17799 , n17798 , n5550 );
and ( n17800 , n17799 , n7702 );
and ( n17801 , n5309 , n7633 );
and ( n17802 , n7711 , n5512 );
nor ( n17803 , n17801 , n17802 );
xnor ( n17804 , n17803 , n5561 );
and ( n17805 , n7702 , n17804 );
and ( n17806 , n17799 , n17804 );
or ( n17807 , n17800 , n17805 , n17806 );
not ( n17808 , n5270 );
and ( n17809 , n5373 , n17808 );
and ( n17810 , n5377 , n5282 );
and ( n17811 , n5393 , n5280 );
nor ( n17812 , n17810 , n17811 );
xnor ( n17813 , n17812 , n5290 );
and ( n17814 , n17808 , n17813 );
and ( n17815 , n5373 , n17813 );
or ( n17816 , n17809 , n17814 , n17815 );
and ( n17817 , n17807 , n17816 );
xor ( n17818 , n17734 , n17737 );
xor ( n17819 , n17818 , n7702 );
and ( n17820 , n17816 , n17819 );
and ( n17821 , n17807 , n17819 );
or ( n17822 , n17817 , n17820 , n17821 );
and ( n17823 , n5408 , n5282 );
and ( n17824 , n5377 , n5280 );
nor ( n17825 , n17823 , n17824 );
xnor ( n17826 , n17825 , n5290 );
and ( n17827 , n5437 , n5540 );
not ( n17828 , n17827 );
xnor ( n17829 , n17828 , n5550 );
and ( n17830 , n17826 , n17829 );
and ( n17831 , n7650 , n5342 );
and ( n17832 , n17829 , n17831 );
and ( n17833 , n17826 , n17831 );
or ( n17834 , n17830 , n17832 , n17833 );
buf ( n17835 , n5373 );
and ( n17836 , n17834 , n17835 );
and ( n17837 , n5296 , n5342 );
and ( n17838 , n17835 , n17837 );
and ( n17839 , n17834 , n17837 );
or ( n17840 , n17836 , n17838 , n17839 );
and ( n17841 , n5393 , n5262 );
not ( n17842 , n17841 );
xnor ( n17843 , n17842 , n5270 );
and ( n17844 , n7711 , n7696 );
not ( n17845 , n17844 );
xnor ( n17846 , n17845 , n7702 );
and ( n17847 , n17843 , n17846 );
and ( n17848 , n5296 , n7633 );
and ( n17849 , n5309 , n5512 );
nor ( n17850 , n17848 , n17849 );
xnor ( n17851 , n17850 , n5561 );
and ( n17852 , n17846 , n17851 );
and ( n17853 , n17843 , n17851 );
or ( n17854 , n17847 , n17852 , n17853 );
xor ( n17855 , n17799 , n7702 );
xor ( n17856 , n17855 , n17804 );
and ( n17857 , n17854 , n17856 );
xor ( n17858 , n5373 , n17808 );
xor ( n17859 , n17858 , n17813 );
and ( n17860 , n17856 , n17859 );
and ( n17861 , n17854 , n17859 );
or ( n17862 , n17857 , n17860 , n17861 );
and ( n17863 , n17840 , n17862 );
xor ( n17864 , n17765 , n17768 );
xor ( n17865 , n17864 , n17770 );
and ( n17866 , n17862 , n17865 );
and ( n17867 , n17840 , n17865 );
or ( n17868 , n17863 , n17866 , n17867 );
and ( n17869 , n17822 , n17868 );
xor ( n17870 , n17773 , n17775 );
xor ( n17871 , n17870 , n17778 );
and ( n17872 , n17868 , n17871 );
and ( n17873 , n17822 , n17871 );
or ( n17874 , n17869 , n17872 , n17873 );
and ( n17875 , n17795 , n17874 );
and ( n17876 , n17793 , n17875 );
xor ( n17877 , n17795 , n17874 );
xor ( n17878 , n17822 , n17868 );
xor ( n17879 , n17878 , n17871 );
and ( n17880 , n5437 , n5282 );
and ( n17881 , n5408 , n5280 );
nor ( n17882 , n17880 , n17881 );
xnor ( n17883 , n17882 , n5290 );
and ( n17884 , n17883 , n5373 );
and ( n17885 , n7647 , n5342 );
and ( n17886 , n5373 , n17885 );
and ( n17887 , n17883 , n17885 );
or ( n17888 , n17884 , n17886 , n17887 );
not ( n17889 , n5251 );
and ( n17890 , n5377 , n5262 );
and ( n17891 , n5393 , n5260 );
nor ( n17892 , n17890 , n17891 );
xnor ( n17893 , n17892 , n5270 );
and ( n17894 , n17889 , n17893 );
and ( n17895 , n5309 , n7696 );
and ( n17896 , n7711 , n7694 );
nor ( n17897 , n17895 , n17896 );
xnor ( n17898 , n17897 , n7702 );
and ( n17899 , n17893 , n17898 );
and ( n17900 , n17889 , n17898 );
or ( n17901 , n17894 , n17899 , n17900 );
and ( n17902 , n17888 , n17901 );
and ( n17903 , n17901 , n17612 );
and ( n17904 , n17888 , n17612 );
or ( n17905 , n17902 , n17903 , n17904 );
and ( n17906 , n5437 , n5280 );
not ( n17907 , n17906 );
xnor ( n17908 , n17907 , n5290 );
buf ( n17909 , n17908 );
and ( n17910 , n17909 , n5550 );
and ( n17911 , n7650 , n7633 );
and ( n17912 , n5296 , n5512 );
nor ( n17913 , n17911 , n17912 );
xnor ( n17914 , n17913 , n5561 );
and ( n17915 , n5550 , n17914 );
and ( n17916 , n17909 , n17914 );
or ( n17917 , n17910 , n17915 , n17916 );
xor ( n17918 , n17843 , n17846 );
xor ( n17919 , n17918 , n17851 );
and ( n17920 , n17917 , n17919 );
xor ( n17921 , n17826 , n17829 );
xor ( n17922 , n17921 , n17831 );
and ( n17923 , n17919 , n17922 );
and ( n17924 , n17917 , n17922 );
or ( n17925 , n17920 , n17923 , n17924 );
and ( n17926 , n17905 , n17925 );
xor ( n17927 , n17834 , n17835 );
xor ( n17928 , n17927 , n17837 );
and ( n17929 , n17925 , n17928 );
and ( n17930 , n17905 , n17928 );
or ( n17931 , n17926 , n17929 , n17930 );
xor ( n17932 , n17807 , n17816 );
xor ( n17933 , n17932 , n17819 );
and ( n17934 , n17931 , n17933 );
xor ( n17935 , n17840 , n17862 );
xor ( n17936 , n17935 , n17865 );
and ( n17937 , n17933 , n17936 );
and ( n17938 , n17931 , n17936 );
or ( n17939 , n17934 , n17937 , n17938 );
and ( n17940 , n17879 , n17939 );
and ( n17941 , n17877 , n17940 );
xor ( n17942 , n17854 , n17856 );
xor ( n17943 , n17942 , n17859 );
xor ( n17944 , n17888 , n17901 );
xor ( n17945 , n17944 , n17612 );
xor ( n17946 , n17883 , n5373 );
xor ( n17947 , n17946 , n17885 );
and ( n17948 , n5393 , n5243 );
not ( n17949 , n17948 );
xnor ( n17950 , n17949 , n5251 );
and ( n17951 , n17950 , n5550 );
and ( n17952 , n7711 , n5365 );
not ( n17953 , n17952 );
xnor ( n17954 , n17953 , n5373 );
and ( n17955 , n5550 , n17954 );
and ( n17956 , n17950 , n17954 );
or ( n17957 , n17951 , n17955 , n17956 );
and ( n17958 , n17947 , n17957 );
and ( n17959 , n17945 , n17958 );
and ( n17960 , n17943 , n17959 );
xor ( n17961 , n17931 , n17933 );
xor ( n17962 , n17961 , n17936 );
and ( n17963 , n17960 , n17962 );
xor ( n17964 , n17879 , n17939 );
and ( n17965 , n17963 , n17964 );
xor ( n17966 , n17943 , n17959 );
xor ( n17967 , n17905 , n17925 );
xor ( n17968 , n17967 , n17928 );
and ( n17969 , n17966 , n17968 );
and ( n17970 , n7647 , n7633 );
and ( n17971 , n7650 , n5512 );
nor ( n17972 , n17970 , n17971 );
xnor ( n17973 , n17972 , n5561 );
not ( n17974 , n17973 );
and ( n17975 , n7716 , n5342 );
and ( n17976 , n17974 , n17975 );
buf ( n17977 , n17973 );
and ( n17978 , n17976 , n17977 );
and ( n17979 , n5377 , n5243 );
and ( n17980 , n5393 , n5241 );
nor ( n17981 , n17979 , n17980 );
xnor ( n17982 , n17981 , n5251 );
and ( n17983 , n17982 , n5550 );
and ( n17984 , n7650 , n7696 );
and ( n17985 , n5296 , n7694 );
nor ( n17986 , n17984 , n17985 );
xnor ( n17987 , n17986 , n7702 );
and ( n17988 , n5550 , n17987 );
and ( n17989 , n17982 , n17987 );
or ( n17990 , n17983 , n17988 , n17989 );
and ( n17991 , n5437 , n5262 );
and ( n17992 , n5408 , n5260 );
nor ( n17993 , n17991 , n17992 );
xnor ( n17994 , n17993 , n5270 );
and ( n17995 , n7716 , n7633 );
and ( n17996 , n7647 , n5512 );
nor ( n17997 , n17995 , n17996 );
xnor ( n17998 , n17997 , n5561 );
and ( n17999 , n17994 , n17998 );
and ( n18000 , n5350 , n5342 );
and ( n18001 , n17998 , n18000 );
and ( n18002 , n17994 , n18000 );
or ( n18003 , n17999 , n18001 , n18002 );
and ( n18004 , n17990 , n18003 );
xor ( n18005 , n17950 , n5550 );
xor ( n18006 , n18005 , n17954 );
and ( n18007 , n18003 , n18006 );
and ( n18008 , n17990 , n18006 );
or ( n18009 , n18004 , n18007 , n18008 );
and ( n18010 , n17977 , n18009 );
and ( n18011 , n17976 , n18009 );
or ( n18012 , n17978 , n18010 , n18011 );
xor ( n18013 , n17945 , n17958 );
and ( n18014 , n18012 , n18013 );
xor ( n18015 , n17917 , n17919 );
xor ( n18016 , n18015 , n17922 );
and ( n18017 , n18013 , n18016 );
and ( n18018 , n18012 , n18016 );
or ( n18019 , n18014 , n18017 , n18018 );
and ( n18020 , n17968 , n18019 );
and ( n18021 , n17966 , n18019 );
or ( n18022 , n17969 , n18020 , n18021 );
not ( n18023 , n5333 );
and ( n18024 , n18023 , n5290 );
and ( n18025 , n5309 , n5365 );
and ( n18026 , n7711 , n5363 );
nor ( n18027 , n18025 , n18026 );
xnor ( n18028 , n18027 , n5373 );
and ( n18029 , n5290 , n18028 );
and ( n18030 , n18023 , n18028 );
or ( n18031 , n18024 , n18029 , n18030 );
and ( n18032 , n5408 , n5262 );
and ( n18033 , n5377 , n5260 );
nor ( n18034 , n18032 , n18033 );
xnor ( n18035 , n18034 , n5270 );
and ( n18036 , n18031 , n18035 );
not ( n18037 , n17908 );
and ( n18038 , n18035 , n18037 );
and ( n18039 , n18031 , n18037 );
or ( n18040 , n18036 , n18038 , n18039 );
xor ( n18041 , n17889 , n17893 );
xor ( n18042 , n18041 , n17898 );
and ( n18043 , n18040 , n18042 );
xor ( n18044 , n17909 , n5550 );
xor ( n18045 , n18044 , n17914 );
and ( n18046 , n18042 , n18045 );
and ( n18047 , n18040 , n18045 );
or ( n18048 , n18043 , n18046 , n18047 );
and ( n18049 , n5296 , n7696 );
and ( n18050 , n5309 , n7694 );
nor ( n18051 , n18049 , n18050 );
xnor ( n18052 , n18051 , n7702 );
xor ( n18053 , n17974 , n17975 );
and ( n18054 , n18052 , n18053 );
xor ( n18055 , n17947 , n17957 );
and ( n18056 , n18054 , n18055 );
and ( n18057 , n5408 , n5243 );
and ( n18058 , n5377 , n5241 );
nor ( n18059 , n18057 , n18058 );
xnor ( n18060 , n18059 , n5251 );
and ( n18061 , n5437 , n5260 );
not ( n18062 , n18061 );
xnor ( n18063 , n18062 , n5270 );
and ( n18064 , n18060 , n18063 );
and ( n18065 , n5350 , n7633 );
and ( n18066 , n7716 , n5512 );
nor ( n18067 , n18065 , n18066 );
xnor ( n18068 , n18067 , n5561 );
and ( n18069 , n18063 , n18068 );
and ( n18070 , n18060 , n18068 );
or ( n18071 , n18064 , n18069 , n18070 );
and ( n18072 , n5393 , n5325 );
not ( n18073 , n18072 );
xnor ( n18074 , n18073 , n5333 );
not ( n18075 , n18074 );
and ( n18076 , n7647 , n7696 );
and ( n18077 , n7650 , n7694 );
nor ( n18078 , n18076 , n18077 );
xnor ( n18079 , n18078 , n7702 );
and ( n18080 , n18075 , n18079 );
and ( n18081 , n5328 , n5342 );
and ( n18082 , n18079 , n18081 );
and ( n18083 , n18075 , n18081 );
or ( n18084 , n18080 , n18082 , n18083 );
and ( n18085 , n18071 , n18084 );
xor ( n18086 , n17994 , n17998 );
xor ( n18087 , n18086 , n18000 );
and ( n18088 , n18084 , n18087 );
and ( n18089 , n18071 , n18087 );
or ( n18090 , n18085 , n18088 , n18089 );
not ( n18091 , n18090 );
xor ( n18092 , n17990 , n18003 );
xor ( n18093 , n18092 , n18006 );
and ( n18094 , n18091 , n18093 );
and ( n18095 , n18055 , n18094 );
and ( n18096 , n18054 , n18094 );
or ( n18097 , n18056 , n18095 , n18096 );
and ( n18098 , n18048 , n18097 );
buf ( n18099 , n18090 );
xor ( n18100 , n18031 , n18035 );
xor ( n18101 , n18100 , n18037 );
and ( n18102 , n7711 , n5542 );
not ( n18103 , n18102 );
xnor ( n18104 , n18103 , n5550 );
and ( n18105 , n5290 , n18104 );
and ( n18106 , n5296 , n5365 );
and ( n18107 , n5309 , n5363 );
nor ( n18108 , n18106 , n18107 );
xnor ( n18109 , n18108 , n5373 );
and ( n18110 , n18104 , n18109 );
and ( n18111 , n5290 , n18109 );
or ( n18112 , n18105 , n18110 , n18111 );
buf ( n18113 , n18074 );
and ( n18114 , n18112 , n18113 );
xor ( n18115 , n18023 , n5290 );
xor ( n18116 , n18115 , n18028 );
and ( n18117 , n18113 , n18116 );
and ( n18118 , n18112 , n18116 );
or ( n18119 , n18114 , n18117 , n18118 );
and ( n18120 , n18101 , n18119 );
xor ( n18121 , n18052 , n18053 );
and ( n18122 , n18119 , n18121 );
and ( n18123 , n18101 , n18121 );
or ( n18124 , n18120 , n18122 , n18123 );
and ( n18125 , n18099 , n18124 );
xor ( n18126 , n17976 , n17977 );
xor ( n18127 , n18126 , n18009 );
and ( n18128 , n18124 , n18127 );
and ( n18129 , n18099 , n18127 );
or ( n18130 , n18125 , n18128 , n18129 );
and ( n18131 , n18097 , n18130 );
and ( n18132 , n18048 , n18130 );
or ( n18133 , n18098 , n18131 , n18132 );
xor ( n18134 , n18040 , n18042 );
xor ( n18135 , n18134 , n18045 );
xor ( n18136 , n18054 , n18055 );
xor ( n18137 , n18136 , n18094 );
and ( n18138 , n18135 , n18137 );
xor ( n18139 , n18099 , n18124 );
xor ( n18140 , n18139 , n18127 );
and ( n18141 , n18137 , n18140 );
and ( n18142 , n18135 , n18140 );
or ( n18143 , n18138 , n18141 , n18142 );
xor ( n18144 , n18012 , n18013 );
xor ( n18145 , n18144 , n18016 );
and ( n18146 , n18143 , n18145 );
xor ( n18147 , n18048 , n18097 );
xor ( n18148 , n18147 , n18130 );
and ( n18149 , n18145 , n18148 );
and ( n18150 , n18143 , n18148 );
or ( n18151 , n18146 , n18149 , n18150 );
and ( n18152 , n18133 , n18151 );
xor ( n18153 , n17966 , n17968 );
xor ( n18154 , n18153 , n18019 );
and ( n18155 , n18151 , n18154 );
and ( n18156 , n18133 , n18154 );
or ( n18157 , n18152 , n18155 , n18156 );
and ( n18158 , n18022 , n18157 );
xor ( n18159 , n17960 , n17962 );
and ( n18160 , n18157 , n18159 );
and ( n18161 , n18022 , n18159 );
or ( n18162 , n18158 , n18160 , n18161 );
and ( n18163 , n17964 , n18162 );
and ( n18164 , n17963 , n18162 );
or ( n18165 , n17965 , n18163 , n18164 );
and ( n18166 , n17940 , n18165 );
and ( n18167 , n17877 , n18165 );
or ( n18168 , n17941 , n18166 , n18167 );
and ( n18169 , n17875 , n18168 );
and ( n18170 , n17793 , n18168 );
or ( n18171 , n17876 , n18169 , n18170 );
and ( n18172 , n17791 , n18171 );
and ( n18173 , n17790 , n18171 );
or ( n18174 , n17792 , n18172 , n18173 );
and ( n18175 , n17761 , n18174 );
and ( n18176 , n17701 , n18174 );
or ( n18177 , n17762 , n18175 , n18176 );
and ( n18178 , n17699 , n18177 );
and ( n18179 , n17663 , n18177 );
or ( n18180 , n17700 , n18178 , n18179 );
and ( n18181 , n17661 , n18180 );
and ( n18182 , n17660 , n18180 );
or ( n18183 , n17662 , n18181 , n18182 );
and ( n18184 , n17634 , n18183 );
and ( n18185 , n17633 , n18183 );
or ( n18186 , n17635 , n18184 , n18185 );
xor ( n18187 , n17608 , n18186 );
xor ( n18188 , n17633 , n17634 );
xor ( n18189 , n18188 , n18183 );
xor ( n18190 , n17660 , n17661 );
xor ( n18191 , n18190 , n18180 );
xor ( n18192 , n17663 , n17699 );
xor ( n18193 , n18192 , n18177 );
xor ( n18194 , n17701 , n17761 );
xor ( n18195 , n18194 , n18174 );
xor ( n18196 , n17790 , n17791 );
xor ( n18197 , n18196 , n18171 );
xor ( n18198 , n17793 , n17875 );
xor ( n18199 , n18198 , n18168 );
xor ( n18200 , n17877 , n17940 );
xor ( n18201 , n18200 , n18165 );
xor ( n18202 , n17963 , n17964 );
xor ( n18203 , n18202 , n18162 );
xor ( n18204 , n18022 , n18157 );
xor ( n18205 , n18204 , n18159 );
xor ( n18206 , n18133 , n18151 );
xor ( n18207 , n18206 , n18154 );
xor ( n18208 , n18143 , n18145 );
xor ( n18209 , n18208 , n18148 );
xor ( n18210 , n18091 , n18093 );
xor ( n18211 , n18101 , n18119 );
xor ( n18212 , n18211 , n18121 );
and ( n18213 , n18210 , n18212 );
and ( n18214 , n5437 , n5243 );
and ( n18215 , n5408 , n5241 );
nor ( n18216 , n18214 , n18215 );
xnor ( n18217 , n18216 , n5251 );
and ( n18218 , n5309 , n5542 );
and ( n18219 , n7711 , n5540 );
nor ( n18220 , n18218 , n18219 );
xnor ( n18221 , n18220 , n5550 );
and ( n18222 , n18217 , n18221 );
and ( n18223 , n5317 , n5342 );
and ( n18224 , n18221 , n18223 );
and ( n18225 , n18217 , n18223 );
or ( n18226 , n18222 , n18224 , n18225 );
and ( n18227 , n5393 , n5499 );
not ( n18228 , n18227 );
xnor ( n18229 , n18228 , n5505 );
buf ( n18230 , n18229 );
not ( n18231 , n5505 );
and ( n18232 , n18230 , n18231 );
and ( n18233 , n5377 , n5325 );
and ( n18234 , n5393 , n5323 );
nor ( n18235 , n18233 , n18234 );
xnor ( n18236 , n18235 , n5333 );
and ( n18237 , n18231 , n18236 );
and ( n18238 , n18230 , n18236 );
or ( n18239 , n18232 , n18237 , n18238 );
and ( n18240 , n18226 , n18239 );
xor ( n18241 , n5290 , n18104 );
xor ( n18242 , n18241 , n18109 );
and ( n18243 , n18239 , n18242 );
and ( n18244 , n18226 , n18242 );
or ( n18245 , n18240 , n18243 , n18244 );
xor ( n18246 , n17982 , n5550 );
xor ( n18247 , n18246 , n17987 );
and ( n18248 , n18245 , n18247 );
xor ( n18249 , n18112 , n18113 );
xor ( n18250 , n18249 , n18116 );
and ( n18251 , n18247 , n18250 );
and ( n18252 , n18245 , n18250 );
or ( n18253 , n18248 , n18251 , n18252 );
and ( n18254 , n18212 , n18253 );
and ( n18255 , n18210 , n18253 );
or ( n18256 , n18213 , n18254 , n18255 );
xor ( n18257 , n18135 , n18137 );
xor ( n18258 , n18257 , n18140 );
and ( n18259 , n18256 , n18258 );
xor ( n18260 , n18210 , n18212 );
xor ( n18261 , n18260 , n18253 );
and ( n18262 , n7650 , n5365 );
and ( n18263 , n5296 , n5363 );
nor ( n18264 , n18262 , n18263 );
xnor ( n18265 , n18264 , n5373 );
and ( n18266 , n5290 , n18265 );
and ( n18267 , n5328 , n7633 );
and ( n18268 , n5350 , n5512 );
nor ( n18269 , n18267 , n18268 );
xnor ( n18270 , n18269 , n5561 );
and ( n18271 , n18265 , n18270 );
and ( n18272 , n5290 , n18270 );
or ( n18273 , n18266 , n18271 , n18272 );
xor ( n18274 , n18060 , n18063 );
xor ( n18275 , n18274 , n18068 );
and ( n18276 , n18273 , n18275 );
xor ( n18277 , n18075 , n18079 );
xor ( n18278 , n18277 , n18081 );
and ( n18279 , n18275 , n18278 );
and ( n18280 , n18273 , n18278 );
or ( n18281 , n18276 , n18279 , n18280 );
and ( n18282 , n7716 , n7696 );
and ( n18283 , n7647 , n7694 );
nor ( n18284 , n18282 , n18283 );
xnor ( n18285 , n18284 , n7702 );
and ( n18286 , n5270 , n18285 );
xor ( n18287 , n18230 , n18231 );
xor ( n18288 , n18287 , n18236 );
and ( n18289 , n18285 , n18288 );
and ( n18290 , n5270 , n18288 );
or ( n18291 , n18286 , n18289 , n18290 );
and ( n18292 , n5393 , n7722 );
not ( n18293 , n18292 );
xnor ( n18294 , n18293 , n7728 );
buf ( n18295 , n18294 );
not ( n18296 , n7728 );
and ( n18297 , n18295 , n18296 );
and ( n18298 , n5377 , n5499 );
and ( n18299 , n5393 , n5497 );
nor ( n18300 , n18298 , n18299 );
xnor ( n18301 , n18300 , n5505 );
and ( n18302 , n18296 , n18301 );
and ( n18303 , n18295 , n18301 );
or ( n18304 , n18297 , n18302 , n18303 );
and ( n18305 , n5437 , n5241 );
not ( n18306 , n18305 );
xnor ( n18307 , n18306 , n5251 );
and ( n18308 , n18304 , n18307 );
and ( n18309 , n7647 , n5365 );
and ( n18310 , n7650 , n5363 );
nor ( n18311 , n18309 , n18310 );
xnor ( n18312 , n18311 , n5373 );
and ( n18313 , n18307 , n18312 );
and ( n18314 , n18304 , n18312 );
or ( n18315 , n18308 , n18313 , n18314 );
not ( n18316 , n18229 );
and ( n18317 , n5408 , n5325 );
and ( n18318 , n5377 , n5323 );
nor ( n18319 , n18317 , n18318 );
xnor ( n18320 , n18319 , n5333 );
and ( n18321 , n18316 , n18320 );
and ( n18322 , n7711 , n5282 );
not ( n18323 , n18322 );
xnor ( n18324 , n18323 , n5290 );
and ( n18325 , n18320 , n18324 );
and ( n18326 , n18316 , n18324 );
or ( n18327 , n18321 , n18325 , n18326 );
and ( n18328 , n18315 , n18327 );
xor ( n18329 , n5290 , n18265 );
xor ( n18330 , n18329 , n18270 );
and ( n18331 , n18327 , n18330 );
and ( n18332 , n18315 , n18330 );
or ( n18333 , n18328 , n18331 , n18332 );
and ( n18334 , n18291 , n18333 );
xor ( n18335 , n18226 , n18239 );
xor ( n18336 , n18335 , n18242 );
and ( n18337 , n18333 , n18336 );
and ( n18338 , n18291 , n18336 );
or ( n18339 , n18334 , n18337 , n18338 );
and ( n18340 , n18281 , n18339 );
xor ( n18341 , n18071 , n18084 );
xor ( n18342 , n18341 , n18087 );
and ( n18343 , n18339 , n18342 );
and ( n18344 , n18281 , n18342 );
or ( n18345 , n18340 , n18343 , n18344 );
and ( n18346 , n18261 , n18345 );
and ( n18347 , n5296 , n5542 );
and ( n18348 , n5309 , n5540 );
nor ( n18349 , n18347 , n18348 );
xnor ( n18350 , n18349 , n5550 );
and ( n18351 , n5350 , n7696 );
and ( n18352 , n7716 , n7694 );
nor ( n18353 , n18351 , n18352 );
xnor ( n18354 , n18353 , n7702 );
and ( n18355 , n18350 , n18354 );
and ( n18356 , n5317 , n7633 );
and ( n18357 , n5328 , n5512 );
nor ( n18358 , n18356 , n18357 );
xnor ( n18359 , n18358 , n5561 );
and ( n18360 , n18354 , n18359 );
and ( n18361 , n18350 , n18359 );
or ( n18362 , n18355 , n18360 , n18361 );
and ( n18363 , n5437 , n5325 );
and ( n18364 , n5408 , n5323 );
nor ( n18365 , n18363 , n18364 );
xnor ( n18366 , n18365 , n5333 );
and ( n18367 , n5309 , n5282 );
and ( n18368 , n7711 , n5280 );
nor ( n18369 , n18367 , n18368 );
xnor ( n18370 , n18369 , n5290 );
and ( n18371 , n18366 , n18370 );
and ( n18372 , n7716 , n5365 );
and ( n18373 , n7647 , n5363 );
nor ( n18374 , n18372 , n18373 );
xnor ( n18375 , n18374 , n5373 );
and ( n18376 , n18370 , n18375 );
and ( n18377 , n18366 , n18375 );
or ( n18378 , n18371 , n18376 , n18377 );
and ( n18379 , n18378 , n5270 );
and ( n18380 , n5246 , n5342 );
and ( n18381 , n5270 , n18380 );
and ( n18382 , n18378 , n18380 );
or ( n18383 , n18379 , n18381 , n18382 );
and ( n18384 , n18362 , n18383 );
xor ( n18385 , n18217 , n18221 );
xor ( n18386 , n18385 , n18223 );
and ( n18387 , n18383 , n18386 );
and ( n18388 , n18362 , n18386 );
or ( n18389 , n18384 , n18387 , n18388 );
and ( n18390 , n5246 , n7633 );
and ( n18391 , n5317 , n5512 );
nor ( n18392 , n18390 , n18391 );
xnor ( n18393 , n18392 , n5561 );
and ( n18394 , n5251 , n18393 );
and ( n18395 , n5233 , n5342 );
and ( n18396 , n18393 , n18395 );
and ( n18397 , n5251 , n18395 );
or ( n18398 , n18394 , n18396 , n18397 );
xor ( n18399 , n18304 , n18307 );
xor ( n18400 , n18399 , n18312 );
and ( n18401 , n18398 , n18400 );
xor ( n18402 , n18316 , n18320 );
xor ( n18403 , n18402 , n18324 );
and ( n18404 , n18400 , n18403 );
and ( n18405 , n18398 , n18403 );
or ( n18406 , n18401 , n18404 , n18405 );
xor ( n18407 , n5270 , n18285 );
xor ( n18408 , n18407 , n18288 );
and ( n18409 , n18406 , n18408 );
xor ( n18410 , n18315 , n18327 );
xor ( n18411 , n18410 , n18330 );
and ( n18412 , n18408 , n18411 );
and ( n18413 , n18406 , n18411 );
or ( n18414 , n18409 , n18412 , n18413 );
and ( n18415 , n18389 , n18414 );
xor ( n18416 , n18273 , n18275 );
xor ( n18417 , n18416 , n18278 );
and ( n18418 , n18414 , n18417 );
and ( n18419 , n18389 , n18417 );
or ( n18420 , n18415 , n18418 , n18419 );
xor ( n18421 , n18245 , n18247 );
xor ( n18422 , n18421 , n18250 );
and ( n18423 , n18420 , n18422 );
xor ( n18424 , n18281 , n18339 );
xor ( n18425 , n18424 , n18342 );
and ( n18426 , n18422 , n18425 );
and ( n18427 , n18420 , n18425 );
or ( n18428 , n18423 , n18426 , n18427 );
and ( n18429 , n18345 , n18428 );
and ( n18430 , n18261 , n18428 );
or ( n18431 , n18346 , n18429 , n18430 );
and ( n18432 , n18258 , n18431 );
and ( n18433 , n18256 , n18431 );
or ( n18434 , n18259 , n18432 , n18433 );
and ( n18435 , n18209 , n18434 );
xor ( n18436 , n18256 , n18258 );
xor ( n18437 , n18436 , n18431 );
xor ( n18438 , n18420 , n18422 );
xor ( n18439 , n18438 , n18425 );
and ( n18440 , n5437 , n5323 );
not ( n18441 , n18440 );
xnor ( n18442 , n18441 , n5333 );
and ( n18443 , n5296 , n5282 );
and ( n18444 , n5309 , n5280 );
nor ( n18445 , n18443 , n18444 );
xnor ( n18446 , n18445 , n5290 );
and ( n18447 , n18442 , n18446 );
and ( n18448 , n5350 , n5365 );
and ( n18449 , n7716 , n5363 );
nor ( n18450 , n18448 , n18449 );
xnor ( n18451 , n18450 , n5373 );
and ( n18452 , n18446 , n18451 );
and ( n18453 , n18442 , n18451 );
or ( n18454 , n18447 , n18452 , n18453 );
and ( n18455 , n18454 , n5270 );
and ( n18456 , n5328 , n7696 );
and ( n18457 , n5350 , n7694 );
nor ( n18458 , n18456 , n18457 );
xnor ( n18459 , n18458 , n7702 );
and ( n18460 , n5270 , n18459 );
and ( n18461 , n18454 , n18459 );
or ( n18462 , n18455 , n18460 , n18461 );
and ( n18463 , n5393 , n5306 );
not ( n18464 , n18463 );
xnor ( n18465 , n18464 , n5314 );
buf ( n18466 , n18465 );
not ( n18467 , n5314 );
and ( n18468 , n18466 , n18467 );
and ( n18469 , n5377 , n7722 );
and ( n18470 , n5393 , n7720 );
nor ( n18471 , n18469 , n18470 );
xnor ( n18472 , n18471 , n7728 );
and ( n18473 , n18467 , n18472 );
and ( n18474 , n18466 , n18472 );
or ( n18475 , n18468 , n18473 , n18474 );
not ( n18476 , n18294 );
and ( n18477 , n18475 , n18476 );
and ( n18478 , n5408 , n5499 );
and ( n18479 , n5377 , n5497 );
nor ( n18480 , n18478 , n18479 );
xnor ( n18481 , n18480 , n5505 );
and ( n18482 , n18476 , n18481 );
and ( n18483 , n18475 , n18481 );
or ( n18484 , n18477 , n18482 , n18483 );
and ( n18485 , n7650 , n5542 );
and ( n18486 , n5296 , n5540 );
nor ( n18487 , n18485 , n18486 );
xnor ( n18488 , n18487 , n5550 );
and ( n18489 , n18484 , n18488 );
xor ( n18490 , n18295 , n18296 );
xor ( n18491 , n18490 , n18301 );
and ( n18492 , n18488 , n18491 );
and ( n18493 , n18484 , n18491 );
or ( n18494 , n18489 , n18492 , n18493 );
and ( n18495 , n18462 , n18494 );
xor ( n18496 , n18350 , n18354 );
xor ( n18497 , n18496 , n18359 );
and ( n18498 , n18494 , n18497 );
and ( n18499 , n18462 , n18497 );
or ( n18500 , n18495 , n18498 , n18499 );
xor ( n18501 , n18362 , n18383 );
xor ( n18502 , n18501 , n18386 );
and ( n18503 , n18500 , n18502 );
xor ( n18504 , n18406 , n18408 );
xor ( n18505 , n18504 , n18411 );
and ( n18506 , n18502 , n18505 );
and ( n18507 , n18500 , n18505 );
or ( n18508 , n18503 , n18506 , n18507 );
xor ( n18509 , n18291 , n18333 );
xor ( n18510 , n18509 , n18336 );
and ( n18511 , n18508 , n18510 );
xor ( n18512 , n18389 , n18414 );
xor ( n18513 , n18512 , n18417 );
and ( n18514 , n18510 , n18513 );
and ( n18515 , n18508 , n18513 );
or ( n18516 , n18511 , n18514 , n18515 );
and ( n18517 , n18439 , n18516 );
xor ( n18518 , n18261 , n18345 );
xor ( n18519 , n18518 , n18428 );
and ( n18520 , n18517 , n18519 );
xor ( n18521 , n18508 , n18510 );
xor ( n18522 , n18521 , n18513 );
and ( n18523 , n7711 , n5262 );
not ( n18524 , n18523 );
xnor ( n18525 , n18524 , n5270 );
and ( n18526 , n5251 , n18525 );
and ( n18527 , n5265 , n5342 );
and ( n18528 , n18525 , n18527 );
and ( n18529 , n5251 , n18527 );
or ( n18530 , n18526 , n18528 , n18529 );
and ( n18531 , n7647 , n5542 );
and ( n18532 , n7650 , n5540 );
nor ( n18533 , n18531 , n18532 );
xnor ( n18534 , n18533 , n5550 );
and ( n18535 , n5233 , n7633 );
and ( n18536 , n5246 , n5512 );
nor ( n18537 , n18535 , n18536 );
xnor ( n18538 , n18537 , n5561 );
and ( n18539 , n18534 , n18538 );
xor ( n18540 , n18475 , n18476 );
xor ( n18541 , n18540 , n18481 );
and ( n18542 , n18538 , n18541 );
and ( n18543 , n18534 , n18541 );
or ( n18544 , n18539 , n18542 , n18543 );
and ( n18545 , n18530 , n18544 );
xor ( n18546 , n18366 , n18370 );
xor ( n18547 , n18546 , n18375 );
and ( n18548 , n18544 , n18547 );
and ( n18549 , n18530 , n18547 );
or ( n18550 , n18545 , n18548 , n18549 );
xor ( n18551 , n18378 , n5270 );
xor ( n18552 , n18551 , n18380 );
and ( n18553 , n18550 , n18552 );
xor ( n18554 , n18398 , n18400 );
xor ( n18555 , n18554 , n18403 );
and ( n18556 , n18552 , n18555 );
and ( n18557 , n18550 , n18555 );
or ( n18558 , n18553 , n18556 , n18557 );
and ( n18559 , n7650 , n5282 );
and ( n18560 , n5296 , n5280 );
nor ( n18561 , n18559 , n18560 );
xnor ( n18562 , n18561 , n5290 );
and ( n18563 , n5333 , n18562 );
and ( n18564 , n5328 , n5365 );
and ( n18565 , n5350 , n5363 );
nor ( n18566 , n18564 , n18565 );
xnor ( n18567 , n18566 , n5373 );
and ( n18568 , n18562 , n18567 );
and ( n18569 , n5333 , n18567 );
or ( n18570 , n18563 , n18568 , n18569 );
and ( n18571 , n5393 , n5487 );
not ( n18572 , n18571 );
xnor ( n18573 , n18572 , n5478 );
buf ( n18574 , n18573 );
not ( n18575 , n5478 );
and ( n18576 , n18574 , n18575 );
and ( n18577 , n5377 , n5306 );
and ( n18578 , n5393 , n5304 );
nor ( n18579 , n18577 , n18578 );
xnor ( n18580 , n18579 , n5314 );
and ( n18581 , n18575 , n18580 );
and ( n18582 , n18574 , n18580 );
or ( n18583 , n18576 , n18581 , n18582 );
not ( n18584 , n18465 );
and ( n18585 , n18583 , n18584 );
and ( n18586 , n5408 , n7722 );
and ( n18587 , n5377 , n7720 );
nor ( n18588 , n18586 , n18587 );
xnor ( n18589 , n18588 , n7728 );
and ( n18590 , n18584 , n18589 );
and ( n18591 , n18583 , n18589 );
or ( n18592 , n18585 , n18590 , n18591 );
and ( n18593 , n5437 , n5499 );
and ( n18594 , n5408 , n5497 );
nor ( n18595 , n18593 , n18594 );
xnor ( n18596 , n18595 , n5505 );
and ( n18597 , n18592 , n18596 );
xor ( n18598 , n18466 , n18467 );
xor ( n18599 , n18598 , n18472 );
and ( n18600 , n18596 , n18599 );
and ( n18601 , n18592 , n18599 );
or ( n18602 , n18597 , n18600 , n18601 );
and ( n18603 , n18570 , n18602 );
and ( n18604 , n5317 , n7696 );
and ( n18605 , n5328 , n7694 );
nor ( n18606 , n18604 , n18605 );
xnor ( n18607 , n18606 , n7702 );
and ( n18608 , n18602 , n18607 );
and ( n18609 , n18570 , n18607 );
or ( n18610 , n18603 , n18608 , n18609 );
xor ( n18611 , n5251 , n18393 );
xor ( n18612 , n18611 , n18395 );
and ( n18613 , n18610 , n18612 );
xor ( n18614 , n18484 , n18488 );
xor ( n18615 , n18614 , n18491 );
and ( n18616 , n18612 , n18615 );
and ( n18617 , n18610 , n18615 );
or ( n18618 , n18613 , n18616 , n18617 );
xor ( n18619 , n18462 , n18494 );
xor ( n18620 , n18619 , n18497 );
and ( n18621 , n18618 , n18620 );
xor ( n18622 , n18550 , n18552 );
xor ( n18623 , n18622 , n18555 );
and ( n18624 , n18620 , n18623 );
and ( n18625 , n18618 , n18623 );
or ( n18626 , n18621 , n18624 , n18625 );
and ( n18627 , n18558 , n18626 );
xor ( n18628 , n18500 , n18502 );
xor ( n18629 , n18628 , n18505 );
and ( n18630 , n18626 , n18629 );
and ( n18631 , n18558 , n18629 );
or ( n18632 , n18627 , n18630 , n18631 );
and ( n18633 , n18522 , n18632 );
xor ( n18634 , n18439 , n18516 );
and ( n18635 , n18633 , n18634 );
xor ( n18636 , n18558 , n18626 );
xor ( n18637 , n18636 , n18629 );
and ( n18638 , n7716 , n5542 );
and ( n18639 , n7647 , n5540 );
nor ( n18640 , n18638 , n18639 );
xnor ( n18641 , n18640 , n5550 );
and ( n18642 , n5265 , n7633 );
and ( n18643 , n5233 , n5512 );
nor ( n18644 , n18642 , n18643 );
xnor ( n18645 , n18644 , n5561 );
and ( n18646 , n18641 , n18645 );
and ( n18647 , n5254 , n5342 );
and ( n18648 , n18645 , n18647 );
and ( n18649 , n18641 , n18647 );
or ( n18650 , n18646 , n18648 , n18649 );
and ( n18651 , n5309 , n5262 );
and ( n18652 , n7711 , n5260 );
nor ( n18653 , n18651 , n18652 );
xnor ( n18654 , n18653 , n5270 );
and ( n18655 , n5251 , n18654 );
and ( n18656 , n5246 , n7696 );
and ( n18657 , n5317 , n7694 );
nor ( n18658 , n18656 , n18657 );
xnor ( n18659 , n18658 , n7702 );
and ( n18660 , n18654 , n18659 );
and ( n18661 , n5251 , n18659 );
or ( n18662 , n18655 , n18660 , n18661 );
and ( n18663 , n18650 , n18662 );
xor ( n18664 , n18442 , n18446 );
xor ( n18665 , n18664 , n18451 );
and ( n18666 , n18662 , n18665 );
and ( n18667 , n18650 , n18665 );
or ( n18668 , n18663 , n18666 , n18667 );
xor ( n18669 , n18454 , n5270 );
xor ( n18670 , n18669 , n18459 );
and ( n18671 , n18668 , n18670 );
xor ( n18672 , n18530 , n18544 );
xor ( n18673 , n18672 , n18547 );
and ( n18674 , n18670 , n18673 );
and ( n18675 , n18668 , n18673 );
or ( n18676 , n18671 , n18674 , n18675 );
and ( n18677 , n7647 , n5282 );
and ( n18678 , n7650 , n5280 );
nor ( n18679 , n18677 , n18678 );
xnor ( n18680 , n18679 , n5290 );
and ( n18681 , n5333 , n18680 );
and ( n18682 , n5317 , n5365 );
and ( n18683 , n5328 , n5363 );
nor ( n18684 , n18682 , n18683 );
xnor ( n18685 , n18684 , n5373 );
and ( n18686 , n18680 , n18685 );
and ( n18687 , n5333 , n18685 );
or ( n18688 , n18681 , n18686 , n18687 );
and ( n18689 , n5437 , n7722 );
and ( n18690 , n5408 , n7720 );
nor ( n18691 , n18689 , n18690 );
xnor ( n18692 , n18691 , n7728 );
and ( n18693 , n18692 , n5505 );
xor ( n18694 , n18574 , n18575 );
xor ( n18695 , n18694 , n18580 );
and ( n18696 , n5505 , n18695 );
and ( n18697 , n18692 , n18695 );
or ( n18698 , n18693 , n18696 , n18697 );
and ( n18699 , n5437 , n5497 );
not ( n18700 , n18699 );
xnor ( n18701 , n18700 , n5505 );
and ( n18702 , n18698 , n18701 );
xor ( n18703 , n18583 , n18584 );
xor ( n18704 , n18703 , n18589 );
and ( n18705 , n18701 , n18704 );
and ( n18706 , n18698 , n18704 );
or ( n18707 , n18702 , n18705 , n18706 );
and ( n18708 , n18688 , n18707 );
xor ( n18709 , n18592 , n18596 );
xor ( n18710 , n18709 , n18599 );
and ( n18711 , n18707 , n18710 );
and ( n18712 , n18688 , n18710 );
or ( n18713 , n18708 , n18711 , n18712 );
xor ( n18714 , n5251 , n18525 );
xor ( n18715 , n18714 , n18527 );
and ( n18716 , n18713 , n18715 );
xor ( n18717 , n18534 , n18538 );
xor ( n18718 , n18717 , n18541 );
and ( n18719 , n18715 , n18718 );
and ( n18720 , n18713 , n18718 );
or ( n18721 , n18716 , n18719 , n18720 );
xor ( n18722 , n18668 , n18670 );
xor ( n18723 , n18722 , n18673 );
and ( n18724 , n18721 , n18723 );
xor ( n18725 , n18610 , n18612 );
xor ( n18726 , n18725 , n18615 );
and ( n18727 , n18723 , n18726 );
and ( n18728 , n18721 , n18726 );
or ( n18729 , n18724 , n18727 , n18728 );
and ( n18730 , n18676 , n18729 );
xor ( n18731 , n18618 , n18620 );
xor ( n18732 , n18731 , n18623 );
and ( n18733 , n18729 , n18732 );
and ( n18734 , n18676 , n18732 );
or ( n18735 , n18730 , n18733 , n18734 );
and ( n18736 , n18637 , n18735 );
xor ( n18737 , n18522 , n18632 );
and ( n18738 , n18736 , n18737 );
and ( n18739 , n5350 , n5542 );
and ( n18740 , n7716 , n5540 );
nor ( n18741 , n18739 , n18740 );
xnor ( n18742 , n18741 , n5550 );
and ( n18743 , n5233 , n7696 );
and ( n18744 , n5246 , n7694 );
nor ( n18745 , n18743 , n18744 );
xnor ( n18746 , n18745 , n7702 );
and ( n18747 , n18742 , n18746 );
and ( n18748 , n5285 , n5342 );
and ( n18749 , n18746 , n18748 );
and ( n18750 , n18742 , n18748 );
or ( n18751 , n18747 , n18749 , n18750 );
and ( n18752 , n7711 , n5243 );
not ( n18753 , n18752 );
xnor ( n18754 , n18753 , n5251 );
and ( n18755 , n5296 , n5262 );
and ( n18756 , n5309 , n5260 );
nor ( n18757 , n18755 , n18756 );
xnor ( n18758 , n18757 , n5270 );
and ( n18759 , n18754 , n18758 );
and ( n18760 , n5254 , n7633 );
and ( n18761 , n5265 , n5512 );
nor ( n18762 , n18760 , n18761 );
xnor ( n18763 , n18762 , n5561 );
and ( n18764 , n18758 , n18763 );
and ( n18765 , n18754 , n18763 );
or ( n18766 , n18759 , n18764 , n18765 );
and ( n18767 , n18751 , n18766 );
xor ( n18768 , n5333 , n18562 );
xor ( n18769 , n18768 , n18567 );
and ( n18770 , n18766 , n18769 );
and ( n18771 , n18751 , n18769 );
or ( n18772 , n18767 , n18770 , n18771 );
xor ( n18773 , n18570 , n18602 );
xor ( n18774 , n18773 , n18607 );
and ( n18775 , n18772 , n18774 );
xor ( n18776 , n18650 , n18662 );
xor ( n18777 , n18776 , n18665 );
and ( n18778 , n18774 , n18777 );
and ( n18779 , n18772 , n18777 );
or ( n18780 , n18775 , n18778 , n18779 );
and ( n18781 , n5393 , n7865 );
not ( n18782 , n18781 );
xnor ( n18783 , n18782 , n5429 );
buf ( n18784 , n18783 );
not ( n18785 , n5429 );
and ( n18786 , n18784 , n18785 );
and ( n18787 , n5377 , n5487 );
and ( n18788 , n5393 , n5485 );
nor ( n18789 , n18787 , n18788 );
xnor ( n18790 , n18789 , n5478 );
and ( n18791 , n18785 , n18790 );
and ( n18792 , n18784 , n18790 );
or ( n18793 , n18786 , n18791 , n18792 );
not ( n18794 , n18573 );
and ( n18795 , n18793 , n18794 );
and ( n18796 , n5408 , n5306 );
and ( n18797 , n5377 , n5304 );
nor ( n18798 , n18796 , n18797 );
xnor ( n18799 , n18798 , n5314 );
and ( n18800 , n18794 , n18799 );
and ( n18801 , n18793 , n18799 );
or ( n18802 , n18795 , n18800 , n18801 );
and ( n18803 , n7716 , n5282 );
and ( n18804 , n7647 , n5280 );
nor ( n18805 , n18803 , n18804 );
xnor ( n18806 , n18805 , n5290 );
and ( n18807 , n18802 , n18806 );
and ( n18808 , n5246 , n5365 );
and ( n18809 , n5317 , n5363 );
nor ( n18810 , n18808 , n18809 );
xnor ( n18811 , n18810 , n5373 );
and ( n18812 , n18806 , n18811 );
and ( n18813 , n18802 , n18811 );
or ( n18814 , n18807 , n18812 , n18813 );
and ( n18815 , n5437 , n7720 );
not ( n18816 , n18815 );
xnor ( n18817 , n18816 , n7728 );
and ( n18818 , n18817 , n5505 );
xor ( n18819 , n18793 , n18794 );
xor ( n18820 , n18819 , n18799 );
and ( n18821 , n5505 , n18820 );
and ( n18822 , n18817 , n18820 );
or ( n18823 , n18818 , n18821 , n18822 );
and ( n18824 , n18823 , n5333 );
xor ( n18825 , n18692 , n5505 );
xor ( n18826 , n18825 , n18695 );
and ( n18827 , n5333 , n18826 );
and ( n18828 , n18823 , n18826 );
or ( n18829 , n18824 , n18827 , n18828 );
and ( n18830 , n18814 , n18829 );
xor ( n18831 , n18698 , n18701 );
xor ( n18832 , n18831 , n18704 );
and ( n18833 , n18829 , n18832 );
and ( n18834 , n18814 , n18832 );
or ( n18835 , n18830 , n18833 , n18834 );
xor ( n18836 , n18641 , n18645 );
xor ( n18837 , n18836 , n18647 );
and ( n18838 , n18835 , n18837 );
xor ( n18839 , n5251 , n18654 );
xor ( n18840 , n18839 , n18659 );
and ( n18841 , n18837 , n18840 );
and ( n18842 , n18835 , n18840 );
or ( n18843 , n18838 , n18841 , n18842 );
xor ( n18844 , n18772 , n18774 );
xor ( n18845 , n18844 , n18777 );
and ( n18846 , n18843 , n18845 );
xor ( n18847 , n18713 , n18715 );
xor ( n18848 , n18847 , n18718 );
and ( n18849 , n18845 , n18848 );
and ( n18850 , n18843 , n18848 );
or ( n18851 , n18846 , n18849 , n18850 );
and ( n18852 , n18780 , n18851 );
xor ( n18853 , n18721 , n18723 );
xor ( n18854 , n18853 , n18726 );
and ( n18855 , n18851 , n18854 );
and ( n18856 , n18780 , n18854 );
or ( n18857 , n18852 , n18855 , n18856 );
xor ( n18858 , n18742 , n18746 );
xor ( n18859 , n18858 , n18748 );
xor ( n18860 , n18754 , n18758 );
xor ( n18861 , n18860 , n18763 );
or ( n18862 , n18859 , n18861 );
xnor ( n18863 , n18859 , n18861 );
and ( n18864 , n5317 , n5542 );
and ( n18865 , n5328 , n5540 );
nor ( n18866 , n18864 , n18865 );
xnor ( n18867 , n18866 , n5550 );
and ( n18868 , n5254 , n7696 );
and ( n18869 , n5265 , n7694 );
nor ( n18870 , n18868 , n18869 );
xnor ( n18871 , n18870 , n7702 );
and ( n18872 , n18867 , n18871 );
and ( n18873 , n5274 , n7633 );
and ( n18874 , n5285 , n5512 );
nor ( n18875 , n18873 , n18874 );
xnor ( n18876 , n18875 , n5561 );
and ( n18877 , n18871 , n18876 );
and ( n18878 , n18867 , n18876 );
or ( n18879 , n18872 , n18877 , n18878 );
xor ( n18880 , n18802 , n18806 );
xor ( n18881 , n18880 , n18811 );
and ( n18882 , n18879 , n18881 );
and ( n18883 , n18863 , n18882 );
and ( n18884 , n18862 , n18883 );
and ( n18885 , n5309 , n5243 );
and ( n18886 , n7711 , n5241 );
nor ( n18887 , n18885 , n18886 );
xnor ( n18888 , n18887 , n5251 );
and ( n18889 , n7650 , n5262 );
and ( n18890 , n5296 , n5260 );
nor ( n18891 , n18889 , n18890 );
xnor ( n18892 , n18891 , n5270 );
and ( n18893 , n18888 , n18892 );
and ( n18894 , n5274 , n5342 );
and ( n18895 , n18892 , n18894 );
and ( n18896 , n18888 , n18894 );
or ( n18897 , n18893 , n18895 , n18896 );
and ( n18898 , n5328 , n5542 );
and ( n18899 , n5350 , n5540 );
nor ( n18900 , n18898 , n18899 );
xnor ( n18901 , n18900 , n5550 );
and ( n18902 , n5265 , n7696 );
and ( n18903 , n5233 , n7694 );
nor ( n18904 , n18902 , n18903 );
xnor ( n18905 , n18904 , n7702 );
and ( n18906 , n18901 , n18905 );
and ( n18907 , n5285 , n7633 );
and ( n18908 , n5254 , n5512 );
nor ( n18909 , n18907 , n18908 );
xnor ( n18910 , n18909 , n5561 );
and ( n18911 , n18905 , n18910 );
and ( n18912 , n18901 , n18910 );
or ( n18913 , n18906 , n18911 , n18912 );
and ( n18914 , n18897 , n18913 );
xor ( n18915 , n5333 , n18680 );
xor ( n18916 , n18915 , n18685 );
and ( n18917 , n18913 , n18916 );
and ( n18918 , n18897 , n18916 );
or ( n18919 , n18914 , n18917 , n18918 );
xor ( n18920 , n18751 , n18766 );
xor ( n18921 , n18920 , n18769 );
and ( n18922 , n18919 , n18921 );
xor ( n18923 , n18688 , n18707 );
xor ( n18924 , n18923 , n18710 );
and ( n18925 , n18921 , n18924 );
and ( n18926 , n18919 , n18924 );
or ( n18927 , n18922 , n18925 , n18926 );
and ( n18928 , n18884 , n18927 );
and ( n18929 , n7650 , n5243 );
and ( n18930 , n5296 , n5241 );
nor ( n18931 , n18929 , n18930 );
xnor ( n18932 , n18931 , n5251 );
and ( n18933 , n5529 , n7633 );
and ( n18934 , n5274 , n5512 );
nor ( n18935 , n18933 , n18934 );
xnor ( n18936 , n18935 , n5561 );
and ( n18937 , n18932 , n18936 );
not ( n18938 , n5405 );
and ( n18939 , n5377 , n7865 );
and ( n18940 , n5393 , n7863 );
nor ( n18941 , n18939 , n18940 );
xnor ( n18942 , n18941 , n5429 );
and ( n18943 , n18938 , n18942 );
and ( n18944 , n5437 , n5487 );
and ( n18945 , n5408 , n5485 );
nor ( n18946 , n18944 , n18945 );
xnor ( n18947 , n18946 , n5478 );
and ( n18948 , n18942 , n18947 );
and ( n18949 , n18938 , n18947 );
or ( n18950 , n18943 , n18948 , n18949 );
not ( n18951 , n18783 );
and ( n18952 , n18950 , n18951 );
and ( n18953 , n5408 , n5487 );
and ( n18954 , n5377 , n5485 );
nor ( n18955 , n18953 , n18954 );
xnor ( n18956 , n18955 , n5478 );
and ( n18957 , n18951 , n18956 );
and ( n18958 , n18950 , n18956 );
or ( n18959 , n18952 , n18957 , n18958 );
and ( n18960 , n5437 , n5304 );
not ( n18961 , n18960 );
xnor ( n18962 , n18961 , n5314 );
and ( n18963 , n18962 , n7728 );
xor ( n18964 , n18950 , n18951 );
xor ( n18965 , n18964 , n18956 );
and ( n18966 , n7728 , n18965 );
and ( n18967 , n18962 , n18965 );
or ( n18968 , n18963 , n18966 , n18967 );
xor ( n18969 , n18959 , n18968 );
xor ( n18970 , n18969 , n5505 );
and ( n18971 , n18936 , n18970 );
and ( n18972 , n18932 , n18970 );
or ( n18973 , n18937 , n18971 , n18972 );
and ( n18974 , n5309 , n5325 );
and ( n18975 , n7711 , n5323 );
nor ( n18976 , n18974 , n18975 );
xnor ( n18977 , n18976 , n5333 );
and ( n18978 , n5328 , n5282 );
and ( n18979 , n5350 , n5280 );
nor ( n18980 , n18978 , n18979 );
xnor ( n18981 , n18980 , n5290 );
and ( n18982 , n18977 , n18981 );
and ( n18983 , n5437 , n5306 );
and ( n18984 , n5408 , n5304 );
nor ( n18985 , n18983 , n18984 );
xnor ( n18986 , n18985 , n5314 );
xor ( n18987 , n18986 , n7728 );
xor ( n18988 , n18784 , n18785 );
xor ( n18989 , n18988 , n18790 );
xor ( n18990 , n18987 , n18989 );
and ( n18991 , n18981 , n18990 );
and ( n18992 , n18977 , n18990 );
or ( n18993 , n18982 , n18991 , n18992 );
and ( n18994 , n18973 , n18993 );
and ( n18995 , n18986 , n7728 );
and ( n18996 , n7728 , n18989 );
and ( n18997 , n18986 , n18989 );
or ( n18998 , n18995 , n18996 , n18997 );
and ( n18999 , n5350 , n5282 );
and ( n19000 , n7716 , n5280 );
nor ( n19001 , n18999 , n19000 );
xnor ( n19002 , n19001 , n5290 );
xor ( n19003 , n18998 , n19002 );
and ( n19004 , n5233 , n5365 );
and ( n19005 , n5246 , n5363 );
nor ( n19006 , n19004 , n19005 );
xnor ( n19007 , n19006 , n5373 );
xor ( n19008 , n19003 , n19007 );
and ( n19009 , n18993 , n19008 );
and ( n19010 , n18973 , n19008 );
or ( n19011 , n18994 , n19009 , n19010 );
xor ( n19012 , n18888 , n18892 );
xor ( n19013 , n19012 , n18894 );
and ( n19014 , n19011 , n19013 );
xor ( n19015 , n18901 , n18905 );
xor ( n19016 , n19015 , n18910 );
and ( n19017 , n19013 , n19016 );
and ( n19018 , n19011 , n19016 );
or ( n19019 , n19014 , n19017 , n19018 );
and ( n19020 , n18959 , n18968 );
and ( n19021 , n18968 , n5505 );
and ( n19022 , n18959 , n5505 );
or ( n19023 , n19020 , n19021 , n19022 );
and ( n19024 , n5296 , n5243 );
and ( n19025 , n5309 , n5241 );
nor ( n19026 , n19024 , n19025 );
xnor ( n19027 , n19026 , n5251 );
and ( n19028 , n19023 , n19027 );
and ( n19029 , n7647 , n5262 );
and ( n19030 , n7650 , n5260 );
nor ( n19031 , n19029 , n19030 );
xnor ( n19032 , n19031 , n5270 );
and ( n19033 , n19027 , n19032 );
and ( n19034 , n19023 , n19032 );
or ( n19035 , n19028 , n19033 , n19034 );
xor ( n19036 , n18867 , n18871 );
xor ( n19037 , n19036 , n18876 );
xor ( n19038 , n19023 , n19027 );
xor ( n19039 , n19038 , n19032 );
and ( n19040 , n19037 , n19039 );
and ( n19041 , n19035 , n19040 );
xor ( n19042 , n18879 , n18881 );
and ( n19043 , n19040 , n19042 );
and ( n19044 , n19035 , n19042 );
or ( n19045 , n19041 , n19043 , n19044 );
and ( n19046 , n19019 , n19045 );
xor ( n19047 , n18863 , n18882 );
and ( n19048 , n19045 , n19047 );
and ( n19049 , n19019 , n19047 );
or ( n19050 , n19046 , n19048 , n19049 );
xor ( n19051 , n18862 , n18883 );
and ( n19052 , n19050 , n19051 );
xor ( n19053 , n18835 , n18837 );
xor ( n19054 , n19053 , n18840 );
and ( n19055 , n19051 , n19054 );
and ( n19056 , n19050 , n19054 );
or ( n19057 , n19052 , n19055 , n19056 );
xor ( n19058 , n18843 , n18845 );
xor ( n19059 , n19058 , n18848 );
and ( n19060 , n19057 , n19059 );
and ( n19061 , n18998 , n19002 );
and ( n19062 , n19002 , n19007 );
and ( n19063 , n18998 , n19007 );
or ( n19064 , n19061 , n19062 , n19063 );
and ( n19065 , n7711 , n5325 );
not ( n19066 , n19065 );
xnor ( n19067 , n19066 , n5333 );
and ( n19068 , n5529 , n5342 );
and ( n19069 , n19067 , n19068 );
xor ( n19070 , n18817 , n5505 );
xor ( n19071 , n19070 , n18820 );
and ( n19072 , n19068 , n19071 );
and ( n19073 , n19067 , n19071 );
or ( n19074 , n19069 , n19072 , n19073 );
and ( n19075 , n19064 , n19074 );
xor ( n19076 , n18823 , n5333 );
xor ( n19077 , n19076 , n18826 );
and ( n19078 , n19074 , n19077 );
and ( n19079 , n19064 , n19077 );
or ( n19080 , n19075 , n19078 , n19079 );
xor ( n19081 , n18897 , n18913 );
xor ( n19082 , n19081 , n18916 );
and ( n19083 , n19080 , n19082 );
xor ( n19084 , n18814 , n18829 );
xor ( n19085 , n19084 , n18832 );
and ( n19086 , n19082 , n19085 );
and ( n19087 , n19080 , n19085 );
or ( n19088 , n19083 , n19086 , n19087 );
xor ( n19089 , n18919 , n18921 );
xor ( n19090 , n19089 , n18924 );
and ( n19091 , n19088 , n19090 );
xor ( n19092 , n19011 , n19013 );
xor ( n19093 , n19092 , n19016 );
and ( n19094 , n7716 , n5262 );
and ( n19095 , n7647 , n5260 );
nor ( n19096 , n19094 , n19095 );
xnor ( n19097 , n19096 , n5270 );
and ( n19098 , n5265 , n5365 );
and ( n19099 , n5233 , n5363 );
nor ( n19100 , n19098 , n19099 );
xnor ( n19101 , n19100 , n5373 );
and ( n19102 , n19097 , n19101 );
and ( n19103 , n5368 , n5342 );
and ( n19104 , n19101 , n19103 );
and ( n19105 , n19097 , n19103 );
or ( n19106 , n19102 , n19104 , n19105 );
and ( n19107 , n5408 , n7865 );
and ( n19108 , n5377 , n7863 );
nor ( n19109 , n19107 , n19108 );
xnor ( n19110 , n19109 , n5429 );
buf ( n19111 , n19110 );
and ( n19112 , n19111 , n5314 );
xor ( n19113 , n18938 , n18942 );
xor ( n19114 , n19113 , n18947 );
and ( n19115 , n5314 , n19114 );
and ( n19116 , n19111 , n19114 );
or ( n19117 , n19112 , n19115 , n19116 );
and ( n19118 , n7711 , n5499 );
not ( n19119 , n19118 );
xnor ( n19120 , n19119 , n5505 );
and ( n19121 , n19117 , n19120 );
xor ( n19122 , n18962 , n7728 );
xor ( n19123 , n19122 , n18965 );
and ( n19124 , n19120 , n19123 );
and ( n19125 , n19117 , n19123 );
or ( n19126 , n19121 , n19124 , n19125 );
and ( n19127 , n5246 , n5542 );
and ( n19128 , n5317 , n5540 );
nor ( n19129 , n19127 , n19128 );
xnor ( n19130 , n19129 , n5550 );
and ( n19131 , n19126 , n19130 );
and ( n19132 , n5285 , n7696 );
and ( n19133 , n5254 , n7694 );
nor ( n19134 , n19132 , n19133 );
xnor ( n19135 , n19134 , n7702 );
and ( n19136 , n19130 , n19135 );
and ( n19137 , n19126 , n19135 );
or ( n19138 , n19131 , n19136 , n19137 );
and ( n19139 , n19106 , n19138 );
xor ( n19140 , n19067 , n19068 );
xor ( n19141 , n19140 , n19071 );
and ( n19142 , n19138 , n19141 );
and ( n19143 , n19106 , n19141 );
or ( n19144 , n19139 , n19142 , n19143 );
and ( n19145 , n19093 , n19144 );
and ( n19146 , n5328 , n5262 );
and ( n19147 , n5350 , n5260 );
nor ( n19148 , n19146 , n19147 );
xnor ( n19149 , n19148 , n5270 );
and ( n19150 , n5265 , n5542 );
and ( n19151 , n5233 , n5540 );
nor ( n19152 , n19150 , n19151 );
xnor ( n19153 , n19152 , n5550 );
and ( n19154 , n19149 , n19153 );
and ( n19155 , n5355 , n7633 );
and ( n19156 , n5368 , n5512 );
nor ( n19157 , n19155 , n19156 );
xnor ( n19158 , n19157 , n5561 );
and ( n19159 , n19153 , n19158 );
and ( n19160 , n19149 , n19158 );
or ( n19161 , n19154 , n19159 , n19160 );
and ( n19162 , n5309 , n5499 );
and ( n19163 , n7711 , n5497 );
nor ( n19164 , n19162 , n19163 );
xnor ( n19165 , n19164 , n5505 );
and ( n19166 , n5246 , n5282 );
and ( n19167 , n5317 , n5280 );
nor ( n19168 , n19166 , n19167 );
xnor ( n19169 , n19168 , n5290 );
and ( n19170 , n19165 , n19169 );
and ( n19171 , n5393 , n5468 );
not ( n19172 , n19171 );
xnor ( n19173 , n19172 , n5405 );
not ( n19174 , n19110 );
and ( n19175 , n19173 , n19174 );
and ( n19176 , n5437 , n5485 );
not ( n19177 , n19176 );
xnor ( n19178 , n19177 , n5478 );
and ( n19179 , n19174 , n19178 );
and ( n19180 , n19173 , n19178 );
or ( n19181 , n19175 , n19179 , n19180 );
not ( n19182 , n5420 );
and ( n19183 , n5437 , n7865 );
and ( n19184 , n5408 , n7863 );
nor ( n19185 , n19183 , n19184 );
xnor ( n19186 , n19185 , n5429 );
and ( n19187 , n19182 , n19186 );
and ( n19188 , n19186 , n5478 );
and ( n19189 , n19182 , n5478 );
or ( n19190 , n19187 , n19188 , n19189 );
and ( n19191 , n19190 , n5314 );
xor ( n19192 , n19173 , n19174 );
xor ( n19193 , n19192 , n19178 );
and ( n19194 , n5314 , n19193 );
and ( n19195 , n19190 , n19193 );
or ( n19196 , n19191 , n19194 , n19195 );
xor ( n19197 , n19181 , n19196 );
xor ( n19198 , n19197 , n7728 );
and ( n19199 , n19169 , n19198 );
and ( n19200 , n19165 , n19198 );
or ( n19201 , n19170 , n19199 , n19200 );
and ( n19202 , n19161 , n19201 );
and ( n19203 , n19181 , n19196 );
and ( n19204 , n19196 , n7728 );
and ( n19205 , n19181 , n7728 );
or ( n19206 , n19203 , n19204 , n19205 );
and ( n19207 , n5296 , n5325 );
and ( n19208 , n5309 , n5323 );
nor ( n19209 , n19207 , n19208 );
xnor ( n19210 , n19209 , n5333 );
xor ( n19211 , n19206 , n19210 );
and ( n19212 , n5254 , n5365 );
and ( n19213 , n5265 , n5363 );
nor ( n19214 , n19212 , n19213 );
xnor ( n19215 , n19214 , n5373 );
xor ( n19216 , n19211 , n19215 );
and ( n19217 , n19201 , n19216 );
and ( n19218 , n19161 , n19216 );
or ( n19219 , n19202 , n19217 , n19218 );
and ( n19220 , n7650 , n5325 );
and ( n19221 , n5296 , n5323 );
nor ( n19222 , n19220 , n19221 );
xnor ( n19223 , n19222 , n5333 );
and ( n19224 , n5285 , n5365 );
and ( n19225 , n5254 , n5363 );
nor ( n19226 , n19224 , n19225 );
xnor ( n19227 , n19226 , n5373 );
and ( n19228 , n19223 , n19227 );
xor ( n19229 , n19111 , n5314 );
xor ( n19230 , n19229 , n19114 );
and ( n19231 , n19227 , n19230 );
and ( n19232 , n19223 , n19230 );
or ( n19233 , n19228 , n19231 , n19232 );
and ( n19234 , n7647 , n5243 );
and ( n19235 , n7650 , n5241 );
nor ( n19236 , n19234 , n19235 );
xnor ( n19237 , n19236 , n5251 );
and ( n19238 , n19233 , n19237 );
xor ( n19239 , n19117 , n19120 );
xor ( n19240 , n19239 , n19123 );
and ( n19241 , n19237 , n19240 );
and ( n19242 , n19233 , n19240 );
or ( n19243 , n19238 , n19241 , n19242 );
and ( n19244 , n19219 , n19243 );
xor ( n19245 , n19126 , n19130 );
xor ( n19246 , n19245 , n19135 );
and ( n19247 , n19243 , n19246 );
and ( n19248 , n19219 , n19246 );
or ( n19249 , n19244 , n19247 , n19248 );
and ( n19250 , n5317 , n5282 );
and ( n19251 , n5328 , n5280 );
nor ( n19252 , n19250 , n19251 );
xnor ( n19253 , n19252 , n5290 );
and ( n19254 , n5233 , n5542 );
and ( n19255 , n5246 , n5540 );
nor ( n19256 , n19254 , n19255 );
xnor ( n19257 , n19256 , n5550 );
and ( n19258 , n19253 , n19257 );
and ( n19259 , n5274 , n7696 );
and ( n19260 , n5285 , n7694 );
nor ( n19261 , n19259 , n19260 );
xnor ( n19262 , n19261 , n7702 );
and ( n19263 , n19257 , n19262 );
and ( n19264 , n19253 , n19262 );
or ( n19265 , n19258 , n19263 , n19264 );
and ( n19266 , n19206 , n19210 );
and ( n19267 , n19210 , n19215 );
and ( n19268 , n19206 , n19215 );
or ( n19269 , n19266 , n19267 , n19268 );
and ( n19270 , n19265 , n19269 );
xor ( n19271 , n18977 , n18981 );
xor ( n19272 , n19271 , n18990 );
and ( n19273 , n19269 , n19272 );
and ( n19274 , n19265 , n19272 );
or ( n19275 , n19270 , n19273 , n19274 );
and ( n19276 , n19249 , n19275 );
xor ( n19277 , n19037 , n19039 );
and ( n19278 , n19275 , n19277 );
and ( n19279 , n19249 , n19277 );
or ( n19280 , n19276 , n19278 , n19279 );
and ( n19281 , n19144 , n19280 );
and ( n19282 , n19093 , n19280 );
or ( n19283 , n19145 , n19281 , n19282 );
xor ( n19284 , n19019 , n19045 );
xor ( n19285 , n19284 , n19047 );
and ( n19286 , n19283 , n19285 );
xor ( n19287 , n19080 , n19082 );
xor ( n19288 , n19287 , n19085 );
and ( n19289 , n19285 , n19288 );
and ( n19290 , n19283 , n19288 );
or ( n19291 , n19286 , n19289 , n19290 );
and ( n19292 , n19090 , n19291 );
and ( n19293 , n19088 , n19291 );
or ( n19294 , n19091 , n19292 , n19293 );
and ( n19295 , n19059 , n19294 );
and ( n19296 , n19057 , n19294 );
or ( n19297 , n19060 , n19295 , n19296 );
and ( n19298 , n18928 , n19297 );
and ( n19299 , n18857 , n19298 );
xor ( n19300 , n18637 , n18735 );
and ( n19301 , n19299 , n19300 );
xor ( n19302 , n18676 , n18729 );
xor ( n19303 , n19302 , n18732 );
xor ( n19304 , n18857 , n19298 );
and ( n19305 , n19303 , n19304 );
xor ( n19306 , n18780 , n18851 );
xor ( n19307 , n19306 , n18854 );
xor ( n19308 , n18928 , n19297 );
and ( n19309 , n19307 , n19308 );
xor ( n19310 , n18884 , n18927 );
xor ( n19311 , n19057 , n19059 );
xor ( n19312 , n19311 , n19294 );
and ( n19313 , n19310 , n19312 );
xor ( n19314 , n19050 , n19051 );
xor ( n19315 , n19314 , n19054 );
xor ( n19316 , n19088 , n19090 );
xor ( n19317 , n19316 , n19291 );
and ( n19318 , n19315 , n19317 );
xor ( n19319 , n19035 , n19040 );
xor ( n19320 , n19319 , n19042 );
xor ( n19321 , n19064 , n19074 );
xor ( n19322 , n19321 , n19077 );
and ( n19323 , n19320 , n19322 );
and ( n19324 , n5350 , n5262 );
and ( n19325 , n7716 , n5260 );
nor ( n19326 , n19324 , n19325 );
xnor ( n19327 , n19326 , n5270 );
and ( n19328 , n5368 , n7633 );
and ( n19329 , n5529 , n5512 );
nor ( n19330 , n19328 , n19329 );
xnor ( n19331 , n19330 , n5561 );
and ( n19332 , n19327 , n19331 );
and ( n19333 , n5355 , n5342 );
and ( n19334 , n19331 , n19333 );
and ( n19335 , n19327 , n19333 );
or ( n19336 , n19332 , n19334 , n19335 );
xor ( n19337 , n19097 , n19101 );
xor ( n19338 , n19337 , n19103 );
and ( n19339 , n19336 , n19338 );
xor ( n19340 , n18932 , n18936 );
xor ( n19341 , n19340 , n18970 );
and ( n19342 , n19338 , n19341 );
and ( n19343 , n19336 , n19341 );
or ( n19344 , n19339 , n19342 , n19343 );
xor ( n19345 , n18973 , n18993 );
xor ( n19346 , n19345 , n19008 );
and ( n19347 , n19344 , n19346 );
xor ( n19348 , n19106 , n19138 );
xor ( n19349 , n19348 , n19141 );
and ( n19350 , n19346 , n19349 );
and ( n19351 , n19344 , n19349 );
or ( n19352 , n19347 , n19350 , n19351 );
and ( n19353 , n19322 , n19352 );
and ( n19354 , n19320 , n19352 );
or ( n19355 , n19323 , n19353 , n19354 );
xor ( n19356 , n19283 , n19285 );
xor ( n19357 , n19356 , n19288 );
and ( n19358 , n19355 , n19357 );
xor ( n19359 , n19093 , n19144 );
xor ( n19360 , n19359 , n19280 );
xor ( n19361 , n19320 , n19322 );
xor ( n19362 , n19361 , n19352 );
and ( n19363 , n19360 , n19362 );
xor ( n19364 , n19149 , n19153 );
xor ( n19365 , n19364 , n19158 );
and ( n19366 , n5393 , n5414 );
not ( n19367 , n19366 );
xnor ( n19368 , n19367 , n5420 );
and ( n19369 , n5437 , n7863 );
not ( n19370 , n19369 );
xnor ( n19371 , n19370 , n5429 );
and ( n19372 , n19368 , n19371 );
and ( n19373 , n19371 , n5478 );
and ( n19374 , n19368 , n5478 );
or ( n19375 , n19372 , n19373 , n19374 );
and ( n19376 , n5408 , n5468 );
and ( n19377 , n5377 , n5438 );
nor ( n19378 , n19376 , n19377 );
xnor ( n19379 , n19378 , n5405 );
buf ( n19380 , n19379 );
and ( n19381 , n19375 , n19380 );
and ( n19382 , n5377 , n5468 );
and ( n19383 , n5393 , n5438 );
nor ( n19384 , n19382 , n19383 );
xnor ( n19385 , n19384 , n5405 );
and ( n19386 , n19380 , n19385 );
and ( n19387 , n19375 , n19385 );
or ( n19388 , n19381 , n19386 , n19387 );
and ( n19389 , n7711 , n7722 );
not ( n19390 , n19389 );
xnor ( n19391 , n19390 , n7728 );
and ( n19392 , n19388 , n19391 );
xor ( n19393 , n19190 , n5314 );
xor ( n19394 , n19393 , n19193 );
and ( n19395 , n19391 , n19394 );
and ( n19396 , n19388 , n19394 );
or ( n19397 , n19392 , n19395 , n19396 );
and ( n19398 , n7716 , n5243 );
and ( n19399 , n7647 , n5241 );
nor ( n19400 , n19398 , n19399 );
xnor ( n19401 , n19400 , n5251 );
xor ( n19402 , n19397 , n19401 );
and ( n19403 , n5545 , n5342 );
xor ( n19404 , n19402 , n19403 );
and ( n19405 , n19365 , n19404 );
xor ( n19406 , n19223 , n19227 );
xor ( n19407 , n19406 , n19230 );
and ( n19408 , n19404 , n19407 );
and ( n19409 , n19365 , n19407 );
or ( n19410 , n19405 , n19408 , n19409 );
xor ( n19411 , n19161 , n19201 );
xor ( n19412 , n19411 , n19216 );
and ( n19413 , n19410 , n19412 );
and ( n19414 , n19397 , n19401 );
and ( n19415 , n19401 , n19403 );
and ( n19416 , n19397 , n19403 );
or ( n19417 , n19414 , n19415 , n19416 );
xor ( n19418 , n19327 , n19331 );
xor ( n19419 , n19418 , n19333 );
xor ( n19420 , n19417 , n19419 );
xor ( n19421 , n19253 , n19257 );
xor ( n19422 , n19421 , n19262 );
xor ( n19423 , n19420 , n19422 );
and ( n19424 , n19412 , n19423 );
and ( n19425 , n19410 , n19423 );
or ( n19426 , n19413 , n19424 , n19425 );
and ( n19427 , n5350 , n5243 );
and ( n19428 , n7716 , n5241 );
nor ( n19429 , n19427 , n19428 );
xnor ( n19430 , n19429 , n5251 );
and ( n19431 , n5368 , n7696 );
and ( n19432 , n5529 , n7694 );
nor ( n19433 , n19431 , n19432 );
xnor ( n19434 , n19433 , n7702 );
and ( n19435 , n19430 , n19434 );
and ( n19436 , n5536 , n5342 );
and ( n19437 , n19434 , n19436 );
and ( n19438 , n19430 , n19436 );
or ( n19439 , n19435 , n19437 , n19438 );
and ( n19440 , n5296 , n5499 );
and ( n19441 , n5309 , n5497 );
nor ( n19442 , n19440 , n19441 );
xnor ( n19443 , n19442 , n5505 );
and ( n19444 , n5233 , n5282 );
and ( n19445 , n5246 , n5280 );
nor ( n19446 , n19444 , n19445 );
xnor ( n19447 , n19446 , n5290 );
and ( n19448 , n19443 , n19447 );
and ( n19449 , n5545 , n7633 );
and ( n19450 , n5355 , n5512 );
nor ( n19451 , n19449 , n19450 );
xnor ( n19452 , n19451 , n5561 );
and ( n19453 , n19447 , n19452 );
and ( n19454 , n19443 , n19452 );
or ( n19455 , n19448 , n19453 , n19454 );
and ( n19456 , n19439 , n19455 );
and ( n19457 , n5317 , n5262 );
and ( n19458 , n5328 , n5260 );
nor ( n19459 , n19457 , n19458 );
xnor ( n19460 , n19459 , n5270 );
and ( n19461 , n5254 , n5542 );
and ( n19462 , n5265 , n5540 );
nor ( n19463 , n19461 , n19462 );
xnor ( n19464 , n19463 , n5550 );
and ( n19465 , n19460 , n19464 );
xor ( n19466 , n19388 , n19391 );
xor ( n19467 , n19466 , n19394 );
and ( n19468 , n19464 , n19467 );
and ( n19469 , n19460 , n19467 );
or ( n19470 , n19465 , n19468 , n19469 );
and ( n19471 , n19455 , n19470 );
and ( n19472 , n19439 , n19470 );
or ( n19473 , n19456 , n19471 , n19472 );
and ( n19474 , n5472 , n5429 );
and ( n19475 , n5429 , n5478 );
and ( n19476 , n5472 , n5478 );
or ( n19477 , n19474 , n19475 , n19476 );
buf ( n19478 , n5463 );
and ( n19479 , n19477 , n19478 );
not ( n19480 , n19379 );
and ( n19481 , n19478 , n19480 );
and ( n19482 , n19477 , n19480 );
or ( n19483 , n19479 , n19481 , n19482 );
and ( n19484 , n19483 , n5314 );
xor ( n19485 , n19182 , n19186 );
xor ( n19486 , n19485 , n5478 );
and ( n19487 , n5314 , n19486 );
and ( n19488 , n19483 , n19486 );
or ( n19489 , n19484 , n19487 , n19488 );
and ( n19490 , n7647 , n5325 );
and ( n19491 , n7650 , n5323 );
nor ( n19492 , n19490 , n19491 );
xnor ( n19493 , n19492 , n5333 );
and ( n19494 , n19489 , n19493 );
and ( n19495 , n5274 , n5365 );
and ( n19496 , n5285 , n5363 );
nor ( n19497 , n19495 , n19496 );
xnor ( n19498 , n19497 , n5373 );
and ( n19499 , n19493 , n19498 );
and ( n19500 , n19489 , n19498 );
or ( n19501 , n19494 , n19499 , n19500 );
and ( n19502 , n5529 , n7696 );
and ( n19503 , n5274 , n7694 );
nor ( n19504 , n19502 , n19503 );
xnor ( n19505 , n19504 , n7702 );
and ( n19506 , n19501 , n19505 );
xor ( n19507 , n19165 , n19169 );
xor ( n19508 , n19507 , n19198 );
and ( n19509 , n19505 , n19508 );
and ( n19510 , n19501 , n19508 );
or ( n19511 , n19506 , n19509 , n19510 );
and ( n19512 , n19473 , n19511 );
xor ( n19513 , n19233 , n19237 );
xor ( n19514 , n19513 , n19240 );
and ( n19515 , n19511 , n19514 );
and ( n19516 , n19473 , n19514 );
or ( n19517 , n19512 , n19515 , n19516 );
and ( n19518 , n19426 , n19517 );
xor ( n19519 , n19219 , n19243 );
xor ( n19520 , n19519 , n19246 );
and ( n19521 , n19517 , n19520 );
and ( n19522 , n19426 , n19520 );
or ( n19523 , n19518 , n19521 , n19522 );
and ( n19524 , n19417 , n19419 );
and ( n19525 , n19419 , n19422 );
and ( n19526 , n19417 , n19422 );
or ( n19527 , n19524 , n19525 , n19526 );
xor ( n19528 , n19336 , n19338 );
xor ( n19529 , n19528 , n19341 );
and ( n19530 , n19527 , n19529 );
xor ( n19531 , n19265 , n19269 );
xor ( n19532 , n19531 , n19272 );
and ( n19533 , n19529 , n19532 );
and ( n19534 , n19527 , n19532 );
or ( n19535 , n19530 , n19533 , n19534 );
or ( n19536 , n19523 , n19535 );
and ( n19537 , n19362 , n19536 );
and ( n19538 , n19360 , n19536 );
or ( n19539 , n19363 , n19537 , n19538 );
and ( n19540 , n19357 , n19539 );
and ( n19541 , n19355 , n19539 );
or ( n19542 , n19358 , n19540 , n19541 );
and ( n19543 , n19317 , n19542 );
and ( n19544 , n19315 , n19542 );
or ( n19545 , n19318 , n19543 , n19544 );
and ( n19546 , n19312 , n19545 );
and ( n19547 , n19310 , n19545 );
or ( n19548 , n19313 , n19546 , n19547 );
and ( n19549 , n19308 , n19548 );
and ( n19550 , n19307 , n19548 );
or ( n19551 , n19309 , n19549 , n19550 );
and ( n19552 , n19304 , n19551 );
and ( n19553 , n19303 , n19551 );
or ( n19554 , n19305 , n19552 , n19553 );
and ( n19555 , n19300 , n19554 );
and ( n19556 , n19299 , n19554 );
or ( n19557 , n19301 , n19555 , n19556 );
and ( n19558 , n18737 , n19557 );
and ( n19559 , n18736 , n19557 );
or ( n19560 , n18738 , n19558 , n19559 );
and ( n19561 , n18634 , n19560 );
and ( n19562 , n18633 , n19560 );
or ( n19563 , n18635 , n19561 , n19562 );
and ( n19564 , n18519 , n19563 );
and ( n19565 , n18517 , n19563 );
or ( n19566 , n18520 , n19564 , n19565 );
and ( n19567 , n18437 , n19566 );
xor ( n19568 , n18517 , n18519 );
xor ( n19569 , n19568 , n19563 );
xor ( n19570 , n18633 , n18634 );
xor ( n19571 , n19570 , n19560 );
xor ( n19572 , n18736 , n18737 );
xor ( n19573 , n19572 , n19557 );
xor ( n19574 , n19299 , n19300 );
xor ( n19575 , n19574 , n19554 );
xor ( n19576 , n19303 , n19304 );
xor ( n19577 , n19576 , n19551 );
xor ( n19578 , n19307 , n19308 );
xor ( n19579 , n19578 , n19548 );
xor ( n19580 , n19310 , n19312 );
xor ( n19581 , n19580 , n19545 );
xor ( n19582 , n19315 , n19317 );
xor ( n19583 , n19582 , n19542 );
xor ( n19584 , n19355 , n19357 );
xor ( n19585 , n19584 , n19539 );
xor ( n19586 , n19249 , n19275 );
xor ( n19587 , n19586 , n19277 );
xor ( n19588 , n19344 , n19346 );
xor ( n19589 , n19588 , n19349 );
and ( n19590 , n19587 , n19589 );
xnor ( n19591 , n19523 , n19535 );
and ( n19592 , n19589 , n19591 );
and ( n19593 , n19587 , n19591 );
or ( n19594 , n19590 , n19592 , n19593 );
xor ( n19595 , n19360 , n19362 );
xor ( n19596 , n19595 , n19536 );
and ( n19597 , n19594 , n19596 );
and ( n19598 , n5265 , n5282 );
and ( n19599 , n5233 , n5280 );
nor ( n19600 , n19598 , n19599 );
xnor ( n19601 , n19600 , n5290 );
and ( n19602 , n5529 , n5365 );
and ( n19603 , n5274 , n5363 );
nor ( n19604 , n19602 , n19603 );
xnor ( n19605 , n19604 , n5373 );
and ( n19606 , n19601 , n19605 );
and ( n19607 , n7660 , n5342 );
and ( n19608 , n19605 , n19607 );
and ( n19609 , n19601 , n19607 );
or ( n19610 , n19606 , n19608 , n19609 );
and ( n19611 , n5246 , n5262 );
and ( n19612 , n5317 , n5260 );
nor ( n19613 , n19611 , n19612 );
xnor ( n19614 , n19613 , n5270 );
and ( n19615 , n5285 , n5542 );
and ( n19616 , n5254 , n5540 );
nor ( n19617 , n19615 , n19616 );
xnor ( n19618 , n19617 , n5550 );
and ( n19619 , n19614 , n19618 );
and ( n19620 , n5536 , n7633 );
and ( n19621 , n5545 , n5512 );
nor ( n19622 , n19620 , n19621 );
xnor ( n19623 , n19622 , n5561 );
and ( n19624 , n19618 , n19623 );
and ( n19625 , n19614 , n19623 );
or ( n19626 , n19619 , n19624 , n19625 );
and ( n19627 , n19610 , n19626 );
xor ( n19628 , n19489 , n19493 );
xor ( n19629 , n19628 , n19498 );
and ( n19630 , n19626 , n19629 );
and ( n19631 , n19610 , n19629 );
or ( n19632 , n19627 , n19630 , n19631 );
and ( n19633 , n5309 , n7722 );
and ( n19634 , n7711 , n7720 );
nor ( n19635 , n19633 , n19634 );
xnor ( n19636 , n19635 , n7728 );
and ( n19637 , n7650 , n5499 );
and ( n19638 , n5296 , n5497 );
nor ( n19639 , n19637 , n19638 );
xnor ( n19640 , n19639 , n5505 );
and ( n19641 , n19636 , n19640 );
and ( n19642 , n7716 , n5325 );
and ( n19643 , n7647 , n5323 );
nor ( n19644 , n19642 , n19643 );
xnor ( n19645 , n19644 , n5333 );
and ( n19646 , n19640 , n19645 );
and ( n19647 , n19636 , n19645 );
or ( n19648 , n19641 , n19646 , n19647 );
and ( n19649 , n5459 , n5464 );
and ( n19650 , n5464 , n5479 );
and ( n19651 , n5459 , n5479 );
or ( n19652 , n19649 , n19650 , n19651 );
xor ( n19653 , n19368 , n19371 );
xor ( n19654 , n19653 , n5478 );
and ( n19655 , n19652 , n19654 );
xor ( n19656 , n19477 , n19478 );
xor ( n19657 , n19656 , n19480 );
and ( n19658 , n19654 , n19657 );
and ( n19659 , n19652 , n19657 );
or ( n19660 , n19655 , n19658 , n19659 );
xor ( n19661 , n19375 , n19380 );
xor ( n19662 , n19661 , n19385 );
and ( n19663 , n19660 , n19662 );
xor ( n19664 , n19483 , n5314 );
xor ( n19665 , n19664 , n19486 );
and ( n19666 , n19662 , n19665 );
and ( n19667 , n19660 , n19665 );
or ( n19668 , n19663 , n19666 , n19667 );
and ( n19669 , n19648 , n19668 );
xor ( n19670 , n19443 , n19447 );
xor ( n19671 , n19670 , n19452 );
and ( n19672 , n19668 , n19671 );
and ( n19673 , n19648 , n19671 );
or ( n19674 , n19669 , n19672 , n19673 );
and ( n19675 , n19632 , n19674 );
xor ( n19676 , n19501 , n19505 );
xor ( n19677 , n19676 , n19508 );
and ( n19678 , n19674 , n19677 );
and ( n19679 , n19632 , n19677 );
or ( n19680 , n19675 , n19678 , n19679 );
and ( n19681 , n5328 , n5243 );
and ( n19682 , n5350 , n5241 );
nor ( n19683 , n19681 , n19682 );
xnor ( n19684 , n19683 , n5251 );
and ( n19685 , n5355 , n7696 );
and ( n19686 , n5368 , n7694 );
nor ( n19687 , n19685 , n19686 );
xnor ( n19688 , n19687 , n7702 );
and ( n19689 , n19684 , n19688 );
xor ( n19690 , n19660 , n19662 );
xor ( n19691 , n19690 , n19665 );
and ( n19692 , n19688 , n19691 );
and ( n19693 , n19684 , n19691 );
or ( n19694 , n19689 , n19692 , n19693 );
xor ( n19695 , n19430 , n19434 );
xor ( n19696 , n19695 , n19436 );
and ( n19697 , n19694 , n19696 );
xor ( n19698 , n19460 , n19464 );
xor ( n19699 , n19698 , n19467 );
and ( n19700 , n19696 , n19699 );
and ( n19701 , n19694 , n19699 );
or ( n19702 , n19697 , n19700 , n19701 );
xor ( n19703 , n19439 , n19455 );
xor ( n19704 , n19703 , n19470 );
and ( n19705 , n19702 , n19704 );
xor ( n19706 , n19365 , n19404 );
xor ( n19707 , n19706 , n19407 );
and ( n19708 , n19704 , n19707 );
and ( n19709 , n19702 , n19707 );
or ( n19710 , n19705 , n19708 , n19709 );
and ( n19711 , n19680 , n19710 );
xor ( n19712 , n19473 , n19511 );
xor ( n19713 , n19712 , n19514 );
and ( n19714 , n19710 , n19713 );
and ( n19715 , n19680 , n19713 );
or ( n19716 , n19711 , n19714 , n19715 );
xor ( n19717 , n19426 , n19517 );
xor ( n19718 , n19717 , n19520 );
and ( n19719 , n19716 , n19718 );
xor ( n19720 , n19527 , n19529 );
xor ( n19721 , n19720 , n19532 );
and ( n19722 , n19718 , n19721 );
and ( n19723 , n19716 , n19721 );
or ( n19724 , n19719 , n19722 , n19723 );
xor ( n19725 , n19716 , n19718 );
xor ( n19726 , n19725 , n19721 );
and ( n19727 , n5233 , n5262 );
and ( n19728 , n5246 , n5260 );
nor ( n19729 , n19727 , n19728 );
xnor ( n19730 , n19729 , n5270 );
and ( n19731 , n7660 , n7633 );
and ( n19732 , n5536 , n5512 );
nor ( n19733 , n19731 , n19732 );
xnor ( n19734 , n19733 , n5561 );
and ( n19735 , n19730 , n19734 );
and ( n19736 , n7690 , n5342 );
and ( n19737 , n19734 , n19736 );
and ( n19738 , n19730 , n19736 );
or ( n19739 , n19735 , n19737 , n19738 );
and ( n19740 , n5432 , n5457 );
and ( n19741 , n5457 , n5480 );
and ( n19742 , n5432 , n5480 );
or ( n19743 , n19740 , n19741 , n19742 );
and ( n19744 , n7647 , n5499 );
and ( n19745 , n7650 , n5497 );
nor ( n19746 , n19744 , n19745 );
xnor ( n19747 , n19746 , n5505 );
and ( n19748 , n19743 , n19747 );
and ( n19749 , n5350 , n5325 );
and ( n19750 , n7716 , n5323 );
nor ( n19751 , n19749 , n19750 );
xnor ( n19752 , n19751 , n5333 );
and ( n19753 , n19747 , n19752 );
and ( n19754 , n19743 , n19752 );
or ( n19755 , n19748 , n19753 , n19754 );
and ( n19756 , n19739 , n19755 );
and ( n19757 , n7711 , n5306 );
not ( n19758 , n19757 );
xnor ( n19759 , n19758 , n5314 );
and ( n19760 , n5296 , n7722 );
and ( n19761 , n5309 , n7720 );
nor ( n19762 , n19760 , n19761 );
xnor ( n19763 , n19762 , n7728 );
and ( n19764 , n19759 , n19763 );
xor ( n19765 , n19652 , n19654 );
xor ( n19766 , n19765 , n19657 );
and ( n19767 , n19763 , n19766 );
and ( n19768 , n19759 , n19766 );
or ( n19769 , n19764 , n19767 , n19768 );
and ( n19770 , n19755 , n19769 );
and ( n19771 , n19739 , n19769 );
or ( n19772 , n19756 , n19770 , n19771 );
and ( n19773 , n5317 , n5243 );
and ( n19774 , n5328 , n5241 );
nor ( n19775 , n19773 , n19774 );
xnor ( n19776 , n19775 , n5251 );
and ( n19777 , n5254 , n5282 );
and ( n19778 , n5265 , n5280 );
nor ( n19779 , n19777 , n19778 );
xnor ( n19780 , n19779 , n5290 );
and ( n19781 , n19776 , n19780 );
and ( n19782 , n5368 , n5365 );
and ( n19783 , n5529 , n5363 );
nor ( n19784 , n19782 , n19783 );
xnor ( n19785 , n19784 , n5373 );
and ( n19786 , n19780 , n19785 );
and ( n19787 , n19776 , n19785 );
or ( n19788 , n19781 , n19786 , n19787 );
xor ( n19789 , n19601 , n19605 );
xor ( n19790 , n19789 , n19607 );
and ( n19791 , n19788 , n19790 );
xor ( n19792 , n19636 , n19640 );
xor ( n19793 , n19792 , n19645 );
and ( n19794 , n19790 , n19793 );
and ( n19795 , n19788 , n19793 );
or ( n19796 , n19791 , n19794 , n19795 );
and ( n19797 , n19772 , n19796 );
xor ( n19798 , n19648 , n19668 );
xor ( n19799 , n19798 , n19671 );
and ( n19800 , n19796 , n19799 );
and ( n19801 , n19772 , n19799 );
or ( n19802 , n19797 , n19800 , n19801 );
and ( n19803 , n5353 , n5374 );
and ( n19804 , n5374 , n5481 );
and ( n19805 , n5353 , n5481 );
or ( n19806 , n19803 , n19804 , n19805 );
and ( n19807 , n5274 , n5542 );
and ( n19808 , n5285 , n5540 );
nor ( n19809 , n19807 , n19808 );
xnor ( n19810 , n19809 , n5550 );
and ( n19811 , n19806 , n19810 );
and ( n19812 , n5545 , n7696 );
and ( n19813 , n5355 , n7694 );
nor ( n19814 , n19812 , n19813 );
xnor ( n19815 , n19814 , n7702 );
and ( n19816 , n19810 , n19815 );
and ( n19817 , n19806 , n19815 );
or ( n19818 , n19811 , n19816 , n19817 );
xor ( n19819 , n19614 , n19618 );
xor ( n19820 , n19819 , n19623 );
and ( n19821 , n19818 , n19820 );
xor ( n19822 , n19684 , n19688 );
xor ( n19823 , n19822 , n19691 );
and ( n19824 , n19820 , n19823 );
and ( n19825 , n19818 , n19823 );
or ( n19826 , n19821 , n19824 , n19825 );
xor ( n19827 , n19610 , n19626 );
xor ( n19828 , n19827 , n19629 );
and ( n19829 , n19826 , n19828 );
xor ( n19830 , n19694 , n19696 );
xor ( n19831 , n19830 , n19699 );
and ( n19832 , n19828 , n19831 );
and ( n19833 , n19826 , n19831 );
or ( n19834 , n19829 , n19832 , n19833 );
and ( n19835 , n19802 , n19834 );
xor ( n19836 , n19632 , n19674 );
xor ( n19837 , n19836 , n19677 );
and ( n19838 , n19834 , n19837 );
and ( n19839 , n19802 , n19837 );
or ( n19840 , n19835 , n19838 , n19839 );
xor ( n19841 , n19410 , n19412 );
xor ( n19842 , n19841 , n19423 );
and ( n19843 , n19840 , n19842 );
xor ( n19844 , n19680 , n19710 );
xor ( n19845 , n19844 , n19713 );
and ( n19846 , n19842 , n19845 );
and ( n19847 , n19840 , n19845 );
or ( n19848 , n19843 , n19846 , n19847 );
and ( n19849 , n19726 , n19848 );
and ( n19850 , n19724 , n19849 );
xor ( n19851 , n19587 , n19589 );
xor ( n19852 , n19851 , n19591 );
and ( n19853 , n19849 , n19852 );
and ( n19854 , n19724 , n19852 );
or ( n19855 , n19850 , n19853 , n19854 );
and ( n19856 , n19596 , n19855 );
and ( n19857 , n19594 , n19855 );
or ( n19858 , n19597 , n19856 , n19857 );
and ( n19859 , n19585 , n19858 );
xor ( n19860 , n19594 , n19596 );
xor ( n19861 , n19860 , n19855 );
xor ( n19862 , n19724 , n19849 );
xor ( n19863 , n19862 , n19852 );
xor ( n19864 , n19788 , n19790 );
xor ( n19865 , n19864 , n19793 );
xor ( n19866 , n19730 , n19734 );
xor ( n19867 , n19866 , n19736 );
and ( n19868 , n8176 , n8180 );
and ( n19869 , n8180 , n8185 );
and ( n19870 , n8176 , n8185 );
or ( n19871 , n19868 , n19869 , n19870 );
and ( n19872 , n19867 , n19871 );
and ( n19873 , n19865 , n19872 );
and ( n19874 , n8191 , n8192 );
and ( n19875 , n8151 , n8165 );
and ( n19876 , n8165 , n8170 );
and ( n19877 , n8151 , n8170 );
or ( n19878 , n19875 , n19876 , n19877 );
and ( n19879 , n19874 , n19878 );
and ( n19880 , n8175 , n8186 );
and ( n19881 , n8186 , n8193 );
and ( n19882 , n8175 , n8193 );
or ( n19883 , n19880 , n19881 , n19882 );
and ( n19884 , n19878 , n19883 );
and ( n19885 , n19874 , n19883 );
or ( n19886 , n19879 , n19884 , n19885 );
xor ( n19887 , n19865 , n19872 );
and ( n19888 , n19886 , n19887 );
xor ( n19889 , n19867 , n19871 );
and ( n19890 , n8118 , n8119 );
and ( n19891 , n8119 , n8121 );
and ( n19892 , n8118 , n8121 );
or ( n19893 , n19890 , n19891 , n19892 );
and ( n19894 , n19889 , n19893 );
xor ( n19895 , n19874 , n19878 );
xor ( n19896 , n19895 , n19883 );
and ( n19897 , n19893 , n19896 );
and ( n19898 , n19889 , n19896 );
or ( n19899 , n19894 , n19897 , n19898 );
and ( n19900 , n19887 , n19899 );
and ( n19901 , n19886 , n19899 );
or ( n19902 , n19888 , n19900 , n19901 );
and ( n19903 , n19873 , n19902 );
xor ( n19904 , n19702 , n19704 );
xor ( n19905 , n19904 , n19707 );
and ( n19906 , n19903 , n19905 );
xor ( n19907 , n19840 , n19842 );
xor ( n19908 , n19907 , n19845 );
and ( n19909 , n19906 , n19908 );
xor ( n19910 , n19726 , n19848 );
and ( n19911 , n19909 , n19910 );
xor ( n19912 , n19873 , n19902 );
xor ( n19913 , n19772 , n19796 );
xor ( n19914 , n19913 , n19799 );
and ( n19915 , n19912 , n19914 );
and ( n19916 , n8171 , n8194 );
and ( n19917 , n8194 , n8199 );
and ( n19918 , n8171 , n8199 );
or ( n19919 , n19916 , n19917 , n19918 );
and ( n19920 , n8109 , n8113 );
and ( n19921 , n8113 , n8122 );
and ( n19922 , n8109 , n8122 );
or ( n19923 , n19920 , n19921 , n19922 );
and ( n19924 , n19919 , n19923 );
xor ( n19925 , n19889 , n19893 );
xor ( n19926 , n19925 , n19896 );
and ( n19927 , n19923 , n19926 );
and ( n19928 , n19919 , n19926 );
or ( n19929 , n19924 , n19927 , n19928 );
xor ( n19930 , n19886 , n19887 );
xor ( n19931 , n19930 , n19899 );
and ( n19932 , n19929 , n19931 );
xor ( n19933 , n19739 , n19755 );
xor ( n19934 , n19933 , n19769 );
and ( n19935 , n19931 , n19934 );
and ( n19936 , n19929 , n19934 );
or ( n19937 , n19932 , n19935 , n19936 );
and ( n19938 , n19914 , n19937 );
and ( n19939 , n19912 , n19937 );
or ( n19940 , n19915 , n19938 , n19939 );
xor ( n19941 , n19802 , n19834 );
xor ( n19942 , n19941 , n19837 );
and ( n19943 , n19940 , n19942 );
and ( n19944 , n8155 , n8159 );
and ( n19945 , n8159 , n8164 );
and ( n19946 , n8155 , n8164 );
or ( n19947 , n19944 , n19945 , n19946 );
xor ( n19948 , n19776 , n19780 );
xor ( n19949 , n19948 , n19785 );
and ( n19950 , n19947 , n19949 );
xor ( n19951 , n19743 , n19747 );
xor ( n19952 , n19951 , n19752 );
and ( n19953 , n19949 , n19952 );
and ( n19954 , n19947 , n19952 );
or ( n19955 , n19950 , n19953 , n19954 );
and ( n19956 , n8141 , n8145 );
and ( n19957 , n8145 , n8150 );
and ( n19958 , n8141 , n8150 );
or ( n19959 , n19956 , n19957 , n19958 );
not ( n19960 , n19959 );
xor ( n19961 , n19759 , n19763 );
xor ( n19962 , n19961 , n19766 );
and ( n19963 , n19960 , n19962 );
and ( n19964 , n19955 , n19963 );
buf ( n19965 , n19959 );
and ( n19966 , n19963 , n19965 );
and ( n19967 , n19955 , n19965 );
or ( n19968 , n19964 , n19966 , n19967 );
xor ( n19969 , n19826 , n19828 );
xor ( n19970 , n19969 , n19831 );
and ( n19971 , n19968 , n19970 );
xor ( n19972 , n19818 , n19820 );
xor ( n19973 , n19972 , n19823 );
and ( n19974 , n8132 , n8136 );
and ( n19975 , n8136 , n8200 );
and ( n19976 , n8132 , n8200 );
or ( n19977 , n19974 , n19975 , n19976 );
xor ( n19978 , n19919 , n19923 );
xor ( n19979 , n19978 , n19926 );
and ( n19980 , n19977 , n19979 );
xor ( n19981 , n19806 , n19810 );
xor ( n19982 , n19981 , n19815 );
and ( n19983 , n19979 , n19982 );
and ( n19984 , n19977 , n19982 );
or ( n19985 , n19980 , n19983 , n19984 );
and ( n19986 , n19973 , n19985 );
xor ( n19987 , n19947 , n19949 );
xor ( n19988 , n19987 , n19952 );
xor ( n19989 , n19960 , n19962 );
and ( n19990 , n19988 , n19989 );
and ( n19991 , n5294 , n5346 );
and ( n19992 , n5346 , n5482 );
and ( n19993 , n5294 , n5482 );
or ( n19994 , n19991 , n19992 , n19993 );
and ( n19995 , n19989 , n19994 );
and ( n19996 , n19988 , n19994 );
or ( n19997 , n19990 , n19995 , n19996 );
and ( n19998 , n19985 , n19997 );
and ( n19999 , n19973 , n19997 );
or ( n20000 , n19986 , n19998 , n19999 );
and ( n20001 , n19970 , n20000 );
and ( n20002 , n19968 , n20000 );
or ( n20003 , n19971 , n20001 , n20002 );
and ( n20004 , n19942 , n20003 );
and ( n20005 , n19940 , n20003 );
or ( n20006 , n19943 , n20004 , n20005 );
xor ( n20007 , n19903 , n19905 );
xor ( n20008 , n19912 , n19914 );
xor ( n20009 , n20008 , n19937 );
xor ( n20010 , n19929 , n19931 );
xor ( n20011 , n20010 , n19934 );
xor ( n20012 , n19955 , n19963 );
xor ( n20013 , n20012 , n19965 );
and ( n20014 , n20011 , n20013 );
and ( n20015 , n8123 , n8127 );
and ( n20016 , n8127 , n8201 );
and ( n20017 , n8123 , n8201 );
or ( n20018 , n20015 , n20016 , n20017 );
and ( n20019 , n5483 , n8104 );
and ( n20020 , n8104 , n8202 );
and ( n20021 , n5483 , n8202 );
or ( n20022 , n20019 , n20020 , n20021 );
and ( n20023 , n20018 , n20022 );
xor ( n20024 , n19977 , n19979 );
xor ( n20025 , n20024 , n19982 );
and ( n20026 , n20022 , n20025 );
and ( n20027 , n20018 , n20025 );
or ( n20028 , n20023 , n20026 , n20027 );
and ( n20029 , n20013 , n20028 );
and ( n20030 , n20011 , n20028 );
or ( n20031 , n20014 , n20029 , n20030 );
and ( n20032 , n20009 , n20031 );
xor ( n20033 , n19968 , n19970 );
xor ( n20034 , n20033 , n20000 );
and ( n20035 , n20031 , n20034 );
and ( n20036 , n20009 , n20034 );
or ( n20037 , n20032 , n20035 , n20036 );
and ( n20038 , n20007 , n20037 );
xor ( n20039 , n19940 , n19942 );
xor ( n20040 , n20039 , n20003 );
and ( n20041 , n20037 , n20040 );
and ( n20042 , n20007 , n20040 );
or ( n20043 , n20038 , n20041 , n20042 );
and ( n20044 , n20006 , n20043 );
xor ( n20045 , n19906 , n19908 );
and ( n20046 , n20043 , n20045 );
and ( n20047 , n20006 , n20045 );
or ( n20048 , n20044 , n20046 , n20047 );
and ( n20049 , n19910 , n20048 );
and ( n20050 , n19909 , n20048 );
or ( n20051 , n19911 , n20049 , n20050 );
and ( n20052 , n19863 , n20051 );
xor ( n20053 , n19909 , n19910 );
xor ( n20054 , n20053 , n20048 );
xor ( n20055 , n20006 , n20043 );
xor ( n20056 , n20055 , n20045 );
xor ( n20057 , n20007 , n20037 );
xor ( n20058 , n20057 , n20040 );
xor ( n20059 , n20009 , n20031 );
xor ( n20060 , n20059 , n20034 );
xor ( n20061 , n19973 , n19985 );
xor ( n20062 , n20061 , n19997 );
xor ( n20063 , n20011 , n20013 );
xor ( n20064 , n20063 , n20028 );
and ( n20065 , n20062 , n20064 );
xor ( n20066 , n19988 , n19989 );
xor ( n20067 , n20066 , n19994 );
xor ( n20068 , n20018 , n20022 );
xor ( n20069 , n20068 , n20025 );
and ( n20070 , n20067 , n20069 );
or ( n20071 , n8203 , n8499 );
and ( n20072 , n20069 , n20071 );
and ( n20073 , n20067 , n20071 );
or ( n20074 , n20070 , n20072 , n20073 );
and ( n20075 , n20064 , n20074 );
and ( n20076 , n20062 , n20074 );
or ( n20077 , n20065 , n20075 , n20076 );
or ( n20078 , n20060 , n20077 );
or ( n20079 , n20058 , n20078 );
or ( n20080 , n20056 , n20079 );
or ( n20081 , n20054 , n20080 );
and ( n20082 , n20051 , n20081 );
and ( n20083 , n19863 , n20081 );
or ( n20084 , n20052 , n20082 , n20083 );
or ( n20085 , n19861 , n20084 );
and ( n20086 , n19858 , n20085 );
and ( n20087 , n19585 , n20085 );
or ( n20088 , n19859 , n20086 , n20087 );
or ( n20089 , n19583 , n20088 );
or ( n20090 , n19581 , n20089 );
or ( n20091 , n19579 , n20090 );
or ( n20092 , n19577 , n20091 );
or ( n20093 , n19575 , n20092 );
or ( n20094 , n19573 , n20093 );
or ( n20095 , n19571 , n20094 );
or ( n20096 , n19569 , n20095 );
and ( n20097 , n19566 , n20096 );
and ( n20098 , n18437 , n20096 );
or ( n20099 , n19567 , n20097 , n20098 );
and ( n20100 , n18434 , n20099 );
and ( n20101 , n18209 , n20099 );
or ( n20102 , n18435 , n20100 , n20101 );
or ( n20103 , n18207 , n20102 );
or ( n20104 , n18205 , n20103 );
or ( n20105 , n18203 , n20104 );
or ( n20106 , n18201 , n20105 );
or ( n20107 , n18199 , n20106 );
or ( n20108 , n18197 , n20107 );
or ( n20109 , n18195 , n20108 );
or ( n20110 , n18193 , n20109 );
or ( n20111 , n18191 , n20110 );
or ( n20112 , n18189 , n20111 );
xnor ( n20113 , n18187 , n20112 );
xnor ( n20114 , n18189 , n20111 );
xnor ( n20115 , n18191 , n20110 );
xnor ( n20116 , n18193 , n20109 );
xnor ( n20117 , n18195 , n20108 );
xnor ( n20118 , n18197 , n20107 );
xnor ( n20119 , n18199 , n20106 );
xnor ( n20120 , n18201 , n20105 );
xnor ( n20121 , n18203 , n20104 );
xnor ( n20122 , n18205 , n20103 );
xnor ( n20123 , n18207 , n20102 );
xor ( n20124 , n18209 , n18434 );
xor ( n20125 , n20124 , n20099 );
not ( n20126 , n20125 );
xor ( n20127 , n18437 , n19566 );
xor ( n20128 , n20127 , n20096 );
xnor ( n20129 , n19569 , n20095 );
xnor ( n20130 , n19571 , n20094 );
xnor ( n20131 , n19573 , n20093 );
xnor ( n20132 , n19575 , n20092 );
xnor ( n20133 , n19577 , n20091 );
xnor ( n20134 , n19579 , n20090 );
xnor ( n20135 , n19581 , n20089 );
xnor ( n20136 , n19583 , n20088 );
xor ( n20137 , n19585 , n19858 );
xor ( n20138 , n20137 , n20085 );
xnor ( n20139 , n19861 , n20084 );
xor ( n20140 , n19863 , n20051 );
xor ( n20141 , n20140 , n20081 );
xnor ( n20142 , n20054 , n20080 );
xnor ( n20143 , n20056 , n20079 );
xnor ( n20144 , n20058 , n20078 );
xnor ( n20145 , n20060 , n20077 );
xor ( n20146 , n20062 , n20064 );
xor ( n20147 , n20146 , n20074 );
not ( n20148 , n20147 );
xor ( n20149 , n20067 , n20069 );
xor ( n20150 , n20149 , n20071 );
and ( n20151 , n8500 , n10627 );
and ( n20152 , n20150 , n20151 );
and ( n20153 , n20148 , n20152 );
or ( n20154 , n20147 , n20153 );
and ( n20155 , n20145 , n20154 );
and ( n20156 , n20144 , n20155 );
and ( n20157 , n20143 , n20156 );
and ( n20158 , n20142 , n20157 );
and ( n20159 , n20141 , n20158 );
and ( n20160 , n20139 , n20159 );
and ( n20161 , n20138 , n20160 );
and ( n20162 , n20136 , n20161 );
and ( n20163 , n20135 , n20162 );
and ( n20164 , n20134 , n20163 );
and ( n20165 , n20133 , n20164 );
and ( n20166 , n20132 , n20165 );
and ( n20167 , n20131 , n20166 );
and ( n20168 , n20130 , n20167 );
and ( n20169 , n20129 , n20168 );
and ( n20170 , n20128 , n20169 );
and ( n20171 , n20126 , n20170 );
or ( n20172 , n20125 , n20171 );
and ( n20173 , n20123 , n20172 );
and ( n20174 , n20122 , n20173 );
and ( n20175 , n20121 , n20174 );
and ( n20176 , n20120 , n20175 );
and ( n20177 , n20119 , n20176 );
and ( n20178 , n20118 , n20177 );
and ( n20179 , n20117 , n20178 );
and ( n20180 , n20116 , n20179 );
and ( n20181 , n20115 , n20180 );
and ( n20182 , n20114 , n20181 );
xor ( n20183 , n20113 , n20182 );
buf ( n20184 , n20183 );
buf ( n20185 , n20184 );
xor ( n20186 , n20114 , n20181 );
buf ( n20187 , n20186 );
buf ( n20188 , n20187 );
xor ( n20189 , n20115 , n20180 );
buf ( n20190 , n20189 );
buf ( n20191 , n20190 );
xor ( n20192 , n20116 , n20179 );
buf ( n20193 , n20192 );
buf ( n20194 , n20193 );
xor ( n20195 , n20117 , n20178 );
buf ( n20196 , n20195 );
buf ( n20197 , n20196 );
xor ( n20198 , n20118 , n20177 );
buf ( n20199 , n20198 );
buf ( n20200 , n20199 );
xor ( n20201 , n20119 , n20176 );
buf ( n20202 , n20201 );
buf ( n20203 , n20202 );
xor ( n20204 , n20120 , n20175 );
buf ( n20205 , n20204 );
buf ( n20206 , n20205 );
xor ( n20207 , n20121 , n20174 );
buf ( n20208 , n20207 );
buf ( n20209 , n20208 );
xor ( n20210 , n20122 , n20173 );
buf ( n20211 , n20210 );
buf ( n20212 , n20211 );
xor ( n20213 , n20123 , n20172 );
buf ( n20214 , n20213 );
buf ( n20215 , n20214 );
xor ( n20216 , n20126 , n20170 );
buf ( n20217 , n20216 );
buf ( n20218 , n20217 );
xor ( n20219 , n20128 , n20169 );
buf ( n20220 , n20219 );
buf ( n20221 , n20220 );
xor ( n20222 , n20129 , n20168 );
buf ( n20223 , n20222 );
buf ( n20224 , n20223 );
xor ( n20225 , n20130 , n20167 );
buf ( n20226 , n20225 );
buf ( n20227 , n20226 );
xor ( n20228 , n20131 , n20166 );
buf ( n20229 , n20228 );
buf ( n20230 , n20229 );
xor ( n20231 , n20132 , n20165 );
buf ( n20232 , n20231 );
buf ( n20233 , n20232 );
xor ( n20234 , n20133 , n20164 );
buf ( n20235 , n20234 );
buf ( n20236 , n20235 );
xor ( n20237 , n20134 , n20163 );
buf ( n20238 , n20237 );
buf ( n20239 , n20238 );
xor ( n20240 , n20135 , n20162 );
buf ( n20241 , n20240 );
buf ( n20242 , n20241 );
xor ( n20243 , n20136 , n20161 );
buf ( n20244 , n20243 );
buf ( n20245 , n20244 );
xor ( n20246 , n20138 , n20160 );
buf ( n20247 , n20246 );
buf ( n20248 , n20247 );
buf ( n20249 , n1103 );
and ( n20250 , n20248 , n20249 );
xor ( n20251 , n20139 , n20159 );
buf ( n20252 , n20251 );
buf ( n20253 , n20252 );
buf ( n20254 , n1273 );
and ( n20255 , n20253 , n20254 );
xor ( n20256 , n20141 , n20158 );
buf ( n20257 , n20256 );
buf ( n20258 , n20257 );
buf ( n20259 , n1310 );
and ( n20260 , n20258 , n20259 );
xor ( n20261 , n20142 , n20157 );
buf ( n20262 , n20261 );
buf ( n20263 , n20262 );
buf ( n20264 , n1346 );
and ( n20265 , n20263 , n20264 );
xor ( n20266 , n20143 , n20156 );
buf ( n20267 , n20266 );
buf ( n20268 , n20267 );
xor ( n20269 , n20144 , n20155 );
buf ( n20270 , n20269 );
buf ( n20271 , n20270 );
xor ( n20272 , n20145 , n20154 );
buf ( n20273 , n20272 );
buf ( n20274 , n20273 );
xor ( n20275 , n20148 , n20152 );
buf ( n20276 , n20275 );
buf ( n20277 , n20276 );
xor ( n20278 , n20150 , n20151 );
buf ( n20279 , n20278 );
buf ( n20280 , n20279 );
buf ( n20281 , n1687 );
and ( n20282 , n20280 , n20281 );
buf ( n20283 , n10629 );
buf ( n20284 , n1717 );
and ( n20285 , n20283 , n20284 );
buf ( n20286 , n10921 );
buf ( n20287 , n1776 );
and ( n20288 , n20286 , n20287 );
buf ( n20289 , n11378 );
buf ( n20290 , n1904 );
and ( n20291 , n20289 , n20290 );
buf ( n20292 , n11708 );
buf ( n20293 , n1988 );
and ( n20294 , n20292 , n20293 );
buf ( n20295 , n11835 );
buf ( n20296 , n2046 );
and ( n20297 , n20295 , n20296 );
buf ( n20298 , n12120 );
buf ( n20299 , n2248 );
and ( n20300 , n20298 , n20299 );
buf ( n20301 , n12619 );
buf ( n20302 , n2302 );
and ( n20303 , n20301 , n20302 );
buf ( n20304 , n12668 );
buf ( n20305 , n2490 );
and ( n20306 , n20304 , n20305 );
buf ( n20307 , n12963 );
buf ( n20308 , n2584 );
and ( n20309 , n20307 , n20308 );
buf ( n20310 , n13411 );
buf ( n20311 , n2716 );
and ( n20312 , n20310 , n20311 );
buf ( n20313 , n13689 );
buf ( n20314 , n2921 );
and ( n20315 , n20313 , n20314 );
buf ( n20316 , n13781 );
buf ( n20317 , n3144 );
and ( n20318 , n20316 , n20317 );
buf ( n20319 , n14265 );
buf ( n20320 , n3286 );
and ( n20321 , n20319 , n20320 );
buf ( n20322 , n14507 );
buf ( n20323 , n3447 );
and ( n20324 , n20322 , n20323 );
buf ( n20325 , n14700 );
buf ( n20326 , n3726 );
and ( n20327 , n20325 , n20326 );
buf ( n20328 , n14989 );
buf ( n20329 , n3890 );
and ( n20330 , n20328 , n20329 );
buf ( n20331 , n15019 );
buf ( n20332 , n4148 );
and ( n20333 , n20331 , n20332 );
buf ( n20334 , n15236 );
buf ( n20335 , n4360 );
and ( n20336 , n20334 , n20335 );
buf ( n20337 , n15630 );
buf ( n20338 , n4732 );
and ( n20339 , n20337 , n20338 );
buf ( n20340 , n15810 );
buf ( n20341 , n4980 );
and ( n20342 , n20340 , n20341 );
buf ( n20343 , n15972 );
buf ( n20344 , n5084 );
and ( n20345 , n20343 , n20344 );
buf ( n20346 , n16248 );
buf ( n20347 , n7637 );
and ( n20348 , n20346 , n20347 );
buf ( n20349 , n16310 );
buf ( n20350 , n5338 );
and ( n20351 , n20349 , n20350 );
and ( n20352 , n20347 , n20351 );
and ( n20353 , n20346 , n20351 );
or ( n20354 , n20348 , n20352 , n20353 );
and ( n20355 , n20344 , n20354 );
and ( n20356 , n20343 , n20354 );
or ( n20357 , n20345 , n20355 , n20356 );
and ( n20358 , n20341 , n20357 );
and ( n20359 , n20340 , n20357 );
or ( n20360 , n20342 , n20358 , n20359 );
and ( n20361 , n20338 , n20360 );
and ( n20362 , n20337 , n20360 );
or ( n20363 , n20339 , n20361 , n20362 );
and ( n20364 , n20335 , n20363 );
and ( n20365 , n20334 , n20363 );
or ( n20366 , n20336 , n20364 , n20365 );
and ( n20367 , n20332 , n20366 );
and ( n20368 , n20331 , n20366 );
or ( n20369 , n20333 , n20367 , n20368 );
and ( n20370 , n20329 , n20369 );
and ( n20371 , n20328 , n20369 );
or ( n20372 , n20330 , n20370 , n20371 );
and ( n20373 , n20326 , n20372 );
and ( n20374 , n20325 , n20372 );
or ( n20375 , n20327 , n20373 , n20374 );
and ( n20376 , n20323 , n20375 );
and ( n20377 , n20322 , n20375 );
or ( n20378 , n20324 , n20376 , n20377 );
and ( n20379 , n20320 , n20378 );
and ( n20380 , n20319 , n20378 );
or ( n20381 , n20321 , n20379 , n20380 );
and ( n20382 , n20317 , n20381 );
and ( n20383 , n20316 , n20381 );
or ( n20384 , n20318 , n20382 , n20383 );
and ( n20385 , n20314 , n20384 );
and ( n20386 , n20313 , n20384 );
or ( n20387 , n20315 , n20385 , n20386 );
and ( n20388 , n20311 , n20387 );
and ( n20389 , n20310 , n20387 );
or ( n20390 , n20312 , n20388 , n20389 );
and ( n20391 , n20308 , n20390 );
and ( n20392 , n20307 , n20390 );
or ( n20393 , n20309 , n20391 , n20392 );
and ( n20394 , n20305 , n20393 );
and ( n20395 , n20304 , n20393 );
or ( n20396 , n20306 , n20394 , n20395 );
and ( n20397 , n20302 , n20396 );
and ( n20398 , n20301 , n20396 );
or ( n20399 , n20303 , n20397 , n20398 );
and ( n20400 , n20299 , n20399 );
and ( n20401 , n20298 , n20399 );
or ( n20402 , n20300 , n20400 , n20401 );
and ( n20403 , n20296 , n20402 );
and ( n20404 , n20295 , n20402 );
or ( n20405 , n20297 , n20403 , n20404 );
and ( n20406 , n20293 , n20405 );
and ( n20407 , n20292 , n20405 );
or ( n20408 , n20294 , n20406 , n20407 );
and ( n20409 , n20290 , n20408 );
and ( n20410 , n20289 , n20408 );
or ( n20411 , n20291 , n20409 , n20410 );
and ( n20412 , n20287 , n20411 );
and ( n20413 , n20286 , n20411 );
or ( n20414 , n20288 , n20412 , n20413 );
and ( n20415 , n20284 , n20414 );
and ( n20416 , n20283 , n20414 );
or ( n20417 , n20285 , n20415 , n20416 );
and ( n20418 , n20281 , n20417 );
and ( n20419 , n20280 , n20417 );
or ( n20420 , n20282 , n20418 , n20419 );
and ( n20421 , n20277 , n20420 );
buf ( n20422 , n20421 );
and ( n20423 , n20274 , n20422 );
buf ( n20424 , n20423 );
and ( n20425 , n20271 , n20424 );
buf ( n20426 , n20425 );
and ( n20427 , n20268 , n20426 );
buf ( n20428 , n20427 );
and ( n20429 , n20264 , n20428 );
and ( n20430 , n20263 , n20428 );
or ( n20431 , n20265 , n20429 , n20430 );
and ( n20432 , n20259 , n20431 );
and ( n20433 , n20258 , n20431 );
or ( n20434 , n20260 , n20432 , n20433 );
and ( n20435 , n20254 , n20434 );
and ( n20436 , n20253 , n20434 );
or ( n20437 , n20255 , n20435 , n20436 );
and ( n20438 , n20249 , n20437 );
and ( n20439 , n20248 , n20437 );
or ( n20440 , n20250 , n20438 , n20439 );
and ( n20441 , n20245 , n20440 );
and ( n20442 , n20242 , n20441 );
and ( n20443 , n20239 , n20442 );
and ( n20444 , n20236 , n20443 );
and ( n20445 , n20233 , n20444 );
and ( n20446 , n20230 , n20445 );
and ( n20447 , n20227 , n20446 );
and ( n20448 , n20224 , n20447 );
and ( n20449 , n20221 , n20448 );
and ( n20450 , n20218 , n20449 );
and ( n20451 , n20215 , n20450 );
and ( n20452 , n20212 , n20451 );
and ( n20453 , n20209 , n20452 );
and ( n20454 , n20206 , n20453 );
and ( n20455 , n20203 , n20454 );
and ( n20456 , n20200 , n20455 );
and ( n20457 , n20197 , n20456 );
and ( n20458 , n20194 , n20457 );
and ( n20459 , n20191 , n20458 );
and ( n20460 , n20188 , n20459 );
and ( n20461 , n20185 , n20460 );
buf ( n20462 , n20461 );
buf ( n20463 , n20462 );
xor ( n20464 , n20185 , n20460 );
buf ( n20465 , n20464 );
buf ( n20466 , n20465 );
xor ( n20467 , n20188 , n20459 );
buf ( n20468 , n20467 );
buf ( n20469 , n20468 );
xor ( n20470 , n20191 , n20458 );
buf ( n20471 , n20470 );
buf ( n20472 , n20471 );
xor ( n20473 , n20194 , n20457 );
buf ( n20474 , n20473 );
buf ( n20475 , n20474 );
xor ( n20476 , n20197 , n20456 );
buf ( n20477 , n20476 );
buf ( n20478 , n20477 );
xor ( n20479 , n20200 , n20455 );
buf ( n20480 , n20479 );
buf ( n20481 , n20480 );
xor ( n20482 , n20203 , n20454 );
buf ( n20483 , n20482 );
buf ( n20484 , n20483 );
xor ( n20485 , n20206 , n20453 );
buf ( n20486 , n20485 );
buf ( n20487 , n20486 );
xor ( n20488 , n20209 , n20452 );
buf ( n20489 , n20488 );
buf ( n20490 , n20489 );
xor ( n20491 , n20212 , n20451 );
buf ( n20492 , n20491 );
buf ( n20493 , n20492 );
xor ( n20494 , n20215 , n20450 );
buf ( n20495 , n20494 );
buf ( n20496 , n20495 );
xor ( n20497 , n20218 , n20449 );
buf ( n20498 , n20497 );
buf ( n20499 , n20498 );
xor ( n20500 , n20221 , n20448 );
buf ( n20501 , n20500 );
buf ( n20502 , n20501 );
xor ( n20503 , n20224 , n20447 );
buf ( n20504 , n20503 );
buf ( n20505 , n20504 );
xor ( n20506 , n20227 , n20446 );
buf ( n20507 , n20506 );
buf ( n20508 , n20507 );
xor ( n20509 , n20230 , n20445 );
buf ( n20510 , n20509 );
buf ( n20511 , n20510 );
xor ( n20512 , n20233 , n20444 );
buf ( n20513 , n20512 );
buf ( n20514 , n20513 );
xor ( n20515 , n20236 , n20443 );
buf ( n20516 , n20515 );
buf ( n20517 , n20516 );
xor ( n20518 , n20239 , n20442 );
buf ( n20519 , n20518 );
buf ( n20520 , n20519 );
xor ( n20521 , n20242 , n20441 );
buf ( n20522 , n20521 );
buf ( n20523 , n20522 );
xor ( n20524 , n20245 , n20440 );
buf ( n20525 , n20524 );
buf ( n20526 , n20525 );
xor ( n20527 , n20248 , n20249 );
xor ( n20528 , n20527 , n20437 );
buf ( n20529 , n20528 );
buf ( n20530 , n20529 );
xor ( n20531 , n20253 , n20254 );
xor ( n20532 , n20531 , n20434 );
buf ( n20533 , n20532 );
buf ( n20534 , n20533 );
xor ( n20535 , n20258 , n20259 );
xor ( n20536 , n20535 , n20431 );
buf ( n20537 , n20536 );
buf ( n20538 , n20537 );
xor ( n20539 , n20263 , n20264 );
xor ( n20540 , n20539 , n20428 );
buf ( n20541 , n20540 );
buf ( n20542 , n20541 );
buf ( n20543 , n20268 );
xor ( n20544 , n20543 , n20426 );
buf ( n20545 , n20544 );
buf ( n20546 , n20545 );
buf ( n20547 , n20271 );
xor ( n20548 , n20547 , n20424 );
buf ( n20549 , n20548 );
buf ( n20550 , n20549 );
buf ( n20551 , n20274 );
xor ( n20552 , n20551 , n20422 );
buf ( n20553 , n20552 );
buf ( n20554 , n20553 );
buf ( n20555 , n20277 );
xor ( n20556 , n20555 , n20420 );
buf ( n20557 , n20556 );
buf ( n20558 , n20557 );
xor ( n20559 , n20280 , n20281 );
xor ( n20560 , n20559 , n20417 );
buf ( n20561 , n20560 );
buf ( n20562 , n20561 );
xor ( n20563 , n20283 , n20284 );
xor ( n20564 , n20563 , n20414 );
buf ( n20565 , n20564 );
buf ( n20566 , n20565 );
xor ( n20567 , n20286 , n20287 );
xor ( n20568 , n20567 , n20411 );
buf ( n20569 , n20568 );
buf ( n20570 , n20569 );
xor ( n20571 , n20289 , n20290 );
xor ( n20572 , n20571 , n20408 );
buf ( n20573 , n20572 );
buf ( n20574 , n20573 );
xor ( n20575 , n20292 , n20293 );
xor ( n20576 , n20575 , n20405 );
buf ( n20577 , n20576 );
buf ( n20578 , n20577 );
xor ( n20579 , n20295 , n20296 );
xor ( n20580 , n20579 , n20402 );
buf ( n20581 , n20580 );
buf ( n20582 , n20581 );
xor ( n20583 , n20298 , n20299 );
xor ( n20584 , n20583 , n20399 );
buf ( n20585 , n20584 );
buf ( n20586 , n20585 );
xor ( n20587 , n20301 , n20302 );
xor ( n20588 , n20587 , n20396 );
buf ( n20589 , n20588 );
buf ( n20590 , n20589 );
xor ( n20591 , n20304 , n20305 );
xor ( n20592 , n20591 , n20393 );
buf ( n20593 , n20592 );
buf ( n20594 , n20593 );
xor ( n20595 , n20307 , n20308 );
xor ( n20596 , n20595 , n20390 );
buf ( n20597 , n20596 );
buf ( n20598 , n20597 );
xor ( n20599 , n20310 , n20311 );
xor ( n20600 , n20599 , n20387 );
buf ( n20601 , n20600 );
buf ( n20602 , n20601 );
xor ( n20603 , n20313 , n20314 );
xor ( n20604 , n20603 , n20384 );
buf ( n20605 , n20604 );
buf ( n20606 , n20605 );
xor ( n20607 , n20316 , n20317 );
xor ( n20608 , n20607 , n20381 );
buf ( n20609 , n20608 );
buf ( n20610 , n20609 );
xor ( n20611 , n20319 , n20320 );
xor ( n20612 , n20611 , n20378 );
buf ( n20613 , n20612 );
buf ( n20614 , n20613 );
xor ( n20615 , n20322 , n20323 );
xor ( n20616 , n20615 , n20375 );
buf ( n20617 , n20616 );
buf ( n20618 , n20617 );
xor ( n20619 , n20325 , n20326 );
xor ( n20620 , n20619 , n20372 );
buf ( n20621 , n20620 );
buf ( n20622 , n20621 );
xor ( n20623 , n20328 , n20329 );
xor ( n20624 , n20623 , n20369 );
buf ( n20625 , n20624 );
buf ( n20626 , n20625 );
xor ( n20627 , n20331 , n20332 );
xor ( n20628 , n20627 , n20366 );
buf ( n20629 , n20628 );
buf ( n20630 , n20629 );
xor ( n20631 , n20334 , n20335 );
xor ( n20632 , n20631 , n20363 );
buf ( n20633 , n20632 );
buf ( n20634 , n20633 );
xor ( n20635 , n20337 , n20338 );
xor ( n20636 , n20635 , n20360 );
buf ( n20637 , n20636 );
buf ( n20638 , n20637 );
xor ( n20639 , n20340 , n20341 );
xor ( n20640 , n20639 , n20357 );
buf ( n20641 , n20640 );
buf ( n20642 , n20641 );
xor ( n20643 , n20343 , n20344 );
xor ( n20644 , n20643 , n20354 );
buf ( n20645 , n20644 );
buf ( n20646 , n20645 );
xor ( n20647 , n20346 , n20347 );
xor ( n20648 , n20647 , n20351 );
buf ( n20649 , n20648 );
buf ( n20650 , n20649 );
xor ( n20651 , n20349 , n20350 );
buf ( n20652 , n20651 );
buf ( n20653 , n20652 );
and ( n20654 , n20650 , n20653 );
or ( n20655 , n20646 , n20654 );
and ( n20656 , n20642 , n20655 );
and ( n20657 , n20638 , n20656 );
and ( n20658 , n20634 , n20657 );
and ( n20659 , n20630 , n20658 );
or ( n20660 , n20626 , n20659 );
or ( n20661 , n20622 , n20660 );
or ( n20662 , n20618 , n20661 );
or ( n20663 , n20614 , n20662 );
or ( n20664 , n20610 , n20663 );
or ( n20665 , n20606 , n20664 );
or ( n20666 , n20602 , n20665 );
or ( n20667 , n20598 , n20666 );
or ( n20668 , n20594 , n20667 );
or ( n20669 , n20590 , n20668 );
or ( n20670 , n20586 , n20669 );
or ( n20671 , n20582 , n20670 );
or ( n20672 , n20578 , n20671 );
or ( n20673 , n20574 , n20672 );
or ( n20674 , n20570 , n20673 );
or ( n20675 , n20566 , n20674 );
or ( n20676 , n20562 , n20675 );
or ( n20677 , n20558 , n20676 );
or ( n20678 , n20554 , n20677 );
or ( n20679 , n20550 , n20678 );
or ( n20680 , n20546 , n20679 );
or ( n20681 , n20542 , n20680 );
or ( n20682 , n20538 , n20681 );
or ( n20683 , n20534 , n20682 );
or ( n20684 , n20530 , n20683 );
or ( n20685 , n20526 , n20684 );
or ( n20686 , n20523 , n20685 );
or ( n20687 , n20520 , n20686 );
or ( n20688 , n20517 , n20687 );
or ( n20689 , n20514 , n20688 );
or ( n20690 , n20511 , n20689 );
or ( n20691 , n20508 , n20690 );
or ( n20692 , n20505 , n20691 );
or ( n20693 , n20502 , n20692 );
or ( n20694 , n20499 , n20693 );
or ( n20695 , n20496 , n20694 );
or ( n20696 , n20493 , n20695 );
or ( n20697 , n20490 , n20696 );
or ( n20698 , n20487 , n20697 );
or ( n20699 , n20484 , n20698 );
or ( n20700 , n20481 , n20699 );
or ( n20701 , n20478 , n20700 );
or ( n20702 , n20475 , n20701 );
or ( n20703 , n20472 , n20702 );
or ( n20704 , n20469 , n20703 );
or ( n20705 , n20466 , n20704 );
or ( n20706 , n20463 , n20705 );
not ( n20707 , n20706 );
buf ( n20708 , n20707 );
xnor ( n20709 , n20463 , n20705 );
buf ( n20710 , n20709 );
xnor ( n20711 , n20466 , n20704 );
buf ( n20712 , n20711 );
xnor ( n20713 , n20469 , n20703 );
buf ( n20714 , n20713 );
xnor ( n20715 , n20472 , n20702 );
buf ( n20716 , n20715 );
xnor ( n20717 , n20475 , n20701 );
buf ( n20718 , n20717 );
xnor ( n20719 , n20478 , n20700 );
buf ( n20720 , n20719 );
xnor ( n20721 , n20481 , n20699 );
buf ( n20722 , n20721 );
xnor ( n20723 , n20484 , n20698 );
buf ( n20724 , n20723 );
xnor ( n20725 , n20487 , n20697 );
buf ( n20726 , n20725 );
xnor ( n20727 , n20490 , n20696 );
buf ( n20728 , n20727 );
xnor ( n20729 , n20493 , n20695 );
buf ( n20730 , n20729 );
xnor ( n20731 , n20496 , n20694 );
buf ( n20732 , n20731 );
xnor ( n20733 , n20499 , n20693 );
buf ( n20734 , n20733 );
xnor ( n20735 , n20502 , n20692 );
buf ( n20736 , n20735 );
xnor ( n20737 , n20505 , n20691 );
buf ( n20738 , n20737 );
xnor ( n20739 , n20508 , n20690 );
buf ( n20740 , n20739 );
xnor ( n20741 , n20511 , n20689 );
buf ( n20742 , n20741 );
xnor ( n20743 , n20514 , n20688 );
buf ( n20744 , n20743 );
xnor ( n20745 , n20517 , n20687 );
buf ( n20746 , n20745 );
xnor ( n20747 , n20520 , n20686 );
buf ( n20748 , n20747 );
xnor ( n20749 , n20523 , n20685 );
buf ( n20750 , n20749 );
xnor ( n20751 , n20526 , n20684 );
buf ( n20752 , n20751 );
xnor ( n20753 , n20530 , n20683 );
buf ( n20754 , n20753 );
xnor ( n20755 , n20534 , n20682 );
buf ( n20756 , n20755 );
xnor ( n20757 , n20538 , n20681 );
buf ( n20758 , n20757 );
xnor ( n20759 , n20542 , n20680 );
buf ( n20760 , n20759 );
xnor ( n20761 , n20546 , n20679 );
buf ( n20762 , n20761 );
xnor ( n20763 , n20550 , n20678 );
buf ( n20764 , n20763 );
xnor ( n20765 , n20554 , n20677 );
buf ( n20766 , n20765 );
xnor ( n20767 , n20558 , n20676 );
buf ( n20768 , n20767 );
xnor ( n20769 , n20562 , n20675 );
buf ( n20770 , n20769 );
xnor ( n20771 , n20566 , n20674 );
buf ( n20772 , n20771 );
xnor ( n20773 , n20570 , n20673 );
buf ( n20774 , n20773 );
xnor ( n20775 , n20574 , n20672 );
buf ( n20776 , n20775 );
xnor ( n20777 , n20578 , n20671 );
buf ( n20778 , n20777 );
xnor ( n20779 , n20582 , n20670 );
buf ( n20780 , n20779 );
xnor ( n20781 , n20586 , n20669 );
buf ( n20782 , n20781 );
xnor ( n20783 , n20590 , n20668 );
buf ( n20784 , n20783 );
xnor ( n20785 , n20594 , n20667 );
buf ( n20786 , n20785 );
xnor ( n20787 , n20598 , n20666 );
buf ( n20788 , n20787 );
xnor ( n20789 , n20602 , n20665 );
buf ( n20790 , n20789 );
xnor ( n20791 , n20606 , n20664 );
buf ( n20792 , n20791 );
xnor ( n20793 , n20610 , n20663 );
buf ( n20794 , n20793 );
xnor ( n20795 , n20614 , n20662 );
buf ( n20796 , n20795 );
xnor ( n20797 , n20618 , n20661 );
buf ( n20798 , n20797 );
xnor ( n20799 , n20622 , n20660 );
buf ( n20800 , n20799 );
xnor ( n20801 , n20626 , n20659 );
buf ( n20802 , n20801 );
xor ( n20803 , n20630 , n20658 );
buf ( n20804 , n20803 );
xor ( n20805 , n20634 , n20657 );
buf ( n20806 , n20805 );
xor ( n20807 , n20638 , n20656 );
buf ( n20808 , n20807 );
xor ( n20809 , n20642 , n20655 );
buf ( n20810 , n20809 );
xnor ( n20811 , n20646 , n20654 );
buf ( n20812 , n20811 );
xor ( n20813 , n20650 , n20653 );
buf ( n20814 , n20813 );
not ( n20815 , n20653 );
buf ( n20816 , n20815 );
buf ( n20817 , n794 );
buf ( n20818 , n795 );
buf ( n20819 , n796 );
buf ( n20820 , n797 );
buf ( n20821 , n798 );
buf ( n20822 , n799 );
buf ( n20823 , n800 );
buf ( n20824 , n801 );
buf ( n20825 , n802 );
buf ( n20826 , n803 );
buf ( n20827 , n804 );
buf ( n20828 , n805 );
buf ( n20829 , n806 );
buf ( n20830 , n807 );
buf ( n20831 , n808 );
buf ( n20832 , n809 );
buf ( n20833 , n17449 );
buf ( n20834 , n20833 );
buf ( n20835 , n17451 );
buf ( n20836 , n20835 );
buf ( n20837 , n17453 );
buf ( n20838 , n20837 );
and ( n20839 , n20836 , n20838 );
not ( n20840 , n20839 );
and ( n20841 , n20834 , n20840 );
not ( n20842 , n20841 );
buf ( n20843 , n20708 );
buf ( n20844 , n20843 );
buf ( n20845 , n17445 );
buf ( n20846 , n20845 );
buf ( n20847 , n17447 );
buf ( n20848 , n20847 );
xor ( n20849 , n20846 , n20848 );
xor ( n20850 , n20848 , n20834 );
not ( n20851 , n20850 );
and ( n20852 , n20849 , n20851 );
and ( n20853 , n20844 , n20852 );
buf ( n20854 , n20708 );
buf ( n20855 , n20854 );
and ( n20856 , n20855 , n20850 );
nor ( n20857 , n20853 , n20856 );
and ( n20858 , n20848 , n20834 );
not ( n20859 , n20858 );
and ( n20860 , n20846 , n20859 );
xnor ( n20861 , n20857 , n20860 );
and ( n20862 , n20842 , n20861 );
buf ( n20863 , n20708 );
buf ( n20864 , n20863 );
and ( n20865 , n20864 , n20846 );
and ( n20866 , n20861 , n20865 );
and ( n20867 , n20842 , n20865 );
or ( n20868 , n20862 , n20866 , n20867 );
and ( n20869 , n20855 , n20852 );
not ( n20870 , n20869 );
xnor ( n20871 , n20870 , n20860 );
and ( n20872 , n20844 , n20846 );
xor ( n20873 , n20871 , n20872 );
buf ( n20874 , n20187 );
buf ( n20875 , n20874 );
buf ( n20876 , n20184 );
buf ( n20877 , n20876 );
and ( n20878 , n20875 , n20877 );
buf ( n20879 , n20184 );
buf ( n20880 , n20879 );
buf ( n20881 , n20880 );
xor ( n20882 , n20878 , n20881 );
buf ( n20883 , n20190 );
buf ( n20884 , n20883 );
and ( n20885 , n20884 , n20877 );
buf ( n20886 , n20193 );
buf ( n20887 , n20886 );
and ( n20888 , n20887 , n20877 );
buf ( n20889 , n20187 );
buf ( n20890 , n20889 );
and ( n20891 , n20884 , n20890 );
and ( n20892 , n20888 , n20891 );
buf ( n20893 , n20875 );
and ( n20894 , n20891 , n20893 );
and ( n20895 , n20888 , n20893 );
or ( n20896 , n20892 , n20894 , n20895 );
and ( n20897 , n20885 , n20896 );
xor ( n20898 , n20888 , n20891 );
xor ( n20899 , n20898 , n20893 );
buf ( n20900 , n20196 );
buf ( n20901 , n20900 );
and ( n20902 , n20901 , n20877 );
and ( n20903 , n20887 , n20890 );
and ( n20904 , n20902 , n20903 );
buf ( n20905 , n20199 );
buf ( n20906 , n20905 );
and ( n20907 , n20906 , n20877 );
buf ( n20908 , n20190 );
buf ( n20909 , n20908 );
and ( n20910 , n20887 , n20909 );
and ( n20911 , n20907 , n20910 );
buf ( n20912 , n20884 );
and ( n20913 , n20910 , n20912 );
and ( n20914 , n20907 , n20912 );
or ( n20915 , n20911 , n20913 , n20914 );
and ( n20916 , n20903 , n20915 );
and ( n20917 , n20902 , n20915 );
or ( n20918 , n20904 , n20916 , n20917 );
and ( n20919 , n20899 , n20918 );
xor ( n20920 , n20902 , n20903 );
xor ( n20921 , n20920 , n20915 );
buf ( n20922 , n20202 );
buf ( n20923 , n20922 );
and ( n20924 , n20923 , n20877 );
and ( n20925 , n20906 , n20890 );
and ( n20926 , n20924 , n20925 );
and ( n20927 , n20901 , n20909 );
and ( n20928 , n20925 , n20927 );
and ( n20929 , n20924 , n20927 );
or ( n20930 , n20926 , n20928 , n20929 );
buf ( n20931 , n20887 );
buf ( n20932 , n20931 );
buf ( n20933 , n20932 );
and ( n20934 , n20930 , n20933 );
and ( n20935 , n20901 , n20890 );
and ( n20936 , n20933 , n20935 );
and ( n20937 , n20930 , n20935 );
or ( n20938 , n20934 , n20936 , n20937 );
and ( n20939 , n20921 , n20938 );
xor ( n20940 , n20907 , n20910 );
xor ( n20941 , n20940 , n20912 );
buf ( n20942 , n20205 );
buf ( n20943 , n20942 );
and ( n20944 , n20943 , n20890 );
buf ( n20945 , n20944 );
and ( n20946 , n20906 , n20909 );
and ( n20947 , n20945 , n20946 );
buf ( n20948 , n20193 );
buf ( n20949 , n20948 );
and ( n20950 , n20901 , n20949 );
and ( n20951 , n20946 , n20950 );
and ( n20952 , n20945 , n20950 );
or ( n20953 , n20947 , n20951 , n20952 );
and ( n20954 , n20943 , n20877 );
and ( n20955 , n20923 , n20890 );
and ( n20956 , n20954 , n20955 );
not ( n20957 , n20931 );
and ( n20958 , n20955 , n20957 );
and ( n20959 , n20954 , n20957 );
or ( n20960 , n20956 , n20958 , n20959 );
and ( n20961 , n20953 , n20960 );
not ( n20962 , n20932 );
and ( n20963 , n20960 , n20962 );
and ( n20964 , n20953 , n20962 );
or ( n20965 , n20961 , n20963 , n20964 );
and ( n20966 , n20941 , n20965 );
xor ( n20967 , n20930 , n20933 );
xor ( n20968 , n20967 , n20935 );
and ( n20969 , n20965 , n20968 );
and ( n20970 , n20941 , n20968 );
or ( n20971 , n20966 , n20969 , n20970 );
and ( n20972 , n20938 , n20971 );
and ( n20973 , n20921 , n20971 );
or ( n20974 , n20939 , n20972 , n20973 );
and ( n20975 , n20918 , n20974 );
and ( n20976 , n20899 , n20974 );
or ( n20977 , n20919 , n20975 , n20976 );
and ( n20978 , n20896 , n20977 );
and ( n20979 , n20885 , n20977 );
or ( n20980 , n20897 , n20978 , n20979 );
xor ( n20981 , n20882 , n20980 );
xor ( n20982 , n20885 , n20896 );
xor ( n20983 , n20982 , n20977 );
xor ( n20984 , n20899 , n20918 );
xor ( n20985 , n20984 , n20974 );
xor ( n20986 , n20921 , n20938 );
xor ( n20987 , n20986 , n20971 );
buf ( n20988 , n20208 );
buf ( n20989 , n20988 );
and ( n20990 , n20989 , n20877 );
and ( n20991 , n20923 , n20909 );
and ( n20992 , n20990 , n20991 );
and ( n20993 , n20906 , n20949 );
and ( n20994 , n20991 , n20993 );
and ( n20995 , n20990 , n20993 );
or ( n20996 , n20992 , n20994 , n20995 );
xor ( n20997 , n20945 , n20946 );
xor ( n20998 , n20997 , n20950 );
and ( n20999 , n20996 , n20998 );
xor ( n21000 , n20954 , n20955 );
xor ( n21001 , n21000 , n20957 );
and ( n21002 , n20998 , n21001 );
and ( n21003 , n20996 , n21001 );
or ( n21004 , n20999 , n21002 , n21003 );
xor ( n21005 , n20924 , n20925 );
xor ( n21006 , n21005 , n20927 );
and ( n21007 , n21004 , n21006 );
xor ( n21008 , n20953 , n20960 );
xor ( n21009 , n21008 , n20962 );
and ( n21010 , n21006 , n21009 );
and ( n21011 , n21004 , n21009 );
or ( n21012 , n21007 , n21010 , n21011 );
xor ( n21013 , n20941 , n20965 );
xor ( n21014 , n21013 , n20968 );
and ( n21015 , n21012 , n21014 );
xor ( n21016 , n21004 , n21006 );
xor ( n21017 , n21016 , n21009 );
buf ( n21018 , n20211 );
buf ( n21019 , n21018 );
and ( n21020 , n21019 , n20877 );
and ( n21021 , n20923 , n20949 );
and ( n21022 , n21020 , n21021 );
buf ( n21023 , n20901 );
and ( n21024 , n21021 , n21023 );
and ( n21025 , n21020 , n21023 );
or ( n21026 , n21022 , n21024 , n21025 );
and ( n21027 , n20943 , n20909 );
buf ( n21028 , n21027 );
and ( n21029 , n21026 , n21028 );
not ( n21030 , n20944 );
and ( n21031 , n21028 , n21030 );
and ( n21032 , n21026 , n21030 );
or ( n21033 , n21029 , n21031 , n21032 );
and ( n21034 , n20943 , n20949 );
buf ( n21035 , n21034 );
and ( n21036 , n20989 , n20890 );
and ( n21037 , n21035 , n21036 );
buf ( n21038 , n20196 );
buf ( n21039 , n21038 );
and ( n21040 , n20906 , n21039 );
and ( n21041 , n21036 , n21040 );
and ( n21042 , n21035 , n21040 );
or ( n21043 , n21037 , n21041 , n21042 );
xor ( n21044 , n20990 , n20991 );
xor ( n21045 , n21044 , n20993 );
and ( n21046 , n21043 , n21045 );
xor ( n21047 , n21026 , n21028 );
xor ( n21048 , n21047 , n21030 );
and ( n21049 , n21045 , n21048 );
and ( n21050 , n21043 , n21048 );
or ( n21051 , n21046 , n21049 , n21050 );
and ( n21052 , n21033 , n21051 );
xor ( n21053 , n20996 , n20998 );
xor ( n21054 , n21053 , n21001 );
and ( n21055 , n21051 , n21054 );
and ( n21056 , n21033 , n21054 );
or ( n21057 , n21052 , n21055 , n21056 );
and ( n21058 , n21017 , n21057 );
buf ( n21059 , n20214 );
buf ( n21060 , n21059 );
and ( n21061 , n21060 , n20877 );
and ( n21062 , n21019 , n20890 );
and ( n21063 , n21061 , n21062 );
and ( n21064 , n20923 , n21039 );
and ( n21065 , n21062 , n21064 );
and ( n21066 , n21061 , n21064 );
or ( n21067 , n21063 , n21065 , n21066 );
buf ( n21068 , n20906 );
buf ( n21069 , n21068 );
and ( n21070 , n20989 , n20909 );
and ( n21071 , n21069 , n21070 );
not ( n21072 , n21034 );
and ( n21073 , n21070 , n21072 );
and ( n21074 , n21069 , n21072 );
or ( n21075 , n21071 , n21073 , n21074 );
and ( n21076 , n21067 , n21075 );
not ( n21077 , n21027 );
and ( n21078 , n21075 , n21077 );
and ( n21079 , n21067 , n21077 );
or ( n21080 , n21076 , n21078 , n21079 );
and ( n21081 , n21060 , n20890 );
and ( n21082 , n21019 , n20909 );
and ( n21083 , n21081 , n21082 );
buf ( n21084 , n20199 );
buf ( n21085 , n21084 );
and ( n21086 , n20923 , n21085 );
and ( n21087 , n21082 , n21086 );
and ( n21088 , n21081 , n21086 );
or ( n21089 , n21083 , n21087 , n21088 );
buf ( n21090 , n20217 );
buf ( n21091 , n21090 );
and ( n21092 , n21091 , n20877 );
and ( n21093 , n20989 , n20949 );
and ( n21094 , n21092 , n21093 );
not ( n21095 , n21068 );
and ( n21096 , n21093 , n21095 );
and ( n21097 , n21092 , n21095 );
or ( n21098 , n21094 , n21096 , n21097 );
and ( n21099 , n21089 , n21098 );
xor ( n21100 , n21061 , n21062 );
xor ( n21101 , n21100 , n21064 );
and ( n21102 , n21098 , n21101 );
and ( n21103 , n21089 , n21101 );
or ( n21104 , n21099 , n21102 , n21103 );
xor ( n21105 , n21020 , n21021 );
xor ( n21106 , n21105 , n21023 );
and ( n21107 , n21104 , n21106 );
xor ( n21108 , n21035 , n21036 );
xor ( n21109 , n21108 , n21040 );
and ( n21110 , n21106 , n21109 );
and ( n21111 , n21104 , n21109 );
or ( n21112 , n21107 , n21110 , n21111 );
and ( n21113 , n21080 , n21112 );
xor ( n21114 , n21043 , n21045 );
xor ( n21115 , n21114 , n21048 );
and ( n21116 , n21112 , n21115 );
and ( n21117 , n21080 , n21115 );
or ( n21118 , n21113 , n21116 , n21117 );
xor ( n21119 , n21033 , n21051 );
xor ( n21120 , n21119 , n21054 );
and ( n21121 , n21118 , n21120 );
buf ( n21122 , n20220 );
buf ( n21123 , n21122 );
and ( n21124 , n21123 , n20877 );
and ( n21125 , n21060 , n20909 );
and ( n21126 , n21124 , n21125 );
and ( n21127 , n20943 , n21085 );
and ( n21128 , n21125 , n21127 );
and ( n21129 , n21124 , n21127 );
or ( n21130 , n21126 , n21128 , n21129 );
and ( n21131 , n21091 , n20890 );
buf ( n21132 , n21131 );
and ( n21133 , n21130 , n21132 );
and ( n21134 , n20943 , n21039 );
and ( n21135 , n21132 , n21134 );
and ( n21136 , n21130 , n21134 );
or ( n21137 , n21133 , n21135 , n21136 );
not ( n21138 , n21131 );
and ( n21139 , n21019 , n20949 );
and ( n21140 , n21138 , n21139 );
and ( n21141 , n20989 , n21039 );
and ( n21142 , n21139 , n21141 );
and ( n21143 , n21138 , n21141 );
or ( n21144 , n21140 , n21142 , n21143 );
xor ( n21145 , n21081 , n21082 );
xor ( n21146 , n21145 , n21086 );
and ( n21147 , n21144 , n21146 );
xor ( n21148 , n21092 , n21093 );
xor ( n21149 , n21148 , n21095 );
and ( n21150 , n21146 , n21149 );
and ( n21151 , n21144 , n21149 );
or ( n21152 , n21147 , n21150 , n21151 );
and ( n21153 , n21137 , n21152 );
xor ( n21154 , n21069 , n21070 );
xor ( n21155 , n21154 , n21072 );
and ( n21156 , n21152 , n21155 );
and ( n21157 , n21137 , n21155 );
or ( n21158 , n21153 , n21156 , n21157 );
xor ( n21159 , n21067 , n21075 );
xor ( n21160 , n21159 , n21077 );
and ( n21161 , n21158 , n21160 );
xor ( n21162 , n21104 , n21106 );
xor ( n21163 , n21162 , n21109 );
and ( n21164 , n21160 , n21163 );
and ( n21165 , n21158 , n21163 );
or ( n21166 , n21161 , n21164 , n21165 );
xor ( n21167 , n21080 , n21112 );
xor ( n21168 , n21167 , n21115 );
and ( n21169 , n21166 , n21168 );
xor ( n21170 , n21158 , n21160 );
xor ( n21171 , n21170 , n21163 );
buf ( n21172 , n20223 );
buf ( n21173 , n21172 );
and ( n21174 , n21173 , n20877 );
and ( n21175 , n21091 , n20909 );
and ( n21176 , n21174 , n21175 );
buf ( n21177 , n20202 );
buf ( n21178 , n21177 );
and ( n21179 , n20943 , n21178 );
and ( n21180 , n21175 , n21179 );
and ( n21181 , n21174 , n21179 );
or ( n21182 , n21176 , n21180 , n21181 );
and ( n21183 , n21091 , n20949 );
buf ( n21184 , n21183 );
and ( n21185 , n21019 , n21039 );
and ( n21186 , n21184 , n21185 );
and ( n21187 , n20989 , n21085 );
and ( n21188 , n21185 , n21187 );
and ( n21189 , n21184 , n21187 );
or ( n21190 , n21186 , n21188 , n21189 );
and ( n21191 , n21182 , n21190 );
buf ( n21192 , n20923 );
buf ( n21193 , n21192 );
and ( n21194 , n21190 , n21193 );
and ( n21195 , n21182 , n21193 );
or ( n21196 , n21191 , n21194 , n21195 );
and ( n21197 , n21123 , n20890 );
and ( n21198 , n21060 , n20949 );
and ( n21199 , n21197 , n21198 );
not ( n21200 , n21192 );
and ( n21201 , n21198 , n21200 );
and ( n21202 , n21197 , n21200 );
or ( n21203 , n21199 , n21201 , n21202 );
xor ( n21204 , n21124 , n21125 );
xor ( n21205 , n21204 , n21127 );
and ( n21206 , n21203 , n21205 );
xor ( n21207 , n21138 , n21139 );
xor ( n21208 , n21207 , n21141 );
and ( n21209 , n21205 , n21208 );
and ( n21210 , n21203 , n21208 );
or ( n21211 , n21206 , n21209 , n21210 );
and ( n21212 , n21196 , n21211 );
xor ( n21213 , n21130 , n21132 );
xor ( n21214 , n21213 , n21134 );
and ( n21215 , n21211 , n21214 );
and ( n21216 , n21196 , n21214 );
or ( n21217 , n21212 , n21215 , n21216 );
xor ( n21218 , n21089 , n21098 );
xor ( n21219 , n21218 , n21101 );
and ( n21220 , n21217 , n21219 );
xor ( n21221 , n21137 , n21152 );
xor ( n21222 , n21221 , n21155 );
and ( n21223 , n21219 , n21222 );
and ( n21224 , n21217 , n21222 );
or ( n21225 , n21220 , n21223 , n21224 );
and ( n21226 , n21171 , n21225 );
xor ( n21227 , n21217 , n21219 );
xor ( n21228 , n21227 , n21222 );
buf ( n21229 , n20943 );
buf ( n21230 , n21229 );
and ( n21231 , n21173 , n20890 );
and ( n21232 , n21230 , n21231 );
and ( n21233 , n21019 , n21085 );
and ( n21234 , n21231 , n21233 );
and ( n21235 , n21230 , n21233 );
or ( n21236 , n21232 , n21234 , n21235 );
buf ( n21237 , n20226 );
buf ( n21238 , n21237 );
and ( n21239 , n21238 , n20877 );
and ( n21240 , n21123 , n20909 );
and ( n21241 , n21239 , n21240 );
not ( n21242 , n21183 );
and ( n21243 , n21240 , n21242 );
and ( n21244 , n21239 , n21242 );
or ( n21245 , n21241 , n21243 , n21244 );
and ( n21246 , n21236 , n21245 );
xor ( n21247 , n21197 , n21198 );
xor ( n21248 , n21247 , n21200 );
and ( n21249 , n21245 , n21248 );
and ( n21250 , n21236 , n21248 );
or ( n21251 , n21246 , n21249 , n21250 );
xor ( n21252 , n21182 , n21190 );
xor ( n21253 , n21252 , n21193 );
and ( n21254 , n21251 , n21253 );
xor ( n21255 , n21203 , n21205 );
xor ( n21256 , n21255 , n21208 );
and ( n21257 , n21253 , n21256 );
and ( n21258 , n21251 , n21256 );
or ( n21259 , n21254 , n21257 , n21258 );
xor ( n21260 , n21144 , n21146 );
xor ( n21261 , n21260 , n21149 );
and ( n21262 , n21259 , n21261 );
xor ( n21263 , n21196 , n21211 );
xor ( n21264 , n21263 , n21214 );
and ( n21265 , n21261 , n21264 );
and ( n21266 , n21259 , n21264 );
or ( n21267 , n21262 , n21265 , n21266 );
and ( n21268 , n21228 , n21267 );
xor ( n21269 , n21259 , n21261 );
xor ( n21270 , n21269 , n21264 );
and ( n21271 , n21238 , n20890 );
and ( n21272 , n21173 , n20909 );
and ( n21273 , n21271 , n21272 );
and ( n21274 , n21060 , n21085 );
and ( n21275 , n21272 , n21274 );
and ( n21276 , n21271 , n21274 );
or ( n21277 , n21273 , n21275 , n21276 );
and ( n21278 , n21060 , n21039 );
and ( n21279 , n21277 , n21278 );
and ( n21280 , n20989 , n21178 );
and ( n21281 , n21278 , n21280 );
and ( n21282 , n21277 , n21280 );
or ( n21283 , n21279 , n21281 , n21282 );
xor ( n21284 , n21174 , n21175 );
xor ( n21285 , n21284 , n21179 );
and ( n21286 , n21283 , n21285 );
xor ( n21287 , n21184 , n21185 );
xor ( n21288 , n21287 , n21187 );
and ( n21289 , n21285 , n21288 );
and ( n21290 , n21283 , n21288 );
or ( n21291 , n21286 , n21289 , n21290 );
and ( n21292 , n21091 , n21039 );
and ( n21293 , n21019 , n21178 );
and ( n21294 , n21292 , n21293 );
buf ( n21295 , n20205 );
buf ( n21296 , n21295 );
and ( n21297 , n20989 , n21296 );
and ( n21298 , n21293 , n21297 );
and ( n21299 , n21292 , n21297 );
or ( n21300 , n21294 , n21298 , n21299 );
buf ( n21301 , n20229 );
buf ( n21302 , n21301 );
and ( n21303 , n21302 , n20877 );
and ( n21304 , n21123 , n20949 );
and ( n21305 , n21303 , n21304 );
not ( n21306 , n21229 );
and ( n21307 , n21304 , n21306 );
and ( n21308 , n21303 , n21306 );
or ( n21309 , n21305 , n21307 , n21308 );
and ( n21310 , n21300 , n21309 );
xor ( n21311 , n21239 , n21240 );
xor ( n21312 , n21311 , n21242 );
and ( n21313 , n21309 , n21312 );
and ( n21314 , n21300 , n21312 );
or ( n21315 , n21310 , n21313 , n21314 );
and ( n21316 , n21302 , n20890 );
and ( n21317 , n21238 , n20909 );
and ( n21318 , n21316 , n21317 );
and ( n21319 , n21019 , n21296 );
and ( n21320 , n21317 , n21319 );
and ( n21321 , n21316 , n21319 );
or ( n21322 , n21318 , n21320 , n21321 );
and ( n21323 , n21173 , n20949 );
buf ( n21324 , n21323 );
and ( n21325 , n21322 , n21324 );
xor ( n21326 , n21271 , n21272 );
xor ( n21327 , n21326 , n21274 );
and ( n21328 , n21324 , n21327 );
and ( n21329 , n21322 , n21327 );
or ( n21330 , n21325 , n21328 , n21329 );
xor ( n21331 , n21230 , n21231 );
xor ( n21332 , n21331 , n21233 );
and ( n21333 , n21330 , n21332 );
xor ( n21334 , n21277 , n21278 );
xor ( n21335 , n21334 , n21280 );
and ( n21336 , n21332 , n21335 );
and ( n21337 , n21330 , n21335 );
or ( n21338 , n21333 , n21336 , n21337 );
and ( n21339 , n21315 , n21338 );
xor ( n21340 , n21236 , n21245 );
xor ( n21341 , n21340 , n21248 );
and ( n21342 , n21338 , n21341 );
and ( n21343 , n21315 , n21341 );
or ( n21344 , n21339 , n21342 , n21343 );
and ( n21345 , n21291 , n21344 );
xor ( n21346 , n21251 , n21253 );
xor ( n21347 , n21346 , n21256 );
and ( n21348 , n21344 , n21347 );
and ( n21349 , n21291 , n21347 );
or ( n21350 , n21345 , n21348 , n21349 );
and ( n21351 , n21270 , n21350 );
xor ( n21352 , n21291 , n21344 );
xor ( n21353 , n21352 , n21347 );
buf ( n21354 , n20232 );
buf ( n21355 , n21354 );
and ( n21356 , n21355 , n20877 );
and ( n21357 , n21091 , n21085 );
and ( n21358 , n21356 , n21357 );
and ( n21359 , n21060 , n21178 );
and ( n21360 , n21357 , n21359 );
and ( n21361 , n21356 , n21359 );
or ( n21362 , n21358 , n21360 , n21361 );
and ( n21363 , n21238 , n20949 );
buf ( n21364 , n21363 );
not ( n21365 , n21323 );
and ( n21366 , n21364 , n21365 );
and ( n21367 , n21123 , n21039 );
and ( n21368 , n21365 , n21367 );
and ( n21369 , n21364 , n21367 );
or ( n21370 , n21366 , n21368 , n21369 );
and ( n21371 , n21362 , n21370 );
xor ( n21372 , n21303 , n21304 );
xor ( n21373 , n21372 , n21306 );
and ( n21374 , n21370 , n21373 );
and ( n21375 , n21362 , n21373 );
or ( n21376 , n21371 , n21374 , n21375 );
and ( n21377 , n21355 , n20890 );
and ( n21378 , n21302 , n20909 );
and ( n21379 , n21377 , n21378 );
and ( n21380 , n21091 , n21178 );
and ( n21381 , n21378 , n21380 );
and ( n21382 , n21377 , n21380 );
or ( n21383 , n21379 , n21381 , n21382 );
buf ( n21384 , n20235 );
buf ( n21385 , n21384 );
and ( n21386 , n21385 , n20877 );
and ( n21387 , n21123 , n21085 );
and ( n21388 , n21386 , n21387 );
buf ( n21389 , n20989 );
and ( n21390 , n21387 , n21389 );
and ( n21391 , n21386 , n21389 );
or ( n21392 , n21388 , n21390 , n21391 );
and ( n21393 , n21383 , n21392 );
xor ( n21394 , n21316 , n21317 );
xor ( n21395 , n21394 , n21319 );
and ( n21396 , n21392 , n21395 );
and ( n21397 , n21383 , n21395 );
or ( n21398 , n21393 , n21396 , n21397 );
xor ( n21399 , n21292 , n21293 );
xor ( n21400 , n21399 , n21297 );
and ( n21401 , n21398 , n21400 );
xor ( n21402 , n21322 , n21324 );
xor ( n21403 , n21402 , n21327 );
and ( n21404 , n21400 , n21403 );
and ( n21405 , n21398 , n21403 );
or ( n21406 , n21401 , n21404 , n21405 );
and ( n21407 , n21376 , n21406 );
xor ( n21408 , n21300 , n21309 );
xor ( n21409 , n21408 , n21312 );
and ( n21410 , n21406 , n21409 );
and ( n21411 , n21376 , n21409 );
or ( n21412 , n21407 , n21410 , n21411 );
xor ( n21413 , n21283 , n21285 );
xor ( n21414 , n21413 , n21288 );
and ( n21415 , n21412 , n21414 );
xor ( n21416 , n21315 , n21338 );
xor ( n21417 , n21416 , n21341 );
and ( n21418 , n21414 , n21417 );
and ( n21419 , n21412 , n21417 );
or ( n21420 , n21415 , n21418 , n21419 );
and ( n21421 , n21353 , n21420 );
xor ( n21422 , n21412 , n21414 );
xor ( n21423 , n21422 , n21417 );
and ( n21424 , n21302 , n20949 );
buf ( n21425 , n21424 );
and ( n21426 , n21060 , n21296 );
and ( n21427 , n21425 , n21426 );
buf ( n21428 , n20208 );
buf ( n21429 , n21428 );
and ( n21430 , n21019 , n21429 );
and ( n21431 , n21426 , n21430 );
and ( n21432 , n21425 , n21430 );
or ( n21433 , n21427 , n21431 , n21432 );
xor ( n21434 , n21356 , n21357 );
xor ( n21435 , n21434 , n21359 );
and ( n21436 , n21433 , n21435 );
xor ( n21437 , n21364 , n21365 );
xor ( n21438 , n21437 , n21367 );
and ( n21439 , n21435 , n21438 );
and ( n21440 , n21433 , n21438 );
or ( n21441 , n21436 , n21439 , n21440 );
and ( n21442 , n21385 , n20890 );
and ( n21443 , n21355 , n20909 );
and ( n21444 , n21442 , n21443 );
and ( n21445 , n21091 , n21296 );
and ( n21446 , n21443 , n21445 );
and ( n21447 , n21442 , n21445 );
or ( n21448 , n21444 , n21446 , n21447 );
not ( n21449 , n21363 );
and ( n21450 , n21448 , n21449 );
and ( n21451 , n21173 , n21039 );
and ( n21452 , n21449 , n21451 );
and ( n21453 , n21448 , n21451 );
or ( n21454 , n21450 , n21452 , n21453 );
buf ( n21455 , n20238 );
buf ( n21456 , n21455 );
and ( n21457 , n21456 , n20877 );
not ( n21458 , n21424 );
and ( n21459 , n21457 , n21458 );
and ( n21460 , n21173 , n21085 );
and ( n21461 , n21458 , n21460 );
and ( n21462 , n21457 , n21460 );
or ( n21463 , n21459 , n21461 , n21462 );
xor ( n21464 , n21377 , n21378 );
xor ( n21465 , n21464 , n21380 );
and ( n21466 , n21463 , n21465 );
xor ( n21467 , n21386 , n21387 );
xor ( n21468 , n21467 , n21389 );
and ( n21469 , n21465 , n21468 );
and ( n21470 , n21463 , n21468 );
or ( n21471 , n21466 , n21469 , n21470 );
and ( n21472 , n21454 , n21471 );
xor ( n21473 , n21383 , n21392 );
xor ( n21474 , n21473 , n21395 );
and ( n21475 , n21471 , n21474 );
and ( n21476 , n21454 , n21474 );
or ( n21477 , n21472 , n21475 , n21476 );
and ( n21478 , n21441 , n21477 );
xor ( n21479 , n21362 , n21370 );
xor ( n21480 , n21479 , n21373 );
and ( n21481 , n21477 , n21480 );
and ( n21482 , n21441 , n21480 );
or ( n21483 , n21478 , n21481 , n21482 );
xor ( n21484 , n21330 , n21332 );
xor ( n21485 , n21484 , n21335 );
and ( n21486 , n21483 , n21485 );
xor ( n21487 , n21376 , n21406 );
xor ( n21488 , n21487 , n21409 );
and ( n21489 , n21485 , n21488 );
and ( n21490 , n21483 , n21488 );
or ( n21491 , n21486 , n21489 , n21490 );
and ( n21492 , n21423 , n21491 );
and ( n21493 , n21238 , n21039 );
and ( n21494 , n21123 , n21178 );
and ( n21495 , n21493 , n21494 );
and ( n21496 , n21060 , n21429 );
and ( n21497 , n21494 , n21496 );
and ( n21498 , n21493 , n21496 );
or ( n21499 , n21495 , n21497 , n21498 );
xor ( n21500 , n21425 , n21426 );
xor ( n21501 , n21500 , n21430 );
and ( n21502 , n21499 , n21501 );
xor ( n21503 , n21448 , n21449 );
xor ( n21504 , n21503 , n21451 );
and ( n21505 , n21501 , n21504 );
and ( n21506 , n21499 , n21504 );
or ( n21507 , n21502 , n21505 , n21506 );
and ( n21508 , n21456 , n20890 );
and ( n21509 , n21385 , n20909 );
and ( n21510 , n21508 , n21509 );
buf ( n21511 , n21019 );
and ( n21512 , n21509 , n21511 );
and ( n21513 , n21508 , n21511 );
or ( n21514 , n21510 , n21512 , n21513 );
and ( n21515 , n21355 , n20949 );
buf ( n21516 , n21515 );
and ( n21517 , n21514 , n21516 );
xor ( n21518 , n21442 , n21443 );
xor ( n21519 , n21518 , n21445 );
and ( n21520 , n21516 , n21519 );
and ( n21521 , n21514 , n21519 );
or ( n21522 , n21517 , n21520 , n21521 );
and ( n21523 , n21173 , n21178 );
and ( n21524 , n21123 , n21296 );
and ( n21525 , n21523 , n21524 );
buf ( n21526 , n20211 );
buf ( n21527 , n21526 );
and ( n21528 , n21060 , n21527 );
and ( n21529 , n21524 , n21528 );
and ( n21530 , n21523 , n21528 );
or ( n21531 , n21525 , n21529 , n21530 );
and ( n21532 , n21385 , n20949 );
buf ( n21533 , n21532 );
buf ( n21534 , n20241 );
buf ( n21535 , n21534 );
and ( n21536 , n21535 , n20877 );
and ( n21537 , n21533 , n21536 );
and ( n21538 , n21238 , n21085 );
and ( n21539 , n21536 , n21538 );
and ( n21540 , n21533 , n21538 );
or ( n21541 , n21537 , n21539 , n21540 );
and ( n21542 , n21531 , n21541 );
xor ( n21543 , n21457 , n21458 );
xor ( n21544 , n21543 , n21460 );
and ( n21545 , n21541 , n21544 );
and ( n21546 , n21531 , n21544 );
or ( n21547 , n21542 , n21545 , n21546 );
and ( n21548 , n21522 , n21547 );
xor ( n21549 , n21463 , n21465 );
xor ( n21550 , n21549 , n21468 );
and ( n21551 , n21547 , n21550 );
and ( n21552 , n21522 , n21550 );
or ( n21553 , n21548 , n21551 , n21552 );
and ( n21554 , n21507 , n21553 );
xor ( n21555 , n21433 , n21435 );
xor ( n21556 , n21555 , n21438 );
and ( n21557 , n21553 , n21556 );
and ( n21558 , n21507 , n21556 );
or ( n21559 , n21554 , n21557 , n21558 );
xor ( n21560 , n21398 , n21400 );
xor ( n21561 , n21560 , n21403 );
and ( n21562 , n21559 , n21561 );
xor ( n21563 , n21441 , n21477 );
xor ( n21564 , n21563 , n21480 );
and ( n21565 , n21561 , n21564 );
and ( n21566 , n21559 , n21564 );
or ( n21567 , n21562 , n21565 , n21566 );
xor ( n21568 , n21483 , n21485 );
xor ( n21569 , n21568 , n21488 );
and ( n21570 , n21567 , n21569 );
xor ( n21571 , n21559 , n21561 );
xor ( n21572 , n21571 , n21564 );
not ( n21573 , n21515 );
and ( n21574 , n21302 , n21039 );
and ( n21575 , n21573 , n21574 );
and ( n21576 , n21091 , n21429 );
and ( n21577 , n21574 , n21576 );
and ( n21578 , n21573 , n21576 );
or ( n21579 , n21575 , n21577 , n21578 );
and ( n21580 , n21535 , n20890 );
and ( n21581 , n21456 , n20909 );
and ( n21582 , n21580 , n21581 );
and ( n21583 , n21173 , n21296 );
and ( n21584 , n21581 , n21583 );
and ( n21585 , n21580 , n21583 );
or ( n21586 , n21582 , n21584 , n21585 );
and ( n21587 , n21456 , n20949 );
buf ( n21588 , n21587 );
and ( n21589 , n21302 , n21085 );
and ( n21590 , n21588 , n21589 );
and ( n21591 , n21091 , n21527 );
and ( n21592 , n21589 , n21591 );
and ( n21593 , n21588 , n21591 );
or ( n21594 , n21590 , n21592 , n21593 );
and ( n21595 , n21586 , n21594 );
xor ( n21596 , n21508 , n21509 );
xor ( n21597 , n21596 , n21511 );
and ( n21598 , n21594 , n21597 );
and ( n21599 , n21586 , n21597 );
or ( n21600 , n21595 , n21598 , n21599 );
and ( n21601 , n21579 , n21600 );
xor ( n21602 , n21493 , n21494 );
xor ( n21603 , n21602 , n21496 );
and ( n21604 , n21600 , n21603 );
and ( n21605 , n21579 , n21603 );
or ( n21606 , n21601 , n21604 , n21605 );
buf ( n21607 , n20244 );
buf ( n21608 , n21607 );
and ( n21609 , n21608 , n20877 );
not ( n21610 , n21532 );
and ( n21611 , n21609 , n21610 );
and ( n21612 , n21238 , n21178 );
and ( n21613 , n21610 , n21612 );
and ( n21614 , n21609 , n21612 );
or ( n21615 , n21611 , n21613 , n21614 );
xor ( n21616 , n21523 , n21524 );
xor ( n21617 , n21616 , n21528 );
and ( n21618 , n21615 , n21617 );
xor ( n21619 , n21533 , n21536 );
xor ( n21620 , n21619 , n21538 );
and ( n21621 , n21617 , n21620 );
and ( n21622 , n21615 , n21620 );
or ( n21623 , n21618 , n21621 , n21622 );
xor ( n21624 , n21514 , n21516 );
xor ( n21625 , n21624 , n21519 );
and ( n21626 , n21623 , n21625 );
xor ( n21627 , n21531 , n21541 );
xor ( n21628 , n21627 , n21544 );
and ( n21629 , n21625 , n21628 );
and ( n21630 , n21623 , n21628 );
or ( n21631 , n21626 , n21629 , n21630 );
and ( n21632 , n21606 , n21631 );
xor ( n21633 , n21499 , n21501 );
xor ( n21634 , n21633 , n21504 );
and ( n21635 , n21631 , n21634 );
and ( n21636 , n21606 , n21634 );
or ( n21637 , n21632 , n21635 , n21636 );
xor ( n21638 , n21454 , n21471 );
xor ( n21639 , n21638 , n21474 );
and ( n21640 , n21637 , n21639 );
xor ( n21641 , n21507 , n21553 );
xor ( n21642 , n21641 , n21556 );
and ( n21643 , n21639 , n21642 );
and ( n21644 , n21637 , n21642 );
or ( n21645 , n21640 , n21643 , n21644 );
and ( n21646 , n21572 , n21645 );
xor ( n21647 , n21637 , n21639 );
xor ( n21648 , n21647 , n21642 );
and ( n21649 , n21535 , n20909 );
and ( n21650 , n21238 , n21296 );
and ( n21651 , n21649 , n21650 );
buf ( n21652 , n21060 );
and ( n21653 , n21650 , n21652 );
and ( n21654 , n21649 , n21652 );
or ( n21655 , n21651 , n21653 , n21654 );
and ( n21656 , n21355 , n21039 );
and ( n21657 , n21655 , n21656 );
and ( n21658 , n21123 , n21429 );
and ( n21659 , n21656 , n21658 );
and ( n21660 , n21655 , n21658 );
or ( n21661 , n21657 , n21659 , n21660 );
and ( n21662 , n21608 , n20890 );
and ( n21663 , n21123 , n21527 );
and ( n21664 , n21662 , n21663 );
buf ( n21665 , n20214 );
buf ( n21666 , n21665 );
and ( n21667 , n21091 , n21666 );
and ( n21668 , n21663 , n21667 );
and ( n21669 , n21662 , n21667 );
or ( n21670 , n21664 , n21668 , n21669 );
buf ( n21671 , n20247 );
buf ( n21672 , n21671 );
and ( n21673 , n21672 , n20877 );
not ( n21674 , n21587 );
and ( n21675 , n21673 , n21674 );
and ( n21676 , n21302 , n21178 );
and ( n21677 , n21674 , n21676 );
and ( n21678 , n21673 , n21676 );
or ( n21679 , n21675 , n21677 , n21678 );
and ( n21680 , n21670 , n21679 );
xor ( n21681 , n21580 , n21581 );
xor ( n21682 , n21681 , n21583 );
and ( n21683 , n21679 , n21682 );
and ( n21684 , n21670 , n21682 );
or ( n21685 , n21680 , n21683 , n21684 );
and ( n21686 , n21661 , n21685 );
xor ( n21687 , n21573 , n21574 );
xor ( n21688 , n21687 , n21576 );
and ( n21689 , n21685 , n21688 );
and ( n21690 , n21661 , n21688 );
or ( n21691 , n21686 , n21689 , n21690 );
and ( n21692 , n21535 , n20949 );
buf ( n21693 , n21692 );
and ( n21694 , n21385 , n21039 );
and ( n21695 , n21693 , n21694 );
and ( n21696 , n21355 , n21085 );
and ( n21697 , n21694 , n21696 );
and ( n21698 , n21693 , n21696 );
or ( n21699 , n21695 , n21697 , n21698 );
xor ( n21700 , n21588 , n21589 );
xor ( n21701 , n21700 , n21591 );
and ( n21702 , n21699 , n21701 );
xor ( n21703 , n21609 , n21610 );
xor ( n21704 , n21703 , n21612 );
and ( n21705 , n21701 , n21704 );
and ( n21706 , n21699 , n21704 );
or ( n21707 , n21702 , n21705 , n21706 );
xor ( n21708 , n21615 , n21617 );
xor ( n21709 , n21708 , n21620 );
and ( n21710 , n21707 , n21709 );
xor ( n21711 , n21586 , n21594 );
xor ( n21712 , n21711 , n21597 );
and ( n21713 , n21709 , n21712 );
and ( n21714 , n21707 , n21712 );
or ( n21715 , n21710 , n21713 , n21714 );
and ( n21716 , n21691 , n21715 );
xor ( n21717 , n21579 , n21600 );
xor ( n21718 , n21717 , n21603 );
and ( n21719 , n21715 , n21718 );
and ( n21720 , n21691 , n21718 );
or ( n21721 , n21716 , n21719 , n21720 );
xor ( n21722 , n21522 , n21547 );
xor ( n21723 , n21722 , n21550 );
and ( n21724 , n21721 , n21723 );
xor ( n21725 , n21606 , n21631 );
xor ( n21726 , n21725 , n21634 );
and ( n21727 , n21723 , n21726 );
and ( n21728 , n21721 , n21726 );
or ( n21729 , n21724 , n21727 , n21728 );
and ( n21730 , n21648 , n21729 );
xor ( n21731 , n21721 , n21723 );
xor ( n21732 , n21731 , n21726 );
and ( n21733 , n21672 , n20890 );
and ( n21734 , n21608 , n20909 );
and ( n21735 , n21733 , n21734 );
and ( n21736 , n21302 , n21296 );
and ( n21737 , n21734 , n21736 );
and ( n21738 , n21733 , n21736 );
or ( n21739 , n21735 , n21737 , n21738 );
and ( n21740 , n21608 , n20949 );
buf ( n21741 , n21740 );
buf ( n21742 , n20252 );
buf ( n21743 , n21742 );
and ( n21744 , n21743 , n20877 );
and ( n21745 , n21741 , n21744 );
and ( n21746 , n21385 , n21085 );
and ( n21747 , n21744 , n21746 );
and ( n21748 , n21741 , n21746 );
or ( n21749 , n21745 , n21747 , n21748 );
and ( n21750 , n21739 , n21749 );
and ( n21751 , n21173 , n21429 );
and ( n21752 , n21749 , n21751 );
and ( n21753 , n21739 , n21751 );
or ( n21754 , n21750 , n21752 , n21753 );
xor ( n21755 , n21655 , n21656 );
xor ( n21756 , n21755 , n21658 );
and ( n21757 , n21754 , n21756 );
xor ( n21758 , n21670 , n21679 );
xor ( n21759 , n21758 , n21682 );
and ( n21760 , n21756 , n21759 );
and ( n21761 , n21754 , n21759 );
or ( n21762 , n21757 , n21760 , n21761 );
not ( n21763 , n21692 );
and ( n21764 , n21456 , n21039 );
and ( n21765 , n21763 , n21764 );
and ( n21766 , n21238 , n21429 );
and ( n21767 , n21764 , n21766 );
and ( n21768 , n21763 , n21766 );
or ( n21769 , n21765 , n21767 , n21768 );
xor ( n21770 , n21662 , n21663 );
xor ( n21771 , n21770 , n21667 );
and ( n21772 , n21769 , n21771 );
xor ( n21773 , n21673 , n21674 );
xor ( n21774 , n21773 , n21676 );
and ( n21775 , n21771 , n21774 );
and ( n21776 , n21769 , n21774 );
or ( n21777 , n21772 , n21775 , n21776 );
and ( n21778 , n21355 , n21178 );
and ( n21779 , n21173 , n21527 );
and ( n21780 , n21778 , n21779 );
and ( n21781 , n21123 , n21666 );
and ( n21782 , n21779 , n21781 );
and ( n21783 , n21778 , n21781 );
or ( n21784 , n21780 , n21782 , n21783 );
xor ( n21785 , n21649 , n21650 );
xor ( n21786 , n21785 , n21652 );
and ( n21787 , n21784 , n21786 );
xor ( n21788 , n21693 , n21694 );
xor ( n21789 , n21788 , n21696 );
and ( n21790 , n21786 , n21789 );
and ( n21791 , n21784 , n21789 );
or ( n21792 , n21787 , n21790 , n21791 );
and ( n21793 , n21777 , n21792 );
xor ( n21794 , n21699 , n21701 );
xor ( n21795 , n21794 , n21704 );
and ( n21796 , n21792 , n21795 );
and ( n21797 , n21777 , n21795 );
or ( n21798 , n21793 , n21796 , n21797 );
and ( n21799 , n21762 , n21798 );
xor ( n21800 , n21661 , n21685 );
xor ( n21801 , n21800 , n21688 );
and ( n21802 , n21798 , n21801 );
and ( n21803 , n21762 , n21801 );
or ( n21804 , n21799 , n21802 , n21803 );
xor ( n21805 , n21623 , n21625 );
xor ( n21806 , n21805 , n21628 );
and ( n21807 , n21804 , n21806 );
xor ( n21808 , n21691 , n21715 );
xor ( n21809 , n21808 , n21718 );
and ( n21810 , n21806 , n21809 );
and ( n21811 , n21804 , n21809 );
or ( n21812 , n21807 , n21810 , n21811 );
and ( n21813 , n21732 , n21812 );
xor ( n21814 , n21804 , n21806 );
xor ( n21815 , n21814 , n21809 );
and ( n21816 , n21743 , n20890 );
and ( n21817 , n21672 , n20909 );
and ( n21818 , n21816 , n21817 );
buf ( n21819 , n21091 );
and ( n21820 , n21817 , n21819 );
and ( n21821 , n21816 , n21819 );
or ( n21822 , n21818 , n21820 , n21821 );
and ( n21823 , n21456 , n21085 );
and ( n21824 , n21173 , n21666 );
and ( n21825 , n21823 , n21824 );
buf ( n21826 , n20217 );
buf ( n21827 , n21826 );
and ( n21828 , n21123 , n21827 );
and ( n21829 , n21824 , n21828 );
and ( n21830 , n21823 , n21828 );
or ( n21831 , n21825 , n21829 , n21830 );
and ( n21832 , n21822 , n21831 );
and ( n21833 , n21672 , n20949 );
buf ( n21834 , n21833 );
buf ( n21835 , n20257 );
buf ( n21836 , n21835 );
and ( n21837 , n21836 , n20877 );
and ( n21838 , n21834 , n21837 );
and ( n21839 , n21385 , n21178 );
and ( n21840 , n21837 , n21839 );
and ( n21841 , n21834 , n21839 );
or ( n21842 , n21838 , n21840 , n21841 );
and ( n21843 , n21831 , n21842 );
and ( n21844 , n21822 , n21842 );
or ( n21845 , n21832 , n21843 , n21844 );
not ( n21846 , n21740 );
and ( n21847 , n21355 , n21296 );
and ( n21848 , n21846 , n21847 );
and ( n21849 , n21238 , n21527 );
and ( n21850 , n21847 , n21849 );
and ( n21851 , n21846 , n21849 );
or ( n21852 , n21848 , n21850 , n21851 );
xor ( n21853 , n21733 , n21734 );
xor ( n21854 , n21853 , n21736 );
and ( n21855 , n21852 , n21854 );
xor ( n21856 , n21741 , n21744 );
xor ( n21857 , n21856 , n21746 );
and ( n21858 , n21854 , n21857 );
and ( n21859 , n21852 , n21857 );
or ( n21860 , n21855 , n21858 , n21859 );
and ( n21861 , n21845 , n21860 );
xor ( n21862 , n21739 , n21749 );
xor ( n21863 , n21862 , n21751 );
and ( n21864 , n21860 , n21863 );
and ( n21865 , n21845 , n21863 );
or ( n21866 , n21861 , n21864 , n21865 );
and ( n21867 , n21743 , n20909 );
and ( n21868 , n21385 , n21296 );
and ( n21869 , n21867 , n21868 );
and ( n21870 , n21173 , n21827 );
and ( n21871 , n21868 , n21870 );
and ( n21872 , n21867 , n21870 );
or ( n21873 , n21869 , n21871 , n21872 );
and ( n21874 , n21535 , n21039 );
and ( n21875 , n21873 , n21874 );
and ( n21876 , n21302 , n21429 );
and ( n21877 , n21874 , n21876 );
and ( n21878 , n21873 , n21876 );
or ( n21879 , n21875 , n21877 , n21878 );
xor ( n21880 , n21778 , n21779 );
xor ( n21881 , n21880 , n21781 );
and ( n21882 , n21879 , n21881 );
xor ( n21883 , n21763 , n21764 );
xor ( n21884 , n21883 , n21766 );
and ( n21885 , n21881 , n21884 );
and ( n21886 , n21879 , n21884 );
or ( n21887 , n21882 , n21885 , n21886 );
xor ( n21888 , n21769 , n21771 );
xor ( n21889 , n21888 , n21774 );
and ( n21890 , n21887 , n21889 );
xor ( n21891 , n21784 , n21786 );
xor ( n21892 , n21891 , n21789 );
and ( n21893 , n21889 , n21892 );
and ( n21894 , n21887 , n21892 );
or ( n21895 , n21890 , n21893 , n21894 );
and ( n21896 , n21866 , n21895 );
xor ( n21897 , n21754 , n21756 );
xor ( n21898 , n21897 , n21759 );
and ( n21899 , n21895 , n21898 );
and ( n21900 , n21866 , n21898 );
or ( n21901 , n21896 , n21899 , n21900 );
xor ( n21902 , n21707 , n21709 );
xor ( n21903 , n21902 , n21712 );
and ( n21904 , n21901 , n21903 );
xor ( n21905 , n21762 , n21798 );
xor ( n21906 , n21905 , n21801 );
and ( n21907 , n21903 , n21906 );
and ( n21908 , n21901 , n21906 );
or ( n21909 , n21904 , n21907 , n21908 );
and ( n21910 , n21815 , n21909 );
xor ( n21911 , n21901 , n21903 );
xor ( n21912 , n21911 , n21906 );
buf ( n21913 , n20262 );
buf ( n21914 , n21913 );
and ( n21915 , n21914 , n20877 );
and ( n21916 , n21456 , n21178 );
and ( n21917 , n21915 , n21916 );
and ( n21918 , n21302 , n21527 );
and ( n21919 , n21916 , n21918 );
and ( n21920 , n21915 , n21918 );
or ( n21921 , n21917 , n21919 , n21920 );
and ( n21922 , n21836 , n20890 );
not ( n21923 , n21833 );
and ( n21924 , n21922 , n21923 );
and ( n21925 , n21238 , n21666 );
and ( n21926 , n21923 , n21925 );
and ( n21927 , n21922 , n21925 );
or ( n21928 , n21924 , n21926 , n21927 );
and ( n21929 , n21921 , n21928 );
xor ( n21930 , n21816 , n21817 );
xor ( n21931 , n21930 , n21819 );
and ( n21932 , n21928 , n21931 );
and ( n21933 , n21921 , n21931 );
or ( n21934 , n21929 , n21932 , n21933 );
xor ( n21935 , n21823 , n21824 );
xor ( n21936 , n21935 , n21828 );
xor ( n21937 , n21834 , n21837 );
xor ( n21938 , n21937 , n21839 );
and ( n21939 , n21936 , n21938 );
xor ( n21940 , n21846 , n21847 );
xor ( n21941 , n21940 , n21849 );
and ( n21942 , n21938 , n21941 );
and ( n21943 , n21936 , n21941 );
or ( n21944 , n21939 , n21942 , n21943 );
and ( n21945 , n21934 , n21944 );
xor ( n21946 , n21852 , n21854 );
xor ( n21947 , n21946 , n21857 );
and ( n21948 , n21944 , n21947 );
and ( n21949 , n21934 , n21947 );
or ( n21950 , n21945 , n21948 , n21949 );
xor ( n21951 , n21845 , n21860 );
xor ( n21952 , n21951 , n21863 );
and ( n21953 , n21950 , n21952 );
xor ( n21954 , n21887 , n21889 );
xor ( n21955 , n21954 , n21892 );
and ( n21956 , n21952 , n21955 );
and ( n21957 , n21950 , n21955 );
or ( n21958 , n21953 , n21956 , n21957 );
xor ( n21959 , n21777 , n21792 );
xor ( n21960 , n21959 , n21795 );
and ( n21961 , n21958 , n21960 );
xor ( n21962 , n21866 , n21895 );
xor ( n21963 , n21962 , n21898 );
and ( n21964 , n21960 , n21963 );
and ( n21965 , n21958 , n21963 );
or ( n21966 , n21961 , n21964 , n21965 );
and ( n21967 , n21912 , n21966 );
xor ( n21968 , n21958 , n21960 );
xor ( n21969 , n21968 , n21963 );
and ( n21970 , n21743 , n20949 );
buf ( n21971 , n21970 );
and ( n21972 , n21608 , n21039 );
and ( n21973 , n21971 , n21972 );
and ( n21974 , n21535 , n21085 );
and ( n21975 , n21972 , n21974 );
and ( n21976 , n21971 , n21974 );
or ( n21977 , n21973 , n21975 , n21976 );
and ( n21978 , n21836 , n20949 );
buf ( n21979 , n21978 );
and ( n21980 , n21608 , n21085 );
and ( n21981 , n21979 , n21980 );
and ( n21982 , n21535 , n21178 );
and ( n21983 , n21980 , n21982 );
and ( n21984 , n21979 , n21982 );
or ( n21985 , n21981 , n21983 , n21984 );
not ( n21986 , n21970 );
and ( n21987 , n21355 , n21527 );
and ( n21988 , n21986 , n21987 );
buf ( n21989 , n20220 );
buf ( n21990 , n21989 );
and ( n21991 , n21173 , n21990 );
and ( n21992 , n21987 , n21991 );
and ( n21993 , n21986 , n21991 );
or ( n21994 , n21988 , n21992 , n21993 );
and ( n21995 , n21985 , n21994 );
xor ( n21996 , n21867 , n21868 );
xor ( n21997 , n21996 , n21870 );
and ( n21998 , n21994 , n21997 );
and ( n21999 , n21985 , n21997 );
or ( n22000 , n21995 , n21998 , n21999 );
and ( n22001 , n21977 , n22000 );
xor ( n22002 , n21873 , n21874 );
xor ( n22003 , n22002 , n21876 );
and ( n22004 , n22000 , n22003 );
and ( n22005 , n21977 , n22003 );
or ( n22006 , n22001 , n22004 , n22005 );
xor ( n22007 , n21822 , n21831 );
xor ( n22008 , n22007 , n21842 );
and ( n22009 , n22006 , n22008 );
xor ( n22010 , n21879 , n21881 );
xor ( n22011 , n22010 , n21884 );
and ( n22012 , n22008 , n22011 );
and ( n22013 , n22006 , n22011 );
or ( n22014 , n22009 , n22012 , n22013 );
and ( n22015 , n21914 , n20890 );
and ( n22016 , n21836 , n20909 );
and ( n22017 , n22015 , n22016 );
buf ( n22018 , n21123 );
and ( n22019 , n22016 , n22018 );
and ( n22020 , n22015 , n22018 );
or ( n22021 , n22017 , n22019 , n22020 );
and ( n22022 , n21456 , n21296 );
and ( n22023 , n21302 , n21666 );
and ( n22024 , n22022 , n22023 );
and ( n22025 , n21238 , n21827 );
and ( n22026 , n22023 , n22025 );
and ( n22027 , n22022 , n22025 );
or ( n22028 , n22024 , n22026 , n22027 );
and ( n22029 , n22021 , n22028 );
and ( n22030 , n21355 , n21429 );
and ( n22031 , n22028 , n22030 );
and ( n22032 , n22021 , n22030 );
or ( n22033 , n22029 , n22031 , n22032 );
buf ( n22034 , n20267 );
buf ( n22035 , n22034 );
and ( n22036 , n22035 , n20877 );
and ( n22037 , n21672 , n21039 );
and ( n22038 , n22036 , n22037 );
and ( n22039 , n21385 , n21429 );
and ( n22040 , n22037 , n22039 );
and ( n22041 , n22036 , n22039 );
or ( n22042 , n22038 , n22040 , n22041 );
xor ( n22043 , n21915 , n21916 );
xor ( n22044 , n22043 , n21918 );
and ( n22045 , n22042 , n22044 );
xor ( n22046 , n21922 , n21923 );
xor ( n22047 , n22046 , n21925 );
and ( n22048 , n22044 , n22047 );
and ( n22049 , n22042 , n22047 );
or ( n22050 , n22045 , n22048 , n22049 );
and ( n22051 , n22033 , n22050 );
xor ( n22052 , n21921 , n21928 );
xor ( n22053 , n22052 , n21931 );
and ( n22054 , n22050 , n22053 );
and ( n22055 , n22033 , n22053 );
or ( n22056 , n22051 , n22054 , n22055 );
and ( n22057 , n22035 , n20890 );
and ( n22058 , n21914 , n20909 );
and ( n22059 , n22057 , n22058 );
and ( n22060 , n21302 , n21827 );
and ( n22061 , n22058 , n22060 );
and ( n22062 , n22057 , n22060 );
or ( n22063 , n22059 , n22061 , n22062 );
and ( n22064 , n21672 , n21085 );
and ( n22065 , n21355 , n21666 );
and ( n22066 , n22064 , n22065 );
and ( n22067 , n21238 , n21990 );
and ( n22068 , n22065 , n22067 );
and ( n22069 , n22064 , n22067 );
or ( n22070 , n22066 , n22068 , n22069 );
and ( n22071 , n22063 , n22070 );
not ( n22072 , n21978 );
and ( n22073 , n21535 , n21296 );
and ( n22074 , n22072 , n22073 );
and ( n22075 , n21385 , n21527 );
and ( n22076 , n22073 , n22075 );
and ( n22077 , n22072 , n22075 );
or ( n22078 , n22074 , n22076 , n22077 );
and ( n22079 , n22070 , n22078 );
and ( n22080 , n22063 , n22078 );
or ( n22081 , n22071 , n22079 , n22080 );
xor ( n22082 , n21971 , n21972 );
xor ( n22083 , n22082 , n21974 );
and ( n22084 , n22081 , n22083 );
xor ( n22085 , n22021 , n22028 );
xor ( n22086 , n22085 , n22030 );
and ( n22087 , n22083 , n22086 );
and ( n22088 , n22081 , n22086 );
or ( n22089 , n22084 , n22087 , n22088 );
xor ( n22090 , n21936 , n21938 );
xor ( n22091 , n22090 , n21941 );
and ( n22092 , n22089 , n22091 );
xor ( n22093 , n21977 , n22000 );
xor ( n22094 , n22093 , n22003 );
and ( n22095 , n22091 , n22094 );
and ( n22096 , n22089 , n22094 );
or ( n22097 , n22092 , n22095 , n22096 );
and ( n22098 , n22056 , n22097 );
xor ( n22099 , n21934 , n21944 );
xor ( n22100 , n22099 , n21947 );
and ( n22101 , n22097 , n22100 );
and ( n22102 , n22056 , n22100 );
or ( n22103 , n22098 , n22101 , n22102 );
and ( n22104 , n22014 , n22103 );
xor ( n22105 , n21950 , n21952 );
xor ( n22106 , n22105 , n21955 );
and ( n22107 , n22103 , n22106 );
and ( n22108 , n22014 , n22106 );
or ( n22109 , n22104 , n22107 , n22108 );
and ( n22110 , n21969 , n22109 );
xor ( n22111 , n22014 , n22103 );
xor ( n22112 , n22111 , n22106 );
buf ( n22113 , n21173 );
buf ( n22114 , n22113 );
buf ( n22115 , n20270 );
buf ( n22116 , n22115 );
and ( n22117 , n22116 , n20877 );
and ( n22118 , n22114 , n22117 );
and ( n22119 , n21608 , n21178 );
and ( n22120 , n22117 , n22119 );
and ( n22121 , n22114 , n22119 );
or ( n22122 , n22118 , n22120 , n22121 );
xor ( n22123 , n22015 , n22016 );
xor ( n22124 , n22123 , n22018 );
and ( n22125 , n22122 , n22124 );
xor ( n22126 , n22022 , n22023 );
xor ( n22127 , n22126 , n22025 );
and ( n22128 , n22124 , n22127 );
and ( n22129 , n22122 , n22127 );
or ( n22130 , n22125 , n22128 , n22129 );
xor ( n22131 , n22042 , n22044 );
xor ( n22132 , n22131 , n22047 );
and ( n22133 , n22130 , n22132 );
xor ( n22134 , n21985 , n21994 );
xor ( n22135 , n22134 , n21997 );
and ( n22136 , n22132 , n22135 );
and ( n22137 , n22130 , n22135 );
or ( n22138 , n22133 , n22136 , n22137 );
xor ( n22139 , n22033 , n22050 );
xor ( n22140 , n22139 , n22053 );
and ( n22141 , n22138 , n22140 );
xor ( n22142 , n22089 , n22091 );
xor ( n22143 , n22142 , n22094 );
and ( n22144 , n22140 , n22143 );
and ( n22145 , n22138 , n22143 );
or ( n22146 , n22141 , n22144 , n22145 );
xor ( n22147 , n22006 , n22008 );
xor ( n22148 , n22147 , n22011 );
and ( n22149 , n22146 , n22148 );
xor ( n22150 , n22056 , n22097 );
xor ( n22151 , n22150 , n22100 );
and ( n22152 , n22148 , n22151 );
and ( n22153 , n22146 , n22151 );
or ( n22154 , n22149 , n22152 , n22153 );
and ( n22155 , n22112 , n22154 );
xor ( n22156 , n22146 , n22148 );
xor ( n22157 , n22156 , n22151 );
xor ( n22158 , n22036 , n22037 );
xor ( n22159 , n22158 , n22039 );
xor ( n22160 , n21979 , n21980 );
xor ( n22161 , n22160 , n21982 );
and ( n22162 , n22159 , n22161 );
xor ( n22163 , n21986 , n21987 );
xor ( n22164 , n22163 , n21991 );
and ( n22165 , n22161 , n22164 );
and ( n22166 , n22159 , n22164 );
or ( n22167 , n22162 , n22165 , n22166 );
and ( n22168 , n21914 , n20949 );
and ( n22169 , n21355 , n21827 );
and ( n22170 , n22168 , n22169 );
buf ( n22171 , n20223 );
buf ( n22172 , n22171 );
and ( n22173 , n21238 , n22172 );
and ( n22174 , n22169 , n22173 );
and ( n22175 , n22168 , n22173 );
or ( n22176 , n22170 , n22174 , n22175 );
and ( n22177 , n21743 , n21039 );
and ( n22178 , n22176 , n22177 );
and ( n22179 , n21456 , n21429 );
and ( n22180 , n22177 , n22179 );
and ( n22181 , n22176 , n22179 );
or ( n22182 , n22178 , n22180 , n22181 );
and ( n22183 , n21743 , n21085 );
and ( n22184 , n21456 , n21527 );
and ( n22185 , n22183 , n22184 );
and ( n22186 , n21385 , n21666 );
and ( n22187 , n22184 , n22186 );
and ( n22188 , n22183 , n22186 );
or ( n22189 , n22185 , n22187 , n22188 );
and ( n22190 , n22116 , n20890 );
and ( n22191 , n22035 , n20909 );
and ( n22192 , n22190 , n22191 );
and ( n22193 , n21608 , n21296 );
and ( n22194 , n22191 , n22193 );
and ( n22195 , n22190 , n22193 );
or ( n22196 , n22192 , n22194 , n22195 );
and ( n22197 , n22189 , n22196 );
and ( n22198 , n22035 , n20949 );
buf ( n22199 , n22198 );
and ( n22200 , n21672 , n21178 );
and ( n22201 , n22199 , n22200 );
not ( n22202 , n22113 );
and ( n22203 , n22200 , n22202 );
and ( n22204 , n22199 , n22202 );
or ( n22205 , n22201 , n22203 , n22204 );
and ( n22206 , n22196 , n22205 );
and ( n22207 , n22189 , n22205 );
or ( n22208 , n22197 , n22206 , n22207 );
and ( n22209 , n22182 , n22208 );
xor ( n22210 , n22122 , n22124 );
xor ( n22211 , n22210 , n22127 );
and ( n22212 , n22208 , n22211 );
and ( n22213 , n22182 , n22211 );
or ( n22214 , n22209 , n22212 , n22213 );
and ( n22215 , n22167 , n22214 );
xor ( n22216 , n22081 , n22083 );
xor ( n22217 , n22216 , n22086 );
and ( n22218 , n22214 , n22217 );
and ( n22219 , n22167 , n22217 );
or ( n22220 , n22215 , n22218 , n22219 );
xor ( n22221 , n22064 , n22065 );
xor ( n22222 , n22221 , n22067 );
xor ( n22223 , n22176 , n22177 );
xor ( n22224 , n22223 , n22179 );
and ( n22225 , n22222 , n22224 );
xor ( n22226 , n22072 , n22073 );
xor ( n22227 , n22226 , n22075 );
and ( n22228 , n22224 , n22227 );
and ( n22229 , n22222 , n22227 );
or ( n22230 , n22225 , n22228 , n22229 );
buf ( n22231 , n20273 );
buf ( n22232 , n22231 );
and ( n22233 , n22232 , n20877 );
and ( n22234 , n21836 , n21039 );
and ( n22235 , n22233 , n22234 );
and ( n22236 , n21302 , n21990 );
and ( n22237 , n22234 , n22236 );
and ( n22238 , n22233 , n22236 );
or ( n22239 , n22235 , n22237 , n22238 );
xor ( n22240 , n22057 , n22058 );
xor ( n22241 , n22240 , n22060 );
and ( n22242 , n22239 , n22241 );
xor ( n22243 , n22114 , n22117 );
xor ( n22244 , n22243 , n22119 );
and ( n22245 , n22241 , n22244 );
and ( n22246 , n22239 , n22244 );
or ( n22247 , n22242 , n22245 , n22246 );
and ( n22248 , n22230 , n22247 );
xor ( n22249 , n22063 , n22070 );
xor ( n22250 , n22249 , n22078 );
and ( n22251 , n22247 , n22250 );
and ( n22252 , n22230 , n22250 );
or ( n22253 , n22248 , n22251 , n22252 );
and ( n22254 , n21672 , n21296 );
and ( n22255 , n21456 , n21666 );
and ( n22256 , n22254 , n22255 );
and ( n22257 , n21385 , n21827 );
and ( n22258 , n22255 , n22257 );
and ( n22259 , n22254 , n22257 );
or ( n22260 , n22256 , n22258 , n22259 );
and ( n22261 , n22232 , n20890 );
and ( n22262 , n22116 , n20909 );
and ( n22263 , n22261 , n22262 );
and ( n22264 , n21302 , n22172 );
and ( n22265 , n22262 , n22264 );
and ( n22266 , n22261 , n22264 );
or ( n22267 , n22263 , n22265 , n22266 );
and ( n22268 , n22260 , n22267 );
and ( n22269 , n21535 , n21429 );
and ( n22270 , n22267 , n22269 );
and ( n22271 , n22260 , n22269 );
or ( n22272 , n22268 , n22270 , n22271 );
buf ( n22273 , n21238 );
buf ( n22274 , n22273 );
and ( n22275 , n21836 , n21085 );
and ( n22276 , n22274 , n22275 );
and ( n22277 , n21743 , n21178 );
and ( n22278 , n22275 , n22277 );
and ( n22279 , n22274 , n22277 );
or ( n22280 , n22276 , n22278 , n22279 );
not ( n22281 , n22198 );
and ( n22282 , n21535 , n21527 );
and ( n22283 , n22281 , n22282 );
and ( n22284 , n21355 , n21990 );
and ( n22285 , n22282 , n22284 );
and ( n22286 , n22281 , n22284 );
or ( n22287 , n22283 , n22285 , n22286 );
and ( n22288 , n22280 , n22287 );
xor ( n22289 , n22190 , n22191 );
xor ( n22290 , n22289 , n22193 );
and ( n22291 , n22287 , n22290 );
and ( n22292 , n22280 , n22290 );
or ( n22293 , n22288 , n22291 , n22292 );
and ( n22294 , n22272 , n22293 );
xor ( n22295 , n22189 , n22196 );
xor ( n22296 , n22295 , n22205 );
and ( n22297 , n22293 , n22296 );
and ( n22298 , n22272 , n22296 );
or ( n22299 , n22294 , n22297 , n22298 );
xor ( n22300 , n22159 , n22161 );
xor ( n22301 , n22300 , n22164 );
and ( n22302 , n22299 , n22301 );
xor ( n22303 , n22182 , n22208 );
xor ( n22304 , n22303 , n22211 );
and ( n22305 , n22301 , n22304 );
and ( n22306 , n22299 , n22304 );
or ( n22307 , n22302 , n22305 , n22306 );
and ( n22308 , n22253 , n22307 );
xor ( n22309 , n22130 , n22132 );
xor ( n22310 , n22309 , n22135 );
and ( n22311 , n22307 , n22310 );
and ( n22312 , n22253 , n22310 );
or ( n22313 , n22308 , n22311 , n22312 );
and ( n22314 , n22220 , n22313 );
xor ( n22315 , n22138 , n22140 );
xor ( n22316 , n22315 , n22143 );
and ( n22317 , n22313 , n22316 );
and ( n22318 , n22220 , n22316 );
or ( n22319 , n22314 , n22317 , n22318 );
and ( n22320 , n22157 , n22319 );
xor ( n22321 , n22220 , n22313 );
xor ( n22322 , n22321 , n22316 );
xor ( n22323 , n22183 , n22184 );
xor ( n22324 , n22323 , n22186 );
xor ( n22325 , n22260 , n22267 );
xor ( n22326 , n22325 , n22269 );
and ( n22327 , n22324 , n22326 );
xor ( n22328 , n22199 , n22200 );
xor ( n22329 , n22328 , n22202 );
and ( n22330 , n22326 , n22329 );
and ( n22331 , n22324 , n22329 );
or ( n22332 , n22327 , n22330 , n22331 );
and ( n22333 , n22116 , n20949 );
and ( n22334 , n21743 , n21296 );
and ( n22335 , n22333 , n22334 );
buf ( n22336 , n20226 );
buf ( n22337 , n22336 );
and ( n22338 , n21302 , n22337 );
and ( n22339 , n22334 , n22338 );
and ( n22340 , n22333 , n22338 );
or ( n22341 , n22335 , n22339 , n22340 );
and ( n22342 , n22232 , n20909 );
and ( n22343 , n21456 , n21827 );
and ( n22344 , n22342 , n22343 );
and ( n22345 , n21355 , n22172 );
and ( n22346 , n22343 , n22345 );
and ( n22347 , n22342 , n22345 );
or ( n22348 , n22344 , n22346 , n22347 );
and ( n22349 , n22341 , n22348 );
buf ( n22350 , n20279 );
buf ( n22351 , n22350 );
and ( n22352 , n22351 , n20877 );
buf ( n22353 , n20276 );
buf ( n22354 , n22353 );
and ( n22355 , n22354 , n20890 );
and ( n22356 , n22352 , n22355 );
not ( n22357 , n22273 );
and ( n22358 , n22355 , n22357 );
and ( n22359 , n22352 , n22357 );
or ( n22360 , n22356 , n22358 , n22359 );
and ( n22361 , n22348 , n22360 );
and ( n22362 , n22341 , n22360 );
or ( n22363 , n22349 , n22361 , n22362 );
and ( n22364 , n21914 , n21085 );
and ( n22365 , n21608 , n21527 );
and ( n22366 , n22364 , n22365 );
and ( n22367 , n21535 , n21666 );
and ( n22368 , n22365 , n22367 );
and ( n22369 , n22364 , n22367 );
or ( n22370 , n22366 , n22368 , n22369 );
and ( n22371 , n22232 , n20949 );
buf ( n22372 , n22371 );
and ( n22373 , n21836 , n21178 );
and ( n22374 , n22372 , n22373 );
and ( n22375 , n21385 , n21990 );
and ( n22376 , n22373 , n22375 );
and ( n22377 , n22372 , n22375 );
or ( n22378 , n22374 , n22376 , n22377 );
and ( n22379 , n22370 , n22378 );
xor ( n22380 , n22254 , n22255 );
xor ( n22381 , n22380 , n22257 );
and ( n22382 , n22378 , n22381 );
and ( n22383 , n22370 , n22381 );
or ( n22384 , n22379 , n22382 , n22383 );
and ( n22385 , n22363 , n22384 );
xor ( n22386 , n22280 , n22287 );
xor ( n22387 , n22386 , n22290 );
and ( n22388 , n22384 , n22387 );
and ( n22389 , n22363 , n22387 );
or ( n22390 , n22385 , n22388 , n22389 );
and ( n22391 , n22332 , n22390 );
xor ( n22392 , n22272 , n22293 );
xor ( n22393 , n22392 , n22296 );
and ( n22394 , n22390 , n22393 );
and ( n22395 , n22332 , n22393 );
or ( n22396 , n22391 , n22394 , n22395 );
and ( n22397 , n22354 , n20877 );
and ( n22398 , n21914 , n21039 );
and ( n22399 , n22397 , n22398 );
and ( n22400 , n21608 , n21429 );
and ( n22401 , n22398 , n22400 );
and ( n22402 , n22397 , n22400 );
or ( n22403 , n22399 , n22401 , n22402 );
xor ( n22404 , n22168 , n22169 );
xor ( n22405 , n22404 , n22173 );
and ( n22406 , n22403 , n22405 );
xor ( n22407 , n22233 , n22234 );
xor ( n22408 , n22407 , n22236 );
and ( n22409 , n22405 , n22408 );
and ( n22410 , n22403 , n22408 );
or ( n22411 , n22406 , n22409 , n22410 );
xor ( n22412 , n22222 , n22224 );
xor ( n22413 , n22412 , n22227 );
and ( n22414 , n22411 , n22413 );
xor ( n22415 , n22239 , n22241 );
xor ( n22416 , n22415 , n22244 );
and ( n22417 , n22413 , n22416 );
and ( n22418 , n22411 , n22416 );
or ( n22419 , n22414 , n22417 , n22418 );
and ( n22420 , n22396 , n22419 );
xor ( n22421 , n22230 , n22247 );
xor ( n22422 , n22421 , n22250 );
and ( n22423 , n22419 , n22422 );
and ( n22424 , n22396 , n22422 );
or ( n22425 , n22420 , n22423 , n22424 );
xor ( n22426 , n22167 , n22214 );
xor ( n22427 , n22426 , n22217 );
and ( n22428 , n22425 , n22427 );
xor ( n22429 , n22253 , n22307 );
xor ( n22430 , n22429 , n22310 );
and ( n22431 , n22427 , n22430 );
and ( n22432 , n22425 , n22430 );
or ( n22433 , n22428 , n22431 , n22432 );
and ( n22434 , n22322 , n22433 );
xor ( n22435 , n22261 , n22262 );
xor ( n22436 , n22435 , n22264 );
xor ( n22437 , n22274 , n22275 );
xor ( n22438 , n22437 , n22277 );
and ( n22439 , n22436 , n22438 );
xor ( n22440 , n22281 , n22282 );
xor ( n22441 , n22440 , n22284 );
and ( n22442 , n22438 , n22441 );
and ( n22443 , n22436 , n22441 );
or ( n22444 , n22439 , n22442 , n22443 );
and ( n22445 , n21836 , n21296 );
and ( n22446 , n21535 , n21827 );
and ( n22447 , n22445 , n22446 );
and ( n22448 , n21385 , n22172 );
and ( n22449 , n22446 , n22448 );
and ( n22450 , n22445 , n22448 );
or ( n22451 , n22447 , n22449 , n22450 );
and ( n22452 , n22035 , n21039 );
and ( n22453 , n22451 , n22452 );
and ( n22454 , n21672 , n21429 );
and ( n22455 , n22452 , n22454 );
and ( n22456 , n22451 , n22454 );
or ( n22457 , n22453 , n22455 , n22456 );
xor ( n22458 , n22397 , n22398 );
xor ( n22459 , n22458 , n22400 );
and ( n22460 , n22457 , n22459 );
xor ( n22461 , n22341 , n22348 );
xor ( n22462 , n22461 , n22360 );
and ( n22463 , n22459 , n22462 );
and ( n22464 , n22457 , n22462 );
or ( n22465 , n22460 , n22463 , n22464 );
and ( n22466 , n22444 , n22465 );
xor ( n22467 , n22403 , n22405 );
xor ( n22468 , n22467 , n22408 );
and ( n22469 , n22465 , n22468 );
and ( n22470 , n22444 , n22468 );
or ( n22471 , n22466 , n22469 , n22470 );
and ( n22472 , n22035 , n21085 );
and ( n22473 , n21672 , n21527 );
and ( n22474 , n22472 , n22473 );
and ( n22475 , n21608 , n21666 );
and ( n22476 , n22473 , n22475 );
and ( n22477 , n22472 , n22475 );
or ( n22478 , n22474 , n22476 , n22477 );
buf ( n22479 , n21302 );
buf ( n22480 , n22479 );
and ( n22481 , n22354 , n20909 );
and ( n22482 , n22480 , n22481 );
and ( n22483 , n21355 , n22337 );
and ( n22484 , n22481 , n22483 );
and ( n22485 , n22480 , n22483 );
or ( n22486 , n22482 , n22484 , n22485 );
and ( n22487 , n22478 , n22486 );
and ( n22488 , n22351 , n20890 );
not ( n22489 , n22371 );
and ( n22490 , n22488 , n22489 );
and ( n22491 , n21914 , n21178 );
and ( n22492 , n22489 , n22491 );
and ( n22493 , n22488 , n22491 );
or ( n22494 , n22490 , n22492 , n22493 );
and ( n22495 , n22486 , n22494 );
and ( n22496 , n22478 , n22494 );
or ( n22497 , n22487 , n22495 , n22496 );
xor ( n22498 , n22364 , n22365 );
xor ( n22499 , n22498 , n22367 );
xor ( n22500 , n22372 , n22373 );
xor ( n22501 , n22500 , n22375 );
and ( n22502 , n22499 , n22501 );
xor ( n22503 , n22352 , n22355 );
xor ( n22504 , n22503 , n22357 );
and ( n22505 , n22501 , n22504 );
and ( n22506 , n22499 , n22504 );
or ( n22507 , n22502 , n22505 , n22506 );
and ( n22508 , n22497 , n22507 );
xor ( n22509 , n22370 , n22378 );
xor ( n22510 , n22509 , n22381 );
and ( n22511 , n22507 , n22510 );
and ( n22512 , n22497 , n22510 );
or ( n22513 , n22508 , n22511 , n22512 );
xor ( n22514 , n22324 , n22326 );
xor ( n22515 , n22514 , n22329 );
and ( n22516 , n22513 , n22515 );
xor ( n22517 , n22363 , n22384 );
xor ( n22518 , n22517 , n22387 );
and ( n22519 , n22515 , n22518 );
and ( n22520 , n22513 , n22518 );
or ( n22521 , n22516 , n22519 , n22520 );
and ( n22522 , n22471 , n22521 );
xor ( n22523 , n22411 , n22413 );
xor ( n22524 , n22523 , n22416 );
and ( n22525 , n22521 , n22524 );
and ( n22526 , n22471 , n22524 );
or ( n22527 , n22522 , n22525 , n22526 );
xor ( n22528 , n22396 , n22419 );
xor ( n22529 , n22528 , n22422 );
and ( n22530 , n22527 , n22529 );
xor ( n22531 , n22299 , n22301 );
xor ( n22532 , n22531 , n22304 );
and ( n22533 , n22529 , n22532 );
and ( n22534 , n22527 , n22532 );
or ( n22535 , n22530 , n22533 , n22534 );
xor ( n22536 , n22425 , n22427 );
xor ( n22537 , n22536 , n22430 );
and ( n22538 , n22535 , n22537 );
xor ( n22539 , n22527 , n22529 );
xor ( n22540 , n22539 , n22532 );
buf ( n22541 , n10629 );
buf ( n22542 , n22541 );
and ( n22543 , n22542 , n20877 );
and ( n22544 , n22116 , n21039 );
and ( n22545 , n22543 , n22544 );
and ( n22546 , n21456 , n21990 );
and ( n22547 , n22544 , n22546 );
and ( n22548 , n22543 , n22546 );
or ( n22549 , n22545 , n22547 , n22548 );
xor ( n22550 , n22333 , n22334 );
xor ( n22551 , n22550 , n22338 );
and ( n22552 , n22549 , n22551 );
xor ( n22553 , n22342 , n22343 );
xor ( n22554 , n22553 , n22345 );
and ( n22555 , n22551 , n22554 );
and ( n22556 , n22549 , n22554 );
or ( n22557 , n22552 , n22555 , n22556 );
and ( n22558 , n22542 , n20890 );
and ( n22559 , n22354 , n20949 );
and ( n22560 , n22558 , n22559 );
buf ( n22561 , n20229 );
buf ( n22562 , n22561 );
and ( n22563 , n21355 , n22562 );
and ( n22564 , n22559 , n22563 );
and ( n22565 , n22558 , n22563 );
or ( n22566 , n22560 , n22564 , n22565 );
and ( n22567 , n21914 , n21296 );
and ( n22568 , n21456 , n22172 );
and ( n22569 , n22567 , n22568 );
not ( n22570 , n22479 );
and ( n22571 , n22568 , n22570 );
and ( n22572 , n22567 , n22570 );
or ( n22573 , n22569 , n22571 , n22572 );
and ( n22574 , n22566 , n22573 );
and ( n22575 , n21743 , n21429 );
and ( n22576 , n22573 , n22575 );
and ( n22577 , n22566 , n22575 );
or ( n22578 , n22574 , n22576 , n22577 );
and ( n22579 , n22351 , n20909 );
and ( n22580 , n21608 , n21827 );
and ( n22581 , n22579 , n22580 );
and ( n22582 , n21385 , n22337 );
and ( n22583 , n22580 , n22582 );
and ( n22584 , n22579 , n22582 );
or ( n22585 , n22581 , n22583 , n22584 );
and ( n22586 , n21385 , n22562 );
buf ( n22587 , n22586 );
buf ( n22588 , n10921 );
buf ( n22589 , n22588 );
and ( n22590 , n22589 , n20877 );
and ( n22591 , n22587 , n22590 );
and ( n22592 , n21743 , n21527 );
and ( n22593 , n22590 , n22592 );
and ( n22594 , n22587 , n22592 );
or ( n22595 , n22591 , n22593 , n22594 );
and ( n22596 , n22585 , n22595 );
xor ( n22597 , n22480 , n22481 );
xor ( n22598 , n22597 , n22483 );
and ( n22599 , n22595 , n22598 );
and ( n22600 , n22585 , n22598 );
or ( n22601 , n22596 , n22599 , n22600 );
and ( n22602 , n22578 , n22601 );
xor ( n22603 , n22451 , n22452 );
xor ( n22604 , n22603 , n22454 );
and ( n22605 , n22601 , n22604 );
and ( n22606 , n22578 , n22604 );
or ( n22607 , n22602 , n22605 , n22606 );
and ( n22608 , n22557 , n22607 );
xor ( n22609 , n22436 , n22438 );
xor ( n22610 , n22609 , n22441 );
and ( n22611 , n22607 , n22610 );
and ( n22612 , n22557 , n22610 );
or ( n22613 , n22608 , n22611 , n22612 );
and ( n22614 , n22116 , n21085 );
and ( n22615 , n22035 , n21178 );
and ( n22616 , n22614 , n22615 );
and ( n22617 , n21535 , n21990 );
and ( n22618 , n22615 , n22617 );
and ( n22619 , n22614 , n22617 );
or ( n22620 , n22616 , n22618 , n22619 );
xor ( n22621 , n22543 , n22544 );
xor ( n22622 , n22621 , n22546 );
and ( n22623 , n22620 , n22622 );
xor ( n22624 , n22445 , n22446 );
xor ( n22625 , n22624 , n22448 );
and ( n22626 , n22622 , n22625 );
and ( n22627 , n22620 , n22625 );
or ( n22628 , n22623 , n22626 , n22627 );
and ( n22629 , n22232 , n21039 );
and ( n22630 , n21836 , n21429 );
and ( n22631 , n22629 , n22630 );
and ( n22632 , n21672 , n21666 );
and ( n22633 , n22630 , n22632 );
and ( n22634 , n22629 , n22632 );
or ( n22635 , n22631 , n22633 , n22634 );
xor ( n22636 , n22472 , n22473 );
xor ( n22637 , n22636 , n22475 );
and ( n22638 , n22635 , n22637 );
xor ( n22639 , n22488 , n22489 );
xor ( n22640 , n22639 , n22491 );
and ( n22641 , n22637 , n22640 );
and ( n22642 , n22635 , n22640 );
or ( n22643 , n22638 , n22641 , n22642 );
and ( n22644 , n22628 , n22643 );
xor ( n22645 , n22549 , n22551 );
xor ( n22646 , n22645 , n22554 );
and ( n22647 , n22643 , n22646 );
and ( n22648 , n22628 , n22646 );
or ( n22649 , n22644 , n22647 , n22648 );
xor ( n22650 , n22457 , n22459 );
xor ( n22651 , n22650 , n22462 );
and ( n22652 , n22649 , n22651 );
xor ( n22653 , n22497 , n22507 );
xor ( n22654 , n22653 , n22510 );
and ( n22655 , n22651 , n22654 );
and ( n22656 , n22649 , n22654 );
or ( n22657 , n22652 , n22655 , n22656 );
and ( n22658 , n22613 , n22657 );
xor ( n22659 , n22444 , n22465 );
xor ( n22660 , n22659 , n22468 );
and ( n22661 , n22657 , n22660 );
and ( n22662 , n22613 , n22660 );
or ( n22663 , n22658 , n22661 , n22662 );
xor ( n22664 , n22332 , n22390 );
xor ( n22665 , n22664 , n22393 );
and ( n22666 , n22663 , n22665 );
xor ( n22667 , n22471 , n22521 );
xor ( n22668 , n22667 , n22524 );
and ( n22669 , n22665 , n22668 );
and ( n22670 , n22663 , n22668 );
or ( n22671 , n22666 , n22669 , n22670 );
and ( n22672 , n22540 , n22671 );
xor ( n22673 , n22663 , n22665 );
xor ( n22674 , n22673 , n22668 );
xor ( n22675 , n22478 , n22486 );
xor ( n22676 , n22675 , n22494 );
xor ( n22677 , n22499 , n22501 );
xor ( n22678 , n22677 , n22504 );
and ( n22679 , n22676 , n22678 );
xor ( n22680 , n22578 , n22601 );
xor ( n22681 , n22680 , n22604 );
and ( n22682 , n22678 , n22681 );
and ( n22683 , n22676 , n22681 );
or ( n22684 , n22679 , n22682 , n22683 );
and ( n22685 , n22232 , n21085 );
and ( n22686 , n21836 , n21527 );
and ( n22687 , n22685 , n22686 );
and ( n22688 , n21743 , n21666 );
and ( n22689 , n22686 , n22688 );
and ( n22690 , n22685 , n22688 );
or ( n22691 , n22687 , n22689 , n22690 );
buf ( n22692 , n21355 );
buf ( n22693 , n22692 );
and ( n22694 , n22116 , n21178 );
and ( n22695 , n22693 , n22694 );
and ( n22696 , n21608 , n21990 );
and ( n22697 , n22694 , n22696 );
and ( n22698 , n22693 , n22696 );
or ( n22699 , n22695 , n22697 , n22698 );
and ( n22700 , n22691 , n22699 );
buf ( n22701 , n11378 );
buf ( n22702 , n22701 );
and ( n22703 , n22702 , n20877 );
and ( n22704 , n22589 , n20890 );
and ( n22705 , n22703 , n22704 );
not ( n22706 , n22586 );
and ( n22707 , n22704 , n22706 );
and ( n22708 , n22703 , n22706 );
or ( n22709 , n22705 , n22707 , n22708 );
and ( n22710 , n22699 , n22709 );
and ( n22711 , n22691 , n22709 );
or ( n22712 , n22700 , n22710 , n22711 );
and ( n22713 , n22351 , n20949 );
and ( n22714 , n22035 , n21296 );
and ( n22715 , n22713 , n22714 );
and ( n22716 , n21456 , n22337 );
and ( n22717 , n22714 , n22716 );
and ( n22718 , n22713 , n22716 );
or ( n22719 , n22715 , n22717 , n22718 );
and ( n22720 , n22542 , n20909 );
and ( n22721 , n21672 , n21827 );
and ( n22722 , n22720 , n22721 );
and ( n22723 , n21535 , n22172 );
and ( n22724 , n22721 , n22723 );
and ( n22725 , n22720 , n22723 );
or ( n22726 , n22722 , n22724 , n22725 );
and ( n22727 , n22719 , n22726 );
xor ( n22728 , n22558 , n22559 );
xor ( n22729 , n22728 , n22563 );
and ( n22730 , n22726 , n22729 );
and ( n22731 , n22719 , n22729 );
or ( n22732 , n22727 , n22730 , n22731 );
and ( n22733 , n22712 , n22732 );
xor ( n22734 , n22566 , n22573 );
xor ( n22735 , n22734 , n22575 );
and ( n22736 , n22732 , n22735 );
and ( n22737 , n22712 , n22735 );
or ( n22738 , n22733 , n22736 , n22737 );
xor ( n22739 , n22579 , n22580 );
xor ( n22740 , n22739 , n22582 );
xor ( n22741 , n22614 , n22615 );
xor ( n22742 , n22741 , n22617 );
and ( n22743 , n22740 , n22742 );
xor ( n22744 , n22567 , n22568 );
xor ( n22745 , n22744 , n22570 );
and ( n22746 , n22742 , n22745 );
and ( n22747 , n22740 , n22745 );
or ( n22748 , n22743 , n22746 , n22747 );
xor ( n22749 , n22620 , n22622 );
xor ( n22750 , n22749 , n22625 );
and ( n22751 , n22748 , n22750 );
xor ( n22752 , n22585 , n22595 );
xor ( n22753 , n22752 , n22598 );
and ( n22754 , n22750 , n22753 );
and ( n22755 , n22748 , n22753 );
or ( n22756 , n22751 , n22754 , n22755 );
and ( n22757 , n22738 , n22756 );
xor ( n22758 , n22628 , n22643 );
xor ( n22759 , n22758 , n22646 );
and ( n22760 , n22756 , n22759 );
and ( n22761 , n22738 , n22759 );
or ( n22762 , n22757 , n22760 , n22761 );
and ( n22763 , n22684 , n22762 );
xor ( n22764 , n22557 , n22607 );
xor ( n22765 , n22764 , n22610 );
and ( n22766 , n22762 , n22765 );
and ( n22767 , n22684 , n22765 );
or ( n22768 , n22763 , n22766 , n22767 );
xor ( n22769 , n22513 , n22515 );
xor ( n22770 , n22769 , n22518 );
and ( n22771 , n22768 , n22770 );
xor ( n22772 , n22613 , n22657 );
xor ( n22773 , n22772 , n22660 );
and ( n22774 , n22770 , n22773 );
and ( n22775 , n22768 , n22773 );
or ( n22776 , n22771 , n22774 , n22775 );
and ( n22777 , n22674 , n22776 );
xor ( n22778 , n22768 , n22770 );
xor ( n22779 , n22778 , n22773 );
and ( n22780 , n22542 , n20949 );
and ( n22781 , n21456 , n22562 );
and ( n22782 , n22780 , n22781 );
buf ( n22783 , n20232 );
buf ( n22784 , n22783 );
and ( n22785 , n21385 , n22784 );
and ( n22786 , n22781 , n22785 );
and ( n22787 , n22780 , n22785 );
or ( n22788 , n22782 , n22786 , n22787 );
and ( n22789 , n22354 , n21039 );
and ( n22790 , n22788 , n22789 );
and ( n22791 , n21914 , n21429 );
and ( n22792 , n22789 , n22791 );
and ( n22793 , n22788 , n22791 );
or ( n22794 , n22790 , n22792 , n22793 );
xor ( n22795 , n22629 , n22630 );
xor ( n22796 , n22795 , n22632 );
and ( n22797 , n22794 , n22796 );
xor ( n22798 , n22587 , n22590 );
xor ( n22799 , n22798 , n22592 );
and ( n22800 , n22796 , n22799 );
and ( n22801 , n22794 , n22799 );
or ( n22802 , n22797 , n22800 , n22801 );
and ( n22803 , n22702 , n20890 );
and ( n22804 , n22589 , n20909 );
and ( n22805 , n22803 , n22804 );
and ( n22806 , n21535 , n22337 );
and ( n22807 , n22804 , n22806 );
and ( n22808 , n22803 , n22806 );
or ( n22809 , n22805 , n22807 , n22808 );
and ( n22810 , n22116 , n21296 );
and ( n22811 , n21743 , n21827 );
and ( n22812 , n22810 , n22811 );
and ( n22813 , n21608 , n22172 );
and ( n22814 , n22811 , n22813 );
and ( n22815 , n22810 , n22813 );
or ( n22816 , n22812 , n22814 , n22815 );
and ( n22817 , n22809 , n22816 );
xor ( n22818 , n22713 , n22714 );
xor ( n22819 , n22818 , n22716 );
and ( n22820 , n22816 , n22819 );
and ( n22821 , n22809 , n22819 );
or ( n22822 , n22817 , n22820 , n22821 );
buf ( n22823 , n11708 );
buf ( n22824 , n22823 );
and ( n22825 , n22824 , n20877 );
and ( n22826 , n21914 , n21527 );
and ( n22827 , n22825 , n22826 );
and ( n22828 , n21836 , n21666 );
and ( n22829 , n22826 , n22828 );
and ( n22830 , n22825 , n22828 );
or ( n22831 , n22827 , n22829 , n22830 );
and ( n22832 , n21535 , n22562 );
buf ( n22833 , n22832 );
and ( n22834 , n22232 , n21178 );
and ( n22835 , n22833 , n22834 );
and ( n22836 , n21672 , n21990 );
and ( n22837 , n22834 , n22836 );
and ( n22838 , n22833 , n22836 );
or ( n22839 , n22835 , n22837 , n22838 );
and ( n22840 , n22831 , n22839 );
xor ( n22841 , n22720 , n22721 );
xor ( n22842 , n22841 , n22723 );
and ( n22843 , n22839 , n22842 );
and ( n22844 , n22831 , n22842 );
or ( n22845 , n22840 , n22843 , n22844 );
and ( n22846 , n22822 , n22845 );
xor ( n22847 , n22719 , n22726 );
xor ( n22848 , n22847 , n22729 );
and ( n22849 , n22845 , n22848 );
and ( n22850 , n22822 , n22848 );
or ( n22851 , n22846 , n22849 , n22850 );
and ( n22852 , n22802 , n22851 );
xor ( n22853 , n22635 , n22637 );
xor ( n22854 , n22853 , n22640 );
and ( n22855 , n22851 , n22854 );
and ( n22856 , n22802 , n22854 );
or ( n22857 , n22852 , n22855 , n22856 );
and ( n22858 , n22354 , n21085 );
and ( n22859 , n22035 , n21429 );
and ( n22860 , n22858 , n22859 );
not ( n22861 , n22692 );
and ( n22862 , n22859 , n22861 );
and ( n22863 , n22858 , n22861 );
or ( n22864 , n22860 , n22862 , n22863 );
xor ( n22865 , n22685 , n22686 );
xor ( n22866 , n22865 , n22688 );
and ( n22867 , n22864 , n22866 );
xor ( n22868 , n22693 , n22694 );
xor ( n22869 , n22868 , n22696 );
and ( n22870 , n22866 , n22869 );
and ( n22871 , n22864 , n22869 );
or ( n22872 , n22867 , n22870 , n22871 );
xor ( n22873 , n22691 , n22699 );
xor ( n22874 , n22873 , n22709 );
and ( n22875 , n22872 , n22874 );
xor ( n22876 , n22740 , n22742 );
xor ( n22877 , n22876 , n22745 );
and ( n22878 , n22874 , n22877 );
and ( n22879 , n22872 , n22877 );
or ( n22880 , n22875 , n22878 , n22879 );
xor ( n22881 , n22712 , n22732 );
xor ( n22882 , n22881 , n22735 );
and ( n22883 , n22880 , n22882 );
xor ( n22884 , n22748 , n22750 );
xor ( n22885 , n22884 , n22753 );
and ( n22886 , n22882 , n22885 );
and ( n22887 , n22880 , n22885 );
or ( n22888 , n22883 , n22886 , n22887 );
and ( n22889 , n22857 , n22888 );
xor ( n22890 , n22676 , n22678 );
xor ( n22891 , n22890 , n22681 );
and ( n22892 , n22888 , n22891 );
and ( n22893 , n22857 , n22891 );
or ( n22894 , n22889 , n22892 , n22893 );
xor ( n22895 , n22649 , n22651 );
xor ( n22896 , n22895 , n22654 );
and ( n22897 , n22894 , n22896 );
xor ( n22898 , n22684 , n22762 );
xor ( n22899 , n22898 , n22765 );
and ( n22900 , n22896 , n22899 );
and ( n22901 , n22894 , n22899 );
or ( n22902 , n22897 , n22900 , n22901 );
and ( n22903 , n22779 , n22902 );
xor ( n22904 , n22894 , n22896 );
xor ( n22905 , n22904 , n22899 );
and ( n22906 , n22824 , n20890 );
and ( n22907 , n22589 , n20949 );
and ( n22908 , n22906 , n22907 );
and ( n22909 , n21456 , n22784 );
and ( n22910 , n22907 , n22909 );
and ( n22911 , n22906 , n22909 );
or ( n22912 , n22908 , n22910 , n22911 );
and ( n22913 , n22351 , n21039 );
and ( n22914 , n22912 , n22913 );
xor ( n22915 , n22780 , n22781 );
xor ( n22916 , n22915 , n22785 );
and ( n22917 , n22913 , n22916 );
and ( n22918 , n22912 , n22916 );
or ( n22919 , n22914 , n22917 , n22918 );
xor ( n22920 , n22788 , n22789 );
xor ( n22921 , n22920 , n22791 );
and ( n22922 , n22919 , n22921 );
xor ( n22923 , n22703 , n22704 );
xor ( n22924 , n22923 , n22706 );
and ( n22925 , n22921 , n22924 );
and ( n22926 , n22919 , n22924 );
or ( n22927 , n22922 , n22925 , n22926 );
and ( n22928 , n22351 , n21085 );
and ( n22929 , n22354 , n21178 );
and ( n22930 , n22928 , n22929 );
and ( n22931 , n21743 , n21990 );
and ( n22932 , n22929 , n22931 );
and ( n22933 , n22928 , n22931 );
or ( n22934 , n22930 , n22932 , n22933 );
buf ( n22935 , n11835 );
buf ( n22936 , n22935 );
and ( n22937 , n22936 , n20877 );
and ( n22938 , n22035 , n21527 );
and ( n22939 , n22937 , n22938 );
not ( n22940 , n22832 );
and ( n22941 , n22938 , n22940 );
and ( n22942 , n22937 , n22940 );
or ( n22943 , n22939 , n22941 , n22942 );
and ( n22944 , n22934 , n22943 );
xor ( n22945 , n22810 , n22811 );
xor ( n22946 , n22945 , n22813 );
and ( n22947 , n22943 , n22946 );
and ( n22948 , n22934 , n22946 );
or ( n22949 , n22944 , n22947 , n22948 );
and ( n22950 , n22702 , n20909 );
and ( n22951 , n21836 , n21827 );
and ( n22952 , n22950 , n22951 );
and ( n22953 , n21608 , n22337 );
and ( n22954 , n22951 , n22953 );
and ( n22955 , n22950 , n22953 );
or ( n22956 , n22952 , n22954 , n22955 );
buf ( n22957 , n21385 );
buf ( n22958 , n22957 );
and ( n22959 , n22232 , n21296 );
and ( n22960 , n22958 , n22959 );
and ( n22961 , n21672 , n22172 );
and ( n22962 , n22959 , n22961 );
and ( n22963 , n22958 , n22961 );
or ( n22964 , n22960 , n22962 , n22963 );
and ( n22965 , n22956 , n22964 );
xor ( n22966 , n22803 , n22804 );
xor ( n22967 , n22966 , n22806 );
and ( n22968 , n22964 , n22967 );
and ( n22969 , n22956 , n22967 );
or ( n22970 , n22965 , n22968 , n22969 );
and ( n22971 , n22949 , n22970 );
xor ( n22972 , n22809 , n22816 );
xor ( n22973 , n22972 , n22819 );
and ( n22974 , n22970 , n22973 );
and ( n22975 , n22949 , n22973 );
or ( n22976 , n22971 , n22974 , n22975 );
and ( n22977 , n22927 , n22976 );
xor ( n22978 , n22794 , n22796 );
xor ( n22979 , n22978 , n22799 );
and ( n22980 , n22976 , n22979 );
and ( n22981 , n22927 , n22979 );
or ( n22982 , n22977 , n22980 , n22981 );
and ( n22983 , n22702 , n20949 );
and ( n22984 , n21608 , n22562 );
and ( n22985 , n22983 , n22984 );
buf ( n22986 , n20235 );
buf ( n22987 , n22986 );
and ( n22988 , n21456 , n22987 );
and ( n22989 , n22984 , n22988 );
and ( n22990 , n22983 , n22988 );
or ( n22991 , n22985 , n22989 , n22990 );
and ( n22992 , n22116 , n21429 );
and ( n22993 , n22991 , n22992 );
and ( n22994 , n21914 , n21666 );
and ( n22995 , n22992 , n22994 );
and ( n22996 , n22991 , n22994 );
or ( n22997 , n22993 , n22995 , n22996 );
xor ( n22998 , n22825 , n22826 );
xor ( n22999 , n22998 , n22828 );
and ( n23000 , n22997 , n22999 );
xor ( n23001 , n22858 , n22859 );
xor ( n23002 , n23001 , n22861 );
and ( n23003 , n22999 , n23002 );
and ( n23004 , n22997 , n23002 );
or ( n23005 , n23000 , n23003 , n23004 );
xor ( n23006 , n22831 , n22839 );
xor ( n23007 , n23006 , n22842 );
and ( n23008 , n23005 , n23007 );
xor ( n23009 , n22864 , n22866 );
xor ( n23010 , n23009 , n22869 );
and ( n23011 , n23007 , n23010 );
and ( n23012 , n23005 , n23010 );
or ( n23013 , n23008 , n23011 , n23012 );
xor ( n23014 , n22822 , n22845 );
xor ( n23015 , n23014 , n22848 );
and ( n23016 , n23013 , n23015 );
xor ( n23017 , n22872 , n22874 );
xor ( n23018 , n23017 , n22877 );
and ( n23019 , n23015 , n23018 );
and ( n23020 , n23013 , n23018 );
or ( n23021 , n23016 , n23019 , n23020 );
and ( n23022 , n22982 , n23021 );
xor ( n23023 , n22802 , n22851 );
xor ( n23024 , n23023 , n22854 );
and ( n23025 , n23021 , n23024 );
and ( n23026 , n22982 , n23024 );
or ( n23027 , n23022 , n23025 , n23026 );
xor ( n23028 , n22738 , n22756 );
xor ( n23029 , n23028 , n22759 );
and ( n23030 , n23027 , n23029 );
xor ( n23031 , n22857 , n22888 );
xor ( n23032 , n23031 , n22891 );
and ( n23033 , n23029 , n23032 );
and ( n23034 , n23027 , n23032 );
or ( n23035 , n23030 , n23033 , n23034 );
and ( n23036 , n22905 , n23035 );
xor ( n23037 , n23027 , n23029 );
xor ( n23038 , n23037 , n23032 );
and ( n23039 , n22936 , n20890 );
and ( n23040 , n22824 , n20909 );
and ( n23041 , n23039 , n23040 );
and ( n23042 , n21914 , n21827 );
and ( n23043 , n23040 , n23042 );
and ( n23044 , n23039 , n23042 );
or ( n23045 , n23041 , n23043 , n23044 );
and ( n23046 , n21672 , n22337 );
and ( n23047 , n21535 , n22784 );
and ( n23048 , n23046 , n23047 );
not ( n23049 , n22957 );
and ( n23050 , n23047 , n23049 );
and ( n23051 , n23046 , n23049 );
or ( n23052 , n23048 , n23050 , n23051 );
and ( n23053 , n23045 , n23052 );
and ( n23054 , n22542 , n21039 );
and ( n23055 , n23052 , n23054 );
and ( n23056 , n23045 , n23054 );
or ( n23057 , n23053 , n23055 , n23056 );
and ( n23058 , n22354 , n21296 );
and ( n23059 , n22035 , n21666 );
and ( n23060 , n23058 , n23059 );
and ( n23061 , n21743 , n22172 );
and ( n23062 , n23059 , n23061 );
and ( n23063 , n23058 , n23061 );
or ( n23064 , n23060 , n23062 , n23063 );
xor ( n23065 , n22906 , n22907 );
xor ( n23066 , n23065 , n22909 );
and ( n23067 , n23064 , n23066 );
xor ( n23068 , n22958 , n22959 );
xor ( n23069 , n23068 , n22961 );
and ( n23070 , n23066 , n23069 );
and ( n23071 , n23064 , n23069 );
or ( n23072 , n23067 , n23070 , n23071 );
and ( n23073 , n23057 , n23072 );
xor ( n23074 , n22833 , n22834 );
xor ( n23075 , n23074 , n22836 );
and ( n23076 , n23072 , n23075 );
and ( n23077 , n23057 , n23075 );
or ( n23078 , n23073 , n23076 , n23077 );
and ( n23079 , n22542 , n21085 );
and ( n23080 , n22351 , n21178 );
and ( n23081 , n23079 , n23080 );
and ( n23082 , n21836 , n21990 );
and ( n23083 , n23080 , n23082 );
and ( n23084 , n23079 , n23082 );
or ( n23085 , n23081 , n23083 , n23084 );
and ( n23086 , n21535 , n22987 );
buf ( n23087 , n23086 );
buf ( n23088 , n12120 );
buf ( n23089 , n23088 );
and ( n23090 , n23089 , n20877 );
and ( n23091 , n23087 , n23090 );
and ( n23092 , n22116 , n21527 );
and ( n23093 , n23090 , n23092 );
and ( n23094 , n23087 , n23092 );
or ( n23095 , n23091 , n23093 , n23094 );
and ( n23096 , n23085 , n23095 );
xor ( n23097 , n22950 , n22951 );
xor ( n23098 , n23097 , n22953 );
and ( n23099 , n23095 , n23098 );
and ( n23100 , n23085 , n23098 );
or ( n23101 , n23096 , n23099 , n23100 );
xor ( n23102 , n22912 , n22913 );
xor ( n23103 , n23102 , n22916 );
and ( n23104 , n23101 , n23103 );
xor ( n23105 , n22956 , n22964 );
xor ( n23106 , n23105 , n22967 );
and ( n23107 , n23103 , n23106 );
and ( n23108 , n23101 , n23106 );
or ( n23109 , n23104 , n23107 , n23108 );
and ( n23110 , n23078 , n23109 );
xor ( n23111 , n22919 , n22921 );
xor ( n23112 , n23111 , n22924 );
and ( n23113 , n23109 , n23112 );
and ( n23114 , n23078 , n23112 );
or ( n23115 , n23110 , n23113 , n23114 );
and ( n23116 , n22589 , n21039 );
and ( n23117 , n22232 , n21429 );
and ( n23118 , n23116 , n23117 );
xor ( n23119 , n22983 , n22984 );
xor ( n23120 , n23119 , n22988 );
and ( n23121 , n23117 , n23120 );
and ( n23122 , n23116 , n23120 );
or ( n23123 , n23118 , n23121 , n23122 );
xor ( n23124 , n22928 , n22929 );
xor ( n23125 , n23124 , n22931 );
and ( n23126 , n23123 , n23125 );
xor ( n23127 , n22937 , n22938 );
xor ( n23128 , n23127 , n22940 );
and ( n23129 , n23125 , n23128 );
and ( n23130 , n23123 , n23128 );
or ( n23131 , n23126 , n23129 , n23130 );
xor ( n23132 , n22934 , n22943 );
xor ( n23133 , n23132 , n22946 );
and ( n23134 , n23131 , n23133 );
xor ( n23135 , n22997 , n22999 );
xor ( n23136 , n23135 , n23002 );
and ( n23137 , n23133 , n23136 );
and ( n23138 , n23131 , n23136 );
or ( n23139 , n23134 , n23137 , n23138 );
xor ( n23140 , n22949 , n22970 );
xor ( n23141 , n23140 , n22973 );
and ( n23142 , n23139 , n23141 );
xor ( n23143 , n23005 , n23007 );
xor ( n23144 , n23143 , n23010 );
and ( n23145 , n23141 , n23144 );
and ( n23146 , n23139 , n23144 );
or ( n23147 , n23142 , n23145 , n23146 );
and ( n23148 , n23115 , n23147 );
xor ( n23149 , n22927 , n22976 );
xor ( n23150 , n23149 , n22979 );
and ( n23151 , n23147 , n23150 );
and ( n23152 , n23115 , n23150 );
or ( n23153 , n23148 , n23151 , n23152 );
xor ( n23154 , n22880 , n22882 );
xor ( n23155 , n23154 , n22885 );
and ( n23156 , n23153 , n23155 );
xor ( n23157 , n22982 , n23021 );
xor ( n23158 , n23157 , n23024 );
and ( n23159 , n23155 , n23158 );
and ( n23160 , n23153 , n23158 );
or ( n23161 , n23156 , n23159 , n23160 );
and ( n23162 , n23038 , n23161 );
xor ( n23163 , n23153 , n23155 );
xor ( n23164 , n23163 , n23158 );
and ( n23165 , n22824 , n20949 );
and ( n23166 , n21672 , n22562 );
and ( n23167 , n23165 , n23166 );
and ( n23168 , n21608 , n22784 );
and ( n23169 , n23166 , n23168 );
and ( n23170 , n23165 , n23168 );
or ( n23171 , n23167 , n23169 , n23170 );
and ( n23172 , n23089 , n20890 );
and ( n23173 , n22936 , n20909 );
and ( n23174 , n23172 , n23173 );
and ( n23175 , n21743 , n22337 );
and ( n23176 , n23173 , n23175 );
and ( n23177 , n23172 , n23175 );
or ( n23178 , n23174 , n23176 , n23177 );
and ( n23179 , n23171 , n23178 );
buf ( n23180 , n21456 );
buf ( n23181 , n23180 );
and ( n23182 , n22351 , n21296 );
and ( n23183 , n23181 , n23182 );
and ( n23184 , n21836 , n22172 );
and ( n23185 , n23182 , n23184 );
and ( n23186 , n23181 , n23184 );
or ( n23187 , n23183 , n23185 , n23186 );
and ( n23188 , n23178 , n23187 );
and ( n23189 , n23171 , n23187 );
or ( n23190 , n23179 , n23188 , n23189 );
xor ( n23191 , n23058 , n23059 );
xor ( n23192 , n23191 , n23061 );
xor ( n23193 , n23039 , n23040 );
xor ( n23194 , n23193 , n23042 );
and ( n23195 , n23192 , n23194 );
xor ( n23196 , n23046 , n23047 );
xor ( n23197 , n23196 , n23049 );
and ( n23198 , n23194 , n23197 );
and ( n23199 , n23192 , n23197 );
or ( n23200 , n23195 , n23198 , n23199 );
and ( n23201 , n23190 , n23200 );
xor ( n23202 , n22991 , n22992 );
xor ( n23203 , n23202 , n22994 );
and ( n23204 , n23200 , n23203 );
and ( n23205 , n23190 , n23203 );
or ( n23206 , n23201 , n23204 , n23205 );
and ( n23207 , n22542 , n21178 );
and ( n23208 , n22232 , n21527 );
and ( n23209 , n23207 , n23208 );
and ( n23210 , n21914 , n21990 );
and ( n23211 , n23208 , n23210 );
and ( n23212 , n23207 , n23210 );
or ( n23213 , n23209 , n23211 , n23212 );
buf ( n23214 , n12619 );
buf ( n23215 , n23214 );
and ( n23216 , n23215 , n20877 );
and ( n23217 , n22116 , n21666 );
and ( n23218 , n23216 , n23217 );
and ( n23219 , n22035 , n21827 );
and ( n23220 , n23217 , n23219 );
and ( n23221 , n23216 , n23219 );
or ( n23222 , n23218 , n23220 , n23221 );
and ( n23223 , n23213 , n23222 );
xor ( n23224 , n23079 , n23080 );
xor ( n23225 , n23224 , n23082 );
and ( n23226 , n23222 , n23225 );
and ( n23227 , n23213 , n23225 );
or ( n23228 , n23223 , n23226 , n23227 );
xor ( n23229 , n23045 , n23052 );
xor ( n23230 , n23229 , n23054 );
and ( n23231 , n23228 , n23230 );
xor ( n23232 , n23085 , n23095 );
xor ( n23233 , n23232 , n23098 );
and ( n23234 , n23230 , n23233 );
and ( n23235 , n23228 , n23233 );
or ( n23236 , n23231 , n23234 , n23235 );
and ( n23237 , n23206 , n23236 );
xor ( n23238 , n23057 , n23072 );
xor ( n23239 , n23238 , n23075 );
and ( n23240 , n23236 , n23239 );
and ( n23241 , n23206 , n23239 );
or ( n23242 , n23237 , n23240 , n23241 );
xor ( n23243 , n23078 , n23109 );
xor ( n23244 , n23243 , n23112 );
and ( n23245 , n23242 , n23244 );
xor ( n23246 , n23139 , n23141 );
xor ( n23247 , n23246 , n23144 );
and ( n23248 , n23244 , n23247 );
and ( n23249 , n23242 , n23247 );
or ( n23250 , n23245 , n23248 , n23249 );
xor ( n23251 , n23013 , n23015 );
xor ( n23252 , n23251 , n23018 );
and ( n23253 , n23250 , n23252 );
xor ( n23254 , n23115 , n23147 );
xor ( n23255 , n23254 , n23150 );
and ( n23256 , n23252 , n23255 );
and ( n23257 , n23250 , n23255 );
or ( n23258 , n23253 , n23256 , n23257 );
and ( n23259 , n23164 , n23258 );
xor ( n23260 , n23250 , n23252 );
xor ( n23261 , n23260 , n23255 );
and ( n23262 , n22589 , n21085 );
and ( n23263 , n22354 , n21429 );
and ( n23264 , n23262 , n23263 );
not ( n23265 , n23086 );
and ( n23266 , n23263 , n23265 );
and ( n23267 , n23262 , n23265 );
or ( n23268 , n23264 , n23266 , n23267 );
xor ( n23269 , n23087 , n23090 );
xor ( n23270 , n23269 , n23092 );
and ( n23271 , n23268 , n23270 );
xor ( n23272 , n23116 , n23117 );
xor ( n23273 , n23272 , n23120 );
and ( n23274 , n23270 , n23273 );
and ( n23275 , n23268 , n23273 );
or ( n23276 , n23271 , n23274 , n23275 );
xor ( n23277 , n23064 , n23066 );
xor ( n23278 , n23277 , n23069 );
and ( n23279 , n23276 , n23278 );
xor ( n23280 , n23123 , n23125 );
xor ( n23281 , n23280 , n23128 );
and ( n23282 , n23278 , n23281 );
and ( n23283 , n23276 , n23281 );
or ( n23284 , n23279 , n23282 , n23283 );
xor ( n23285 , n23101 , n23103 );
xor ( n23286 , n23285 , n23106 );
and ( n23287 , n23284 , n23286 );
xor ( n23288 , n23131 , n23133 );
xor ( n23289 , n23288 , n23136 );
and ( n23290 , n23286 , n23289 );
and ( n23291 , n23284 , n23289 );
or ( n23292 , n23287 , n23290 , n23291 );
and ( n23293 , n22542 , n21296 );
and ( n23294 , n21914 , n22172 );
and ( n23295 , n23293 , n23294 );
and ( n23296 , n21836 , n22337 );
and ( n23297 , n23294 , n23296 );
and ( n23298 , n23293 , n23296 );
or ( n23299 , n23295 , n23297 , n23298 );
and ( n23300 , n22116 , n21827 );
and ( n23301 , n21672 , n22784 );
and ( n23302 , n23300 , n23301 );
and ( n23303 , n21608 , n22987 );
and ( n23304 , n23301 , n23303 );
and ( n23305 , n23300 , n23303 );
or ( n23306 , n23302 , n23304 , n23305 );
and ( n23307 , n23299 , n23306 );
and ( n23308 , n23215 , n20890 );
and ( n23309 , n23089 , n20909 );
and ( n23310 , n23308 , n23309 );
not ( n23311 , n23180 );
and ( n23312 , n23309 , n23311 );
and ( n23313 , n23308 , n23311 );
or ( n23314 , n23310 , n23312 , n23313 );
and ( n23315 , n23306 , n23314 );
and ( n23316 , n23299 , n23314 );
or ( n23317 , n23307 , n23315 , n23316 );
and ( n23318 , n22936 , n20949 );
and ( n23319 , n21743 , n22562 );
and ( n23320 , n23318 , n23319 );
buf ( n23321 , n20238 );
buf ( n23322 , n23321 );
and ( n23323 , n21535 , n23322 );
and ( n23324 , n23319 , n23323 );
and ( n23325 , n23318 , n23323 );
or ( n23326 , n23320 , n23324 , n23325 );
and ( n23327 , n22702 , n21039 );
and ( n23328 , n23326 , n23327 );
xor ( n23329 , n23165 , n23166 );
xor ( n23330 , n23329 , n23168 );
and ( n23331 , n23327 , n23330 );
and ( n23332 , n23326 , n23330 );
or ( n23333 , n23328 , n23331 , n23332 );
and ( n23334 , n23317 , n23333 );
buf ( n23335 , n12668 );
buf ( n23336 , n23335 );
and ( n23337 , n23336 , n20877 );
and ( n23338 , n22232 , n21666 );
and ( n23339 , n23337 , n23338 );
and ( n23340 , n22035 , n21990 );
and ( n23341 , n23338 , n23340 );
and ( n23342 , n23337 , n23340 );
or ( n23343 , n23339 , n23341 , n23342 );
xor ( n23344 , n23172 , n23173 );
xor ( n23345 , n23344 , n23175 );
and ( n23346 , n23343 , n23345 );
xor ( n23347 , n23181 , n23182 );
xor ( n23348 , n23347 , n23184 );
and ( n23349 , n23345 , n23348 );
and ( n23350 , n23343 , n23348 );
or ( n23351 , n23346 , n23349 , n23350 );
and ( n23352 , n23333 , n23351 );
and ( n23353 , n23317 , n23351 );
or ( n23354 , n23334 , n23352 , n23353 );
and ( n23355 , n21608 , n23322 );
buf ( n23356 , n23355 );
and ( n23357 , n22589 , n21178 );
and ( n23358 , n23356 , n23357 );
and ( n23359 , n22354 , n21527 );
and ( n23360 , n23357 , n23359 );
and ( n23361 , n23356 , n23359 );
or ( n23362 , n23358 , n23360 , n23361 );
and ( n23363 , n23089 , n20949 );
and ( n23364 , n21836 , n22562 );
and ( n23365 , n23363 , n23364 );
and ( n23366 , n21672 , n22987 );
and ( n23367 , n23364 , n23366 );
and ( n23368 , n23363 , n23366 );
or ( n23369 , n23365 , n23367 , n23368 );
and ( n23370 , n22824 , n21039 );
and ( n23371 , n23369 , n23370 );
and ( n23372 , n22702 , n21085 );
and ( n23373 , n23370 , n23372 );
and ( n23374 , n23369 , n23372 );
or ( n23375 , n23371 , n23373 , n23374 );
and ( n23376 , n23362 , n23375 );
xor ( n23377 , n23262 , n23263 );
xor ( n23378 , n23377 , n23265 );
and ( n23379 , n23375 , n23378 );
and ( n23380 , n23362 , n23378 );
or ( n23381 , n23376 , n23379 , n23380 );
xor ( n23382 , n23171 , n23178 );
xor ( n23383 , n23382 , n23187 );
and ( n23384 , n23381 , n23383 );
xor ( n23385 , n23213 , n23222 );
xor ( n23386 , n23385 , n23225 );
and ( n23387 , n23383 , n23386 );
and ( n23388 , n23381 , n23386 );
or ( n23389 , n23384 , n23387 , n23388 );
and ( n23390 , n23354 , n23389 );
xor ( n23391 , n23190 , n23200 );
xor ( n23392 , n23391 , n23203 );
and ( n23393 , n23389 , n23392 );
and ( n23394 , n23354 , n23392 );
or ( n23395 , n23390 , n23393 , n23394 );
xor ( n23396 , n23206 , n23236 );
xor ( n23397 , n23396 , n23239 );
and ( n23398 , n23395 , n23397 );
xor ( n23399 , n23284 , n23286 );
xor ( n23400 , n23399 , n23289 );
and ( n23401 , n23397 , n23400 );
and ( n23402 , n23395 , n23400 );
or ( n23403 , n23398 , n23401 , n23402 );
and ( n23404 , n23292 , n23403 );
xor ( n23405 , n23242 , n23244 );
xor ( n23406 , n23405 , n23247 );
and ( n23407 , n23403 , n23406 );
and ( n23408 , n23292 , n23406 );
or ( n23409 , n23404 , n23407 , n23408 );
and ( n23410 , n23261 , n23409 );
xor ( n23411 , n23292 , n23403 );
xor ( n23412 , n23411 , n23406 );
xor ( n23413 , n23207 , n23208 );
xor ( n23414 , n23413 , n23210 );
xor ( n23415 , n23216 , n23217 );
xor ( n23416 , n23415 , n23219 );
and ( n23417 , n23414 , n23416 );
xor ( n23418 , n23326 , n23327 );
xor ( n23419 , n23418 , n23330 );
and ( n23420 , n23416 , n23419 );
and ( n23421 , n23414 , n23419 );
or ( n23422 , n23417 , n23420 , n23421 );
xor ( n23423 , n23192 , n23194 );
xor ( n23424 , n23423 , n23197 );
and ( n23425 , n23422 , n23424 );
xor ( n23426 , n23268 , n23270 );
xor ( n23427 , n23426 , n23273 );
and ( n23428 , n23424 , n23427 );
and ( n23429 , n23422 , n23427 );
or ( n23430 , n23425 , n23428 , n23429 );
xor ( n23431 , n23228 , n23230 );
xor ( n23432 , n23431 , n23233 );
and ( n23433 , n23430 , n23432 );
xor ( n23434 , n23276 , n23278 );
xor ( n23435 , n23434 , n23281 );
and ( n23436 , n23432 , n23435 );
and ( n23437 , n23430 , n23435 );
or ( n23438 , n23433 , n23436 , n23437 );
and ( n23439 , n22589 , n21296 );
and ( n23440 , n22354 , n21666 );
and ( n23441 , n23439 , n23440 );
and ( n23442 , n22035 , n22172 );
and ( n23443 , n23440 , n23442 );
and ( n23444 , n23439 , n23442 );
or ( n23445 , n23441 , n23443 , n23444 );
xor ( n23446 , n23293 , n23294 );
xor ( n23447 , n23446 , n23296 );
and ( n23448 , n23445 , n23447 );
xor ( n23449 , n23300 , n23301 );
xor ( n23450 , n23449 , n23303 );
and ( n23451 , n23447 , n23450 );
and ( n23452 , n23445 , n23450 );
or ( n23453 , n23448 , n23451 , n23452 );
buf ( n23454 , n21535 );
buf ( n23455 , n23454 );
and ( n23456 , n23215 , n20909 );
and ( n23457 , n23455 , n23456 );
and ( n23458 , n22232 , n21827 );
and ( n23459 , n23456 , n23458 );
and ( n23460 , n23455 , n23458 );
or ( n23461 , n23457 , n23459 , n23460 );
and ( n23462 , n22351 , n21429 );
and ( n23463 , n23461 , n23462 );
xor ( n23464 , n23318 , n23319 );
xor ( n23465 , n23464 , n23323 );
and ( n23466 , n23462 , n23465 );
and ( n23467 , n23461 , n23465 );
or ( n23468 , n23463 , n23466 , n23467 );
and ( n23469 , n23453 , n23468 );
xor ( n23470 , n23299 , n23306 );
xor ( n23471 , n23470 , n23314 );
and ( n23472 , n23468 , n23471 );
and ( n23473 , n23453 , n23471 );
or ( n23474 , n23469 , n23472 , n23473 );
and ( n23475 , n23336 , n20890 );
and ( n23476 , n21914 , n22337 );
and ( n23477 , n23475 , n23476 );
and ( n23478 , n21743 , n22784 );
and ( n23479 , n23476 , n23478 );
and ( n23480 , n23475 , n23478 );
or ( n23481 , n23477 , n23479 , n23480 );
buf ( n23482 , n12963 );
buf ( n23483 , n23482 );
and ( n23484 , n23483 , n20877 );
and ( n23485 , n22351 , n21527 );
and ( n23486 , n23484 , n23485 );
not ( n23487 , n23355 );
and ( n23488 , n23485 , n23487 );
and ( n23489 , n23484 , n23487 );
or ( n23490 , n23486 , n23488 , n23489 );
and ( n23491 , n23481 , n23490 );
xor ( n23492 , n23308 , n23309 );
xor ( n23493 , n23492 , n23311 );
and ( n23494 , n23490 , n23493 );
and ( n23495 , n23481 , n23493 );
or ( n23496 , n23491 , n23494 , n23495 );
and ( n23497 , n22824 , n21085 );
and ( n23498 , n22702 , n21178 );
and ( n23499 , n23497 , n23498 );
and ( n23500 , n22116 , n21990 );
and ( n23501 , n23498 , n23500 );
and ( n23502 , n23497 , n23500 );
or ( n23503 , n23499 , n23501 , n23502 );
and ( n23504 , n23215 , n20949 );
and ( n23505 , n21743 , n22987 );
and ( n23506 , n23504 , n23505 );
buf ( n23507 , n20241 );
buf ( n23508 , n23507 );
and ( n23509 , n21608 , n23508 );
and ( n23510 , n23505 , n23509 );
and ( n23511 , n23504 , n23509 );
or ( n23512 , n23506 , n23510 , n23511 );
and ( n23513 , n21914 , n22562 );
and ( n23514 , n21672 , n23322 );
and ( n23515 , n23513 , n23514 );
not ( n23516 , n23454 );
and ( n23517 , n23514 , n23516 );
and ( n23518 , n23513 , n23516 );
or ( n23519 , n23515 , n23517 , n23518 );
and ( n23520 , n23512 , n23519 );
and ( n23521 , n22542 , n21429 );
and ( n23522 , n23519 , n23521 );
and ( n23523 , n23512 , n23521 );
or ( n23524 , n23520 , n23522 , n23523 );
and ( n23525 , n23503 , n23524 );
xor ( n23526 , n23356 , n23357 );
xor ( n23527 , n23526 , n23359 );
and ( n23528 , n23524 , n23527 );
and ( n23529 , n23503 , n23527 );
or ( n23530 , n23525 , n23528 , n23529 );
and ( n23531 , n23496 , n23530 );
xor ( n23532 , n23343 , n23345 );
xor ( n23533 , n23532 , n23348 );
and ( n23534 , n23530 , n23533 );
and ( n23535 , n23496 , n23533 );
or ( n23536 , n23531 , n23534 , n23535 );
and ( n23537 , n23474 , n23536 );
xor ( n23538 , n23317 , n23333 );
xor ( n23539 , n23538 , n23351 );
and ( n23540 , n23536 , n23539 );
and ( n23541 , n23474 , n23539 );
or ( n23542 , n23537 , n23540 , n23541 );
and ( n23543 , n23483 , n20890 );
and ( n23544 , n23336 , n20909 );
and ( n23545 , n23543 , n23544 );
and ( n23546 , n22116 , n22172 );
and ( n23547 , n23544 , n23546 );
and ( n23548 , n23543 , n23546 );
or ( n23549 , n23545 , n23547 , n23548 );
and ( n23550 , n22936 , n21039 );
and ( n23551 , n23549 , n23550 );
xor ( n23552 , n23363 , n23364 );
xor ( n23553 , n23552 , n23366 );
and ( n23554 , n23550 , n23553 );
and ( n23555 , n23549 , n23553 );
or ( n23556 , n23551 , n23554 , n23555 );
xor ( n23557 , n23337 , n23338 );
xor ( n23558 , n23557 , n23340 );
and ( n23559 , n23556 , n23558 );
xor ( n23560 , n23369 , n23370 );
xor ( n23561 , n23560 , n23372 );
and ( n23562 , n23558 , n23561 );
and ( n23563 , n23556 , n23561 );
or ( n23564 , n23559 , n23562 , n23563 );
xor ( n23565 , n23362 , n23375 );
xor ( n23566 , n23565 , n23378 );
and ( n23567 , n23564 , n23566 );
xor ( n23568 , n23414 , n23416 );
xor ( n23569 , n23568 , n23419 );
and ( n23570 , n23566 , n23569 );
and ( n23571 , n23564 , n23569 );
or ( n23572 , n23567 , n23570 , n23571 );
xor ( n23573 , n23381 , n23383 );
xor ( n23574 , n23573 , n23386 );
and ( n23575 , n23572 , n23574 );
xor ( n23576 , n23422 , n23424 );
xor ( n23577 , n23576 , n23427 );
and ( n23578 , n23574 , n23577 );
and ( n23579 , n23572 , n23577 );
or ( n23580 , n23575 , n23578 , n23579 );
and ( n23581 , n23542 , n23580 );
xor ( n23582 , n23354 , n23389 );
xor ( n23583 , n23582 , n23392 );
and ( n23584 , n23580 , n23583 );
and ( n23585 , n23542 , n23583 );
or ( n23586 , n23581 , n23584 , n23585 );
and ( n23587 , n23438 , n23586 );
xor ( n23588 , n23395 , n23397 );
xor ( n23589 , n23588 , n23400 );
and ( n23590 , n23586 , n23589 );
and ( n23591 , n23438 , n23589 );
or ( n23592 , n23587 , n23590 , n23591 );
and ( n23593 , n23412 , n23592 );
xor ( n23594 , n23438 , n23586 );
xor ( n23595 , n23594 , n23589 );
and ( n23596 , n23089 , n21039 );
and ( n23597 , n22824 , n21178 );
and ( n23598 , n23596 , n23597 );
and ( n23599 , n22542 , n21527 );
and ( n23600 , n23597 , n23599 );
and ( n23601 , n23596 , n23599 );
or ( n23602 , n23598 , n23600 , n23601 );
xor ( n23603 , n23497 , n23498 );
xor ( n23604 , n23603 , n23500 );
and ( n23605 , n23602 , n23604 );
xor ( n23606 , n23484 , n23485 );
xor ( n23607 , n23606 , n23487 );
and ( n23608 , n23604 , n23607 );
and ( n23609 , n23602 , n23607 );
or ( n23610 , n23605 , n23608 , n23609 );
xor ( n23611 , n23481 , n23490 );
xor ( n23612 , n23611 , n23493 );
and ( n23613 , n23610 , n23612 );
xor ( n23614 , n23445 , n23447 );
xor ( n23615 , n23614 , n23450 );
and ( n23616 , n23612 , n23615 );
and ( n23617 , n23610 , n23615 );
or ( n23618 , n23613 , n23616 , n23617 );
buf ( n23619 , n13411 );
buf ( n23620 , n23619 );
and ( n23621 , n23620 , n20877 );
and ( n23622 , n22351 , n21666 );
and ( n23623 , n23621 , n23622 );
and ( n23624 , n22232 , n21990 );
and ( n23625 , n23622 , n23624 );
and ( n23626 , n23621 , n23624 );
or ( n23627 , n23623 , n23625 , n23626 );
and ( n23628 , n21672 , n23508 );
buf ( n23629 , n23628 );
and ( n23630 , n22354 , n21827 );
and ( n23631 , n23629 , n23630 );
and ( n23632 , n21836 , n22784 );
and ( n23633 , n23630 , n23632 );
and ( n23634 , n23629 , n23632 );
or ( n23635 , n23631 , n23633 , n23634 );
and ( n23636 , n23627 , n23635 );
xor ( n23637 , n23475 , n23476 );
xor ( n23638 , n23637 , n23478 );
and ( n23639 , n23635 , n23638 );
and ( n23640 , n23627 , n23638 );
or ( n23641 , n23636 , n23639 , n23640 );
and ( n23642 , n22936 , n21085 );
and ( n23643 , n22702 , n21296 );
and ( n23644 , n23642 , n23643 );
and ( n23645 , n22035 , n22337 );
and ( n23646 , n23643 , n23645 );
and ( n23647 , n23642 , n23645 );
or ( n23648 , n23644 , n23646 , n23647 );
xor ( n23649 , n23439 , n23440 );
xor ( n23650 , n23649 , n23442 );
and ( n23651 , n23648 , n23650 );
xor ( n23652 , n23455 , n23456 );
xor ( n23653 , n23652 , n23458 );
and ( n23654 , n23650 , n23653 );
and ( n23655 , n23648 , n23653 );
or ( n23656 , n23651 , n23654 , n23655 );
and ( n23657 , n23641 , n23656 );
xor ( n23658 , n23461 , n23462 );
xor ( n23659 , n23658 , n23465 );
and ( n23660 , n23656 , n23659 );
and ( n23661 , n23641 , n23659 );
or ( n23662 , n23657 , n23660 , n23661 );
and ( n23663 , n23618 , n23662 );
xor ( n23664 , n23453 , n23468 );
xor ( n23665 , n23664 , n23471 );
and ( n23666 , n23662 , n23665 );
and ( n23667 , n23618 , n23665 );
or ( n23668 , n23663 , n23666 , n23667 );
xor ( n23669 , n23474 , n23536 );
xor ( n23670 , n23669 , n23539 );
and ( n23671 , n23668 , n23670 );
xor ( n23672 , n23572 , n23574 );
xor ( n23673 , n23672 , n23577 );
and ( n23674 , n23670 , n23673 );
and ( n23675 , n23668 , n23673 );
or ( n23676 , n23671 , n23674 , n23675 );
xor ( n23677 , n23430 , n23432 );
xor ( n23678 , n23677 , n23435 );
and ( n23679 , n23676 , n23678 );
xor ( n23680 , n23542 , n23580 );
xor ( n23681 , n23680 , n23583 );
and ( n23682 , n23678 , n23681 );
and ( n23683 , n23676 , n23681 );
or ( n23684 , n23679 , n23682 , n23683 );
and ( n23685 , n23595 , n23684 );
xor ( n23686 , n23676 , n23678 );
xor ( n23687 , n23686 , n23681 );
and ( n23688 , n23483 , n20949 );
and ( n23689 , n21836 , n23322 );
and ( n23690 , n23688 , n23689 );
and ( n23691 , n21743 , n23508 );
and ( n23692 , n23689 , n23691 );
and ( n23693 , n23688 , n23691 );
or ( n23694 , n23690 , n23692 , n23693 );
and ( n23695 , n23215 , n21039 );
and ( n23696 , n23694 , n23695 );
and ( n23697 , n23089 , n21085 );
and ( n23698 , n23695 , n23697 );
and ( n23699 , n23694 , n23697 );
or ( n23700 , n23696 , n23698 , n23699 );
xor ( n23701 , n23621 , n23622 );
xor ( n23702 , n23701 , n23624 );
and ( n23703 , n23700 , n23702 );
xor ( n23704 , n23596 , n23597 );
xor ( n23705 , n23704 , n23599 );
and ( n23706 , n23702 , n23705 );
and ( n23707 , n23700 , n23705 );
or ( n23708 , n23703 , n23706 , n23707 );
xor ( n23709 , n23627 , n23635 );
xor ( n23710 , n23709 , n23638 );
and ( n23711 , n23708 , n23710 );
xor ( n23712 , n23648 , n23650 );
xor ( n23713 , n23712 , n23653 );
and ( n23714 , n23710 , n23713 );
and ( n23715 , n23708 , n23713 );
or ( n23716 , n23711 , n23714 , n23715 );
xor ( n23717 , n23556 , n23558 );
xor ( n23718 , n23717 , n23561 );
and ( n23719 , n23716 , n23718 );
xor ( n23720 , n23641 , n23656 );
xor ( n23721 , n23720 , n23659 );
and ( n23722 , n23718 , n23721 );
and ( n23723 , n23716 , n23721 );
or ( n23724 , n23719 , n23722 , n23723 );
and ( n23725 , n23620 , n20909 );
and ( n23726 , n22354 , n22172 );
and ( n23727 , n23725 , n23726 );
and ( n23728 , n22232 , n22337 );
and ( n23729 , n23726 , n23728 );
and ( n23730 , n23725 , n23728 );
or ( n23731 , n23727 , n23729 , n23730 );
and ( n23732 , n21836 , n23508 );
buf ( n23733 , n23732 );
and ( n23734 , n22936 , n21296 );
and ( n23735 , n23733 , n23734 );
and ( n23736 , n22035 , n22784 );
and ( n23737 , n23734 , n23736 );
and ( n23738 , n23733 , n23736 );
or ( n23739 , n23735 , n23737 , n23738 );
and ( n23740 , n23731 , n23739 );
buf ( n23741 , n13689 );
buf ( n23742 , n23741 );
and ( n23743 , n23742 , n20890 );
and ( n23744 , n22542 , n21827 );
and ( n23745 , n23743 , n23744 );
buf ( n23746 , n21608 );
not ( n23747 , n23746 );
and ( n23748 , n23744 , n23747 );
and ( n23749 , n23743 , n23747 );
or ( n23750 , n23745 , n23748 , n23749 );
and ( n23751 , n23739 , n23750 );
and ( n23752 , n23731 , n23750 );
or ( n23753 , n23740 , n23751 , n23752 );
and ( n23754 , n22116 , n22562 );
and ( n23755 , n21914 , n22987 );
and ( n23756 , n23754 , n23755 );
buf ( n23757 , n20244 );
buf ( n23758 , n23757 );
and ( n23759 , n21672 , n23758 );
and ( n23760 , n23755 , n23759 );
and ( n23761 , n23754 , n23759 );
or ( n23762 , n23756 , n23760 , n23761 );
and ( n23763 , n22702 , n21429 );
and ( n23764 , n23762 , n23763 );
and ( n23765 , n23336 , n20949 );
and ( n23766 , n22035 , n22562 );
xor ( n23767 , n23765 , n23766 );
and ( n23768 , n21743 , n23322 );
xor ( n23769 , n23767 , n23768 );
and ( n23770 , n23763 , n23769 );
and ( n23771 , n23762 , n23769 );
or ( n23772 , n23764 , n23770 , n23771 );
and ( n23773 , n23753 , n23772 );
and ( n23774 , n23765 , n23766 );
and ( n23775 , n23766 , n23768 );
and ( n23776 , n23765 , n23768 );
or ( n23777 , n23774 , n23775 , n23776 );
buf ( n23778 , n23746 );
and ( n23779 , n22824 , n21296 );
and ( n23780 , n23778 , n23779 );
and ( n23781 , n22116 , n22337 );
and ( n23782 , n23779 , n23781 );
and ( n23783 , n23778 , n23781 );
or ( n23784 , n23780 , n23782 , n23783 );
xor ( n23785 , n23777 , n23784 );
and ( n23786 , n22589 , n21429 );
xor ( n23787 , n23785 , n23786 );
and ( n23788 , n23772 , n23787 );
and ( n23789 , n23753 , n23787 );
or ( n23790 , n23773 , n23788 , n23789 );
xor ( n23791 , n23602 , n23604 );
xor ( n23792 , n23791 , n23607 );
and ( n23793 , n23790 , n23792 );
and ( n23794 , n23777 , n23784 );
and ( n23795 , n23784 , n23786 );
and ( n23796 , n23777 , n23786 );
or ( n23797 , n23794 , n23795 , n23796 );
and ( n23798 , n22351 , n21827 );
and ( n23799 , n21914 , n22784 );
and ( n23800 , n23798 , n23799 );
and ( n23801 , n21836 , n22987 );
and ( n23802 , n23799 , n23801 );
and ( n23803 , n23798 , n23801 );
or ( n23804 , n23800 , n23802 , n23803 );
xor ( n23805 , n23504 , n23505 );
xor ( n23806 , n23805 , n23509 );
and ( n23807 , n23804 , n23806 );
xor ( n23808 , n23513 , n23514 );
xor ( n23809 , n23808 , n23516 );
and ( n23810 , n23806 , n23809 );
and ( n23811 , n23804 , n23809 );
or ( n23812 , n23807 , n23810 , n23811 );
xor ( n23813 , n23797 , n23812 );
xor ( n23814 , n23512 , n23519 );
xor ( n23815 , n23814 , n23521 );
xor ( n23816 , n23813 , n23815 );
and ( n23817 , n23792 , n23816 );
and ( n23818 , n23790 , n23816 );
or ( n23819 , n23793 , n23817 , n23818 );
xor ( n23820 , n23610 , n23612 );
xor ( n23821 , n23820 , n23615 );
and ( n23822 , n23819 , n23821 );
and ( n23823 , n23797 , n23812 );
and ( n23824 , n23812 , n23815 );
and ( n23825 , n23797 , n23815 );
or ( n23826 , n23823 , n23824 , n23825 );
and ( n23827 , n23742 , n20877 );
and ( n23828 , n22936 , n21178 );
and ( n23829 , n23827 , n23828 );
and ( n23830 , n22589 , n21527 );
and ( n23831 , n23828 , n23830 );
and ( n23832 , n23827 , n23830 );
or ( n23833 , n23829 , n23831 , n23832 );
and ( n23834 , n22542 , n21666 );
and ( n23835 , n22354 , n21990 );
and ( n23836 , n23834 , n23835 );
and ( n23837 , n22232 , n22172 );
and ( n23838 , n23835 , n23837 );
and ( n23839 , n23834 , n23837 );
or ( n23840 , n23836 , n23838 , n23839 );
and ( n23841 , n23833 , n23840 );
xor ( n23842 , n23543 , n23544 );
xor ( n23843 , n23842 , n23546 );
and ( n23844 , n23840 , n23843 );
and ( n23845 , n23833 , n23843 );
or ( n23846 , n23841 , n23844 , n23845 );
and ( n23847 , n23620 , n20890 );
and ( n23848 , n23483 , n20909 );
and ( n23849 , n23847 , n23848 );
not ( n23850 , n23628 );
and ( n23851 , n23848 , n23850 );
and ( n23852 , n23847 , n23850 );
or ( n23853 , n23849 , n23851 , n23852 );
xor ( n23854 , n23642 , n23643 );
xor ( n23855 , n23854 , n23645 );
and ( n23856 , n23853 , n23855 );
xor ( n23857 , n23629 , n23630 );
xor ( n23858 , n23857 , n23632 );
and ( n23859 , n23855 , n23858 );
and ( n23860 , n23853 , n23858 );
or ( n23861 , n23856 , n23859 , n23860 );
and ( n23862 , n23846 , n23861 );
xor ( n23863 , n23549 , n23550 );
xor ( n23864 , n23863 , n23553 );
and ( n23865 , n23861 , n23864 );
and ( n23866 , n23846 , n23864 );
or ( n23867 , n23862 , n23865 , n23866 );
xor ( n23868 , n23826 , n23867 );
xor ( n23869 , n23503 , n23524 );
xor ( n23870 , n23869 , n23527 );
xor ( n23871 , n23868 , n23870 );
and ( n23872 , n23821 , n23871 );
and ( n23873 , n23819 , n23871 );
or ( n23874 , n23822 , n23872 , n23873 );
and ( n23875 , n23724 , n23874 );
xor ( n23876 , n23618 , n23662 );
xor ( n23877 , n23876 , n23665 );
and ( n23878 , n23874 , n23877 );
and ( n23879 , n23724 , n23877 );
or ( n23880 , n23875 , n23878 , n23879 );
and ( n23881 , n23826 , n23867 );
and ( n23882 , n23867 , n23870 );
and ( n23883 , n23826 , n23870 );
or ( n23884 , n23881 , n23882 , n23883 );
xor ( n23885 , n23496 , n23530 );
xor ( n23886 , n23885 , n23533 );
and ( n23887 , n23884 , n23886 );
xor ( n23888 , n23564 , n23566 );
xor ( n23889 , n23888 , n23569 );
and ( n23890 , n23886 , n23889 );
and ( n23891 , n23884 , n23889 );
or ( n23892 , n23887 , n23890 , n23891 );
and ( n23893 , n23880 , n23892 );
xor ( n23894 , n23668 , n23670 );
xor ( n23895 , n23894 , n23673 );
and ( n23896 , n23892 , n23895 );
and ( n23897 , n23880 , n23895 );
or ( n23898 , n23893 , n23896 , n23897 );
and ( n23899 , n23687 , n23898 );
xor ( n23900 , n23880 , n23892 );
xor ( n23901 , n23900 , n23895 );
buf ( n23902 , n13781 );
buf ( n23903 , n23902 );
and ( n23904 , n23903 , n20877 );
and ( n23905 , n23215 , n21085 );
and ( n23906 , n23904 , n23905 );
and ( n23907 , n23089 , n21178 );
and ( n23908 , n23905 , n23907 );
and ( n23909 , n23904 , n23907 );
or ( n23910 , n23906 , n23908 , n23909 );
and ( n23911 , n22702 , n21527 );
and ( n23912 , n22589 , n21666 );
and ( n23913 , n23911 , n23912 );
and ( n23914 , n22351 , n21990 );
and ( n23915 , n23912 , n23914 );
and ( n23916 , n23911 , n23914 );
or ( n23917 , n23913 , n23915 , n23916 );
and ( n23918 , n23910 , n23917 );
xor ( n23919 , n23834 , n23835 );
xor ( n23920 , n23919 , n23837 );
and ( n23921 , n23917 , n23920 );
and ( n23922 , n23910 , n23920 );
or ( n23923 , n23918 , n23921 , n23922 );
xor ( n23924 , n23798 , n23799 );
xor ( n23925 , n23924 , n23801 );
xor ( n23926 , n23778 , n23779 );
xor ( n23927 , n23926 , n23781 );
and ( n23928 , n23925 , n23927 );
xor ( n23929 , n23847 , n23848 );
xor ( n23930 , n23929 , n23850 );
and ( n23931 , n23927 , n23930 );
and ( n23932 , n23925 , n23930 );
or ( n23933 , n23928 , n23931 , n23932 );
and ( n23934 , n23923 , n23933 );
xor ( n23935 , n23804 , n23806 );
xor ( n23936 , n23935 , n23809 );
and ( n23937 , n23933 , n23936 );
and ( n23938 , n23923 , n23936 );
or ( n23939 , n23934 , n23937 , n23938 );
xor ( n23940 , n23833 , n23840 );
xor ( n23941 , n23940 , n23843 );
xor ( n23942 , n23853 , n23855 );
xor ( n23943 , n23942 , n23858 );
and ( n23944 , n23941 , n23943 );
xor ( n23945 , n23700 , n23702 );
xor ( n23946 , n23945 , n23705 );
and ( n23947 , n23943 , n23946 );
and ( n23948 , n23941 , n23946 );
or ( n23949 , n23944 , n23947 , n23948 );
and ( n23950 , n23939 , n23949 );
xor ( n23951 , n23846 , n23861 );
xor ( n23952 , n23951 , n23864 );
and ( n23953 , n23949 , n23952 );
and ( n23954 , n23939 , n23952 );
or ( n23955 , n23950 , n23953 , n23954 );
and ( n23956 , n23620 , n20949 );
and ( n23957 , n22035 , n22987 );
and ( n23958 , n23956 , n23957 );
and ( n23959 , n21743 , n23758 );
and ( n23960 , n23957 , n23959 );
and ( n23961 , n23956 , n23959 );
or ( n23962 , n23958 , n23960 , n23961 );
buf ( n23963 , n21672 );
buf ( n23964 , n23963 );
and ( n23965 , n22232 , n22562 );
and ( n23966 , n23964 , n23965 );
and ( n23967 , n21914 , n23322 );
and ( n23968 , n23965 , n23967 );
and ( n23969 , n23964 , n23967 );
or ( n23970 , n23966 , n23968 , n23969 );
and ( n23971 , n23962 , n23970 );
and ( n23972 , n23336 , n21039 );
and ( n23973 , n23970 , n23972 );
and ( n23974 , n23962 , n23972 );
or ( n23975 , n23971 , n23973 , n23974 );
xor ( n23976 , n23827 , n23828 );
xor ( n23977 , n23976 , n23830 );
and ( n23978 , n23975 , n23977 );
xor ( n23979 , n23694 , n23695 );
xor ( n23980 , n23979 , n23697 );
and ( n23981 , n23977 , n23980 );
and ( n23982 , n23975 , n23980 );
or ( n23983 , n23978 , n23981 , n23982 );
and ( n23984 , n22824 , n21429 );
xor ( n23985 , n23688 , n23689 );
xor ( n23986 , n23985 , n23691 );
and ( n23987 , n23984 , n23986 );
xor ( n23988 , n23754 , n23755 );
xor ( n23989 , n23988 , n23759 );
and ( n23990 , n23986 , n23989 );
and ( n23991 , n23984 , n23989 );
or ( n23992 , n23987 , n23990 , n23991 );
and ( n23993 , n23336 , n21085 );
and ( n23994 , n23089 , n21296 );
and ( n23995 , n23993 , n23994 );
and ( n23996 , n22354 , n22337 );
and ( n23997 , n23994 , n23996 );
and ( n23998 , n23993 , n23996 );
or ( n23999 , n23995 , n23997 , n23998 );
xor ( n24000 , n23725 , n23726 );
xor ( n24001 , n24000 , n23728 );
and ( n24002 , n23999 , n24001 );
xor ( n24003 , n23743 , n23744 );
xor ( n24004 , n24003 , n23747 );
and ( n24005 , n24001 , n24004 );
and ( n24006 , n23999 , n24004 );
or ( n24007 , n24002 , n24005 , n24006 );
and ( n24008 , n23992 , n24007 );
xor ( n24009 , n23762 , n23763 );
xor ( n24010 , n24009 , n23769 );
and ( n24011 , n24007 , n24010 );
and ( n24012 , n23992 , n24010 );
or ( n24013 , n24008 , n24011 , n24012 );
and ( n24014 , n23983 , n24013 );
xor ( n24015 , n23753 , n23772 );
xor ( n24016 , n24015 , n23787 );
and ( n24017 , n24013 , n24016 );
and ( n24018 , n23983 , n24016 );
or ( n24019 , n24014 , n24017 , n24018 );
xor ( n24020 , n23708 , n23710 );
xor ( n24021 , n24020 , n23713 );
and ( n24022 , n24019 , n24021 );
xor ( n24023 , n23790 , n23792 );
xor ( n24024 , n24023 , n23816 );
and ( n24025 , n24021 , n24024 );
and ( n24026 , n24019 , n24024 );
or ( n24027 , n24022 , n24025 , n24026 );
and ( n24028 , n23955 , n24027 );
xor ( n24029 , n23716 , n23718 );
xor ( n24030 , n24029 , n23721 );
and ( n24031 , n24027 , n24030 );
and ( n24032 , n23955 , n24030 );
or ( n24033 , n24028 , n24031 , n24032 );
xor ( n24034 , n23724 , n23874 );
xor ( n24035 , n24034 , n23877 );
and ( n24036 , n24033 , n24035 );
xor ( n24037 , n23884 , n23886 );
xor ( n24038 , n24037 , n23889 );
and ( n24039 , n24035 , n24038 );
and ( n24040 , n24033 , n24038 );
or ( n24041 , n24036 , n24039 , n24040 );
and ( n24042 , n23901 , n24041 );
xor ( n24043 , n24033 , n24035 );
xor ( n24044 , n24043 , n24038 );
xor ( n24045 , n23819 , n23821 );
xor ( n24046 , n24045 , n23871 );
xor ( n24047 , n23955 , n24027 );
xor ( n24048 , n24047 , n24030 );
and ( n24049 , n24046 , n24048 );
and ( n24050 , n24044 , n24049 );
buf ( n24051 , n14265 );
buf ( n24052 , n24051 );
and ( n24053 , n24052 , n20877 );
and ( n24054 , n22702 , n21666 );
and ( n24055 , n24053 , n24054 );
and ( n24056 , n22542 , n21990 );
and ( n24057 , n24054 , n24056 );
and ( n24058 , n24053 , n24056 );
or ( n24059 , n24055 , n24057 , n24058 );
and ( n24060 , n22354 , n22562 );
and ( n24061 , n21914 , n23508 );
and ( n24062 , n24060 , n24061 );
buf ( n24063 , n20247 );
buf ( n24064 , n24063 );
and ( n24065 , n21743 , n24064 );
and ( n24066 , n24061 , n24065 );
and ( n24067 , n24060 , n24065 );
or ( n24068 , n24062 , n24066 , n24067 );
and ( n24069 , n23742 , n20949 );
and ( n24070 , n22035 , n23322 );
and ( n24071 , n24069 , n24070 );
not ( n24072 , n23963 );
and ( n24073 , n24070 , n24072 );
and ( n24074 , n24069 , n24072 );
or ( n24075 , n24071 , n24073 , n24074 );
and ( n24076 , n24068 , n24075 );
and ( n24077 , n22936 , n21429 );
and ( n24078 , n24075 , n24077 );
and ( n24079 , n24068 , n24077 );
or ( n24080 , n24076 , n24078 , n24079 );
and ( n24081 , n24059 , n24080 );
xor ( n24082 , n23904 , n23905 );
xor ( n24083 , n24082 , n23907 );
and ( n24084 , n24080 , n24083 );
and ( n24085 , n24059 , n24083 );
or ( n24086 , n24081 , n24084 , n24085 );
and ( n24087 , n23742 , n20909 );
and ( n24088 , n22589 , n21827 );
and ( n24089 , n24087 , n24088 );
and ( n24090 , n22351 , n22172 );
and ( n24091 , n24088 , n24090 );
and ( n24092 , n24087 , n24090 );
or ( n24093 , n24089 , n24091 , n24092 );
and ( n24094 , n23903 , n20890 );
and ( n24095 , n22116 , n22784 );
and ( n24096 , n24094 , n24095 );
not ( n24097 , n23732 );
and ( n24098 , n24095 , n24097 );
and ( n24099 , n24094 , n24097 );
or ( n24100 , n24096 , n24098 , n24099 );
and ( n24101 , n24093 , n24100 );
xor ( n24102 , n23733 , n23734 );
xor ( n24103 , n24102 , n23736 );
and ( n24104 , n24100 , n24103 );
and ( n24105 , n24093 , n24103 );
or ( n24106 , n24101 , n24104 , n24105 );
and ( n24107 , n24086 , n24106 );
xor ( n24108 , n23731 , n23739 );
xor ( n24109 , n24108 , n23750 );
and ( n24110 , n24106 , n24109 );
and ( n24111 , n24086 , n24109 );
or ( n24112 , n24107 , n24110 , n24111 );
xor ( n24113 , n23923 , n23933 );
xor ( n24114 , n24113 , n23936 );
and ( n24115 , n24112 , n24114 );
xor ( n24116 , n23941 , n23943 );
xor ( n24117 , n24116 , n23946 );
and ( n24118 , n24114 , n24117 );
and ( n24119 , n24112 , n24117 );
or ( n24120 , n24115 , n24118 , n24119 );
xor ( n24121 , n23939 , n23949 );
xor ( n24122 , n24121 , n23952 );
and ( n24123 , n24120 , n24122 );
xor ( n24124 , n24019 , n24021 );
xor ( n24125 , n24124 , n24024 );
xor ( n24126 , n24120 , n24122 );
and ( n24127 , n24125 , n24126 );
xor ( n24128 , n23983 , n24013 );
xor ( n24129 , n24128 , n24016 );
xor ( n24130 , n24112 , n24114 );
xor ( n24131 , n24130 , n24117 );
and ( n24132 , n24129 , n24131 );
and ( n24133 , n23483 , n21039 );
and ( n24134 , n23215 , n21178 );
and ( n24135 , n24133 , n24134 );
and ( n24136 , n22824 , n21527 );
and ( n24137 , n24134 , n24136 );
and ( n24138 , n24133 , n24136 );
or ( n24139 , n24135 , n24137 , n24138 );
xor ( n24140 , n23911 , n23912 );
xor ( n24141 , n24140 , n23914 );
and ( n24142 , n24139 , n24141 );
xor ( n24143 , n23962 , n23970 );
xor ( n24144 , n24143 , n23972 );
and ( n24145 , n24141 , n24144 );
and ( n24146 , n24139 , n24144 );
or ( n24147 , n24142 , n24145 , n24146 );
xor ( n24148 , n23910 , n23917 );
xor ( n24149 , n24148 , n23920 );
and ( n24150 , n24147 , n24149 );
xor ( n24151 , n23925 , n23927 );
xor ( n24152 , n24151 , n23930 );
and ( n24153 , n24149 , n24152 );
and ( n24154 , n24147 , n24152 );
or ( n24155 , n24150 , n24153 , n24154 );
and ( n24156 , n24131 , n24155 );
and ( n24157 , n24129 , n24155 );
or ( n24158 , n24132 , n24156 , n24157 );
and ( n24159 , n24126 , n24158 );
and ( n24160 , n24125 , n24158 );
or ( n24161 , n24127 , n24159 , n24160 );
and ( n24162 , n24123 , n24161 );
xor ( n24163 , n24046 , n24048 );
and ( n24164 , n24161 , n24163 );
and ( n24165 , n24123 , n24163 );
or ( n24166 , n24162 , n24164 , n24165 );
and ( n24167 , n24049 , n24166 );
and ( n24168 , n24044 , n24166 );
or ( n24169 , n24050 , n24167 , n24168 );
and ( n24170 , n24041 , n24169 );
and ( n24171 , n23901 , n24169 );
or ( n24172 , n24042 , n24170 , n24171 );
and ( n24173 , n23898 , n24172 );
and ( n24174 , n23687 , n24172 );
or ( n24175 , n23899 , n24173 , n24174 );
and ( n24176 , n23684 , n24175 );
and ( n24177 , n23595 , n24175 );
or ( n24178 , n23685 , n24176 , n24177 );
and ( n24179 , n23592 , n24178 );
and ( n24180 , n23412 , n24178 );
or ( n24181 , n23593 , n24179 , n24180 );
and ( n24182 , n23409 , n24181 );
and ( n24183 , n23261 , n24181 );
or ( n24184 , n23410 , n24182 , n24183 );
and ( n24185 , n23258 , n24184 );
and ( n24186 , n23164 , n24184 );
or ( n24187 , n23259 , n24185 , n24186 );
and ( n24188 , n23161 , n24187 );
and ( n24189 , n23038 , n24187 );
or ( n24190 , n23162 , n24188 , n24189 );
and ( n24191 , n23035 , n24190 );
and ( n24192 , n22905 , n24190 );
or ( n24193 , n23036 , n24191 , n24192 );
and ( n24194 , n22902 , n24193 );
and ( n24195 , n22779 , n24193 );
or ( n24196 , n22903 , n24194 , n24195 );
and ( n24197 , n22776 , n24196 );
and ( n24198 , n22674 , n24196 );
or ( n24199 , n22777 , n24197 , n24198 );
and ( n24200 , n22671 , n24199 );
and ( n24201 , n22540 , n24199 );
or ( n24202 , n22672 , n24200 , n24201 );
and ( n24203 , n22537 , n24202 );
and ( n24204 , n22535 , n24202 );
or ( n24205 , n22538 , n24203 , n24204 );
and ( n24206 , n22433 , n24205 );
and ( n24207 , n22322 , n24205 );
or ( n24208 , n22434 , n24206 , n24207 );
and ( n24209 , n22319 , n24208 );
and ( n24210 , n22157 , n24208 );
or ( n24211 , n22320 , n24209 , n24210 );
and ( n24212 , n22154 , n24211 );
and ( n24213 , n22112 , n24211 );
or ( n24214 , n22155 , n24212 , n24213 );
and ( n24215 , n22109 , n24214 );
and ( n24216 , n21969 , n24214 );
or ( n24217 , n22110 , n24215 , n24216 );
and ( n24218 , n21966 , n24217 );
and ( n24219 , n21912 , n24217 );
or ( n24220 , n21967 , n24218 , n24219 );
and ( n24221 , n21909 , n24220 );
and ( n24222 , n21815 , n24220 );
or ( n24223 , n21910 , n24221 , n24222 );
and ( n24224 , n21812 , n24223 );
and ( n24225 , n21732 , n24223 );
or ( n24226 , n21813 , n24224 , n24225 );
and ( n24227 , n21729 , n24226 );
and ( n24228 , n21648 , n24226 );
or ( n24229 , n21730 , n24227 , n24228 );
and ( n24230 , n21645 , n24229 );
and ( n24231 , n21572 , n24229 );
or ( n24232 , n21646 , n24230 , n24231 );
and ( n24233 , n21569 , n24232 );
and ( n24234 , n21567 , n24232 );
or ( n24235 , n21570 , n24233 , n24234 );
and ( n24236 , n21491 , n24235 );
and ( n24237 , n21423 , n24235 );
or ( n24238 , n21492 , n24236 , n24237 );
and ( n24239 , n21420 , n24238 );
and ( n24240 , n21353 , n24238 );
or ( n24241 , n21421 , n24239 , n24240 );
and ( n24242 , n21350 , n24241 );
and ( n24243 , n21270 , n24241 );
or ( n24244 , n21351 , n24242 , n24243 );
and ( n24245 , n21267 , n24244 );
and ( n24246 , n21228 , n24244 );
or ( n24247 , n21268 , n24245 , n24246 );
and ( n24248 , n21225 , n24247 );
and ( n24249 , n21171 , n24247 );
or ( n24250 , n21226 , n24248 , n24249 );
and ( n24251 , n21168 , n24250 );
and ( n24252 , n21166 , n24250 );
or ( n24253 , n21169 , n24251 , n24252 );
and ( n24254 , n21120 , n24253 );
and ( n24255 , n21118 , n24253 );
or ( n24256 , n21121 , n24254 , n24255 );
and ( n24257 , n21057 , n24256 );
and ( n24258 , n21017 , n24256 );
or ( n24259 , n21058 , n24257 , n24258 );
and ( n24260 , n21014 , n24259 );
and ( n24261 , n21012 , n24259 );
or ( n24262 , n21015 , n24260 , n24261 );
or ( n24263 , n20987 , n24262 );
or ( n24264 , n20985 , n24263 );
or ( n24265 , n20983 , n24264 );
xnor ( n24266 , n20981 , n24265 );
xnor ( n24267 , n20983 , n24264 );
xnor ( n24268 , n20985 , n24263 );
xnor ( n24269 , n20987 , n24262 );
xor ( n24270 , n21012 , n21014 );
xor ( n24271 , n24270 , n24259 );
xor ( n24272 , n21017 , n21057 );
xor ( n24273 , n24272 , n24256 );
xor ( n24274 , n21118 , n21120 );
xor ( n24275 , n24274 , n24253 );
xor ( n24276 , n21166 , n21168 );
xor ( n24277 , n24276 , n24250 );
xor ( n24278 , n21171 , n21225 );
xor ( n24279 , n24278 , n24247 );
xor ( n24280 , n21228 , n21267 );
xor ( n24281 , n24280 , n24244 );
xor ( n24282 , n21270 , n21350 );
xor ( n24283 , n24282 , n24241 );
xor ( n24284 , n21353 , n21420 );
xor ( n24285 , n24284 , n24238 );
xor ( n24286 , n21423 , n21491 );
xor ( n24287 , n24286 , n24235 );
xor ( n24288 , n21567 , n21569 );
xor ( n24289 , n24288 , n24232 );
xor ( n24290 , n21572 , n21645 );
xor ( n24291 , n24290 , n24229 );
xor ( n24292 , n21648 , n21729 );
xor ( n24293 , n24292 , n24226 );
xor ( n24294 , n21732 , n21812 );
xor ( n24295 , n24294 , n24223 );
xor ( n24296 , n21815 , n21909 );
xor ( n24297 , n24296 , n24220 );
xor ( n24298 , n21912 , n21966 );
xor ( n24299 , n24298 , n24217 );
xor ( n24300 , n21969 , n22109 );
xor ( n24301 , n24300 , n24214 );
xor ( n24302 , n22112 , n22154 );
xor ( n24303 , n24302 , n24211 );
xor ( n24304 , n22157 , n22319 );
xor ( n24305 , n24304 , n24208 );
xor ( n24306 , n22322 , n22433 );
xor ( n24307 , n24306 , n24205 );
xor ( n24308 , n22535 , n22537 );
xor ( n24309 , n24308 , n24202 );
xor ( n24310 , n22540 , n22671 );
xor ( n24311 , n24310 , n24199 );
xor ( n24312 , n22674 , n22776 );
xor ( n24313 , n24312 , n24196 );
xor ( n24314 , n22779 , n22902 );
xor ( n24315 , n24314 , n24193 );
xor ( n24316 , n22905 , n23035 );
xor ( n24317 , n24316 , n24190 );
xor ( n24318 , n23038 , n23161 );
xor ( n24319 , n24318 , n24187 );
xor ( n24320 , n23164 , n23258 );
xor ( n24321 , n24320 , n24184 );
xor ( n24322 , n23261 , n23409 );
xor ( n24323 , n24322 , n24181 );
xor ( n24324 , n23412 , n23592 );
xor ( n24325 , n24324 , n24178 );
xor ( n24326 , n23595 , n23684 );
xor ( n24327 , n24326 , n24175 );
xor ( n24328 , n23687 , n23898 );
xor ( n24329 , n24328 , n24172 );
xor ( n24330 , n23901 , n24041 );
xor ( n24331 , n24330 , n24169 );
xor ( n24332 , n24044 , n24049 );
xor ( n24333 , n24332 , n24166 );
xor ( n24334 , n23992 , n24007 );
xor ( n24335 , n24334 , n24010 );
buf ( n24336 , n14507 );
buf ( n24337 , n24336 );
and ( n24338 , n24337 , n20877 );
and ( n24339 , n23336 , n21178 );
and ( n24340 , n24338 , n24339 );
and ( n24341 , n22232 , n22784 );
and ( n24342 , n24339 , n24341 );
and ( n24343 , n24338 , n24341 );
or ( n24344 , n24340 , n24342 , n24343 );
xor ( n24345 , n24087 , n24088 );
xor ( n24346 , n24345 , n24090 );
and ( n24347 , n24344 , n24346 );
xor ( n24348 , n24094 , n24095 );
xor ( n24349 , n24348 , n24097 );
and ( n24350 , n24346 , n24349 );
and ( n24351 , n24344 , n24349 );
or ( n24352 , n24347 , n24350 , n24351 );
xor ( n24353 , n23984 , n23986 );
xor ( n24354 , n24353 , n23989 );
and ( n24355 , n24352 , n24354 );
and ( n24356 , n24335 , n24355 );
xor ( n24357 , n24086 , n24106 );
xor ( n24358 , n24357 , n24109 );
and ( n24359 , n24355 , n24358 );
and ( n24360 , n24335 , n24358 );
or ( n24361 , n24356 , n24359 , n24360 );
xor ( n24362 , n23975 , n23977 );
xor ( n24363 , n24362 , n23980 );
and ( n24364 , n23215 , n21296 );
and ( n24365 , n22116 , n22987 );
and ( n24366 , n24364 , n24365 );
and ( n24367 , n21836 , n23758 );
and ( n24368 , n24365 , n24367 );
and ( n24369 , n24364 , n24367 );
or ( n24370 , n24366 , n24368 , n24369 );
xor ( n24371 , n23956 , n23957 );
xor ( n24372 , n24371 , n23959 );
and ( n24373 , n24370 , n24372 );
xor ( n24374 , n23964 , n23965 );
xor ( n24375 , n24374 , n23967 );
and ( n24376 , n24372 , n24375 );
and ( n24377 , n24370 , n24375 );
or ( n24378 , n24373 , n24376 , n24377 );
xor ( n24379 , n24093 , n24100 );
xor ( n24380 , n24379 , n24103 );
and ( n24381 , n24378 , n24380 );
and ( n24382 , n24363 , n24381 );
and ( n24383 , n23483 , n21085 );
and ( n24384 , n22824 , n21666 );
and ( n24385 , n24383 , n24384 );
and ( n24386 , n22589 , n21990 );
and ( n24387 , n24384 , n24386 );
and ( n24388 , n24383 , n24386 );
or ( n24389 , n24385 , n24387 , n24388 );
xor ( n24390 , n24053 , n24054 );
xor ( n24391 , n24390 , n24056 );
or ( n24392 , n24389 , n24391 );
xor ( n24393 , n24133 , n24134 );
xor ( n24394 , n24393 , n24136 );
xor ( n24395 , n23993 , n23994 );
xor ( n24396 , n24395 , n23996 );
and ( n24397 , n24394 , n24396 );
and ( n24398 , n23903 , n20909 );
and ( n24399 , n22542 , n22172 );
and ( n24400 , n24398 , n24399 );
and ( n24401 , n22351 , n22337 );
and ( n24402 , n24399 , n24401 );
and ( n24403 , n24398 , n24401 );
or ( n24404 , n24400 , n24402 , n24403 );
and ( n24405 , n24396 , n24404 );
and ( n24406 , n24394 , n24404 );
or ( n24407 , n24397 , n24405 , n24406 );
and ( n24408 , n24392 , n24407 );
xor ( n24409 , n24059 , n24080 );
xor ( n24410 , n24409 , n24083 );
and ( n24411 , n24407 , n24410 );
and ( n24412 , n24392 , n24410 );
or ( n24413 , n24408 , n24411 , n24412 );
and ( n24414 , n24381 , n24413 );
and ( n24415 , n24363 , n24413 );
or ( n24416 , n24382 , n24414 , n24415 );
and ( n24417 , n24361 , n24416 );
xor ( n24418 , n24352 , n24354 );
and ( n24419 , n24052 , n20890 );
and ( n24420 , n23089 , n21429 );
and ( n24421 , n24419 , n24420 );
and ( n24422 , n22702 , n21827 );
and ( n24423 , n24420 , n24422 );
and ( n24424 , n24419 , n24422 );
or ( n24425 , n24421 , n24423 , n24424 );
xor ( n24426 , n24068 , n24075 );
xor ( n24427 , n24426 , n24077 );
and ( n24428 , n24425 , n24427 );
xor ( n24429 , n24344 , n24346 );
xor ( n24430 , n24429 , n24349 );
and ( n24431 , n24427 , n24430 );
and ( n24432 , n24425 , n24430 );
or ( n24433 , n24428 , n24431 , n24432 );
and ( n24434 , n24418 , n24433 );
xnor ( n24435 , n24389 , n24391 );
and ( n24436 , n23620 , n21039 );
and ( n24437 , n22936 , n21527 );
and ( n24438 , n24436 , n24437 );
xor ( n24439 , n24060 , n24061 );
xor ( n24440 , n24439 , n24065 );
and ( n24441 , n24437 , n24440 );
and ( n24442 , n24436 , n24440 );
or ( n24443 , n24438 , n24441 , n24442 );
and ( n24444 , n24435 , n24443 );
and ( n24445 , n23620 , n21085 );
and ( n24446 , n23483 , n21178 );
and ( n24447 , n24445 , n24446 );
and ( n24448 , n22702 , n21990 );
and ( n24449 , n24446 , n24448 );
and ( n24450 , n24445 , n24448 );
or ( n24451 , n24447 , n24449 , n24450 );
xor ( n24452 , n24398 , n24399 );
xor ( n24453 , n24452 , n24401 );
or ( n24454 , n24451 , n24453 );
and ( n24455 , n24443 , n24454 );
and ( n24456 , n24435 , n24454 );
or ( n24457 , n24444 , n24455 , n24456 );
and ( n24458 , n24433 , n24457 );
and ( n24459 , n24418 , n24457 );
or ( n24460 , n24434 , n24458 , n24459 );
xor ( n24461 , n24147 , n24149 );
xor ( n24462 , n24461 , n24152 );
and ( n24463 , n24460 , n24462 );
xor ( n24464 , n23999 , n24001 );
xor ( n24465 , n24464 , n24004 );
xor ( n24466 , n24139 , n24141 );
xor ( n24467 , n24466 , n24144 );
or ( n24468 , n24465 , n24467 );
and ( n24469 , n24462 , n24468 );
and ( n24470 , n24460 , n24468 );
or ( n24471 , n24463 , n24469 , n24470 );
and ( n24472 , n24416 , n24471 );
and ( n24473 , n24361 , n24471 );
or ( n24474 , n24417 , n24472 , n24473 );
xor ( n24475 , n24125 , n24126 );
xor ( n24476 , n24475 , n24158 );
and ( n24477 , n24474 , n24476 );
xor ( n24478 , n24364 , n24365 );
xor ( n24479 , n24478 , n24367 );
xor ( n24480 , n24069 , n24070 );
xor ( n24481 , n24480 , n24072 );
and ( n24482 , n24479 , n24481 );
and ( n24483 , n23903 , n20949 );
and ( n24484 , n22116 , n23322 );
and ( n24485 , n24483 , n24484 );
and ( n24486 , n22035 , n23508 );
and ( n24487 , n24484 , n24486 );
and ( n24488 , n24483 , n24486 );
or ( n24489 , n24485 , n24487 , n24488 );
and ( n24490 , n24481 , n24489 );
and ( n24491 , n24479 , n24489 );
or ( n24492 , n24482 , n24490 , n24491 );
and ( n24493 , n22351 , n22562 );
and ( n24494 , n22232 , n22987 );
and ( n24495 , n24493 , n24494 );
and ( n24496 , n21914 , n23758 );
and ( n24497 , n24494 , n24496 );
and ( n24498 , n24493 , n24496 );
or ( n24499 , n24495 , n24497 , n24498 );
and ( n24500 , n23215 , n21429 );
and ( n24501 , n22542 , n22337 );
and ( n24502 , n24500 , n24501 );
and ( n24503 , n21836 , n24064 );
and ( n24504 , n24501 , n24503 );
and ( n24505 , n24500 , n24503 );
or ( n24506 , n24502 , n24504 , n24505 );
and ( n24507 , n24499 , n24506 );
xor ( n24508 , n24419 , n24420 );
xor ( n24509 , n24508 , n24422 );
and ( n24510 , n24506 , n24509 );
and ( n24511 , n24499 , n24509 );
or ( n24512 , n24507 , n24510 , n24511 );
and ( n24513 , n24492 , n24512 );
xor ( n24514 , n24394 , n24396 );
xor ( n24515 , n24514 , n24404 );
and ( n24516 , n24512 , n24515 );
and ( n24517 , n24492 , n24515 );
or ( n24518 , n24513 , n24516 , n24517 );
xor ( n24519 , n24378 , n24380 );
and ( n24520 , n24518 , n24519 );
and ( n24521 , n24337 , n20890 );
and ( n24522 , n24052 , n20909 );
and ( n24523 , n24521 , n24522 );
and ( n24524 , n22589 , n22172 );
and ( n24525 , n24522 , n24524 );
and ( n24526 , n24521 , n24524 );
or ( n24527 , n24523 , n24525 , n24526 );
and ( n24528 , n23336 , n21296 );
and ( n24529 , n22824 , n21827 );
and ( n24530 , n24528 , n24529 );
and ( n24531 , n22354 , n22784 );
and ( n24532 , n24529 , n24531 );
and ( n24533 , n24528 , n24531 );
or ( n24534 , n24530 , n24532 , n24533 );
and ( n24535 , n24527 , n24534 );
and ( n24536 , n22116 , n23508 );
and ( n24537 , n21914 , n24064 );
and ( n24538 , n24536 , n24537 );
buf ( n24539 , n20252 );
buf ( n24540 , n24539 );
and ( n24541 , n21836 , n24540 );
and ( n24542 , n24537 , n24541 );
and ( n24543 , n24536 , n24541 );
or ( n24544 , n24538 , n24542 , n24543 );
buf ( n24545 , n14700 );
buf ( n24546 , n24545 );
and ( n24547 , n24546 , n20877 );
and ( n24548 , n24544 , n24547 );
and ( n24549 , n22936 , n21666 );
and ( n24550 , n24547 , n24549 );
and ( n24551 , n24544 , n24549 );
or ( n24552 , n24548 , n24550 , n24551 );
and ( n24553 , n24534 , n24552 );
and ( n24554 , n24527 , n24552 );
or ( n24555 , n24535 , n24553 , n24554 );
and ( n24556 , n24052 , n20949 );
and ( n24557 , n22542 , n22562 );
and ( n24558 , n24556 , n24557 );
and ( n24559 , n22035 , n23758 );
and ( n24560 , n24557 , n24559 );
and ( n24561 , n24556 , n24559 );
or ( n24562 , n24558 , n24560 , n24561 );
and ( n24563 , n23742 , n21039 );
and ( n24564 , n24562 , n24563 );
and ( n24565 , n23089 , n21527 );
and ( n24566 , n24563 , n24565 );
and ( n24567 , n24562 , n24565 );
or ( n24568 , n24564 , n24566 , n24567 );
xor ( n24569 , n24338 , n24339 );
xor ( n24570 , n24569 , n24341 );
and ( n24571 , n24568 , n24570 );
xor ( n24572 , n24383 , n24384 );
xor ( n24573 , n24572 , n24386 );
and ( n24574 , n24570 , n24573 );
and ( n24575 , n24568 , n24573 );
or ( n24576 , n24571 , n24574 , n24575 );
and ( n24577 , n24555 , n24576 );
xor ( n24578 , n24370 , n24372 );
xor ( n24579 , n24578 , n24375 );
and ( n24580 , n24576 , n24579 );
and ( n24581 , n24555 , n24579 );
or ( n24582 , n24577 , n24580 , n24581 );
and ( n24583 , n24519 , n24582 );
and ( n24584 , n24518 , n24582 );
or ( n24585 , n24520 , n24583 , n24584 );
xor ( n24586 , n24436 , n24437 );
xor ( n24587 , n24586 , n24440 );
xnor ( n24588 , n24451 , n24453 );
and ( n24589 , n24587 , n24588 );
xor ( n24590 , n24483 , n24484 );
xor ( n24591 , n24590 , n24486 );
xor ( n24592 , n24493 , n24494 );
xor ( n24593 , n24592 , n24496 );
and ( n24594 , n24591 , n24593 );
and ( n24595 , n24337 , n20909 );
and ( n24596 , n22702 , n22172 );
and ( n24597 , n24595 , n24596 );
and ( n24598 , n22589 , n22337 );
and ( n24599 , n24596 , n24598 );
and ( n24600 , n24595 , n24598 );
or ( n24601 , n24597 , n24599 , n24600 );
and ( n24602 , n24593 , n24601 );
and ( n24603 , n24591 , n24601 );
or ( n24604 , n24594 , n24602 , n24603 );
and ( n24605 , n24588 , n24604 );
and ( n24606 , n24587 , n24604 );
or ( n24607 , n24589 , n24605 , n24606 );
and ( n24608 , n24546 , n20890 );
and ( n24609 , n23620 , n21178 );
and ( n24610 , n24608 , n24609 );
and ( n24611 , n22936 , n21827 );
and ( n24612 , n24609 , n24611 );
and ( n24613 , n24608 , n24611 );
or ( n24614 , n24610 , n24612 , n24613 );
and ( n24615 , n23483 , n21296 );
and ( n24616 , n22351 , n22784 );
and ( n24617 , n24615 , n24616 );
and ( n24618 , n22354 , n22987 );
and ( n24619 , n24616 , n24618 );
and ( n24620 , n24615 , n24618 );
or ( n24621 , n24617 , n24619 , n24620 );
and ( n24622 , n24614 , n24621 );
buf ( n24623 , n14989 );
buf ( n24624 , n24623 );
and ( n24625 , n24624 , n20877 );
and ( n24626 , n23742 , n21085 );
and ( n24627 , n24625 , n24626 );
and ( n24628 , n22824 , n21990 );
and ( n24629 , n24626 , n24628 );
and ( n24630 , n24625 , n24628 );
or ( n24631 , n24627 , n24629 , n24630 );
and ( n24632 , n24621 , n24631 );
and ( n24633 , n24614 , n24631 );
or ( n24634 , n24622 , n24632 , n24633 );
xor ( n24635 , n24479 , n24481 );
xor ( n24636 , n24635 , n24489 );
and ( n24637 , n24634 , n24636 );
xor ( n24638 , n24499 , n24506 );
xor ( n24639 , n24638 , n24509 );
and ( n24640 , n24636 , n24639 );
and ( n24641 , n24634 , n24639 );
or ( n24642 , n24637 , n24640 , n24641 );
and ( n24643 , n24607 , n24642 );
xor ( n24644 , n24425 , n24427 );
xor ( n24645 , n24644 , n24430 );
and ( n24646 , n24642 , n24645 );
and ( n24647 , n24607 , n24645 );
or ( n24648 , n24643 , n24646 , n24647 );
xor ( n24649 , n24392 , n24407 );
xor ( n24650 , n24649 , n24410 );
and ( n24651 , n24648 , n24650 );
xor ( n24652 , n24418 , n24433 );
xor ( n24653 , n24652 , n24457 );
and ( n24654 , n24650 , n24653 );
and ( n24655 , n24648 , n24653 );
or ( n24656 , n24651 , n24654 , n24655 );
and ( n24657 , n24585 , n24656 );
xor ( n24658 , n24335 , n24355 );
xor ( n24659 , n24658 , n24358 );
and ( n24660 , n24656 , n24659 );
and ( n24661 , n24585 , n24659 );
or ( n24662 , n24657 , n24660 , n24661 );
xor ( n24663 , n24129 , n24131 );
xor ( n24664 , n24663 , n24155 );
and ( n24665 , n24662 , n24664 );
xor ( n24666 , n24363 , n24381 );
xor ( n24667 , n24666 , n24413 );
xnor ( n24668 , n24465 , n24467 );
xor ( n24669 , n24435 , n24443 );
xor ( n24670 , n24669 , n24454 );
xor ( n24671 , n24492 , n24512 );
xor ( n24672 , n24671 , n24515 );
and ( n24673 , n24670 , n24672 );
xor ( n24674 , n24555 , n24576 );
xor ( n24675 , n24674 , n24579 );
and ( n24676 , n24672 , n24675 );
and ( n24677 , n24670 , n24675 );
or ( n24678 , n24673 , n24676 , n24677 );
and ( n24679 , n24668 , n24678 );
xor ( n24680 , n24527 , n24534 );
xor ( n24681 , n24680 , n24552 );
xor ( n24682 , n24568 , n24570 );
xor ( n24683 , n24682 , n24573 );
and ( n24684 , n24681 , n24683 );
and ( n24685 , n22232 , n23508 );
and ( n24686 , n22035 , n24064 );
and ( n24687 , n24685 , n24686 );
and ( n24688 , n21914 , n24540 );
and ( n24689 , n24686 , n24688 );
and ( n24690 , n24685 , n24688 );
or ( n24691 , n24687 , n24689 , n24690 );
and ( n24692 , n23215 , n21527 );
and ( n24693 , n24691 , n24692 );
and ( n24694 , n23089 , n21666 );
and ( n24695 , n24692 , n24694 );
and ( n24696 , n24691 , n24694 );
or ( n24697 , n24693 , n24695 , n24696 );
xor ( n24698 , n24521 , n24522 );
xor ( n24699 , n24698 , n24524 );
and ( n24700 , n24697 , n24699 );
xor ( n24701 , n24528 , n24529 );
xor ( n24702 , n24701 , n24531 );
and ( n24703 , n24699 , n24702 );
and ( n24704 , n24697 , n24702 );
or ( n24705 , n24700 , n24703 , n24704 );
and ( n24706 , n24683 , n24705 );
and ( n24707 , n24681 , n24705 );
or ( n24708 , n24684 , n24706 , n24707 );
and ( n24709 , n23903 , n21039 );
and ( n24710 , n23336 , n21429 );
and ( n24711 , n24709 , n24710 );
xor ( n24712 , n24536 , n24537 );
xor ( n24713 , n24712 , n24541 );
and ( n24714 , n24710 , n24713 );
and ( n24715 , n24709 , n24713 );
or ( n24716 , n24711 , n24714 , n24715 );
xor ( n24717 , n24445 , n24446 );
xor ( n24718 , n24717 , n24448 );
and ( n24719 , n24716 , n24718 );
xor ( n24720 , n24544 , n24547 );
xor ( n24721 , n24720 , n24549 );
and ( n24722 , n24718 , n24721 );
and ( n24723 , n24716 , n24721 );
or ( n24724 , n24719 , n24722 , n24723 );
xor ( n24725 , n24500 , n24501 );
xor ( n24726 , n24725 , n24503 );
xor ( n24727 , n24562 , n24563 );
xor ( n24728 , n24727 , n24565 );
and ( n24729 , n24726 , n24728 );
buf ( n24730 , n15019 );
buf ( n24731 , n24730 );
and ( n24732 , n24731 , n20877 );
and ( n24733 , n23215 , n21666 );
and ( n24734 , n24732 , n24733 );
and ( n24735 , n22936 , n21990 );
and ( n24736 , n24733 , n24735 );
and ( n24737 , n24732 , n24735 );
or ( n24738 , n24734 , n24736 , n24737 );
and ( n24739 , n23903 , n21085 );
and ( n24740 , n23742 , n21178 );
and ( n24741 , n24739 , n24740 );
and ( n24742 , n22542 , n22784 );
and ( n24743 , n24740 , n24742 );
and ( n24744 , n24739 , n24742 );
or ( n24745 , n24741 , n24743 , n24744 );
and ( n24746 , n24738 , n24745 );
xor ( n24747 , n24595 , n24596 );
xor ( n24748 , n24747 , n24598 );
and ( n24749 , n24745 , n24748 );
and ( n24750 , n24738 , n24748 );
or ( n24751 , n24746 , n24749 , n24750 );
and ( n24752 , n24728 , n24751 );
and ( n24753 , n24726 , n24751 );
or ( n24754 , n24729 , n24752 , n24753 );
and ( n24755 , n24724 , n24754 );
and ( n24756 , n22232 , n23322 );
buf ( n24757 , n21743 );
and ( n24758 , n24756 , n24757 );
xor ( n24759 , n24556 , n24557 );
xor ( n24760 , n24759 , n24559 );
and ( n24761 , n24757 , n24760 );
and ( n24762 , n24756 , n24760 );
or ( n24763 , n24758 , n24761 , n24762 );
and ( n24764 , n24337 , n20949 );
and ( n24765 , n22589 , n22562 );
and ( n24766 , n24764 , n24765 );
and ( n24767 , n22354 , n23322 );
and ( n24768 , n24765 , n24767 );
and ( n24769 , n24764 , n24767 );
or ( n24770 , n24766 , n24768 , n24769 );
and ( n24771 , n24624 , n20890 );
and ( n24772 , n24546 , n20909 );
and ( n24773 , n24771 , n24772 );
and ( n24774 , n22824 , n22172 );
and ( n24775 , n24772 , n24774 );
and ( n24776 , n24771 , n24774 );
or ( n24777 , n24773 , n24775 , n24776 );
and ( n24778 , n24770 , n24777 );
and ( n24779 , n23620 , n21296 );
and ( n24780 , n23089 , n21827 );
and ( n24781 , n24779 , n24780 );
and ( n24782 , n22702 , n22337 );
and ( n24783 , n24780 , n24782 );
and ( n24784 , n24779 , n24782 );
or ( n24785 , n24781 , n24783 , n24784 );
and ( n24786 , n24777 , n24785 );
and ( n24787 , n24770 , n24785 );
or ( n24788 , n24778 , n24786 , n24787 );
and ( n24789 , n24763 , n24788 );
xor ( n24790 , n24591 , n24593 );
xor ( n24791 , n24790 , n24601 );
and ( n24792 , n24788 , n24791 );
and ( n24793 , n24763 , n24791 );
or ( n24794 , n24789 , n24792 , n24793 );
and ( n24795 , n24754 , n24794 );
and ( n24796 , n24724 , n24794 );
or ( n24797 , n24755 , n24795 , n24796 );
and ( n24798 , n24708 , n24797 );
xor ( n24799 , n24607 , n24642 );
xor ( n24800 , n24799 , n24645 );
and ( n24801 , n24797 , n24800 );
and ( n24802 , n24708 , n24800 );
or ( n24803 , n24798 , n24801 , n24802 );
and ( n24804 , n24678 , n24803 );
and ( n24805 , n24668 , n24803 );
or ( n24806 , n24679 , n24804 , n24805 );
and ( n24807 , n24667 , n24806 );
xor ( n24808 , n24460 , n24462 );
xor ( n24809 , n24808 , n24468 );
and ( n24810 , n24806 , n24809 );
and ( n24811 , n24667 , n24809 );
or ( n24812 , n24807 , n24810 , n24811 );
and ( n24813 , n24664 , n24812 );
and ( n24814 , n24662 , n24812 );
or ( n24815 , n24665 , n24813 , n24814 );
and ( n24816 , n24476 , n24815 );
and ( n24817 , n24474 , n24815 );
or ( n24818 , n24477 , n24816 , n24817 );
xor ( n24819 , n24123 , n24161 );
xor ( n24820 , n24819 , n24163 );
and ( n24821 , n24818 , n24820 );
xor ( n24822 , n24361 , n24416 );
xor ( n24823 , n24822 , n24471 );
xor ( n24824 , n24585 , n24656 );
xor ( n24825 , n24824 , n24659 );
xor ( n24826 , n24518 , n24519 );
xor ( n24827 , n24826 , n24582 );
xor ( n24828 , n24648 , n24650 );
xor ( n24829 , n24828 , n24653 );
and ( n24830 , n24827 , n24829 );
xor ( n24831 , n24587 , n24588 );
xor ( n24832 , n24831 , n24604 );
xor ( n24833 , n24634 , n24636 );
xor ( n24834 , n24833 , n24639 );
and ( n24835 , n24832 , n24834 );
xor ( n24836 , n24697 , n24699 );
xor ( n24837 , n24836 , n24702 );
xor ( n24838 , n24716 , n24718 );
xor ( n24839 , n24838 , n24721 );
and ( n24840 , n24837 , n24839 );
and ( n24841 , n24834 , n24840 );
and ( n24842 , n24832 , n24840 );
or ( n24843 , n24835 , n24841 , n24842 );
xor ( n24844 , n24614 , n24621 );
xor ( n24845 , n24844 , n24631 );
xor ( n24846 , n24608 , n24609 );
xor ( n24847 , n24846 , n24611 );
xor ( n24848 , n24615 , n24616 );
xor ( n24849 , n24848 , n24618 );
and ( n24850 , n24847 , n24849 );
xor ( n24851 , n24691 , n24692 );
xor ( n24852 , n24851 , n24694 );
and ( n24853 , n24849 , n24852 );
and ( n24854 , n24847 , n24852 );
or ( n24855 , n24850 , n24853 , n24854 );
and ( n24856 , n24845 , n24855 );
and ( n24857 , n22542 , n22987 );
and ( n24858 , n22354 , n23508 );
and ( n24859 , n24857 , n24858 );
and ( n24860 , n22035 , n24540 );
and ( n24861 , n24858 , n24860 );
and ( n24862 , n24857 , n24860 );
or ( n24863 , n24859 , n24861 , n24862 );
and ( n24864 , n24546 , n20949 );
and ( n24865 , n22702 , n22562 );
and ( n24866 , n24864 , n24865 );
and ( n24867 , n22232 , n23758 );
and ( n24868 , n24865 , n24867 );
and ( n24869 , n24864 , n24867 );
or ( n24870 , n24866 , n24868 , n24869 );
and ( n24871 , n24863 , n24870 );
xor ( n24872 , n24685 , n24686 );
xor ( n24873 , n24872 , n24688 );
and ( n24874 , n24870 , n24873 );
and ( n24875 , n24863 , n24873 );
or ( n24876 , n24871 , n24874 , n24875 );
xor ( n24877 , n24625 , n24626 );
xor ( n24878 , n24877 , n24628 );
or ( n24879 , n24876 , n24878 );
and ( n24880 , n24855 , n24879 );
and ( n24881 , n24845 , n24879 );
or ( n24882 , n24856 , n24880 , n24881 );
and ( n24883 , n24052 , n21039 );
and ( n24884 , n23483 , n21429 );
and ( n24885 , n24883 , n24884 );
and ( n24886 , n23336 , n21527 );
and ( n24887 , n24884 , n24886 );
and ( n24888 , n24883 , n24886 );
or ( n24889 , n24885 , n24887 , n24888 );
xor ( n24890 , n24709 , n24710 );
xor ( n24891 , n24890 , n24713 );
and ( n24892 , n24889 , n24891 );
xor ( n24893 , n24738 , n24745 );
xor ( n24894 , n24893 , n24748 );
and ( n24895 , n24891 , n24894 );
and ( n24896 , n24889 , n24894 );
or ( n24897 , n24892 , n24895 , n24896 );
and ( n24898 , n24337 , n21039 );
and ( n24899 , n23620 , n21429 );
and ( n24900 , n24898 , n24899 );
and ( n24901 , n23336 , n21666 );
and ( n24902 , n24899 , n24901 );
and ( n24903 , n24898 , n24901 );
or ( n24904 , n24900 , n24902 , n24903 );
xor ( n24905 , n24779 , n24780 );
xor ( n24906 , n24905 , n24782 );
or ( n24907 , n24904 , n24906 );
and ( n24908 , n22351 , n22987 );
and ( n24909 , n22116 , n23758 );
and ( n24910 , n24908 , n24909 );
xor ( n24911 , n24764 , n24765 );
xor ( n24912 , n24911 , n24767 );
and ( n24913 , n24909 , n24912 );
and ( n24914 , n24908 , n24912 );
or ( n24915 , n24910 , n24913 , n24914 );
and ( n24916 , n24907 , n24915 );
xor ( n24917 , n24732 , n24733 );
xor ( n24918 , n24917 , n24735 );
xor ( n24919 , n24739 , n24740 );
xor ( n24920 , n24919 , n24742 );
and ( n24921 , n24918 , n24920 );
and ( n24922 , n22116 , n24064 );
buf ( n24923 , n21836 );
or ( n24924 , n24922 , n24923 );
and ( n24925 , n24920 , n24924 );
and ( n24926 , n24918 , n24924 );
or ( n24927 , n24921 , n24925 , n24926 );
and ( n24928 , n24915 , n24927 );
and ( n24929 , n24907 , n24927 );
or ( n24930 , n24916 , n24928 , n24929 );
and ( n24931 , n24897 , n24930 );
xor ( n24932 , n24726 , n24728 );
xor ( n24933 , n24932 , n24751 );
and ( n24934 , n24930 , n24933 );
and ( n24935 , n24897 , n24933 );
or ( n24936 , n24931 , n24934 , n24935 );
and ( n24937 , n24882 , n24936 );
xor ( n24938 , n24681 , n24683 );
xor ( n24939 , n24938 , n24705 );
and ( n24940 , n24936 , n24939 );
and ( n24941 , n24882 , n24939 );
or ( n24942 , n24937 , n24940 , n24941 );
and ( n24943 , n24843 , n24942 );
xor ( n24944 , n24670 , n24672 );
xor ( n24945 , n24944 , n24675 );
and ( n24946 , n24942 , n24945 );
and ( n24947 , n24843 , n24945 );
or ( n24948 , n24943 , n24946 , n24947 );
and ( n24949 , n24829 , n24948 );
and ( n24950 , n24827 , n24948 );
or ( n24951 , n24830 , n24949 , n24950 );
and ( n24952 , n24825 , n24951 );
xor ( n24953 , n24667 , n24806 );
xor ( n24954 , n24953 , n24809 );
and ( n24955 , n24951 , n24954 );
and ( n24956 , n24825 , n24954 );
or ( n24957 , n24952 , n24955 , n24956 );
and ( n24958 , n24823 , n24957 );
xor ( n24959 , n24662 , n24664 );
xor ( n24960 , n24959 , n24812 );
and ( n24961 , n24957 , n24960 );
and ( n24962 , n24823 , n24960 );
or ( n24963 , n24958 , n24961 , n24962 );
xor ( n24964 , n24474 , n24476 );
xor ( n24965 , n24964 , n24815 );
and ( n24966 , n24963 , n24965 );
xor ( n24967 , n24668 , n24678 );
xor ( n24968 , n24967 , n24803 );
xor ( n24969 , n24708 , n24797 );
xor ( n24970 , n24969 , n24800 );
xor ( n24971 , n24724 , n24754 );
xor ( n24972 , n24971 , n24794 );
xor ( n24973 , n24763 , n24788 );
xor ( n24974 , n24973 , n24791 );
xor ( n24975 , n24837 , n24839 );
and ( n24976 , n24974 , n24975 );
xor ( n24977 , n24756 , n24757 );
xor ( n24978 , n24977 , n24760 );
xor ( n24979 , n24770 , n24777 );
xor ( n24980 , n24979 , n24785 );
and ( n24981 , n24978 , n24980 );
xor ( n24982 , n24847 , n24849 );
xor ( n24983 , n24982 , n24852 );
and ( n24984 , n24980 , n24983 );
and ( n24985 , n24978 , n24983 );
or ( n24986 , n24981 , n24984 , n24985 );
and ( n24987 , n24975 , n24986 );
and ( n24988 , n24974 , n24986 );
or ( n24989 , n24976 , n24987 , n24988 );
and ( n24990 , n24972 , n24989 );
xnor ( n24991 , n24876 , n24878 );
buf ( n24992 , n15236 );
buf ( n24993 , n24992 );
and ( n24994 , n24993 , n20877 );
and ( n24995 , n23903 , n21178 );
and ( n24996 , n24994 , n24995 );
and ( n24997 , n23483 , n21527 );
and ( n24998 , n24995 , n24997 );
and ( n24999 , n24994 , n24997 );
or ( n25000 , n24996 , n24998 , n24999 );
and ( n25001 , n22351 , n23508 );
and ( n25002 , n22232 , n24064 );
and ( n25003 , n25001 , n25002 );
and ( n25004 , n22116 , n24540 );
and ( n25005 , n25002 , n25004 );
and ( n25006 , n25001 , n25004 );
or ( n25007 , n25003 , n25005 , n25006 );
and ( n25008 , n24052 , n21085 );
and ( n25009 , n25007 , n25008 );
and ( n25010 , n23089 , n21990 );
and ( n25011 , n25008 , n25010 );
and ( n25012 , n25007 , n25010 );
or ( n25013 , n25009 , n25011 , n25012 );
and ( n25014 , n25000 , n25013 );
xor ( n25015 , n24771 , n24772 );
xor ( n25016 , n25015 , n24774 );
and ( n25017 , n25013 , n25016 );
and ( n25018 , n25000 , n25016 );
or ( n25019 , n25014 , n25017 , n25018 );
and ( n25020 , n24991 , n25019 );
xor ( n25021 , n24883 , n24884 );
xor ( n25022 , n25021 , n24886 );
xnor ( n25023 , n24904 , n24906 );
and ( n25024 , n25022 , n25023 );
buf ( n25025 , n20257 );
buf ( n25026 , n25025 );
and ( n25027 , n21914 , n25026 );
xor ( n25028 , n24857 , n24858 );
xor ( n25029 , n25028 , n24860 );
and ( n25030 , n25027 , n25029 );
xor ( n25031 , n24898 , n24899 );
xor ( n25032 , n25031 , n24901 );
and ( n25033 , n25029 , n25032 );
and ( n25034 , n25027 , n25032 );
or ( n25035 , n25030 , n25033 , n25034 );
and ( n25036 , n25023 , n25035 );
and ( n25037 , n25022 , n25035 );
or ( n25038 , n25024 , n25036 , n25037 );
and ( n25039 , n25019 , n25038 );
and ( n25040 , n24991 , n25038 );
or ( n25041 , n25020 , n25039 , n25040 );
xnor ( n25042 , n24922 , n24923 );
and ( n25043 , n24624 , n20949 );
and ( n25044 , n22824 , n22562 );
and ( n25045 , n25043 , n25044 );
and ( n25046 , n22354 , n23758 );
and ( n25047 , n25044 , n25046 );
and ( n25048 , n25043 , n25046 );
or ( n25049 , n25045 , n25047 , n25048 );
and ( n25050 , n25042 , n25049 );
and ( n25051 , n24546 , n21039 );
and ( n25052 , n23742 , n21429 );
and ( n25053 , n25051 , n25052 );
and ( n25054 , n23620 , n21527 );
and ( n25055 , n25052 , n25054 );
and ( n25056 , n25051 , n25054 );
or ( n25057 , n25053 , n25055 , n25056 );
and ( n25058 , n25049 , n25057 );
and ( n25059 , n25042 , n25057 );
or ( n25060 , n25050 , n25058 , n25059 );
xor ( n25061 , n24908 , n24909 );
xor ( n25062 , n25061 , n24912 );
and ( n25063 , n25060 , n25062 );
xor ( n25064 , n24918 , n24920 );
xor ( n25065 , n25064 , n24924 );
and ( n25066 , n25062 , n25065 );
and ( n25067 , n25060 , n25065 );
or ( n25068 , n25063 , n25066 , n25067 );
xor ( n25069 , n24889 , n24891 );
xor ( n25070 , n25069 , n24894 );
and ( n25071 , n25068 , n25070 );
xor ( n25072 , n24907 , n24915 );
xor ( n25073 , n25072 , n24927 );
and ( n25074 , n25070 , n25073 );
and ( n25075 , n25068 , n25073 );
or ( n25076 , n25071 , n25074 , n25075 );
and ( n25077 , n25041 , n25076 );
xor ( n25078 , n24845 , n24855 );
xor ( n25079 , n25078 , n24879 );
and ( n25080 , n25076 , n25079 );
and ( n25081 , n25041 , n25079 );
or ( n25082 , n25077 , n25080 , n25081 );
and ( n25083 , n24989 , n25082 );
and ( n25084 , n24972 , n25082 );
or ( n25085 , n24990 , n25083 , n25084 );
and ( n25086 , n24970 , n25085 );
xor ( n25087 , n24843 , n24942 );
xor ( n25088 , n25087 , n24945 );
and ( n25089 , n25085 , n25088 );
and ( n25090 , n24970 , n25088 );
or ( n25091 , n25086 , n25089 , n25090 );
and ( n25092 , n24968 , n25091 );
xor ( n25093 , n24827 , n24829 );
xor ( n25094 , n25093 , n24948 );
and ( n25095 , n25091 , n25094 );
and ( n25096 , n24968 , n25094 );
or ( n25097 , n25092 , n25095 , n25096 );
xor ( n25098 , n24825 , n24951 );
xor ( n25099 , n25098 , n24954 );
or ( n25100 , n25097 , n25099 );
xor ( n25101 , n24823 , n24957 );
xor ( n25102 , n25101 , n24960 );
or ( n25103 , n25100 , n25102 );
and ( n25104 , n24965 , n25103 );
and ( n25105 , n24963 , n25103 );
or ( n25106 , n24966 , n25104 , n25105 );
and ( n25107 , n24820 , n25106 );
and ( n25108 , n24818 , n25106 );
or ( n25109 , n24821 , n25107 , n25108 );
or ( n25110 , n24333 , n25109 );
or ( n25111 , n24331 , n25110 );
or ( n25112 , n24329 , n25111 );
or ( n25113 , n24327 , n25112 );
or ( n25114 , n24325 , n25113 );
or ( n25115 , n24323 , n25114 );
or ( n25116 , n24321 , n25115 );
or ( n25117 , n24319 , n25116 );
or ( n25118 , n24317 , n25117 );
or ( n25119 , n24315 , n25118 );
or ( n25120 , n24313 , n25119 );
or ( n25121 , n24311 , n25120 );
or ( n25122 , n24309 , n25121 );
or ( n25123 , n24307 , n25122 );
or ( n25124 , n24305 , n25123 );
or ( n25125 , n24303 , n25124 );
or ( n25126 , n24301 , n25125 );
or ( n25127 , n24299 , n25126 );
or ( n25128 , n24297 , n25127 );
or ( n25129 , n24295 , n25128 );
or ( n25130 , n24293 , n25129 );
or ( n25131 , n24291 , n25130 );
or ( n25132 , n24289 , n25131 );
or ( n25133 , n24287 , n25132 );
or ( n25134 , n24285 , n25133 );
or ( n25135 , n24283 , n25134 );
or ( n25136 , n24281 , n25135 );
or ( n25137 , n24279 , n25136 );
or ( n25138 , n24277 , n25137 );
or ( n25139 , n24275 , n25138 );
or ( n25140 , n24273 , n25139 );
and ( n25141 , n24271 , n25140 );
xor ( n25142 , n24271 , n25140 );
xnor ( n25143 , n24273 , n25139 );
xnor ( n25144 , n24275 , n25138 );
xnor ( n25145 , n24277 , n25137 );
xnor ( n25146 , n24279 , n25136 );
xnor ( n25147 , n24281 , n25135 );
xnor ( n25148 , n24283 , n25134 );
xnor ( n25149 , n24285 , n25133 );
xnor ( n25150 , n24287 , n25132 );
xnor ( n25151 , n24289 , n25131 );
xnor ( n25152 , n24291 , n25130 );
xnor ( n25153 , n24293 , n25129 );
xnor ( n25154 , n24295 , n25128 );
xnor ( n25155 , n24297 , n25127 );
xnor ( n25156 , n24299 , n25126 );
xnor ( n25157 , n24301 , n25125 );
xnor ( n25158 , n24303 , n25124 );
xnor ( n25159 , n24305 , n25123 );
xnor ( n25160 , n24307 , n25122 );
xnor ( n25161 , n24309 , n25121 );
xnor ( n25162 , n24311 , n25120 );
xnor ( n25163 , n24313 , n25119 );
xnor ( n25164 , n24315 , n25118 );
xnor ( n25165 , n24317 , n25117 );
xnor ( n25166 , n24319 , n25116 );
xnor ( n25167 , n24321 , n25115 );
xnor ( n25168 , n24323 , n25114 );
xnor ( n25169 , n24325 , n25113 );
xnor ( n25170 , n24327 , n25112 );
xnor ( n25171 , n24329 , n25111 );
xnor ( n25172 , n24331 , n25110 );
xnor ( n25173 , n24333 , n25109 );
xor ( n25174 , n24818 , n24820 );
xor ( n25175 , n25174 , n25106 );
not ( n25176 , n25175 );
xor ( n25177 , n24963 , n24965 );
xor ( n25178 , n25177 , n25103 );
not ( n25179 , n25178 );
xnor ( n25180 , n25100 , n25102 );
xnor ( n25181 , n25097 , n25099 );
xor ( n25182 , n24968 , n25091 );
xor ( n25183 , n25182 , n25094 );
xor ( n25184 , n24832 , n24834 );
xor ( n25185 , n25184 , n24840 );
xor ( n25186 , n24882 , n24936 );
xor ( n25187 , n25186 , n24939 );
and ( n25188 , n25185 , n25187 );
xor ( n25189 , n24897 , n24930 );
xor ( n25190 , n25189 , n24933 );
and ( n25191 , n24624 , n20909 );
and ( n25192 , n23742 , n21296 );
and ( n25193 , n25191 , n25192 );
and ( n25194 , n22824 , n22337 );
and ( n25195 , n25192 , n25194 );
and ( n25196 , n25191 , n25194 );
or ( n25197 , n25193 , n25195 , n25196 );
and ( n25198 , n24731 , n20890 );
and ( n25199 , n23215 , n21827 );
and ( n25200 , n25198 , n25199 );
and ( n25201 , n22936 , n22172 );
and ( n25202 , n25199 , n25201 );
and ( n25203 , n25198 , n25201 );
or ( n25204 , n25200 , n25202 , n25203 );
and ( n25205 , n25197 , n25204 );
and ( n25206 , n22035 , n25026 );
buf ( n25207 , n25206 );
and ( n25208 , n22589 , n22784 );
and ( n25209 , n25207 , n25208 );
and ( n25210 , n22351 , n23322 );
and ( n25211 , n25208 , n25210 );
and ( n25212 , n25207 , n25210 );
or ( n25213 , n25209 , n25211 , n25212 );
and ( n25214 , n25204 , n25213 );
and ( n25215 , n25197 , n25213 );
or ( n25216 , n25205 , n25214 , n25215 );
xor ( n25217 , n25000 , n25013 );
xor ( n25218 , n25217 , n25016 );
buf ( n25219 , n15630 );
buf ( n25220 , n25219 );
and ( n25221 , n25220 , n20877 );
and ( n25222 , n24337 , n21085 );
and ( n25223 , n25221 , n25222 );
and ( n25224 , n24052 , n21178 );
and ( n25225 , n25222 , n25224 );
and ( n25226 , n25221 , n25224 );
or ( n25227 , n25223 , n25225 , n25226 );
xor ( n25228 , n25191 , n25192 );
xor ( n25229 , n25228 , n25194 );
xor ( n25230 , n25227 , n25229 );
xor ( n25231 , n25198 , n25199 );
xor ( n25232 , n25231 , n25201 );
xor ( n25233 , n25230 , n25232 );
and ( n25234 , n23903 , n21296 );
and ( n25235 , n22702 , n22784 );
xor ( n25236 , n25234 , n25235 );
and ( n25237 , n22589 , n22987 );
xor ( n25238 , n25236 , n25237 );
and ( n25239 , n24731 , n20909 );
and ( n25240 , n23089 , n22172 );
xor ( n25241 , n25239 , n25240 );
and ( n25242 , n22936 , n22337 );
xor ( n25243 , n25241 , n25242 );
and ( n25244 , n25238 , n25243 );
and ( n25245 , n24993 , n20890 );
and ( n25246 , n23336 , n21827 );
xor ( n25247 , n25245 , n25246 );
and ( n25248 , n23215 , n21990 );
xor ( n25249 , n25247 , n25248 );
and ( n25250 , n25243 , n25249 );
and ( n25251 , n25238 , n25249 );
or ( n25252 , n25244 , n25250 , n25251 );
and ( n25253 , n25233 , n25252 );
and ( n25254 , n22936 , n22562 );
and ( n25255 , n22702 , n22987 );
and ( n25256 , n25254 , n25255 );
and ( n25257 , n22589 , n23322 );
and ( n25258 , n25255 , n25257 );
and ( n25259 , n25254 , n25257 );
or ( n25260 , n25256 , n25258 , n25259 );
and ( n25261 , n24731 , n20949 );
and ( n25262 , n22351 , n23758 );
and ( n25263 , n25261 , n25262 );
buf ( n25264 , n21914 );
not ( n25265 , n25264 );
and ( n25266 , n25262 , n25265 );
and ( n25267 , n25261 , n25265 );
or ( n25268 , n25263 , n25266 , n25267 );
and ( n25269 , n25260 , n25268 );
xor ( n25270 , n25001 , n25002 );
xor ( n25271 , n25270 , n25004 );
and ( n25272 , n25268 , n25271 );
and ( n25273 , n25260 , n25271 );
or ( n25274 , n25269 , n25272 , n25273 );
and ( n25275 , n25252 , n25274 );
and ( n25276 , n25233 , n25274 );
or ( n25277 , n25253 , n25275 , n25276 );
and ( n25278 , n25218 , n25277 );
and ( n25279 , n23483 , n21666 );
and ( n25280 , n22232 , n24540 );
and ( n25281 , n22116 , n25026 );
and ( n25282 , n25280 , n25281 );
buf ( n25283 , n20262 );
buf ( n25284 , n25283 );
and ( n25285 , n22035 , n25284 );
and ( n25286 , n25281 , n25285 );
and ( n25287 , n25280 , n25285 );
or ( n25288 , n25282 , n25286 , n25287 );
and ( n25289 , n25279 , n25288 );
and ( n25290 , n24624 , n21039 );
and ( n25291 , n23903 , n21429 );
and ( n25292 , n25290 , n25291 );
and ( n25293 , n23336 , n21990 );
and ( n25294 , n25291 , n25293 );
and ( n25295 , n25290 , n25293 );
or ( n25296 , n25292 , n25294 , n25295 );
and ( n25297 , n25288 , n25296 );
and ( n25298 , n25279 , n25296 );
or ( n25299 , n25289 , n25297 , n25298 );
xor ( n25300 , n25027 , n25029 );
xor ( n25301 , n25300 , n25032 );
and ( n25302 , n25299 , n25301 );
xor ( n25303 , n25042 , n25049 );
xor ( n25304 , n25303 , n25057 );
and ( n25305 , n25301 , n25304 );
and ( n25306 , n25299 , n25304 );
or ( n25307 , n25302 , n25305 , n25306 );
and ( n25308 , n25277 , n25307 );
and ( n25309 , n25218 , n25307 );
or ( n25310 , n25278 , n25308 , n25309 );
and ( n25311 , n25216 , n25310 );
xor ( n25312 , n24978 , n24980 );
xor ( n25313 , n25312 , n24983 );
and ( n25314 , n25310 , n25313 );
and ( n25315 , n25216 , n25313 );
or ( n25316 , n25311 , n25314 , n25315 );
and ( n25317 , n25190 , n25316 );
xor ( n25318 , n24974 , n24975 );
xor ( n25319 , n25318 , n24986 );
and ( n25320 , n25316 , n25319 );
and ( n25321 , n25190 , n25319 );
or ( n25322 , n25317 , n25320 , n25321 );
and ( n25323 , n25187 , n25322 );
and ( n25324 , n25185 , n25322 );
or ( n25325 , n25188 , n25323 , n25324 );
xor ( n25326 , n24970 , n25085 );
xor ( n25327 , n25326 , n25088 );
and ( n25328 , n25325 , n25327 );
xor ( n25329 , n24972 , n24989 );
xor ( n25330 , n25329 , n25082 );
xor ( n25331 , n25041 , n25076 );
xor ( n25332 , n25331 , n25079 );
xor ( n25333 , n24991 , n25019 );
xor ( n25334 , n25333 , n25038 );
xor ( n25335 , n25068 , n25070 );
xor ( n25336 , n25335 , n25073 );
and ( n25337 , n25334 , n25336 );
and ( n25338 , n25227 , n25229 );
and ( n25339 , n25229 , n25232 );
and ( n25340 , n25227 , n25232 );
or ( n25341 , n25338 , n25339 , n25340 );
and ( n25342 , n25239 , n25240 );
and ( n25343 , n25240 , n25242 );
and ( n25344 , n25239 , n25242 );
or ( n25345 , n25342 , n25343 , n25344 );
buf ( n25346 , n25264 );
and ( n25347 , n22542 , n23322 );
and ( n25348 , n25346 , n25347 );
not ( n25349 , n25206 );
and ( n25350 , n25347 , n25349 );
and ( n25351 , n25346 , n25349 );
or ( n25352 , n25348 , n25350 , n25351 );
and ( n25353 , n25345 , n25352 );
xor ( n25354 , n25207 , n25208 );
xor ( n25355 , n25354 , n25210 );
and ( n25356 , n25352 , n25355 );
and ( n25357 , n25345 , n25355 );
or ( n25358 , n25353 , n25356 , n25357 );
and ( n25359 , n25341 , n25358 );
xor ( n25360 , n24863 , n24870 );
xor ( n25361 , n25360 , n24873 );
and ( n25362 , n25358 , n25361 );
and ( n25363 , n25341 , n25361 );
or ( n25364 , n25359 , n25362 , n25363 );
and ( n25365 , n25336 , n25364 );
and ( n25366 , n25334 , n25364 );
or ( n25367 , n25337 , n25365 , n25366 );
and ( n25368 , n25332 , n25367 );
and ( n25369 , n25234 , n25235 );
and ( n25370 , n25235 , n25237 );
and ( n25371 , n25234 , n25237 );
or ( n25372 , n25369 , n25370 , n25371 );
and ( n25373 , n25245 , n25246 );
and ( n25374 , n25246 , n25248 );
and ( n25375 , n25245 , n25248 );
or ( n25376 , n25373 , n25374 , n25375 );
and ( n25377 , n25372 , n25376 );
xor ( n25378 , n24864 , n24865 );
xor ( n25379 , n25378 , n24867 );
and ( n25380 , n25376 , n25379 );
and ( n25381 , n25372 , n25379 );
or ( n25382 , n25377 , n25380 , n25381 );
not ( n25383 , n25382 );
xor ( n25384 , n25197 , n25204 );
xor ( n25385 , n25384 , n25213 );
and ( n25386 , n25383 , n25385 );
buf ( n25387 , n25382 );
and ( n25388 , n25386 , n25387 );
xor ( n25389 , n25022 , n25023 );
xor ( n25390 , n25389 , n25035 );
xor ( n25391 , n25060 , n25062 );
xor ( n25392 , n25391 , n25065 );
and ( n25393 , n25390 , n25392 );
and ( n25394 , n25220 , n20890 );
and ( n25395 , n24993 , n20909 );
and ( n25396 , n25394 , n25395 );
and ( n25397 , n23215 , n22172 );
and ( n25398 , n25395 , n25397 );
and ( n25399 , n25394 , n25397 );
or ( n25400 , n25396 , n25398 , n25399 );
xor ( n25401 , n25043 , n25044 );
xor ( n25402 , n25401 , n25046 );
and ( n25403 , n25400 , n25402 );
xor ( n25404 , n25346 , n25347 );
xor ( n25405 , n25404 , n25349 );
and ( n25406 , n25402 , n25405 );
and ( n25407 , n25400 , n25405 );
or ( n25408 , n25403 , n25406 , n25407 );
xor ( n25409 , n24994 , n24995 );
xor ( n25410 , n25409 , n24997 );
and ( n25411 , n25408 , n25410 );
xor ( n25412 , n25007 , n25008 );
xor ( n25413 , n25412 , n25010 );
and ( n25414 , n25410 , n25413 );
and ( n25415 , n25408 , n25413 );
or ( n25416 , n25411 , n25414 , n25415 );
and ( n25417 , n25392 , n25416 );
and ( n25418 , n25390 , n25416 );
or ( n25419 , n25393 , n25417 , n25418 );
and ( n25420 , n25387 , n25419 );
and ( n25421 , n25386 , n25419 );
or ( n25422 , n25388 , n25420 , n25421 );
and ( n25423 , n25367 , n25422 );
and ( n25424 , n25332 , n25422 );
or ( n25425 , n25368 , n25423 , n25424 );
and ( n25426 , n25330 , n25425 );
xor ( n25427 , n25185 , n25187 );
xor ( n25428 , n25427 , n25322 );
and ( n25429 , n25425 , n25428 );
and ( n25430 , n25330 , n25428 );
or ( n25431 , n25426 , n25429 , n25430 );
and ( n25432 , n25327 , n25431 );
and ( n25433 , n25325 , n25431 );
or ( n25434 , n25328 , n25432 , n25433 );
and ( n25435 , n25183 , n25434 );
xor ( n25436 , n25183 , n25434 );
xor ( n25437 , n25325 , n25327 );
xor ( n25438 , n25437 , n25431 );
xor ( n25439 , n25190 , n25316 );
xor ( n25440 , n25439 , n25319 );
xor ( n25441 , n25216 , n25310 );
xor ( n25442 , n25441 , n25313 );
and ( n25443 , n25220 , n20909 );
and ( n25444 , n24337 , n21296 );
and ( n25445 , n25443 , n25444 );
and ( n25446 , n23215 , n22337 );
and ( n25447 , n25444 , n25446 );
and ( n25448 , n25443 , n25446 );
or ( n25449 , n25445 , n25447 , n25448 );
buf ( n25450 , n15810 );
buf ( n25451 , n25450 );
and ( n25452 , n25451 , n20890 );
and ( n25453 , n23620 , n21827 );
and ( n25454 , n25452 , n25453 );
and ( n25455 , n23336 , n22172 );
and ( n25456 , n25453 , n25455 );
and ( n25457 , n25452 , n25455 );
or ( n25458 , n25454 , n25456 , n25457 );
and ( n25459 , n25449 , n25458 );
xor ( n25460 , n25261 , n25262 );
xor ( n25461 , n25460 , n25265 );
and ( n25462 , n25458 , n25461 );
and ( n25463 , n25449 , n25461 );
or ( n25464 , n25459 , n25462 , n25463 );
xor ( n25465 , n25221 , n25222 );
xor ( n25466 , n25465 , n25224 );
and ( n25467 , n25464 , n25466 );
xor ( n25468 , n25260 , n25268 );
xor ( n25469 , n25468 , n25271 );
and ( n25470 , n25466 , n25469 );
and ( n25471 , n25464 , n25469 );
or ( n25472 , n25467 , n25470 , n25471 );
xor ( n25473 , n25238 , n25243 );
xor ( n25474 , n25473 , n25249 );
and ( n25475 , n22542 , n23508 );
and ( n25476 , n22354 , n24064 );
and ( n25477 , n25475 , n25476 );
and ( n25478 , n25451 , n20877 );
and ( n25479 , n23620 , n21666 );
xor ( n25480 , n25478 , n25479 );
and ( n25481 , n23483 , n21827 );
xor ( n25482 , n25480 , n25481 );
and ( n25483 , n25476 , n25482 );
and ( n25484 , n25475 , n25482 );
or ( n25485 , n25477 , n25483 , n25484 );
and ( n25486 , n25474 , n25485 );
and ( n25487 , n22351 , n24064 );
and ( n25488 , n22354 , n24540 );
and ( n25489 , n25487 , n25488 );
and ( n25490 , n22116 , n25284 );
and ( n25491 , n25488 , n25490 );
and ( n25492 , n25487 , n25490 );
or ( n25493 , n25489 , n25491 , n25492 );
and ( n25494 , n24731 , n21039 );
and ( n25495 , n22589 , n23508 );
and ( n25496 , n25494 , n25495 );
and ( n25497 , n22232 , n25026 );
and ( n25498 , n25495 , n25497 );
and ( n25499 , n25494 , n25497 );
or ( n25500 , n25496 , n25498 , n25499 );
and ( n25501 , n25493 , n25500 );
xor ( n25502 , n25290 , n25291 );
xor ( n25503 , n25502 , n25293 );
and ( n25504 , n25500 , n25503 );
and ( n25505 , n25493 , n25503 );
or ( n25506 , n25501 , n25504 , n25505 );
and ( n25507 , n25485 , n25506 );
and ( n25508 , n25474 , n25506 );
or ( n25509 , n25486 , n25507 , n25508 );
and ( n25510 , n25472 , n25509 );
xor ( n25511 , n25233 , n25252 );
xor ( n25512 , n25511 , n25274 );
and ( n25513 , n25509 , n25512 );
and ( n25514 , n25472 , n25512 );
or ( n25515 , n25510 , n25513 , n25514 );
xor ( n25516 , n25218 , n25277 );
xor ( n25517 , n25516 , n25307 );
and ( n25518 , n25515 , n25517 );
xor ( n25519 , n25341 , n25358 );
xor ( n25520 , n25519 , n25361 );
and ( n25521 , n25517 , n25520 );
and ( n25522 , n25515 , n25520 );
or ( n25523 , n25518 , n25521 , n25522 );
and ( n25524 , n25442 , n25523 );
xor ( n25525 , n25383 , n25385 );
and ( n25526 , n24052 , n21296 );
and ( n25527 , n23089 , n22337 );
and ( n25528 , n25526 , n25527 );
and ( n25529 , n22824 , n22784 );
and ( n25530 , n25527 , n25529 );
and ( n25531 , n25526 , n25529 );
or ( n25532 , n25528 , n25530 , n25531 );
and ( n25533 , n25478 , n25479 );
and ( n25534 , n25479 , n25481 );
and ( n25535 , n25478 , n25481 );
or ( n25536 , n25533 , n25534 , n25535 );
and ( n25537 , n25532 , n25536 );
and ( n25538 , n24546 , n21085 );
and ( n25539 , n24337 , n21178 );
and ( n25540 , n25538 , n25539 );
and ( n25541 , n23742 , n21527 );
and ( n25542 , n25539 , n25541 );
and ( n25543 , n25538 , n25541 );
or ( n25544 , n25540 , n25542 , n25543 );
and ( n25545 , n25536 , n25544 );
and ( n25546 , n25532 , n25544 );
or ( n25547 , n25537 , n25545 , n25546 );
xor ( n25548 , n25372 , n25376 );
xor ( n25549 , n25548 , n25379 );
and ( n25550 , n25547 , n25549 );
xor ( n25551 , n25345 , n25352 );
xor ( n25552 , n25551 , n25355 );
and ( n25553 , n25549 , n25552 );
and ( n25554 , n25547 , n25552 );
or ( n25555 , n25550 , n25553 , n25554 );
and ( n25556 , n25525 , n25555 );
xor ( n25557 , n25299 , n25301 );
xor ( n25558 , n25557 , n25304 );
xor ( n25559 , n25408 , n25410 );
xor ( n25560 , n25559 , n25413 );
and ( n25561 , n25558 , n25560 );
and ( n25562 , n23089 , n22562 );
and ( n25563 , n22824 , n22987 );
and ( n25564 , n25562 , n25563 );
and ( n25565 , n22542 , n23758 );
and ( n25566 , n25563 , n25565 );
and ( n25567 , n25562 , n25565 );
or ( n25568 , n25564 , n25566 , n25567 );
and ( n25569 , n24993 , n20949 );
and ( n25570 , n22936 , n22784 );
and ( n25571 , n25569 , n25570 );
and ( n25572 , n22702 , n23322 );
and ( n25573 , n25570 , n25572 );
and ( n25574 , n25569 , n25572 );
or ( n25575 , n25571 , n25573 , n25574 );
and ( n25576 , n25568 , n25575 );
xor ( n25577 , n25280 , n25281 );
xor ( n25578 , n25577 , n25285 );
and ( n25579 , n25575 , n25578 );
and ( n25580 , n25568 , n25578 );
or ( n25581 , n25576 , n25579 , n25580 );
xor ( n25582 , n25051 , n25052 );
xor ( n25583 , n25582 , n25054 );
and ( n25584 , n25581 , n25583 );
xor ( n25585 , n25400 , n25402 );
xor ( n25586 , n25585 , n25405 );
and ( n25587 , n25583 , n25586 );
and ( n25588 , n25581 , n25586 );
or ( n25589 , n25584 , n25587 , n25588 );
and ( n25590 , n25560 , n25589 );
and ( n25591 , n25558 , n25589 );
or ( n25592 , n25561 , n25590 , n25591 );
and ( n25593 , n25555 , n25592 );
and ( n25594 , n25525 , n25592 );
or ( n25595 , n25556 , n25593 , n25594 );
and ( n25596 , n25523 , n25595 );
and ( n25597 , n25442 , n25595 );
or ( n25598 , n25524 , n25596 , n25597 );
and ( n25599 , n25440 , n25598 );
xor ( n25600 , n25332 , n25367 );
xor ( n25601 , n25600 , n25422 );
and ( n25602 , n25598 , n25601 );
and ( n25603 , n25440 , n25601 );
or ( n25604 , n25599 , n25602 , n25603 );
xor ( n25605 , n25330 , n25425 );
xor ( n25606 , n25605 , n25428 );
and ( n25607 , n25604 , n25606 );
xor ( n25608 , n25334 , n25336 );
xor ( n25609 , n25608 , n25364 );
xor ( n25610 , n25386 , n25387 );
xor ( n25611 , n25610 , n25419 );
and ( n25612 , n25609 , n25611 );
and ( n25613 , n22702 , n23508 );
and ( n25614 , n22354 , n25026 );
and ( n25615 , n25613 , n25614 );
buf ( n25616 , n20267 );
buf ( n25617 , n25616 );
and ( n25618 , n22116 , n25617 );
and ( n25619 , n25614 , n25618 );
and ( n25620 , n25613 , n25618 );
or ( n25621 , n25615 , n25619 , n25620 );
buf ( n25622 , n15972 );
buf ( n25623 , n25622 );
and ( n25624 , n25623 , n20877 );
and ( n25625 , n25621 , n25624 );
and ( n25626 , n24624 , n21085 );
and ( n25627 , n25624 , n25626 );
and ( n25628 , n25621 , n25626 );
or ( n25629 , n25625 , n25627 , n25628 );
xor ( n25630 , n25394 , n25395 );
xor ( n25631 , n25630 , n25397 );
and ( n25632 , n25629 , n25631 );
xor ( n25633 , n25254 , n25255 );
xor ( n25634 , n25633 , n25257 );
and ( n25635 , n25631 , n25634 );
and ( n25636 , n25629 , n25634 );
or ( n25637 , n25632 , n25635 , n25636 );
xor ( n25638 , n25532 , n25536 );
xor ( n25639 , n25638 , n25544 );
or ( n25640 , n25637 , n25639 );
xor ( n25641 , n25279 , n25288 );
xor ( n25642 , n25641 , n25296 );
and ( n25643 , n24546 , n21178 );
and ( n25644 , n23903 , n21527 );
and ( n25645 , n25643 , n25644 );
and ( n25646 , n23483 , n21990 );
and ( n25647 , n25644 , n25646 );
and ( n25648 , n25643 , n25646 );
or ( n25649 , n25645 , n25647 , n25648 );
and ( n25650 , n22542 , n24064 );
and ( n25651 , n22351 , n24540 );
and ( n25652 , n25650 , n25651 );
buf ( n25653 , n22035 );
not ( n25654 , n25653 );
and ( n25655 , n25651 , n25654 );
and ( n25656 , n25650 , n25654 );
or ( n25657 , n25652 , n25655 , n25656 );
and ( n25658 , n24052 , n21429 );
and ( n25659 , n25657 , n25658 );
and ( n25660 , n23742 , n21666 );
and ( n25661 , n25658 , n25660 );
and ( n25662 , n25657 , n25660 );
or ( n25663 , n25659 , n25661 , n25662 );
and ( n25664 , n25649 , n25663 );
xor ( n25665 , n25526 , n25527 );
xor ( n25666 , n25665 , n25529 );
and ( n25667 , n25663 , n25666 );
and ( n25668 , n25649 , n25666 );
or ( n25669 , n25664 , n25667 , n25668 );
and ( n25670 , n25642 , n25669 );
xor ( n25671 , n25568 , n25575 );
xor ( n25672 , n25671 , n25578 );
xor ( n25673 , n25449 , n25458 );
xor ( n25674 , n25673 , n25461 );
and ( n25675 , n25672 , n25674 );
and ( n25676 , n25669 , n25675 );
and ( n25677 , n25642 , n25675 );
or ( n25678 , n25670 , n25676 , n25677 );
and ( n25679 , n25640 , n25678 );
xor ( n25680 , n25472 , n25509 );
xor ( n25681 , n25680 , n25512 );
and ( n25682 , n25678 , n25681 );
and ( n25683 , n25640 , n25681 );
or ( n25684 , n25679 , n25682 , n25683 );
xor ( n25685 , n25390 , n25392 );
xor ( n25686 , n25685 , n25416 );
and ( n25687 , n25684 , n25686 );
xor ( n25688 , n25547 , n25549 );
xor ( n25689 , n25688 , n25552 );
and ( n25690 , n25220 , n20949 );
and ( n25691 , n23215 , n22562 );
and ( n25692 , n25690 , n25691 );
and ( n25693 , n22936 , n22987 );
and ( n25694 , n25691 , n25693 );
and ( n25695 , n25690 , n25693 );
or ( n25696 , n25692 , n25694 , n25695 );
and ( n25697 , n24546 , n21296 );
and ( n25698 , n23742 , n21827 );
and ( n25699 , n25697 , n25698 );
and ( n25700 , n22589 , n23758 );
and ( n25701 , n25698 , n25700 );
and ( n25702 , n25697 , n25700 );
or ( n25703 , n25699 , n25701 , n25702 );
and ( n25704 , n25696 , n25703 );
and ( n25705 , n22351 , n25026 );
buf ( n25706 , n25705 );
and ( n25707 , n22824 , n23322 );
and ( n25708 , n25706 , n25707 );
and ( n25709 , n22232 , n25284 );
and ( n25710 , n25707 , n25709 );
and ( n25711 , n25706 , n25709 );
or ( n25712 , n25708 , n25710 , n25711 );
and ( n25713 , n25703 , n25712 );
and ( n25714 , n25696 , n25712 );
or ( n25715 , n25704 , n25713 , n25714 );
and ( n25716 , n25623 , n20890 );
and ( n25717 , n25451 , n20909 );
and ( n25718 , n25716 , n25717 );
and ( n25719 , n23089 , n22784 );
and ( n25720 , n25717 , n25719 );
and ( n25721 , n25716 , n25719 );
or ( n25722 , n25718 , n25720 , n25721 );
xor ( n25723 , n25562 , n25563 );
xor ( n25724 , n25723 , n25565 );
and ( n25725 , n25722 , n25724 );
xor ( n25726 , n25569 , n25570 );
xor ( n25727 , n25726 , n25572 );
and ( n25728 , n25724 , n25727 );
and ( n25729 , n25722 , n25727 );
or ( n25730 , n25725 , n25728 , n25729 );
and ( n25731 , n25715 , n25730 );
xor ( n25732 , n25538 , n25539 );
xor ( n25733 , n25732 , n25541 );
and ( n25734 , n25730 , n25733 );
and ( n25735 , n25715 , n25733 );
or ( n25736 , n25731 , n25734 , n25735 );
xor ( n25737 , n25581 , n25583 );
xor ( n25738 , n25737 , n25586 );
or ( n25739 , n25736 , n25738 );
and ( n25740 , n25689 , n25739 );
buf ( n25741 , n16248 );
buf ( n25742 , n25741 );
and ( n25743 , n25742 , n20877 );
and ( n25744 , n24624 , n21178 );
and ( n25745 , n25743 , n25744 );
and ( n25746 , n24052 , n21527 );
and ( n25747 , n25744 , n25746 );
and ( n25748 , n25743 , n25746 );
or ( n25749 , n25745 , n25747 , n25748 );
xor ( n25750 , n25443 , n25444 );
xor ( n25751 , n25750 , n25446 );
and ( n25752 , n25749 , n25751 );
xor ( n25753 , n25657 , n25658 );
xor ( n25754 , n25753 , n25660 );
and ( n25755 , n25751 , n25754 );
and ( n25756 , n25749 , n25754 );
or ( n25757 , n25752 , n25755 , n25756 );
and ( n25758 , n23903 , n21666 );
and ( n25759 , n23483 , n22172 );
and ( n25760 , n25758 , n25759 );
and ( n25761 , n23336 , n22337 );
and ( n25762 , n25759 , n25761 );
and ( n25763 , n25758 , n25761 );
or ( n25764 , n25760 , n25762 , n25763 );
and ( n25765 , n24731 , n21085 );
and ( n25766 , n23620 , n21990 );
and ( n25767 , n25765 , n25766 );
xor ( n25768 , n25613 , n25614 );
xor ( n25769 , n25768 , n25618 );
and ( n25770 , n25766 , n25769 );
and ( n25771 , n25765 , n25769 );
or ( n25772 , n25767 , n25770 , n25771 );
and ( n25773 , n25764 , n25772 );
xor ( n25774 , n25452 , n25453 );
xor ( n25775 , n25774 , n25455 );
and ( n25776 , n25772 , n25775 );
and ( n25777 , n25764 , n25775 );
or ( n25778 , n25773 , n25776 , n25777 );
and ( n25779 , n25757 , n25778 );
xor ( n25780 , n25649 , n25663 );
xor ( n25781 , n25780 , n25666 );
and ( n25782 , n25778 , n25781 );
and ( n25783 , n25757 , n25781 );
or ( n25784 , n25779 , n25782 , n25783 );
xor ( n25785 , n25464 , n25466 );
xor ( n25786 , n25785 , n25469 );
and ( n25787 , n25784 , n25786 );
and ( n25788 , n25739 , n25787 );
and ( n25789 , n25689 , n25787 );
or ( n25790 , n25740 , n25788 , n25789 );
and ( n25791 , n25686 , n25790 );
and ( n25792 , n25684 , n25790 );
or ( n25793 , n25687 , n25791 , n25792 );
and ( n25794 , n25611 , n25793 );
and ( n25795 , n25609 , n25793 );
or ( n25796 , n25612 , n25794 , n25795 );
xor ( n25797 , n25440 , n25598 );
xor ( n25798 , n25797 , n25601 );
and ( n25799 , n25796 , n25798 );
xor ( n25800 , n25487 , n25488 );
xor ( n25801 , n25800 , n25490 );
xor ( n25802 , n25643 , n25644 );
xor ( n25803 , n25802 , n25646 );
and ( n25804 , n25801 , n25803 );
buf ( n25805 , n25653 );
and ( n25806 , n25803 , n25805 );
and ( n25807 , n25801 , n25805 );
or ( n25808 , n25804 , n25806 , n25807 );
xor ( n25809 , n25475 , n25476 );
xor ( n25810 , n25809 , n25482 );
and ( n25811 , n25808 , n25810 );
xor ( n25812 , n25493 , n25500 );
xor ( n25813 , n25812 , n25503 );
and ( n25814 , n25810 , n25813 );
and ( n25815 , n25808 , n25813 );
or ( n25816 , n25811 , n25814 , n25815 );
xor ( n25817 , n25474 , n25485 );
xor ( n25818 , n25817 , n25506 );
and ( n25819 , n25816 , n25818 );
xnor ( n25820 , n25637 , n25639 );
and ( n25821 , n25818 , n25820 );
and ( n25822 , n25816 , n25820 );
or ( n25823 , n25819 , n25821 , n25822 );
xor ( n25824 , n25558 , n25560 );
xor ( n25825 , n25824 , n25589 );
and ( n25826 , n25823 , n25825 );
xor ( n25827 , n25640 , n25678 );
xor ( n25828 , n25827 , n25681 );
and ( n25829 , n25825 , n25828 );
and ( n25830 , n25823 , n25828 );
or ( n25831 , n25826 , n25829 , n25830 );
xor ( n25832 , n25515 , n25517 );
xor ( n25833 , n25832 , n25520 );
and ( n25834 , n25831 , n25833 );
xor ( n25835 , n25525 , n25555 );
xor ( n25836 , n25835 , n25592 );
and ( n25837 , n25833 , n25836 );
and ( n25838 , n25831 , n25836 );
or ( n25839 , n25834 , n25837 , n25838 );
xor ( n25840 , n25442 , n25523 );
xor ( n25841 , n25840 , n25595 );
and ( n25842 , n25839 , n25841 );
xor ( n25843 , n25629 , n25631 );
xor ( n25844 , n25843 , n25634 );
xor ( n25845 , n25672 , n25674 );
and ( n25846 , n25844 , n25845 );
xor ( n25847 , n25494 , n25495 );
xor ( n25848 , n25847 , n25497 );
xor ( n25849 , n25621 , n25624 );
xor ( n25850 , n25849 , n25626 );
and ( n25851 , n25848 , n25850 );
xor ( n25852 , n25722 , n25724 );
xor ( n25853 , n25852 , n25727 );
and ( n25854 , n25850 , n25853 );
and ( n25855 , n25848 , n25853 );
or ( n25856 , n25851 , n25854 , n25855 );
and ( n25857 , n25845 , n25856 );
and ( n25858 , n25844 , n25856 );
or ( n25859 , n25846 , n25857 , n25858 );
xor ( n25860 , n25642 , n25669 );
xor ( n25861 , n25860 , n25675 );
and ( n25862 , n25859 , n25861 );
xnor ( n25863 , n25736 , n25738 );
and ( n25864 , n25861 , n25863 );
and ( n25865 , n25859 , n25863 );
or ( n25866 , n25862 , n25864 , n25865 );
xor ( n25867 , n25784 , n25786 );
and ( n25868 , n25451 , n20949 );
and ( n25869 , n23336 , n22562 );
and ( n25870 , n25868 , n25869 );
and ( n25871 , n22702 , n23758 );
and ( n25872 , n25869 , n25871 );
and ( n25873 , n25868 , n25871 );
or ( n25874 , n25870 , n25872 , n25873 );
and ( n25875 , n24993 , n21039 );
and ( n25876 , n25874 , n25875 );
and ( n25877 , n24337 , n21429 );
and ( n25878 , n25875 , n25877 );
and ( n25879 , n25874 , n25877 );
or ( n25880 , n25876 , n25878 , n25879 );
and ( n25881 , n25742 , n20890 );
and ( n25882 , n25623 , n20909 );
and ( n25883 , n25881 , n25882 );
and ( n25884 , n23620 , n22172 );
and ( n25885 , n25882 , n25884 );
and ( n25886 , n25881 , n25884 );
or ( n25887 , n25883 , n25885 , n25886 );
xor ( n25888 , n25690 , n25691 );
xor ( n25889 , n25888 , n25693 );
or ( n25890 , n25887 , n25889 );
and ( n25891 , n25880 , n25890 );
and ( n25892 , n22542 , n24540 );
and ( n25893 , n22354 , n25284 );
and ( n25894 , n25892 , n25893 );
and ( n25895 , n22232 , n25617 );
and ( n25896 , n25893 , n25895 );
and ( n25897 , n25892 , n25895 );
or ( n25898 , n25894 , n25896 , n25897 );
and ( n25899 , n22824 , n23508 );
and ( n25900 , n22589 , n24064 );
and ( n25901 , n25899 , n25900 );
not ( n25902 , n25705 );
and ( n25903 , n25900 , n25902 );
and ( n25904 , n25899 , n25902 );
or ( n25905 , n25901 , n25903 , n25904 );
and ( n25906 , n25898 , n25905 );
and ( n25907 , n25890 , n25906 );
and ( n25908 , n25880 , n25906 );
or ( n25909 , n25891 , n25907 , n25908 );
xor ( n25910 , n25808 , n25810 );
xor ( n25911 , n25910 , n25813 );
and ( n25912 , n25909 , n25911 );
xor ( n25913 , n25715 , n25730 );
xor ( n25914 , n25913 , n25733 );
and ( n25915 , n25911 , n25914 );
and ( n25916 , n25909 , n25914 );
or ( n25917 , n25912 , n25915 , n25916 );
and ( n25918 , n25867 , n25917 );
xor ( n25919 , n25757 , n25778 );
xor ( n25920 , n25919 , n25781 );
xor ( n25921 , n25697 , n25698 );
xor ( n25922 , n25921 , n25700 );
and ( n25923 , n24993 , n21085 );
and ( n25924 , n24731 , n21178 );
and ( n25925 , n25923 , n25924 );
and ( n25926 , n24337 , n21527 );
and ( n25927 , n25924 , n25926 );
and ( n25928 , n25923 , n25926 );
or ( n25929 , n25925 , n25927 , n25928 );
and ( n25930 , n25922 , n25929 );
and ( n25931 , n24052 , n21666 );
and ( n25932 , n23903 , n21827 );
or ( n25933 , n25931 , n25932 );
and ( n25934 , n25929 , n25933 );
and ( n25935 , n25922 , n25933 );
or ( n25936 , n25930 , n25934 , n25935 );
xor ( n25937 , n25801 , n25803 );
xor ( n25938 , n25937 , n25805 );
and ( n25939 , n25936 , n25938 );
xor ( n25940 , n25696 , n25703 );
xor ( n25941 , n25940 , n25712 );
and ( n25942 , n25938 , n25941 );
and ( n25943 , n25936 , n25941 );
or ( n25944 , n25939 , n25942 , n25943 );
and ( n25945 , n25920 , n25944 );
xor ( n25946 , n25749 , n25751 );
xor ( n25947 , n25946 , n25754 );
xor ( n25948 , n25764 , n25772 );
xor ( n25949 , n25948 , n25775 );
and ( n25950 , n25947 , n25949 );
and ( n25951 , n22936 , n23508 );
and ( n25952 , n22589 , n24540 );
and ( n25953 , n25951 , n25952 );
and ( n25954 , n22351 , n25284 );
and ( n25955 , n25952 , n25954 );
and ( n25956 , n25951 , n25954 );
or ( n25957 , n25953 , n25955 , n25956 );
buf ( n25958 , n16310 );
buf ( n25959 , n25958 );
and ( n25960 , n25959 , n20877 );
and ( n25961 , n25957 , n25960 );
and ( n25962 , n23742 , n21990 );
and ( n25963 , n25960 , n25962 );
and ( n25964 , n25957 , n25962 );
or ( n25965 , n25961 , n25963 , n25964 );
xor ( n25966 , n25758 , n25759 );
xor ( n25967 , n25966 , n25761 );
and ( n25968 , n25965 , n25967 );
xor ( n25969 , n25716 , n25717 );
xor ( n25970 , n25969 , n25719 );
and ( n25971 , n25967 , n25970 );
and ( n25972 , n25965 , n25970 );
or ( n25973 , n25968 , n25971 , n25972 );
and ( n25974 , n25949 , n25973 );
and ( n25975 , n25947 , n25973 );
or ( n25976 , n25950 , n25974 , n25975 );
and ( n25977 , n25944 , n25976 );
and ( n25978 , n25920 , n25976 );
or ( n25979 , n25945 , n25977 , n25978 );
and ( n25980 , n25917 , n25979 );
and ( n25981 , n25867 , n25979 );
or ( n25982 , n25918 , n25980 , n25981 );
and ( n25983 , n25866 , n25982 );
xor ( n25984 , n25689 , n25739 );
xor ( n25985 , n25984 , n25787 );
and ( n25986 , n25982 , n25985 );
and ( n25987 , n25866 , n25985 );
or ( n25988 , n25983 , n25986 , n25987 );
xor ( n25989 , n25684 , n25686 );
xor ( n25990 , n25989 , n25790 );
and ( n25991 , n25988 , n25990 );
xor ( n25992 , n25831 , n25833 );
xor ( n25993 , n25992 , n25836 );
and ( n25994 , n25990 , n25993 );
and ( n25995 , n25988 , n25993 );
or ( n25996 , n25991 , n25994 , n25995 );
and ( n25997 , n25841 , n25996 );
and ( n25998 , n25839 , n25996 );
or ( n25999 , n25842 , n25997 , n25998 );
and ( n26000 , n25798 , n25999 );
and ( n26001 , n25796 , n25999 );
or ( n26002 , n25799 , n26000 , n26001 );
and ( n26003 , n25606 , n26002 );
and ( n26004 , n25604 , n26002 );
or ( n26005 , n25607 , n26003 , n26004 );
and ( n26006 , n25438 , n26005 );
xor ( n26007 , n25438 , n26005 );
xor ( n26008 , n25604 , n25606 );
xor ( n26009 , n26008 , n26002 );
not ( n26010 , n26009 );
xor ( n26011 , n25796 , n25798 );
xor ( n26012 , n26011 , n25999 );
xor ( n26013 , n25609 , n25611 );
xor ( n26014 , n26013 , n25793 );
xor ( n26015 , n25839 , n25841 );
xor ( n26016 , n26015 , n25996 );
and ( n26017 , n26014 , n26016 );
xor ( n26018 , n25823 , n25825 );
xor ( n26019 , n26018 , n25828 );
and ( n26020 , n24624 , n21296 );
and ( n26021 , n23483 , n22337 );
and ( n26022 , n26020 , n26021 );
and ( n26023 , n23215 , n22784 );
and ( n26024 , n26021 , n26023 );
and ( n26025 , n26020 , n26023 );
or ( n26026 , n26022 , n26024 , n26025 );
xor ( n26027 , n25706 , n25707 );
xor ( n26028 , n26027 , n25709 );
and ( n26029 , n26026 , n26028 );
xor ( n26030 , n25650 , n25651 );
xor ( n26031 , n26030 , n25654 );
and ( n26032 , n26028 , n26031 );
and ( n26033 , n26026 , n26031 );
or ( n26034 , n26029 , n26032 , n26033 );
and ( n26035 , n25220 , n21039 );
and ( n26036 , n24546 , n21429 );
and ( n26037 , n26035 , n26036 );
xor ( n26038 , n25892 , n25893 );
xor ( n26039 , n26038 , n25895 );
and ( n26040 , n26036 , n26039 );
and ( n26041 , n26035 , n26039 );
or ( n26042 , n26037 , n26040 , n26041 );
xor ( n26043 , n25765 , n25766 );
xor ( n26044 , n26043 , n25769 );
and ( n26045 , n26042 , n26044 );
and ( n26046 , n26034 , n26045 );
xnor ( n26047 , n25887 , n25889 );
xor ( n26048 , n25898 , n25905 );
and ( n26049 , n26047 , n26048 );
and ( n26050 , n25742 , n20909 );
and ( n26051 , n24731 , n21296 );
and ( n26052 , n26050 , n26051 );
and ( n26053 , n23336 , n22784 );
and ( n26054 , n26051 , n26053 );
and ( n26055 , n26050 , n26053 );
or ( n26056 , n26052 , n26054 , n26055 );
and ( n26057 , n25623 , n20949 );
and ( n26058 , n24052 , n21827 );
and ( n26059 , n26057 , n26058 );
and ( n26060 , n23483 , n22562 );
and ( n26061 , n26058 , n26060 );
and ( n26062 , n26057 , n26060 );
or ( n26063 , n26059 , n26061 , n26062 );
and ( n26064 , n26056 , n26063 );
and ( n26065 , n25959 , n20890 );
and ( n26066 , n23742 , n22172 );
and ( n26067 , n26065 , n26066 );
and ( n26068 , n23620 , n22337 );
and ( n26069 , n26066 , n26068 );
and ( n26070 , n26065 , n26068 );
or ( n26071 , n26067 , n26069 , n26070 );
and ( n26072 , n26063 , n26071 );
and ( n26073 , n26056 , n26071 );
or ( n26074 , n26064 , n26072 , n26073 );
and ( n26075 , n26048 , n26074 );
and ( n26076 , n26047 , n26074 );
or ( n26077 , n26049 , n26075 , n26076 );
and ( n26078 , n26045 , n26077 );
and ( n26079 , n26034 , n26077 );
or ( n26080 , n26046 , n26078 , n26079 );
and ( n26081 , n25220 , n21085 );
and ( n26082 , n24993 , n21178 );
and ( n26083 , n26081 , n26082 );
and ( n26084 , n24546 , n21527 );
and ( n26085 , n26082 , n26084 );
and ( n26086 , n26081 , n26084 );
or ( n26087 , n26083 , n26085 , n26086 );
xor ( n26088 , n25881 , n25882 );
xor ( n26089 , n26088 , n25884 );
and ( n26090 , n26087 , n26089 );
and ( n26091 , n23215 , n22987 );
and ( n26092 , n23089 , n23322 );
and ( n26093 , n26091 , n26092 );
and ( n26094 , n22824 , n23758 );
and ( n26095 , n26092 , n26094 );
and ( n26096 , n26091 , n26094 );
or ( n26097 , n26093 , n26095 , n26096 );
xor ( n26098 , n25899 , n25900 );
xor ( n26099 , n26098 , n25902 );
and ( n26100 , n26097 , n26099 );
and ( n26101 , n26090 , n26100 );
and ( n26102 , n23089 , n22987 );
and ( n26103 , n22936 , n23322 );
and ( n26104 , n26102 , n26103 );
xor ( n26105 , n25868 , n25869 );
xor ( n26106 , n26105 , n25871 );
and ( n26107 , n26103 , n26106 );
and ( n26108 , n26102 , n26106 );
or ( n26109 , n26104 , n26107 , n26108 );
and ( n26110 , n26100 , n26109 );
and ( n26111 , n26090 , n26109 );
or ( n26112 , n26101 , n26110 , n26111 );
xor ( n26113 , n25848 , n25850 );
xor ( n26114 , n26113 , n25853 );
and ( n26115 , n26112 , n26114 );
xor ( n26116 , n25880 , n25890 );
xor ( n26117 , n26116 , n25906 );
and ( n26118 , n26114 , n26117 );
and ( n26119 , n26112 , n26117 );
or ( n26120 , n26115 , n26118 , n26119 );
and ( n26121 , n26080 , n26120 );
xor ( n26122 , n25844 , n25845 );
xor ( n26123 , n26122 , n25856 );
and ( n26124 , n26120 , n26123 );
and ( n26125 , n26080 , n26123 );
or ( n26126 , n26121 , n26124 , n26125 );
xor ( n26127 , n25816 , n25818 );
xor ( n26128 , n26127 , n25820 );
and ( n26129 , n26126 , n26128 );
xor ( n26130 , n25743 , n25744 );
xor ( n26131 , n26130 , n25746 );
xor ( n26132 , n25874 , n25875 );
xor ( n26133 , n26132 , n25877 );
and ( n26134 , n26131 , n26133 );
xor ( n26135 , n26026 , n26028 );
xor ( n26136 , n26135 , n26031 );
and ( n26137 , n26133 , n26136 );
and ( n26138 , n26131 , n26136 );
or ( n26139 , n26134 , n26137 , n26138 );
and ( n26140 , n23089 , n23508 );
and ( n26141 , n22824 , n24064 );
and ( n26142 , n26140 , n26141 );
and ( n26143 , n22702 , n24540 );
and ( n26144 , n26141 , n26143 );
and ( n26145 , n26140 , n26143 );
or ( n26146 , n26142 , n26144 , n26145 );
buf ( n26147 , n16538 );
buf ( n26148 , n26147 );
and ( n26149 , n26148 , n20877 );
and ( n26150 , n26146 , n26149 );
and ( n26151 , n24337 , n21666 );
and ( n26152 , n26149 , n26151 );
and ( n26153 , n26146 , n26151 );
or ( n26154 , n26150 , n26152 , n26153 );
xor ( n26155 , n26020 , n26021 );
xor ( n26156 , n26155 , n26023 );
and ( n26157 , n26154 , n26156 );
xor ( n26158 , n25957 , n25960 );
xor ( n26159 , n26158 , n25962 );
and ( n26160 , n26156 , n26159 );
and ( n26161 , n26154 , n26159 );
or ( n26162 , n26157 , n26160 , n26161 );
xor ( n26163 , n25965 , n25967 );
xor ( n26164 , n26163 , n25970 );
and ( n26165 , n26162 , n26164 );
and ( n26166 , n26139 , n26165 );
xor ( n26167 , n25923 , n25924 );
xor ( n26168 , n26167 , n25926 );
xnor ( n26169 , n25931 , n25932 );
and ( n26170 , n26168 , n26169 );
and ( n26171 , n25451 , n21039 );
and ( n26172 , n24624 , n21429 );
and ( n26173 , n26171 , n26172 );
and ( n26174 , n23903 , n21990 );
and ( n26175 , n26172 , n26174 );
and ( n26176 , n26171 , n26174 );
or ( n26177 , n26173 , n26175 , n26176 );
and ( n26178 , n26169 , n26177 );
and ( n26179 , n26168 , n26177 );
or ( n26180 , n26170 , n26178 , n26179 );
xor ( n26181 , n25922 , n25929 );
xor ( n26182 , n26181 , n25933 );
and ( n26183 , n26180 , n26182 );
xor ( n26184 , n26042 , n26044 );
and ( n26185 , n26182 , n26184 );
and ( n26186 , n26180 , n26184 );
or ( n26187 , n26183 , n26185 , n26186 );
and ( n26188 , n26165 , n26187 );
and ( n26189 , n26139 , n26187 );
or ( n26190 , n26166 , n26188 , n26189 );
and ( n26191 , n22702 , n24064 );
and ( n26192 , n22542 , n25026 );
and ( n26193 , n26191 , n26192 );
and ( n26194 , n22354 , n25617 );
and ( n26195 , n26192 , n26194 );
and ( n26196 , n26191 , n26194 );
or ( n26197 , n26193 , n26195 , n26196 );
xor ( n26198 , n26056 , n26063 );
xor ( n26199 , n26198 , n26071 );
and ( n26200 , n26197 , n26199 );
xor ( n26201 , n26035 , n26036 );
xor ( n26202 , n26201 , n26039 );
and ( n26203 , n26199 , n26202 );
and ( n26204 , n26197 , n26202 );
or ( n26205 , n26200 , n26203 , n26204 );
xor ( n26206 , n26087 , n26089 );
xor ( n26207 , n26097 , n26099 );
and ( n26208 , n26206 , n26207 );
and ( n26209 , n25451 , n21085 );
and ( n26210 , n25220 , n21178 );
and ( n26211 , n26209 , n26210 );
and ( n26212 , n24624 , n21527 );
and ( n26213 , n26210 , n26212 );
and ( n26214 , n26209 , n26212 );
or ( n26215 , n26211 , n26213 , n26214 );
xor ( n26216 , n26057 , n26058 );
xor ( n26217 , n26216 , n26060 );
and ( n26218 , n26215 , n26217 );
xor ( n26219 , n26091 , n26092 );
xor ( n26220 , n26219 , n26094 );
and ( n26221 , n26217 , n26220 );
and ( n26222 , n26215 , n26220 );
or ( n26223 , n26218 , n26221 , n26222 );
and ( n26224 , n26207 , n26223 );
and ( n26225 , n26206 , n26223 );
or ( n26226 , n26208 , n26224 , n26225 );
and ( n26227 , n26205 , n26226 );
buf ( n26228 , n20270 );
buf ( n26229 , n26228 );
and ( n26230 , n22232 , n26229 );
buf ( n26231 , n22116 );
and ( n26232 , n26230 , n26231 );
xor ( n26233 , n25951 , n25952 );
xor ( n26234 , n26233 , n25954 );
and ( n26235 , n26231 , n26234 );
and ( n26236 , n26230 , n26234 );
or ( n26237 , n26232 , n26235 , n26236 );
xor ( n26238 , n26081 , n26082 );
xor ( n26239 , n26238 , n26084 );
xor ( n26240 , n26050 , n26051 );
xor ( n26241 , n26240 , n26053 );
and ( n26242 , n26239 , n26241 );
and ( n26243 , n25742 , n20949 );
and ( n26244 , n23620 , n22562 );
and ( n26245 , n26243 , n26244 );
and ( n26246 , n23336 , n22987 );
and ( n26247 , n26244 , n26246 );
and ( n26248 , n26243 , n26246 );
or ( n26249 , n26245 , n26247 , n26248 );
and ( n26250 , n26241 , n26249 );
and ( n26251 , n26239 , n26249 );
or ( n26252 , n26242 , n26250 , n26251 );
and ( n26253 , n26237 , n26252 );
and ( n26254 , n22589 , n25026 );
and ( n26255 , n22351 , n25617 );
and ( n26256 , n26254 , n26255 );
and ( n26257 , n22354 , n26229 );
and ( n26258 , n26255 , n26257 );
and ( n26259 , n26254 , n26257 );
or ( n26260 , n26256 , n26258 , n26259 );
and ( n26261 , n25623 , n21039 );
and ( n26262 , n24546 , n21666 );
and ( n26263 , n26261 , n26262 );
and ( n26264 , n23215 , n23322 );
and ( n26265 , n26262 , n26264 );
and ( n26266 , n26261 , n26264 );
or ( n26267 , n26263 , n26265 , n26266 );
and ( n26268 , n26260 , n26267 );
xor ( n26269 , n26171 , n26172 );
xor ( n26270 , n26269 , n26174 );
and ( n26271 , n26267 , n26270 );
and ( n26272 , n26260 , n26270 );
or ( n26273 , n26268 , n26271 , n26272 );
and ( n26274 , n26252 , n26273 );
and ( n26275 , n26237 , n26273 );
or ( n26276 , n26253 , n26274 , n26275 );
and ( n26277 , n26226 , n26276 );
and ( n26278 , n26205 , n26276 );
or ( n26279 , n26227 , n26277 , n26278 );
xor ( n26280 , n25936 , n25938 );
xor ( n26281 , n26280 , n25941 );
and ( n26282 , n26279 , n26281 );
xor ( n26283 , n25947 , n25949 );
xor ( n26284 , n26283 , n25973 );
and ( n26285 , n26281 , n26284 );
and ( n26286 , n26279 , n26284 );
or ( n26287 , n26282 , n26285 , n26286 );
and ( n26288 , n26190 , n26287 );
xor ( n26289 , n25909 , n25911 );
xor ( n26290 , n26289 , n25914 );
and ( n26291 , n26287 , n26290 );
and ( n26292 , n26190 , n26290 );
or ( n26293 , n26288 , n26291 , n26292 );
and ( n26294 , n26128 , n26293 );
and ( n26295 , n26126 , n26293 );
or ( n26296 , n26129 , n26294 , n26295 );
and ( n26297 , n26019 , n26296 );
xor ( n26298 , n25866 , n25982 );
xor ( n26299 , n26298 , n25985 );
and ( n26300 , n26296 , n26299 );
and ( n26301 , n26019 , n26299 );
or ( n26302 , n26297 , n26300 , n26301 );
xor ( n26303 , n25988 , n25990 );
xor ( n26304 , n26303 , n25993 );
and ( n26305 , n26302 , n26304 );
xor ( n26306 , n25859 , n25861 );
xor ( n26307 , n26306 , n25863 );
xor ( n26308 , n25867 , n25917 );
xor ( n26309 , n26308 , n25979 );
and ( n26310 , n26307 , n26309 );
xor ( n26311 , n25920 , n25944 );
xor ( n26312 , n26311 , n25976 );
xor ( n26313 , n26080 , n26120 );
xor ( n26314 , n26313 , n26123 );
and ( n26315 , n26312 , n26314 );
xor ( n26316 , n26034 , n26045 );
xor ( n26317 , n26316 , n26077 );
xor ( n26318 , n26112 , n26114 );
xor ( n26319 , n26318 , n26117 );
and ( n26320 , n26317 , n26319 );
xor ( n26321 , n26047 , n26048 );
xor ( n26322 , n26321 , n26074 );
xor ( n26323 , n26090 , n26100 );
xor ( n26324 , n26323 , n26109 );
and ( n26325 , n26322 , n26324 );
xor ( n26326 , n26131 , n26133 );
xor ( n26327 , n26326 , n26136 );
and ( n26328 , n26324 , n26327 );
and ( n26329 , n26322 , n26327 );
or ( n26330 , n26325 , n26328 , n26329 );
and ( n26331 , n26319 , n26330 );
and ( n26332 , n26317 , n26330 );
or ( n26333 , n26320 , n26331 , n26332 );
and ( n26334 , n26314 , n26333 );
and ( n26335 , n26312 , n26333 );
or ( n26336 , n26315 , n26334 , n26335 );
and ( n26337 , n26309 , n26336 );
and ( n26338 , n26307 , n26336 );
or ( n26339 , n26310 , n26337 , n26338 );
xor ( n26340 , n26019 , n26296 );
xor ( n26341 , n26340 , n26299 );
and ( n26342 , n26339 , n26341 );
xor ( n26343 , n26126 , n26128 );
xor ( n26344 , n26343 , n26293 );
xor ( n26345 , n26162 , n26164 );
xor ( n26346 , n26102 , n26103 );
xor ( n26347 , n26346 , n26106 );
xor ( n26348 , n26168 , n26169 );
xor ( n26349 , n26348 , n26177 );
and ( n26350 , n26347 , n26349 );
xor ( n26351 , n26154 , n26156 );
xor ( n26352 , n26351 , n26159 );
and ( n26353 , n26349 , n26352 );
and ( n26354 , n26347 , n26352 );
or ( n26355 , n26350 , n26353 , n26354 );
and ( n26356 , n26345 , n26355 );
and ( n26357 , n25959 , n20909 );
and ( n26358 , n24993 , n21296 );
and ( n26359 , n26357 , n26358 );
and ( n26360 , n23483 , n22784 );
and ( n26361 , n26358 , n26360 );
and ( n26362 , n26357 , n26360 );
or ( n26363 , n26359 , n26361 , n26362 );
and ( n26364 , n24337 , n21827 );
and ( n26365 , n23903 , n22172 );
and ( n26366 , n26364 , n26365 );
and ( n26367 , n22936 , n23758 );
and ( n26368 , n26365 , n26367 );
and ( n26369 , n26364 , n26367 );
or ( n26370 , n26366 , n26368 , n26369 );
and ( n26371 , n26363 , n26370 );
and ( n26372 , n22702 , n25026 );
and ( n26373 , n22542 , n25617 );
and ( n26374 , n26372 , n26373 );
buf ( n26375 , n20273 );
buf ( n26376 , n26375 );
and ( n26377 , n22354 , n26376 );
and ( n26378 , n26373 , n26377 );
and ( n26379 , n26372 , n26377 );
or ( n26380 , n26374 , n26378 , n26379 );
and ( n26381 , n26148 , n20890 );
and ( n26382 , n26380 , n26381 );
and ( n26383 , n23742 , n22337 );
and ( n26384 , n26381 , n26383 );
and ( n26385 , n26380 , n26383 );
or ( n26386 , n26382 , n26384 , n26385 );
and ( n26387 , n26370 , n26386 );
and ( n26388 , n26363 , n26386 );
or ( n26389 , n26371 , n26387 , n26388 );
and ( n26390 , n22936 , n24064 );
and ( n26391 , n22351 , n26229 );
and ( n26392 , n26390 , n26391 );
buf ( n26393 , n22232 );
not ( n26394 , n26393 );
and ( n26395 , n26391 , n26394 );
and ( n26396 , n26390 , n26394 );
or ( n26397 , n26392 , n26395 , n26396 );
buf ( n26398 , n16732 );
buf ( n26399 , n26398 );
and ( n26400 , n26399 , n20877 );
and ( n26401 , n26397 , n26400 );
and ( n26402 , n24052 , n21990 );
and ( n26403 , n26400 , n26402 );
and ( n26404 , n26397 , n26402 );
or ( n26405 , n26401 , n26403 , n26404 );
xor ( n26406 , n26065 , n26066 );
xor ( n26407 , n26406 , n26068 );
and ( n26408 , n26405 , n26407 );
and ( n26409 , n26389 , n26408 );
xor ( n26410 , n26191 , n26192 );
xor ( n26411 , n26410 , n26194 );
xor ( n26412 , n26146 , n26149 );
xor ( n26413 , n26412 , n26151 );
and ( n26414 , n26411 , n26413 );
and ( n26415 , n22542 , n25284 );
xor ( n26416 , n26140 , n26141 );
xor ( n26417 , n26416 , n26143 );
and ( n26418 , n26415 , n26417 );
xor ( n26419 , n26209 , n26210 );
xor ( n26420 , n26419 , n26212 );
and ( n26421 , n26417 , n26420 );
and ( n26422 , n26415 , n26420 );
or ( n26423 , n26418 , n26421 , n26422 );
and ( n26424 , n26413 , n26423 );
and ( n26425 , n26411 , n26423 );
or ( n26426 , n26414 , n26424 , n26425 );
and ( n26427 , n26408 , n26426 );
and ( n26428 , n26389 , n26426 );
or ( n26429 , n26409 , n26427 , n26428 );
and ( n26430 , n26355 , n26429 );
and ( n26431 , n26345 , n26429 );
or ( n26432 , n26356 , n26430 , n26431 );
xor ( n26433 , n26254 , n26255 );
xor ( n26434 , n26433 , n26257 );
and ( n26435 , n23215 , n23508 );
and ( n26436 , n22824 , n24540 );
and ( n26437 , n26435 , n26436 );
and ( n26438 , n22589 , n25284 );
and ( n26439 , n26436 , n26438 );
and ( n26440 , n26435 , n26438 );
or ( n26441 , n26437 , n26439 , n26440 );
and ( n26442 , n26434 , n26441 );
buf ( n26443 , n26393 );
and ( n26444 , n26441 , n26443 );
and ( n26445 , n26434 , n26443 );
or ( n26446 , n26442 , n26444 , n26445 );
xor ( n26447 , n26230 , n26231 );
xor ( n26448 , n26447 , n26234 );
and ( n26449 , n26446 , n26448 );
xor ( n26450 , n26239 , n26241 );
xor ( n26451 , n26450 , n26249 );
and ( n26452 , n26448 , n26451 );
and ( n26453 , n26446 , n26451 );
or ( n26454 , n26449 , n26452 , n26453 );
xor ( n26455 , n26197 , n26199 );
xor ( n26456 , n26455 , n26202 );
and ( n26457 , n26454 , n26456 );
xor ( n26458 , n26206 , n26207 );
xor ( n26459 , n26458 , n26223 );
and ( n26460 , n26456 , n26459 );
and ( n26461 , n26454 , n26459 );
or ( n26462 , n26457 , n26460 , n26461 );
xor ( n26463 , n26180 , n26182 );
xor ( n26464 , n26463 , n26184 );
and ( n26465 , n26462 , n26464 );
xor ( n26466 , n26205 , n26226 );
xor ( n26467 , n26466 , n26276 );
and ( n26468 , n26464 , n26467 );
and ( n26469 , n26462 , n26467 );
or ( n26470 , n26465 , n26468 , n26469 );
and ( n26471 , n26432 , n26470 );
xor ( n26472 , n26139 , n26165 );
xor ( n26473 , n26472 , n26187 );
and ( n26474 , n26470 , n26473 );
and ( n26475 , n26432 , n26473 );
or ( n26476 , n26471 , n26474 , n26475 );
xor ( n26477 , n26190 , n26287 );
xor ( n26478 , n26477 , n26290 );
and ( n26479 , n26476 , n26478 );
xor ( n26480 , n26279 , n26281 );
xor ( n26481 , n26480 , n26284 );
xor ( n26482 , n26237 , n26252 );
xor ( n26483 , n26482 , n26273 );
and ( n26484 , n25623 , n21085 );
and ( n26485 , n25451 , n21178 );
and ( n26486 , n26484 , n26485 );
xor ( n26487 , n26372 , n26373 );
xor ( n26488 , n26487 , n26377 );
and ( n26489 , n26485 , n26488 );
and ( n26490 , n26484 , n26488 );
or ( n26491 , n26486 , n26489 , n26490 );
xor ( n26492 , n26357 , n26358 );
xor ( n26493 , n26492 , n26360 );
and ( n26494 , n26491 , n26493 );
xor ( n26495 , n26380 , n26381 );
xor ( n26496 , n26495 , n26383 );
and ( n26497 , n26493 , n26496 );
and ( n26498 , n26491 , n26496 );
or ( n26499 , n26494 , n26497 , n26498 );
xor ( n26500 , n26363 , n26370 );
xor ( n26501 , n26500 , n26386 );
and ( n26502 , n26499 , n26501 );
xor ( n26503 , n26215 , n26217 );
xor ( n26504 , n26503 , n26220 );
and ( n26505 , n26501 , n26504 );
and ( n26506 , n26499 , n26504 );
or ( n26507 , n26502 , n26505 , n26506 );
and ( n26508 , n26483 , n26507 );
xor ( n26509 , n26260 , n26267 );
xor ( n26510 , n26509 , n26270 );
xor ( n26511 , n26405 , n26407 );
and ( n26512 , n26510 , n26511 );
and ( n26513 , n26148 , n20909 );
and ( n26514 , n25220 , n21296 );
and ( n26515 , n26513 , n26514 );
and ( n26516 , n23620 , n22784 );
and ( n26517 , n26514 , n26516 );
and ( n26518 , n26513 , n26516 );
or ( n26519 , n26515 , n26517 , n26518 );
and ( n26520 , n22589 , n25617 );
and ( n26521 , n22542 , n26229 );
and ( n26522 , n26520 , n26521 );
and ( n26523 , n22351 , n26376 );
and ( n26524 , n26521 , n26523 );
and ( n26525 , n26520 , n26523 );
or ( n26526 , n26522 , n26524 , n26525 );
and ( n26527 , n24546 , n21827 );
and ( n26528 , n26526 , n26527 );
and ( n26529 , n24052 , n22172 );
and ( n26530 , n26527 , n26529 );
and ( n26531 , n26526 , n26529 );
or ( n26532 , n26528 , n26530 , n26531 );
and ( n26533 , n26519 , n26532 );
xor ( n26534 , n26243 , n26244 );
xor ( n26535 , n26534 , n26246 );
and ( n26536 , n26532 , n26535 );
and ( n26537 , n26519 , n26535 );
or ( n26538 , n26533 , n26536 , n26537 );
and ( n26539 , n26511 , n26538 );
and ( n26540 , n26510 , n26538 );
or ( n26541 , n26512 , n26539 , n26540 );
and ( n26542 , n26507 , n26541 );
and ( n26543 , n26483 , n26541 );
or ( n26544 , n26508 , n26542 , n26543 );
and ( n26545 , n23620 , n22987 );
and ( n26546 , n23483 , n23322 );
and ( n26547 , n26545 , n26546 );
and ( n26548 , n23215 , n23758 );
and ( n26549 , n26546 , n26548 );
and ( n26550 , n26545 , n26548 );
or ( n26551 , n26547 , n26549 , n26550 );
and ( n26552 , n25742 , n21039 );
and ( n26553 , n26551 , n26552 );
and ( n26554 , n24993 , n21429 );
and ( n26555 , n26552 , n26554 );
and ( n26556 , n26551 , n26554 );
or ( n26557 , n26553 , n26555 , n26556 );
and ( n26558 , n26399 , n20890 );
and ( n26559 , n23903 , n22337 );
and ( n26560 , n26558 , n26559 );
xor ( n26561 , n26390 , n26391 );
xor ( n26562 , n26561 , n26394 );
and ( n26563 , n26559 , n26562 );
and ( n26564 , n26558 , n26562 );
or ( n26565 , n26560 , n26563 , n26564 );
and ( n26566 , n26557 , n26565 );
xor ( n26567 , n26397 , n26400 );
xor ( n26568 , n26567 , n26402 );
and ( n26569 , n26565 , n26568 );
and ( n26570 , n26557 , n26568 );
or ( n26571 , n26566 , n26569 , n26570 );
xor ( n26572 , n26261 , n26262 );
xor ( n26573 , n26572 , n26264 );
xor ( n26574 , n26415 , n26417 );
xor ( n26575 , n26574 , n26420 );
and ( n26576 , n26573 , n26575 );
xor ( n26577 , n26434 , n26441 );
xor ( n26578 , n26577 , n26443 );
and ( n26579 , n26575 , n26578 );
and ( n26580 , n26573 , n26578 );
or ( n26581 , n26576 , n26579 , n26580 );
and ( n26582 , n26571 , n26581 );
xor ( n26583 , n26411 , n26413 );
xor ( n26584 , n26583 , n26423 );
and ( n26585 , n26581 , n26584 );
and ( n26586 , n26571 , n26584 );
or ( n26587 , n26582 , n26585 , n26586 );
xor ( n26588 , n26347 , n26349 );
xor ( n26589 , n26588 , n26352 );
and ( n26590 , n26587 , n26589 );
xor ( n26591 , n26389 , n26408 );
xor ( n26592 , n26591 , n26426 );
and ( n26593 , n26589 , n26592 );
and ( n26594 , n26587 , n26592 );
or ( n26595 , n26590 , n26593 , n26594 );
and ( n26596 , n26544 , n26595 );
xor ( n26597 , n26322 , n26324 );
xor ( n26598 , n26597 , n26327 );
and ( n26599 , n26595 , n26598 );
and ( n26600 , n26544 , n26598 );
or ( n26601 , n26596 , n26599 , n26600 );
and ( n26602 , n26481 , n26601 );
xor ( n26603 , n26317 , n26319 );
xor ( n26604 , n26603 , n26330 );
and ( n26605 , n26601 , n26604 );
and ( n26606 , n26481 , n26604 );
or ( n26607 , n26602 , n26605 , n26606 );
and ( n26608 , n26478 , n26607 );
and ( n26609 , n26476 , n26607 );
or ( n26610 , n26479 , n26608 , n26609 );
and ( n26611 , n26344 , n26610 );
xor ( n26612 , n26307 , n26309 );
xor ( n26613 , n26612 , n26336 );
and ( n26614 , n26610 , n26613 );
and ( n26615 , n26344 , n26613 );
or ( n26616 , n26611 , n26614 , n26615 );
and ( n26617 , n26341 , n26616 );
and ( n26618 , n26339 , n26616 );
or ( n26619 , n26342 , n26617 , n26618 );
and ( n26620 , n26304 , n26619 );
and ( n26621 , n26302 , n26619 );
or ( n26622 , n26305 , n26620 , n26621 );
and ( n26623 , n26016 , n26622 );
and ( n26624 , n26014 , n26622 );
or ( n26625 , n26017 , n26623 , n26624 );
and ( n26626 , n26012 , n26625 );
xor ( n26627 , n26012 , n26625 );
xor ( n26628 , n26014 , n26016 );
xor ( n26629 , n26628 , n26622 );
not ( n26630 , n26629 );
xor ( n26631 , n26302 , n26304 );
xor ( n26632 , n26631 , n26619 );
xor ( n26633 , n26339 , n26341 );
xor ( n26634 , n26633 , n26616 );
not ( n26635 , n26634 );
xor ( n26636 , n26312 , n26314 );
xor ( n26637 , n26636 , n26333 );
xor ( n26638 , n26432 , n26470 );
xor ( n26639 , n26638 , n26473 );
xor ( n26640 , n26345 , n26355 );
xor ( n26641 , n26640 , n26429 );
xor ( n26642 , n26462 , n26464 );
xor ( n26643 , n26642 , n26467 );
and ( n26644 , n26641 , n26643 );
xor ( n26645 , n26454 , n26456 );
xor ( n26646 , n26645 , n26459 );
xor ( n26647 , n26446 , n26448 );
xor ( n26648 , n26647 , n26451 );
and ( n26649 , n25959 , n20949 );
and ( n26650 , n23742 , n22562 );
and ( n26651 , n26649 , n26650 );
and ( n26652 , n23483 , n22987 );
and ( n26653 , n26650 , n26652 );
and ( n26654 , n26649 , n26652 );
or ( n26655 , n26651 , n26653 , n26654 );
and ( n26656 , n22824 , n25026 );
buf ( n26657 , n26656 );
and ( n26658 , n23336 , n23322 );
and ( n26659 , n26657 , n26658 );
and ( n26660 , n23089 , n23758 );
and ( n26661 , n26658 , n26660 );
and ( n26662 , n26657 , n26660 );
or ( n26663 , n26659 , n26661 , n26662 );
and ( n26664 , n26655 , n26663 );
and ( n26665 , n24731 , n21429 );
and ( n26666 , n26663 , n26665 );
and ( n26667 , n26655 , n26665 );
or ( n26668 , n26664 , n26666 , n26667 );
and ( n26669 , n26648 , n26668 );
and ( n26670 , n23336 , n23508 );
and ( n26671 , n22936 , n24540 );
and ( n26672 , n26670 , n26671 );
and ( n26673 , n22702 , n25284 );
and ( n26674 , n26671 , n26673 );
and ( n26675 , n26670 , n26673 );
or ( n26676 , n26672 , n26674 , n26675 );
buf ( n26677 , n16750 );
buf ( n26678 , n26677 );
and ( n26679 , n26678 , n20877 );
and ( n26680 , n26676 , n26679 );
and ( n26681 , n24337 , n21990 );
and ( n26682 , n26679 , n26681 );
and ( n26683 , n26676 , n26681 );
or ( n26684 , n26680 , n26682 , n26683 );
buf ( n26685 , n22354 );
buf ( n26686 , n26685 );
and ( n26687 , n23089 , n24064 );
and ( n26688 , n26686 , n26687 );
not ( n26689 , n26656 );
and ( n26690 , n26687 , n26689 );
and ( n26691 , n26686 , n26689 );
or ( n26692 , n26688 , n26690 , n26691 );
and ( n26693 , n24731 , n21527 );
and ( n26694 , n26692 , n26693 );
and ( n26695 , n24624 , n21666 );
and ( n26696 , n26693 , n26695 );
and ( n26697 , n26692 , n26695 );
or ( n26698 , n26694 , n26696 , n26697 );
and ( n26699 , n26684 , n26698 );
xor ( n26700 , n26364 , n26365 );
xor ( n26701 , n26700 , n26367 );
and ( n26702 , n26698 , n26701 );
and ( n26703 , n26684 , n26701 );
or ( n26704 , n26699 , n26702 , n26703 );
and ( n26705 , n26668 , n26704 );
and ( n26706 , n26648 , n26704 );
or ( n26707 , n26669 , n26705 , n26706 );
and ( n26708 , n26646 , n26707 );
xor ( n26709 , n26519 , n26532 );
xor ( n26710 , n26709 , n26535 );
xor ( n26711 , n26557 , n26565 );
xor ( n26712 , n26711 , n26568 );
and ( n26713 , n26710 , n26712 );
xor ( n26714 , n26513 , n26514 );
xor ( n26715 , n26714 , n26516 );
xor ( n26716 , n26526 , n26527 );
xor ( n26717 , n26716 , n26529 );
and ( n26718 , n26715 , n26717 );
xor ( n26719 , n26558 , n26559 );
xor ( n26720 , n26719 , n26562 );
and ( n26721 , n26717 , n26720 );
and ( n26722 , n26715 , n26720 );
or ( n26723 , n26718 , n26721 , n26722 );
and ( n26724 , n26712 , n26723 );
and ( n26725 , n26710 , n26723 );
or ( n26726 , n26713 , n26724 , n26725 );
xor ( n26727 , n26510 , n26511 );
xor ( n26728 , n26727 , n26538 );
and ( n26729 , n26726 , n26728 );
xor ( n26730 , n26571 , n26581 );
xor ( n26731 , n26730 , n26584 );
and ( n26732 , n26728 , n26731 );
and ( n26733 , n26726 , n26731 );
or ( n26734 , n26729 , n26732 , n26733 );
and ( n26735 , n26707 , n26734 );
and ( n26736 , n26646 , n26734 );
or ( n26737 , n26708 , n26735 , n26736 );
and ( n26738 , n26643 , n26737 );
and ( n26739 , n26641 , n26737 );
or ( n26740 , n26644 , n26738 , n26739 );
and ( n26741 , n26639 , n26740 );
xor ( n26742 , n26481 , n26601 );
xor ( n26743 , n26742 , n26604 );
and ( n26744 , n26740 , n26743 );
and ( n26745 , n26639 , n26743 );
or ( n26746 , n26741 , n26744 , n26745 );
and ( n26747 , n26637 , n26746 );
xor ( n26748 , n26476 , n26478 );
xor ( n26749 , n26748 , n26607 );
and ( n26750 , n26746 , n26749 );
and ( n26751 , n26637 , n26749 );
or ( n26752 , n26747 , n26750 , n26751 );
xor ( n26753 , n26344 , n26610 );
xor ( n26754 , n26753 , n26613 );
and ( n26755 , n26752 , n26754 );
xor ( n26756 , n26752 , n26754 );
xor ( n26757 , n26637 , n26746 );
xor ( n26758 , n26757 , n26749 );
xor ( n26759 , n26544 , n26595 );
xor ( n26760 , n26759 , n26598 );
xor ( n26761 , n26483 , n26507 );
xor ( n26762 , n26761 , n26541 );
xor ( n26763 , n26587 , n26589 );
xor ( n26764 , n26763 , n26592 );
and ( n26765 , n26762 , n26764 );
and ( n26766 , n26399 , n20949 );
and ( n26767 , n23742 , n22987 );
and ( n26768 , n26766 , n26767 );
and ( n26769 , n23620 , n23322 );
and ( n26770 , n26767 , n26769 );
and ( n26771 , n26766 , n26769 );
or ( n26772 , n26768 , n26770 , n26771 );
and ( n26773 , n23336 , n23758 );
and ( n26774 , n22824 , n25284 );
and ( n26775 , n26773 , n26774 );
not ( n26776 , n26685 );
and ( n26777 , n26774 , n26776 );
and ( n26778 , n26773 , n26776 );
or ( n26779 , n26775 , n26777 , n26778 );
and ( n26780 , n26772 , n26779 );
buf ( n26781 , n16870 );
buf ( n26782 , n26781 );
and ( n26783 , n26782 , n20877 );
and ( n26784 , n26779 , n26783 );
and ( n26785 , n26772 , n26783 );
or ( n26786 , n26780 , n26784 , n26785 );
and ( n26787 , n25959 , n21039 );
and ( n26788 , n25220 , n21429 );
and ( n26789 , n26787 , n26788 );
xor ( n26790 , n26686 , n26687 );
xor ( n26791 , n26790 , n26689 );
and ( n26792 , n26788 , n26791 );
and ( n26793 , n26787 , n26791 );
or ( n26794 , n26789 , n26792 , n26793 );
and ( n26795 , n26786 , n26794 );
xor ( n26796 , n26484 , n26485 );
xor ( n26797 , n26796 , n26488 );
and ( n26798 , n26794 , n26797 );
and ( n26799 , n26786 , n26797 );
or ( n26800 , n26795 , n26798 , n26799 );
xor ( n26801 , n26491 , n26493 );
xor ( n26802 , n26801 , n26496 );
and ( n26803 , n26800 , n26802 );
xor ( n26804 , n26684 , n26698 );
xor ( n26805 , n26804 , n26701 );
and ( n26806 , n26802 , n26805 );
and ( n26807 , n26800 , n26805 );
or ( n26808 , n26803 , n26806 , n26807 );
xor ( n26809 , n26499 , n26501 );
xor ( n26810 , n26809 , n26504 );
and ( n26811 , n26808 , n26810 );
and ( n26812 , n26764 , n26811 );
and ( n26813 , n26762 , n26811 );
or ( n26814 , n26765 , n26812 , n26813 );
and ( n26815 , n26760 , n26814 );
xor ( n26816 , n26641 , n26643 );
xor ( n26817 , n26816 , n26737 );
and ( n26818 , n26814 , n26817 );
and ( n26819 , n26760 , n26817 );
or ( n26820 , n26815 , n26818 , n26819 );
xor ( n26821 , n26639 , n26740 );
xor ( n26822 , n26821 , n26743 );
and ( n26823 , n26820 , n26822 );
and ( n26824 , n26148 , n20949 );
and ( n26825 , n24624 , n21827 );
and ( n26826 , n26824 , n26825 );
and ( n26827 , n23903 , n22562 );
and ( n26828 , n26825 , n26827 );
and ( n26829 , n26824 , n26827 );
or ( n26830 , n26826 , n26828 , n26829 );
and ( n26831 , n26399 , n20909 );
and ( n26832 , n25451 , n21296 );
and ( n26833 , n26831 , n26832 );
and ( n26834 , n23742 , n22784 );
and ( n26835 , n26832 , n26834 );
and ( n26836 , n26831 , n26834 );
or ( n26837 , n26833 , n26835 , n26836 );
and ( n26838 , n26830 , n26837 );
xor ( n26839 , n26435 , n26436 );
xor ( n26840 , n26839 , n26438 );
and ( n26841 , n26837 , n26840 );
and ( n26842 , n26830 , n26840 );
or ( n26843 , n26838 , n26841 , n26842 );
and ( n26844 , n26678 , n20890 );
and ( n26845 , n24337 , n22172 );
and ( n26846 , n26844 , n26845 );
and ( n26847 , n24052 , n22337 );
and ( n26848 , n26845 , n26847 );
and ( n26849 , n26844 , n26847 );
or ( n26850 , n26846 , n26848 , n26849 );
xor ( n26851 , n26649 , n26650 );
xor ( n26852 , n26851 , n26652 );
and ( n26853 , n26850 , n26852 );
xor ( n26854 , n26657 , n26658 );
xor ( n26855 , n26854 , n26660 );
and ( n26856 , n26852 , n26855 );
and ( n26857 , n26850 , n26855 );
or ( n26858 , n26853 , n26856 , n26857 );
and ( n26859 , n26843 , n26858 );
xor ( n26860 , n26655 , n26663 );
xor ( n26861 , n26860 , n26665 );
and ( n26862 , n26858 , n26861 );
and ( n26863 , n26843 , n26861 );
or ( n26864 , n26859 , n26862 , n26863 );
and ( n26865 , n25742 , n21085 );
and ( n26866 , n25623 , n21178 );
and ( n26867 , n26865 , n26866 );
and ( n26868 , n24993 , n21527 );
and ( n26869 , n26866 , n26868 );
and ( n26870 , n26865 , n26868 );
or ( n26871 , n26867 , n26869 , n26870 );
and ( n26872 , n22936 , n25026 );
and ( n26873 , n22542 , n26376 );
and ( n26874 , n26872 , n26873 );
buf ( n26875 , n20276 );
buf ( n26876 , n26875 );
and ( n26877 , n22351 , n26876 );
and ( n26878 , n26873 , n26877 );
and ( n26879 , n26872 , n26877 );
or ( n26880 , n26874 , n26878 , n26879 );
and ( n26881 , n24546 , n21990 );
and ( n26882 , n26880 , n26881 );
xor ( n26883 , n26520 , n26521 );
xor ( n26884 , n26883 , n26523 );
and ( n26885 , n26881 , n26884 );
and ( n26886 , n26880 , n26884 );
or ( n26887 , n26882 , n26885 , n26886 );
and ( n26888 , n26871 , n26887 );
xor ( n26889 , n26573 , n26575 );
xor ( n26890 , n26889 , n26578 );
and ( n26891 , n26888 , n26890 );
xor ( n26892 , n26676 , n26679 );
xor ( n26893 , n26892 , n26681 );
xor ( n26894 , n26551 , n26552 );
xor ( n26895 , n26894 , n26554 );
and ( n26896 , n26893 , n26895 );
xor ( n26897 , n26692 , n26693 );
xor ( n26898 , n26897 , n26695 );
and ( n26899 , n26895 , n26898 );
and ( n26900 , n26893 , n26898 );
or ( n26901 , n26896 , n26899 , n26900 );
and ( n26902 , n26890 , n26901 );
and ( n26903 , n26888 , n26901 );
or ( n26904 , n26891 , n26902 , n26903 );
and ( n26905 , n26864 , n26904 );
and ( n26906 , n24731 , n21666 );
and ( n26907 , n23089 , n24540 );
and ( n26908 , n22702 , n25617 );
and ( n26909 , n26907 , n26908 );
and ( n26910 , n22589 , n26229 );
and ( n26911 , n26908 , n26910 );
and ( n26912 , n26907 , n26910 );
or ( n26913 , n26909 , n26911 , n26912 );
and ( n26914 , n26906 , n26913 );
and ( n26915 , n25959 , n21085 );
and ( n26916 , n25742 , n21178 );
and ( n26917 , n26915 , n26916 );
and ( n26918 , n25220 , n21527 );
and ( n26919 , n26916 , n26918 );
and ( n26920 , n26915 , n26918 );
or ( n26921 , n26917 , n26919 , n26920 );
and ( n26922 , n26913 , n26921 );
and ( n26923 , n26906 , n26921 );
or ( n26924 , n26914 , n26922 , n26923 );
xor ( n26925 , n26715 , n26717 );
xor ( n26926 , n26925 , n26720 );
and ( n26927 , n26924 , n26926 );
xor ( n26928 , n26871 , n26887 );
and ( n26929 , n26926 , n26928 );
and ( n26930 , n26924 , n26928 );
or ( n26931 , n26927 , n26929 , n26930 );
buf ( n26932 , n16981 );
buf ( n26933 , n26932 );
and ( n26934 , n26933 , n20877 );
and ( n26935 , n26782 , n20890 );
and ( n26936 , n26934 , n26935 );
and ( n26937 , n23483 , n23508 );
and ( n26938 , n26935 , n26937 );
and ( n26939 , n26934 , n26937 );
or ( n26940 , n26936 , n26938 , n26939 );
xor ( n26941 , n26880 , n26881 );
xor ( n26942 , n26941 , n26884 );
and ( n26943 , n26940 , n26942 );
xor ( n26944 , n26831 , n26832 );
xor ( n26945 , n26944 , n26834 );
xor ( n26946 , n26844 , n26845 );
xor ( n26947 , n26946 , n26847 );
xor ( n26948 , n26945 , n26947 );
xor ( n26949 , n26865 , n26866 );
xor ( n26950 , n26949 , n26868 );
xor ( n26951 , n26948 , n26950 );
and ( n26952 , n26942 , n26951 );
and ( n26953 , n26940 , n26951 );
or ( n26954 , n26943 , n26952 , n26953 );
and ( n26955 , n24993 , n21666 );
and ( n26956 , n24624 , n21990 );
and ( n26957 , n26955 , n26956 );
xor ( n26958 , n26907 , n26908 );
xor ( n26959 , n26958 , n26910 );
and ( n26960 , n26956 , n26959 );
and ( n26961 , n26955 , n26959 );
or ( n26962 , n26957 , n26960 , n26961 );
and ( n26963 , n26148 , n21039 );
and ( n26964 , n25451 , n21429 );
and ( n26965 , n26963 , n26964 );
xor ( n26966 , n26773 , n26774 );
xor ( n26967 , n26966 , n26776 );
and ( n26968 , n26964 , n26967 );
and ( n26969 , n26963 , n26967 );
or ( n26970 , n26965 , n26968 , n26969 );
and ( n26971 , n26962 , n26970 );
and ( n26972 , n26933 , n20890 );
and ( n26973 , n26782 , n20909 );
and ( n26974 , n26972 , n26973 );
and ( n26975 , n24052 , n22784 );
and ( n26976 , n26973 , n26975 );
and ( n26977 , n26972 , n26975 );
or ( n26978 , n26974 , n26976 , n26977 );
buf ( n26979 , n17035 );
buf ( n26980 , n26979 );
and ( n26981 , n26980 , n20877 );
and ( n26982 , n26148 , n21085 );
and ( n26983 , n26981 , n26982 );
and ( n26984 , n25959 , n21178 );
and ( n26985 , n26982 , n26984 );
and ( n26986 , n26981 , n26984 );
or ( n26987 , n26983 , n26985 , n26986 );
and ( n26988 , n26978 , n26987 );
xor ( n26989 , n26766 , n26767 );
xor ( n26990 , n26989 , n26769 );
and ( n26991 , n26987 , n26990 );
and ( n26992 , n26978 , n26990 );
or ( n26993 , n26988 , n26991 , n26992 );
and ( n26994 , n26970 , n26993 );
and ( n26995 , n26962 , n26993 );
or ( n26996 , n26971 , n26994 , n26995 );
and ( n26997 , n26954 , n26996 );
and ( n26998 , n23215 , n24064 );
and ( n26999 , n26678 , n20909 );
and ( n27000 , n25623 , n21296 );
xor ( n27001 , n26999 , n27000 );
and ( n27002 , n23903 , n22784 );
xor ( n27003 , n27001 , n27002 );
and ( n27004 , n26998 , n27003 );
and ( n27005 , n23620 , n23508 );
and ( n27006 , n23215 , n24540 );
and ( n27007 , n27005 , n27006 );
and ( n27008 , n22936 , n25284 );
and ( n27009 , n27006 , n27008 );
and ( n27010 , n27005 , n27008 );
or ( n27011 , n27007 , n27009 , n27010 );
and ( n27012 , n27003 , n27011 );
and ( n27013 , n26998 , n27011 );
or ( n27014 , n27004 , n27012 , n27013 );
and ( n27015 , n26678 , n20949 );
and ( n27016 , n23903 , n22987 );
and ( n27017 , n27015 , n27016 );
and ( n27018 , n23742 , n23322 );
and ( n27019 , n27016 , n27018 );
and ( n27020 , n27015 , n27018 );
or ( n27021 , n27017 , n27019 , n27020 );
and ( n27022 , n24624 , n22172 );
and ( n27023 , n24546 , n22337 );
and ( n27024 , n27022 , n27023 );
and ( n27025 , n24337 , n22562 );
and ( n27026 , n27023 , n27025 );
and ( n27027 , n27022 , n27025 );
or ( n27028 , n27024 , n27026 , n27027 );
and ( n27029 , n27021 , n27028 );
and ( n27030 , n25451 , n21527 );
and ( n27031 , n25220 , n21666 );
and ( n27032 , n27030 , n27031 );
and ( n27033 , n24731 , n21990 );
and ( n27034 , n27031 , n27033 );
and ( n27035 , n27030 , n27033 );
or ( n27036 , n27032 , n27034 , n27035 );
and ( n27037 , n27028 , n27036 );
and ( n27038 , n27021 , n27036 );
or ( n27039 , n27029 , n27037 , n27038 );
and ( n27040 , n27014 , n27039 );
xor ( n27041 , n26906 , n26913 );
xor ( n27042 , n27041 , n26921 );
and ( n27043 , n27039 , n27042 );
and ( n27044 , n27014 , n27042 );
or ( n27045 , n27040 , n27043 , n27044 );
and ( n27046 , n26996 , n27045 );
and ( n27047 , n26954 , n27045 );
or ( n27048 , n26997 , n27046 , n27047 );
and ( n27049 , n26931 , n27048 );
xor ( n27050 , n26710 , n26712 );
xor ( n27051 , n27050 , n26723 );
and ( n27052 , n27048 , n27051 );
and ( n27053 , n26931 , n27051 );
or ( n27054 , n27049 , n27052 , n27053 );
and ( n27055 , n26904 , n27054 );
and ( n27056 , n26864 , n27054 );
or ( n27057 , n26905 , n27055 , n27056 );
xor ( n27058 , n26646 , n26707 );
xor ( n27059 , n27058 , n26734 );
and ( n27060 , n27057 , n27059 );
xor ( n27061 , n26648 , n26668 );
xor ( n27062 , n27061 , n26704 );
xor ( n27063 , n26726 , n26728 );
xor ( n27064 , n27063 , n26731 );
and ( n27065 , n27062 , n27064 );
xor ( n27066 , n26808 , n26810 );
and ( n27067 , n27064 , n27066 );
and ( n27068 , n27062 , n27066 );
or ( n27069 , n27065 , n27067 , n27068 );
and ( n27070 , n27059 , n27069 );
and ( n27071 , n27057 , n27069 );
or ( n27072 , n27060 , n27070 , n27071 );
xor ( n27073 , n26760 , n26814 );
xor ( n27074 , n27073 , n26817 );
and ( n27075 , n27072 , n27074 );
and ( n27076 , n26999 , n27000 );
and ( n27077 , n27000 , n27002 );
and ( n27078 , n26999 , n27002 );
or ( n27079 , n27076 , n27077 , n27078 );
xor ( n27080 , n26824 , n26825 );
xor ( n27081 , n27080 , n26827 );
and ( n27082 , n27079 , n27081 );
xor ( n27083 , n26545 , n26546 );
xor ( n27084 , n27083 , n26548 );
and ( n27085 , n27081 , n27084 );
and ( n27086 , n27079 , n27084 );
or ( n27087 , n27082 , n27085 , n27086 );
and ( n27088 , n23089 , n25026 );
and ( n27089 , n22824 , n25617 );
and ( n27090 , n27088 , n27089 );
and ( n27091 , n22542 , n26876 );
and ( n27092 , n27089 , n27091 );
and ( n27093 , n27088 , n27091 );
or ( n27094 , n27090 , n27092 , n27093 );
and ( n27095 , n24731 , n21827 );
and ( n27096 , n27094 , n27095 );
and ( n27097 , n24546 , n22172 );
and ( n27098 , n27095 , n27097 );
and ( n27099 , n27094 , n27097 );
or ( n27100 , n27096 , n27098 , n27099 );
and ( n27101 , n24337 , n22337 );
and ( n27102 , n24052 , n22562 );
and ( n27103 , n27101 , n27102 );
xor ( n27104 , n26872 , n26873 );
xor ( n27105 , n27104 , n26877 );
and ( n27106 , n27102 , n27105 );
and ( n27107 , n27101 , n27105 );
or ( n27108 , n27103 , n27106 , n27107 );
and ( n27109 , n27100 , n27108 );
xor ( n27110 , n26670 , n26671 );
xor ( n27111 , n27110 , n26673 );
and ( n27112 , n27108 , n27111 );
and ( n27113 , n27100 , n27111 );
or ( n27114 , n27109 , n27112 , n27113 );
and ( n27115 , n27087 , n27114 );
xor ( n27116 , n26830 , n26837 );
xor ( n27117 , n27116 , n26840 );
and ( n27118 , n27114 , n27117 );
and ( n27119 , n27087 , n27117 );
or ( n27120 , n27115 , n27118 , n27119 );
xor ( n27121 , n26843 , n26858 );
xor ( n27122 , n27121 , n26861 );
and ( n27123 , n27120 , n27122 );
xor ( n27124 , n26800 , n26802 );
xor ( n27125 , n27124 , n26805 );
and ( n27126 , n26945 , n26947 );
and ( n27127 , n26947 , n26950 );
and ( n27128 , n26945 , n26950 );
or ( n27129 , n27126 , n27127 , n27128 );
xor ( n27130 , n26850 , n26852 );
xor ( n27131 , n27130 , n26855 );
and ( n27132 , n27129 , n27131 );
and ( n27133 , n27125 , n27132 );
xor ( n27134 , n26893 , n26895 );
xor ( n27135 , n27134 , n26898 );
xor ( n27136 , n26786 , n26794 );
xor ( n27137 , n27136 , n26797 );
and ( n27138 , n27135 , n27137 );
xor ( n27139 , n27087 , n27114 );
xor ( n27140 , n27139 , n27117 );
and ( n27141 , n27137 , n27140 );
and ( n27142 , n27135 , n27140 );
or ( n27143 , n27138 , n27141 , n27142 );
and ( n27144 , n27132 , n27143 );
and ( n27145 , n27125 , n27143 );
or ( n27146 , n27133 , n27144 , n27145 );
and ( n27147 , n27123 , n27146 );
xor ( n27148 , n26772 , n26779 );
xor ( n27149 , n27148 , n26783 );
xor ( n27150 , n27079 , n27081 );
xor ( n27151 , n27150 , n27084 );
and ( n27152 , n27149 , n27151 );
xor ( n27153 , n27100 , n27108 );
xor ( n27154 , n27153 , n27111 );
and ( n27155 , n27151 , n27154 );
and ( n27156 , n27149 , n27154 );
or ( n27157 , n27152 , n27155 , n27156 );
xor ( n27158 , n26787 , n26788 );
xor ( n27159 , n27158 , n26791 );
xor ( n27160 , n26915 , n26916 );
xor ( n27161 , n27160 , n26918 );
xor ( n27162 , n27094 , n27095 );
xor ( n27163 , n27162 , n27097 );
and ( n27164 , n27161 , n27163 );
xor ( n27165 , n27101 , n27102 );
xor ( n27166 , n27165 , n27105 );
and ( n27167 , n27163 , n27166 );
and ( n27168 , n27161 , n27166 );
or ( n27169 , n27164 , n27167 , n27168 );
and ( n27170 , n27159 , n27169 );
and ( n27171 , n23483 , n23758 );
and ( n27172 , n23336 , n24064 );
and ( n27173 , n27171 , n27172 );
and ( n27174 , n22702 , n26229 );
and ( n27175 , n27172 , n27174 );
and ( n27176 , n27171 , n27174 );
or ( n27177 , n27173 , n27175 , n27176 );
xor ( n27178 , n26934 , n26935 );
xor ( n27179 , n27178 , n26937 );
and ( n27180 , n27177 , n27179 );
xor ( n27181 , n26955 , n26956 );
xor ( n27182 , n27181 , n26959 );
and ( n27183 , n27179 , n27182 );
and ( n27184 , n27177 , n27182 );
or ( n27185 , n27180 , n27183 , n27184 );
and ( n27186 , n27169 , n27185 );
and ( n27187 , n27159 , n27185 );
or ( n27188 , n27170 , n27186 , n27187 );
and ( n27189 , n27157 , n27188 );
xor ( n27190 , n26963 , n26964 );
xor ( n27191 , n27190 , n26967 );
xor ( n27192 , n26978 , n26987 );
xor ( n27193 , n27192 , n26990 );
and ( n27194 , n27191 , n27193 );
and ( n27195 , n22936 , n25617 );
and ( n27196 , n22824 , n26229 );
and ( n27197 , n27195 , n27196 );
and ( n27198 , n22589 , n26876 );
and ( n27199 , n27196 , n27198 );
and ( n27200 , n27195 , n27198 );
or ( n27201 , n27197 , n27199 , n27200 );
and ( n27202 , n25742 , n21296 );
and ( n27203 , n27201 , n27202 );
and ( n27204 , n24993 , n21827 );
and ( n27205 , n27202 , n27204 );
and ( n27206 , n27201 , n27204 );
or ( n27207 , n27203 , n27205 , n27206 );
and ( n27208 , n27193 , n27207 );
and ( n27209 , n27191 , n27207 );
or ( n27210 , n27194 , n27208 , n27209 );
and ( n27211 , n24546 , n22562 );
and ( n27212 , n23903 , n23322 );
and ( n27213 , n27211 , n27212 );
and ( n27214 , n23620 , n23758 );
and ( n27215 , n27212 , n27214 );
and ( n27216 , n27211 , n27214 );
or ( n27217 , n27213 , n27215 , n27216 );
xor ( n27218 , n27088 , n27089 );
xor ( n27219 , n27218 , n27091 );
and ( n27220 , n27217 , n27219 );
xor ( n27221 , n27005 , n27006 );
xor ( n27222 , n27221 , n27008 );
and ( n27223 , n27219 , n27222 );
and ( n27224 , n27217 , n27222 );
or ( n27225 , n27220 , n27223 , n27224 );
and ( n27226 , n26399 , n21039 );
and ( n27227 , n25623 , n21429 );
and ( n27228 , n27226 , n27227 );
xor ( n27229 , n27015 , n27016 );
xor ( n27230 , n27229 , n27018 );
and ( n27231 , n27227 , n27230 );
and ( n27232 , n27226 , n27230 );
or ( n27233 , n27228 , n27231 , n27232 );
and ( n27234 , n27225 , n27233 );
and ( n27235 , n22589 , n26376 );
and ( n27236 , n23742 , n23508 );
and ( n27237 , n23483 , n24064 );
and ( n27238 , n27236 , n27237 );
and ( n27239 , n23089 , n25284 );
and ( n27240 , n27237 , n27239 );
and ( n27241 , n27236 , n27239 );
or ( n27242 , n27238 , n27240 , n27241 );
and ( n27243 , n27235 , n27242 );
and ( n27244 , n22702 , n26376 );
buf ( n27245 , n20279 );
buf ( n27246 , n27245 );
and ( n27247 , n22542 , n27246 );
or ( n27248 , n27244 , n27247 );
and ( n27249 , n27242 , n27248 );
and ( n27250 , n27235 , n27248 );
or ( n27251 , n27243 , n27249 , n27250 );
and ( n27252 , n27233 , n27251 );
and ( n27253 , n27225 , n27251 );
or ( n27254 , n27234 , n27252 , n27253 );
and ( n27255 , n27210 , n27254 );
and ( n27256 , n26678 , n21039 );
and ( n27257 , n25959 , n21296 );
and ( n27258 , n27256 , n27257 );
and ( n27259 , n25220 , n21827 );
and ( n27260 , n27257 , n27259 );
and ( n27261 , n27256 , n27259 );
or ( n27262 , n27258 , n27260 , n27261 );
and ( n27263 , n23336 , n24540 );
and ( n27264 , n23215 , n25026 );
and ( n27265 , n27263 , n27264 );
buf ( n27266 , n22351 );
and ( n27267 , n27264 , n27266 );
and ( n27268 , n27263 , n27266 );
or ( n27269 , n27265 , n27267 , n27268 );
and ( n27270 , n27262 , n27269 );
xor ( n27271 , n27030 , n27031 );
xor ( n27272 , n27271 , n27033 );
and ( n27273 , n27269 , n27272 );
and ( n27274 , n27262 , n27272 );
or ( n27275 , n27270 , n27273 , n27274 );
xor ( n27276 , n26998 , n27003 );
xor ( n27277 , n27276 , n27011 );
and ( n27278 , n27275 , n27277 );
xor ( n27279 , n27021 , n27028 );
xor ( n27280 , n27279 , n27036 );
and ( n27281 , n27277 , n27280 );
and ( n27282 , n27275 , n27280 );
or ( n27283 , n27278 , n27281 , n27282 );
and ( n27284 , n27254 , n27283 );
and ( n27285 , n27210 , n27283 );
or ( n27286 , n27255 , n27284 , n27285 );
and ( n27287 , n27188 , n27286 );
and ( n27288 , n27157 , n27286 );
or ( n27289 , n27189 , n27287 , n27288 );
xor ( n27290 , n26940 , n26942 );
xor ( n27291 , n27290 , n26951 );
xor ( n27292 , n26962 , n26970 );
xor ( n27293 , n27292 , n26993 );
and ( n27294 , n27291 , n27293 );
xor ( n27295 , n27014 , n27039 );
xor ( n27296 , n27295 , n27042 );
and ( n27297 , n27293 , n27296 );
and ( n27298 , n27291 , n27296 );
or ( n27299 , n27294 , n27297 , n27298 );
xor ( n27300 , n26924 , n26926 );
xor ( n27301 , n27300 , n26928 );
and ( n27302 , n27299 , n27301 );
xor ( n27303 , n26954 , n26996 );
xor ( n27304 , n27303 , n27045 );
and ( n27305 , n27301 , n27304 );
and ( n27306 , n27299 , n27304 );
or ( n27307 , n27302 , n27305 , n27306 );
and ( n27308 , n27289 , n27307 );
xor ( n27309 , n26888 , n26890 );
xor ( n27310 , n27309 , n26901 );
and ( n27311 , n27307 , n27310 );
and ( n27312 , n27289 , n27310 );
or ( n27313 , n27308 , n27311 , n27312 );
and ( n27314 , n27146 , n27313 );
and ( n27315 , n27123 , n27313 );
or ( n27316 , n27147 , n27314 , n27315 );
xor ( n27317 , n26762 , n26764 );
xor ( n27318 , n27317 , n26811 );
and ( n27319 , n27316 , n27318 );
xor ( n27320 , n26864 , n26904 );
xor ( n27321 , n27320 , n27054 );
xor ( n27322 , n26931 , n27048 );
xor ( n27323 , n27322 , n27051 );
xor ( n27324 , n27120 , n27122 );
and ( n27325 , n27323 , n27324 );
xor ( n27326 , n27129 , n27131 );
xor ( n27327 , n27149 , n27151 );
xor ( n27328 , n27327 , n27154 );
and ( n27329 , n26399 , n21085 );
and ( n27330 , n26148 , n21178 );
and ( n27331 , n27329 , n27330 );
xor ( n27332 , n27236 , n27237 );
xor ( n27333 , n27332 , n27239 );
and ( n27334 , n27330 , n27333 );
and ( n27335 , n27329 , n27333 );
or ( n27336 , n27331 , n27334 , n27335 );
xor ( n27337 , n27022 , n27023 );
xor ( n27338 , n27337 , n27025 );
and ( n27339 , n27336 , n27338 );
xor ( n27340 , n26981 , n26982 );
xor ( n27341 , n27340 , n26984 );
and ( n27342 , n27338 , n27341 );
and ( n27343 , n27336 , n27341 );
or ( n27344 , n27339 , n27342 , n27343 );
not ( n27345 , n27344 );
xor ( n27346 , n27161 , n27163 );
xor ( n27347 , n27346 , n27166 );
and ( n27348 , n27345 , n27347 );
and ( n27349 , n27328 , n27348 );
buf ( n27350 , n27344 );
and ( n27351 , n27348 , n27350 );
and ( n27352 , n27328 , n27350 );
or ( n27353 , n27349 , n27351 , n27352 );
and ( n27354 , n27326 , n27353 );
and ( n27355 , n25623 , n21527 );
and ( n27356 , n25451 , n21666 );
and ( n27357 , n27355 , n27356 );
and ( n27358 , n24993 , n21990 );
and ( n27359 , n27356 , n27358 );
and ( n27360 , n27355 , n27358 );
or ( n27361 , n27357 , n27359 , n27360 );
xor ( n27362 , n26972 , n26973 );
xor ( n27363 , n27362 , n26975 );
and ( n27364 , n27361 , n27363 );
xor ( n27365 , n27201 , n27202 );
xor ( n27366 , n27365 , n27204 );
and ( n27367 , n27363 , n27366 );
and ( n27368 , n27361 , n27366 );
or ( n27369 , n27364 , n27367 , n27368 );
xor ( n27370 , n27171 , n27172 );
xor ( n27371 , n27370 , n27174 );
xor ( n27372 , n27217 , n27219 );
xor ( n27373 , n27372 , n27222 );
and ( n27374 , n27371 , n27373 );
xor ( n27375 , n27226 , n27227 );
xor ( n27376 , n27375 , n27230 );
and ( n27377 , n27373 , n27376 );
and ( n27378 , n27371 , n27376 );
or ( n27379 , n27374 , n27377 , n27378 );
and ( n27380 , n27369 , n27379 );
and ( n27381 , n23903 , n23508 );
and ( n27382 , n23620 , n24064 );
and ( n27383 , n27381 , n27382 );
and ( n27384 , n23483 , n24540 );
and ( n27385 , n27382 , n27384 );
and ( n27386 , n27381 , n27384 );
or ( n27387 , n27383 , n27385 , n27386 );
buf ( n27388 , n17176 );
buf ( n27389 , n27388 );
and ( n27390 , n27389 , n20877 );
and ( n27391 , n27387 , n27390 );
xor ( n27392 , n27195 , n27196 );
xor ( n27393 , n27392 , n27198 );
and ( n27394 , n27390 , n27393 );
and ( n27395 , n27387 , n27393 );
or ( n27396 , n27391 , n27394 , n27395 );
xor ( n27397 , n27355 , n27356 );
xor ( n27398 , n27397 , n27358 );
xnor ( n27399 , n27244 , n27247 );
and ( n27400 , n27398 , n27399 );
and ( n27401 , n26933 , n20949 );
and ( n27402 , n24731 , n22337 );
and ( n27403 , n27401 , n27402 );
and ( n27404 , n24624 , n22562 );
and ( n27405 , n27402 , n27404 );
and ( n27406 , n27401 , n27404 );
or ( n27407 , n27403 , n27405 , n27406 );
and ( n27408 , n27399 , n27407 );
and ( n27409 , n27398 , n27407 );
or ( n27410 , n27400 , n27408 , n27409 );
and ( n27411 , n27396 , n27410 );
xor ( n27412 , n27235 , n27242 );
xor ( n27413 , n27412 , n27248 );
and ( n27414 , n27410 , n27413 );
and ( n27415 , n27396 , n27413 );
or ( n27416 , n27411 , n27414 , n27415 );
and ( n27417 , n27379 , n27416 );
and ( n27418 , n27369 , n27416 );
or ( n27419 , n27380 , n27417 , n27418 );
xor ( n27420 , n27177 , n27179 );
xor ( n27421 , n27420 , n27182 );
xor ( n27422 , n27191 , n27193 );
xor ( n27423 , n27422 , n27207 );
and ( n27424 , n27421 , n27423 );
xor ( n27425 , n27225 , n27233 );
xor ( n27426 , n27425 , n27251 );
and ( n27427 , n27423 , n27426 );
and ( n27428 , n27421 , n27426 );
or ( n27429 , n27424 , n27427 , n27428 );
and ( n27430 , n27419 , n27429 );
xor ( n27431 , n27159 , n27169 );
xor ( n27432 , n27431 , n27185 );
and ( n27433 , n27429 , n27432 );
and ( n27434 , n27419 , n27432 );
or ( n27435 , n27430 , n27433 , n27434 );
and ( n27436 , n27353 , n27435 );
and ( n27437 , n27326 , n27435 );
or ( n27438 , n27354 , n27436 , n27437 );
and ( n27439 , n27324 , n27438 );
and ( n27440 , n27323 , n27438 );
or ( n27441 , n27325 , n27439 , n27440 );
and ( n27442 , n27321 , n27441 );
xor ( n27443 , n27135 , n27137 );
xor ( n27444 , n27443 , n27140 );
xor ( n27445 , n27157 , n27188 );
xor ( n27446 , n27445 , n27286 );
and ( n27447 , n27444 , n27446 );
xor ( n27448 , n27299 , n27301 );
xor ( n27449 , n27448 , n27304 );
and ( n27450 , n27446 , n27449 );
and ( n27451 , n27444 , n27449 );
or ( n27452 , n27447 , n27450 , n27451 );
xor ( n27453 , n27125 , n27132 );
xor ( n27454 , n27453 , n27143 );
and ( n27455 , n27452 , n27454 );
xor ( n27456 , n27289 , n27307 );
xor ( n27457 , n27456 , n27310 );
and ( n27458 , n27454 , n27457 );
and ( n27459 , n27452 , n27457 );
or ( n27460 , n27455 , n27458 , n27459 );
and ( n27461 , n27441 , n27460 );
and ( n27462 , n27321 , n27460 );
or ( n27463 , n27442 , n27461 , n27462 );
and ( n27464 , n27318 , n27463 );
and ( n27465 , n27316 , n27463 );
or ( n27466 , n27319 , n27464 , n27465 );
and ( n27467 , n27074 , n27466 );
and ( n27468 , n27072 , n27466 );
or ( n27469 , n27075 , n27467 , n27468 );
and ( n27470 , n26822 , n27469 );
and ( n27471 , n26820 , n27469 );
or ( n27472 , n26823 , n27470 , n27471 );
and ( n27473 , n26758 , n27472 );
xor ( n27474 , n26758 , n27472 );
xor ( n27475 , n26820 , n26822 );
xor ( n27476 , n27475 , n27469 );
xor ( n27477 , n27057 , n27059 );
xor ( n27478 , n27477 , n27069 );
xor ( n27479 , n27062 , n27064 );
xor ( n27480 , n27479 , n27066 );
xor ( n27481 , n27123 , n27146 );
xor ( n27482 , n27481 , n27313 );
and ( n27483 , n27480 , n27482 );
xor ( n27484 , n27210 , n27254 );
xor ( n27485 , n27484 , n27283 );
xor ( n27486 , n27291 , n27293 );
xor ( n27487 , n27486 , n27296 );
and ( n27488 , n27485 , n27487 );
xor ( n27489 , n27275 , n27277 );
xor ( n27490 , n27489 , n27280 );
xor ( n27491 , n27345 , n27347 );
and ( n27492 , n27490 , n27491 );
and ( n27493 , n26782 , n20949 );
and ( n27494 , n24624 , n22337 );
and ( n27495 , n27493 , n27494 );
and ( n27496 , n24052 , n22987 );
and ( n27497 , n27494 , n27496 );
and ( n27498 , n27493 , n27496 );
or ( n27499 , n27495 , n27497 , n27498 );
and ( n27500 , n26980 , n20890 );
and ( n27501 , n26933 , n20909 );
and ( n27502 , n27500 , n27501 );
and ( n27503 , n24337 , n22784 );
and ( n27504 , n27501 , n27503 );
and ( n27505 , n27500 , n27503 );
or ( n27506 , n27502 , n27504 , n27505 );
and ( n27507 , n27499 , n27506 );
and ( n27508 , n23336 , n25026 );
and ( n27509 , n22824 , n26376 );
and ( n27510 , n27508 , n27509 );
and ( n27511 , n22702 , n26876 );
and ( n27512 , n27509 , n27511 );
and ( n27513 , n27508 , n27511 );
or ( n27514 , n27510 , n27512 , n27513 );
buf ( n27515 , n22542 );
buf ( n27516 , n27515 );
and ( n27517 , n23089 , n25617 );
and ( n27518 , n27516 , n27517 );
and ( n27519 , n22936 , n26229 );
and ( n27520 , n27517 , n27519 );
and ( n27521 , n27516 , n27519 );
or ( n27522 , n27518 , n27520 , n27521 );
and ( n27523 , n27514 , n27522 );
and ( n27524 , n24731 , n22172 );
and ( n27525 , n27522 , n27524 );
and ( n27526 , n27514 , n27524 );
or ( n27527 , n27523 , n27525 , n27526 );
and ( n27528 , n27506 , n27527 );
and ( n27529 , n27499 , n27527 );
or ( n27530 , n27507 , n27528 , n27529 );
and ( n27531 , n27491 , n27530 );
and ( n27532 , n27490 , n27530 );
or ( n27533 , n27492 , n27531 , n27532 );
and ( n27534 , n27487 , n27533 );
and ( n27535 , n27485 , n27533 );
or ( n27536 , n27488 , n27534 , n27535 );
xor ( n27537 , n27262 , n27269 );
xor ( n27538 , n27537 , n27272 );
xor ( n27539 , n27361 , n27363 );
xor ( n27540 , n27539 , n27366 );
and ( n27541 , n27538 , n27540 );
xor ( n27542 , n27336 , n27338 );
xor ( n27543 , n27542 , n27341 );
and ( n27544 , n27540 , n27543 );
and ( n27545 , n27538 , n27543 );
or ( n27546 , n27541 , n27544 , n27545 );
and ( n27547 , n24337 , n22987 );
and ( n27548 , n24052 , n23322 );
and ( n27549 , n27547 , n27548 );
and ( n27550 , n23742 , n23758 );
and ( n27551 , n27548 , n27550 );
and ( n27552 , n27547 , n27550 );
or ( n27553 , n27549 , n27551 , n27552 );
and ( n27554 , n23483 , n25026 );
and ( n27555 , n22936 , n26376 );
and ( n27556 , n27554 , n27555 );
buf ( n27557 , n10629 );
buf ( n27558 , n27557 );
and ( n27559 , n22589 , n27558 );
and ( n27560 , n27555 , n27559 );
and ( n27561 , n27554 , n27559 );
or ( n27562 , n27556 , n27560 , n27561 );
and ( n27563 , n23215 , n25284 );
and ( n27564 , n27562 , n27563 );
and ( n27565 , n22589 , n27246 );
not ( n27566 , n27565 );
and ( n27567 , n27563 , n27566 );
and ( n27568 , n27562 , n27566 );
or ( n27569 , n27564 , n27567 , n27568 );
and ( n27570 , n27553 , n27569 );
and ( n27571 , n25742 , n21429 );
and ( n27572 , n27569 , n27571 );
and ( n27573 , n27553 , n27571 );
or ( n27574 , n27570 , n27572 , n27573 );
xor ( n27575 , n27256 , n27257 );
xor ( n27576 , n27575 , n27259 );
xor ( n27577 , n27263 , n27264 );
xor ( n27578 , n27577 , n27266 );
and ( n27579 , n27576 , n27578 );
xor ( n27580 , n27387 , n27390 );
xor ( n27581 , n27580 , n27393 );
and ( n27582 , n27578 , n27581 );
and ( n27583 , n27576 , n27581 );
or ( n27584 , n27579 , n27582 , n27583 );
and ( n27585 , n27574 , n27584 );
xor ( n27586 , n27329 , n27330 );
xor ( n27587 , n27586 , n27333 );
buf ( n27588 , n27565 );
and ( n27589 , n27587 , n27588 );
buf ( n27590 , n17217 );
buf ( n27591 , n27590 );
and ( n27592 , n27591 , n20877 );
and ( n27593 , n26678 , n21085 );
and ( n27594 , n27592 , n27593 );
and ( n27595 , n25451 , n21990 );
and ( n27596 , n24731 , n22562 );
and ( n27597 , n27595 , n27596 );
and ( n27598 , n23903 , n23758 );
and ( n27599 , n27596 , n27598 );
and ( n27600 , n27595 , n27598 );
or ( n27601 , n27597 , n27599 , n27600 );
and ( n27602 , n27593 , n27601 );
and ( n27603 , n27592 , n27601 );
or ( n27604 , n27594 , n27602 , n27603 );
and ( n27605 , n27588 , n27604 );
and ( n27606 , n27587 , n27604 );
or ( n27607 , n27589 , n27605 , n27606 );
and ( n27608 , n27584 , n27607 );
and ( n27609 , n27574 , n27607 );
or ( n27610 , n27585 , n27608 , n27609 );
and ( n27611 , n27546 , n27610 );
xor ( n27612 , n27369 , n27379 );
xor ( n27613 , n27612 , n27416 );
and ( n27614 , n27610 , n27613 );
and ( n27615 , n27546 , n27613 );
or ( n27616 , n27611 , n27614 , n27615 );
xor ( n27617 , n27328 , n27348 );
xor ( n27618 , n27617 , n27350 );
and ( n27619 , n27616 , n27618 );
xor ( n27620 , n27419 , n27429 );
xor ( n27621 , n27620 , n27432 );
and ( n27622 , n27618 , n27621 );
and ( n27623 , n27616 , n27621 );
or ( n27624 , n27619 , n27622 , n27623 );
and ( n27625 , n27536 , n27624 );
xor ( n27626 , n27326 , n27353 );
xor ( n27627 , n27626 , n27435 );
and ( n27628 , n27624 , n27627 );
and ( n27629 , n27536 , n27627 );
or ( n27630 , n27625 , n27628 , n27629 );
xor ( n27631 , n27323 , n27324 );
xor ( n27632 , n27631 , n27438 );
and ( n27633 , n27630 , n27632 );
xor ( n27634 , n27452 , n27454 );
xor ( n27635 , n27634 , n27457 );
and ( n27636 , n27632 , n27635 );
and ( n27637 , n27630 , n27635 );
or ( n27638 , n27633 , n27636 , n27637 );
and ( n27639 , n27482 , n27638 );
and ( n27640 , n27480 , n27638 );
or ( n27641 , n27483 , n27639 , n27640 );
and ( n27642 , n27478 , n27641 );
xor ( n27643 , n27316 , n27318 );
xor ( n27644 , n27643 , n27463 );
and ( n27645 , n27641 , n27644 );
and ( n27646 , n27478 , n27644 );
or ( n27647 , n27642 , n27645 , n27646 );
xor ( n27648 , n27072 , n27074 );
xor ( n27649 , n27648 , n27466 );
and ( n27650 , n27647 , n27649 );
xor ( n27651 , n27478 , n27641 );
xor ( n27652 , n27651 , n27644 );
xor ( n27653 , n27321 , n27441 );
xor ( n27654 , n27653 , n27460 );
xor ( n27655 , n27480 , n27482 );
xor ( n27656 , n27655 , n27638 );
and ( n27657 , n27654 , n27656 );
xor ( n27658 , n27444 , n27446 );
xor ( n27659 , n27658 , n27449 );
xor ( n27660 , n27421 , n27423 );
xor ( n27661 , n27660 , n27426 );
and ( n27662 , n26980 , n20909 );
and ( n27663 , n26148 , n21296 );
and ( n27664 , n27662 , n27663 );
and ( n27665 , n24546 , n22784 );
and ( n27666 , n27663 , n27665 );
and ( n27667 , n27662 , n27665 );
or ( n27668 , n27664 , n27666 , n27667 );
and ( n27669 , n22824 , n26876 );
and ( n27670 , n22702 , n27246 );
and ( n27671 , n27669 , n27670 );
not ( n27672 , n27515 );
and ( n27673 , n27670 , n27672 );
and ( n27674 , n27669 , n27672 );
or ( n27675 , n27671 , n27673 , n27674 );
and ( n27676 , n25451 , n21827 );
and ( n27677 , n27675 , n27676 );
and ( n27678 , n24993 , n22172 );
and ( n27679 , n27676 , n27678 );
and ( n27680 , n27675 , n27678 );
or ( n27681 , n27677 , n27679 , n27680 );
and ( n27682 , n27668 , n27681 );
xor ( n27683 , n27493 , n27494 );
xor ( n27684 , n27683 , n27496 );
and ( n27685 , n27681 , n27684 );
and ( n27686 , n27668 , n27684 );
or ( n27687 , n27682 , n27685 , n27686 );
and ( n27688 , n24052 , n23508 );
and ( n27689 , n23742 , n24064 );
and ( n27690 , n27688 , n27689 );
and ( n27691 , n23620 , n24540 );
and ( n27692 , n27689 , n27691 );
and ( n27693 , n27688 , n27691 );
or ( n27694 , n27690 , n27692 , n27693 );
and ( n27695 , n25220 , n21990 );
and ( n27696 , n27694 , n27695 );
xor ( n27697 , n27516 , n27517 );
xor ( n27698 , n27697 , n27519 );
and ( n27699 , n27695 , n27698 );
and ( n27700 , n27694 , n27698 );
or ( n27701 , n27696 , n27699 , n27700 );
xor ( n27702 , n27211 , n27212 );
xor ( n27703 , n27702 , n27214 );
and ( n27704 , n27701 , n27703 );
xor ( n27705 , n27500 , n27501 );
xor ( n27706 , n27705 , n27503 );
and ( n27707 , n27703 , n27706 );
and ( n27708 , n27701 , n27706 );
or ( n27709 , n27704 , n27707 , n27708 );
and ( n27710 , n27687 , n27709 );
xor ( n27711 , n27499 , n27506 );
xor ( n27712 , n27711 , n27527 );
and ( n27713 , n27709 , n27712 );
and ( n27714 , n27687 , n27712 );
or ( n27715 , n27710 , n27713 , n27714 );
and ( n27716 , n27661 , n27715 );
xor ( n27717 , n27371 , n27373 );
xor ( n27718 , n27717 , n27376 );
xor ( n27719 , n27396 , n27410 );
xor ( n27720 , n27719 , n27413 );
and ( n27721 , n27718 , n27720 );
and ( n27722 , n26399 , n21178 );
and ( n27723 , n25742 , n21527 );
and ( n27724 , n27722 , n27723 );
and ( n27725 , n25623 , n21666 );
and ( n27726 , n27723 , n27725 );
and ( n27727 , n27722 , n27725 );
or ( n27728 , n27724 , n27726 , n27727 );
and ( n27729 , n23336 , n25284 );
and ( n27730 , n23215 , n25617 );
and ( n27731 , n27729 , n27730 );
and ( n27732 , n23089 , n26229 );
and ( n27733 , n27730 , n27732 );
and ( n27734 , n27729 , n27732 );
or ( n27735 , n27731 , n27733 , n27734 );
and ( n27736 , n27389 , n20890 );
and ( n27737 , n27735 , n27736 );
xor ( n27738 , n27508 , n27509 );
xor ( n27739 , n27738 , n27511 );
and ( n27740 , n27736 , n27739 );
and ( n27741 , n27735 , n27739 );
or ( n27742 , n27737 , n27740 , n27741 );
and ( n27743 , n27728 , n27742 );
xor ( n27744 , n27514 , n27522 );
xor ( n27745 , n27744 , n27524 );
and ( n27746 , n27742 , n27745 );
and ( n27747 , n27728 , n27745 );
or ( n27748 , n27743 , n27746 , n27747 );
and ( n27749 , n27720 , n27748 );
and ( n27750 , n27718 , n27748 );
or ( n27751 , n27721 , n27749 , n27750 );
and ( n27752 , n27715 , n27751 );
and ( n27753 , n27661 , n27751 );
or ( n27754 , n27716 , n27752 , n27753 );
and ( n27755 , n27591 , n20890 );
and ( n27756 , n27389 , n20909 );
and ( n27757 , n27755 , n27756 );
and ( n27758 , n26399 , n21296 );
and ( n27759 , n27756 , n27758 );
and ( n27760 , n27755 , n27758 );
or ( n27761 , n27757 , n27759 , n27760 );
and ( n27762 , n25623 , n21827 );
and ( n27763 , n25220 , n22172 );
and ( n27764 , n27762 , n27763 );
and ( n27765 , n24993 , n22337 );
and ( n27766 , n27763 , n27765 );
and ( n27767 , n27762 , n27765 );
or ( n27768 , n27764 , n27766 , n27767 );
and ( n27769 , n27761 , n27768 );
xor ( n27770 , n27401 , n27402 );
xor ( n27771 , n27770 , n27404 );
and ( n27772 , n27768 , n27771 );
and ( n27773 , n27761 , n27771 );
or ( n27774 , n27769 , n27772 , n27773 );
and ( n27775 , n26782 , n21085 );
and ( n27776 , n26678 , n21178 );
and ( n27777 , n27775 , n27776 );
xor ( n27778 , n27669 , n27670 );
xor ( n27779 , n27778 , n27672 );
and ( n27780 , n27776 , n27779 );
and ( n27781 , n27775 , n27779 );
or ( n27782 , n27777 , n27780 , n27781 );
xor ( n27783 , n27662 , n27663 );
xor ( n27784 , n27783 , n27665 );
and ( n27785 , n27782 , n27784 );
xor ( n27786 , n27675 , n27676 );
xor ( n27787 , n27786 , n27678 );
and ( n27788 , n27784 , n27787 );
and ( n27789 , n27782 , n27787 );
or ( n27790 , n27785 , n27788 , n27789 );
and ( n27791 , n27774 , n27790 );
xor ( n27792 , n27668 , n27681 );
xor ( n27793 , n27792 , n27684 );
and ( n27794 , n27790 , n27793 );
and ( n27795 , n27774 , n27793 );
or ( n27796 , n27791 , n27794 , n27795 );
xor ( n27797 , n27398 , n27399 );
xor ( n27798 , n27797 , n27407 );
xor ( n27799 , n27553 , n27569 );
xor ( n27800 , n27799 , n27571 );
and ( n27801 , n27798 , n27800 );
and ( n27802 , n26980 , n20949 );
and ( n27803 , n24546 , n22987 );
and ( n27804 , n27802 , n27803 );
and ( n27805 , n24337 , n23322 );
and ( n27806 , n27803 , n27805 );
and ( n27807 , n27802 , n27805 );
or ( n27808 , n27804 , n27806 , n27807 );
and ( n27809 , n25959 , n21429 );
and ( n27810 , n27808 , n27809 );
xor ( n27811 , n27562 , n27563 );
xor ( n27812 , n27811 , n27566 );
and ( n27813 , n27809 , n27812 );
and ( n27814 , n27808 , n27812 );
or ( n27815 , n27810 , n27813 , n27814 );
and ( n27816 , n27800 , n27815 );
and ( n27817 , n27798 , n27815 );
or ( n27818 , n27801 , n27816 , n27817 );
and ( n27819 , n27796 , n27818 );
and ( n27820 , n23620 , n25026 );
and ( n27821 , n23215 , n26229 );
and ( n27822 , n27820 , n27821 );
and ( n27823 , n23089 , n26376 );
and ( n27824 , n27821 , n27823 );
and ( n27825 , n27820 , n27823 );
or ( n27826 , n27822 , n27824 , n27825 );
and ( n27827 , n24624 , n22784 );
and ( n27828 , n27826 , n27827 );
xor ( n27829 , n27554 , n27555 );
xor ( n27830 , n27829 , n27559 );
and ( n27831 , n27827 , n27830 );
and ( n27832 , n27826 , n27830 );
or ( n27833 , n27828 , n27831 , n27832 );
and ( n27834 , n26782 , n21039 );
and ( n27835 , n27833 , n27834 );
xor ( n27836 , n27381 , n27382 );
xor ( n27837 , n27836 , n27384 );
and ( n27838 , n27834 , n27837 );
and ( n27839 , n27833 , n27837 );
or ( n27840 , n27835 , n27838 , n27839 );
xor ( n27841 , n27547 , n27548 );
xor ( n27842 , n27841 , n27550 );
xor ( n27843 , n27735 , n27736 );
xor ( n27844 , n27843 , n27739 );
or ( n27845 , n27842 , n27844 );
and ( n27846 , n27840 , n27845 );
xor ( n27847 , n27761 , n27768 );
xor ( n27848 , n27847 , n27771 );
and ( n27849 , n26782 , n21178 );
and ( n27850 , n26148 , n21527 );
and ( n27851 , n27849 , n27850 );
and ( n27852 , n25959 , n21666 );
and ( n27853 , n27850 , n27852 );
and ( n27854 , n27849 , n27852 );
or ( n27855 , n27851 , n27853 , n27854 );
xor ( n27856 , n27755 , n27756 );
xor ( n27857 , n27856 , n27758 );
and ( n27858 , n27855 , n27857 );
and ( n27859 , n27848 , n27858 );
xor ( n27860 , n27802 , n27803 );
xor ( n27861 , n27860 , n27805 );
buf ( n27862 , n17247 );
buf ( n27863 , n27862 );
and ( n27864 , n27863 , n20877 );
and ( n27865 , n25959 , n21527 );
xor ( n27866 , n27864 , n27865 );
and ( n27867 , n25742 , n21666 );
xor ( n27868 , n27866 , n27867 );
and ( n27869 , n27861 , n27868 );
and ( n27870 , n24337 , n23508 );
and ( n27871 , n23903 , n24064 );
and ( n27872 , n27870 , n27871 );
and ( n27873 , n23742 , n24540 );
and ( n27874 , n27871 , n27873 );
and ( n27875 , n27870 , n27873 );
or ( n27876 , n27872 , n27874 , n27875 );
and ( n27877 , n27868 , n27876 );
and ( n27878 , n27861 , n27876 );
or ( n27879 , n27869 , n27877 , n27878 );
and ( n27880 , n27858 , n27879 );
and ( n27881 , n27848 , n27879 );
or ( n27882 , n27859 , n27880 , n27881 );
and ( n27883 , n27845 , n27882 );
and ( n27884 , n27840 , n27882 );
or ( n27885 , n27846 , n27883 , n27884 );
and ( n27886 , n27818 , n27885 );
and ( n27887 , n27796 , n27885 );
or ( n27888 , n27819 , n27886 , n27887 );
xor ( n27889 , n27490 , n27491 );
xor ( n27890 , n27889 , n27530 );
and ( n27891 , n27888 , n27890 );
xor ( n27892 , n27546 , n27610 );
xor ( n27893 , n27892 , n27613 );
and ( n27894 , n27890 , n27893 );
and ( n27895 , n27888 , n27893 );
or ( n27896 , n27891 , n27894 , n27895 );
and ( n27897 , n27754 , n27896 );
xor ( n27898 , n27485 , n27487 );
xor ( n27899 , n27898 , n27533 );
and ( n27900 , n27896 , n27899 );
and ( n27901 , n27754 , n27899 );
or ( n27902 , n27897 , n27900 , n27901 );
and ( n27903 , n27659 , n27902 );
xor ( n27904 , n27536 , n27624 );
xor ( n27905 , n27904 , n27627 );
and ( n27906 , n27902 , n27905 );
and ( n27907 , n27659 , n27905 );
or ( n27908 , n27903 , n27906 , n27907 );
xor ( n27909 , n27630 , n27632 );
xor ( n27910 , n27909 , n27635 );
and ( n27911 , n27908 , n27910 );
xor ( n27912 , n27616 , n27618 );
xor ( n27913 , n27912 , n27621 );
xor ( n27914 , n27538 , n27540 );
xor ( n27915 , n27914 , n27543 );
xor ( n27916 , n27574 , n27584 );
xor ( n27917 , n27916 , n27607 );
and ( n27918 , n27915 , n27917 );
xor ( n27919 , n27687 , n27709 );
xor ( n27920 , n27919 , n27712 );
and ( n27921 , n27917 , n27920 );
and ( n27922 , n27915 , n27920 );
or ( n27923 , n27918 , n27921 , n27922 );
and ( n27924 , n24624 , n22987 );
and ( n27925 , n24546 , n23322 );
and ( n27926 , n27924 , n27925 );
and ( n27927 , n24052 , n23758 );
and ( n27928 , n27925 , n27927 );
and ( n27929 , n27924 , n27927 );
or ( n27930 , n27926 , n27928 , n27929 );
and ( n27931 , n26933 , n21039 );
and ( n27932 , n27930 , n27931 );
and ( n27933 , n26148 , n21429 );
and ( n27934 , n27931 , n27933 );
and ( n27935 , n27930 , n27933 );
or ( n27936 , n27932 , n27934 , n27935 );
xor ( n27937 , n27722 , n27723 );
xor ( n27938 , n27937 , n27725 );
and ( n27939 , n27936 , n27938 );
xor ( n27940 , n27694 , n27695 );
xor ( n27941 , n27940 , n27698 );
and ( n27942 , n27938 , n27941 );
and ( n27943 , n27936 , n27941 );
or ( n27944 , n27939 , n27942 , n27943 );
xor ( n27945 , n27728 , n27742 );
xor ( n27946 , n27945 , n27745 );
or ( n27947 , n27944 , n27946 );
xor ( n27948 , n27576 , n27578 );
xor ( n27949 , n27948 , n27581 );
xor ( n27950 , n27587 , n27588 );
xor ( n27951 , n27950 , n27604 );
and ( n27952 , n27949 , n27951 );
xor ( n27953 , n27701 , n27703 );
xor ( n27954 , n27953 , n27706 );
and ( n27955 , n27951 , n27954 );
and ( n27956 , n27949 , n27954 );
or ( n27957 , n27952 , n27955 , n27956 );
and ( n27958 , n27947 , n27957 );
xor ( n27959 , n27774 , n27790 );
xor ( n27960 , n27959 , n27793 );
buf ( n27961 , n17268 );
buf ( n27962 , n27961 );
and ( n27963 , n27962 , n20877 );
and ( n27964 , n26933 , n21085 );
and ( n27965 , n27963 , n27964 );
xor ( n27966 , n27870 , n27871 );
xor ( n27967 , n27966 , n27873 );
and ( n27968 , n27964 , n27967 );
and ( n27969 , n27963 , n27967 );
or ( n27970 , n27965 , n27968 , n27969 );
xor ( n27971 , n27762 , n27763 );
xor ( n27972 , n27971 , n27765 );
and ( n27973 , n27970 , n27972 );
xor ( n27974 , n27826 , n27827 );
xor ( n27975 , n27974 , n27830 );
and ( n27976 , n27972 , n27975 );
and ( n27977 , n27970 , n27975 );
or ( n27978 , n27973 , n27976 , n27977 );
xor ( n27979 , n27782 , n27784 );
xor ( n27980 , n27979 , n27787 );
and ( n27981 , n27978 , n27980 );
and ( n27982 , n27960 , n27981 );
and ( n27983 , n27864 , n27865 );
and ( n27984 , n27865 , n27867 );
and ( n27985 , n27864 , n27867 );
or ( n27986 , n27983 , n27984 , n27985 );
and ( n27987 , n23742 , n25026 );
and ( n27988 , n22936 , n27246 );
and ( n27989 , n27987 , n27988 );
and ( n27990 , n22824 , n27558 );
and ( n27991 , n27988 , n27990 );
and ( n27992 , n27987 , n27990 );
or ( n27993 , n27989 , n27991 , n27992 );
and ( n27994 , n24993 , n22562 );
and ( n27995 , n27993 , n27994 );
and ( n27996 , n23483 , n25284 );
and ( n27997 , n27994 , n27996 );
and ( n27998 , n27993 , n27996 );
or ( n27999 , n27995 , n27997 , n27998 );
xor ( n28000 , n27688 , n27689 );
xor ( n28001 , n28000 , n27691 );
and ( n28002 , n27999 , n28001 );
xor ( n28003 , n27729 , n27730 );
xor ( n28004 , n28003 , n27732 );
and ( n28005 , n28001 , n28004 );
and ( n28006 , n27999 , n28004 );
or ( n28007 , n28002 , n28005 , n28006 );
and ( n28008 , n27986 , n28007 );
and ( n28009 , n27981 , n28008 );
and ( n28010 , n27960 , n28008 );
or ( n28011 , n27982 , n28009 , n28010 );
and ( n28012 , n27957 , n28011 );
and ( n28013 , n27947 , n28011 );
or ( n28014 , n27958 , n28012 , n28013 );
and ( n28015 , n27923 , n28014 );
and ( n28016 , n27591 , n20909 );
and ( n28017 , n26678 , n21296 );
and ( n28018 , n28016 , n28017 );
and ( n28019 , n24731 , n22784 );
and ( n28020 , n28017 , n28019 );
and ( n28021 , n28016 , n28019 );
or ( n28022 , n28018 , n28020 , n28021 );
and ( n28023 , n27863 , n20890 );
and ( n28024 , n27389 , n20949 );
and ( n28025 , n28023 , n28024 );
and ( n28026 , n25623 , n21990 );
and ( n28027 , n28024 , n28026 );
and ( n28028 , n28023 , n28026 );
or ( n28029 , n28025 , n28027 , n28028 );
and ( n28030 , n28022 , n28029 );
and ( n28031 , n25220 , n22337 );
and ( n28032 , n23336 , n25617 );
and ( n28033 , n28031 , n28032 );
and ( n28034 , n22936 , n26876 );
and ( n28035 , n28032 , n28034 );
and ( n28036 , n28031 , n28034 );
or ( n28037 , n28033 , n28035 , n28036 );
and ( n28038 , n28029 , n28037 );
and ( n28039 , n28022 , n28037 );
or ( n28040 , n28030 , n28038 , n28039 );
xor ( n28041 , n27592 , n27593 );
xor ( n28042 , n28041 , n27601 );
and ( n28043 , n28040 , n28042 );
xor ( n28044 , n27808 , n27809 );
xor ( n28045 , n28044 , n27812 );
and ( n28046 , n28042 , n28045 );
and ( n28047 , n28040 , n28045 );
or ( n28048 , n28043 , n28046 , n28047 );
xor ( n28049 , n27833 , n27834 );
xor ( n28050 , n28049 , n27837 );
xnor ( n28051 , n27842 , n27844 );
and ( n28052 , n28050 , n28051 );
xor ( n28053 , n27595 , n27596 );
xor ( n28054 , n28053 , n27598 );
xor ( n28055 , n27775 , n27776 );
xor ( n28056 , n28055 , n27779 );
and ( n28057 , n28054 , n28056 );
xor ( n28058 , n27855 , n27857 );
and ( n28059 , n28056 , n28058 );
and ( n28060 , n28054 , n28058 );
or ( n28061 , n28057 , n28059 , n28060 );
and ( n28062 , n28051 , n28061 );
and ( n28063 , n28050 , n28061 );
or ( n28064 , n28052 , n28062 , n28063 );
and ( n28065 , n28048 , n28064 );
xor ( n28066 , n27798 , n27800 );
xor ( n28067 , n28066 , n27815 );
and ( n28068 , n28064 , n28067 );
and ( n28069 , n28048 , n28067 );
or ( n28070 , n28065 , n28068 , n28069 );
xor ( n28071 , n27718 , n27720 );
xor ( n28072 , n28071 , n27748 );
and ( n28073 , n28070 , n28072 );
xor ( n28074 , n27796 , n27818 );
xor ( n28075 , n28074 , n27885 );
and ( n28076 , n28072 , n28075 );
and ( n28077 , n28070 , n28075 );
or ( n28078 , n28073 , n28076 , n28077 );
and ( n28079 , n28014 , n28078 );
and ( n28080 , n27923 , n28078 );
or ( n28081 , n28015 , n28079 , n28080 );
and ( n28082 , n27913 , n28081 );
xor ( n28083 , n27754 , n27896 );
xor ( n28084 , n28083 , n27899 );
and ( n28085 , n28081 , n28084 );
and ( n28086 , n27913 , n28084 );
or ( n28087 , n28082 , n28085 , n28086 );
xor ( n28088 , n27659 , n27902 );
xor ( n28089 , n28088 , n27905 );
and ( n28090 , n28087 , n28089 );
xor ( n28091 , n27661 , n27715 );
xor ( n28092 , n28091 , n27751 );
xor ( n28093 , n27888 , n27890 );
xor ( n28094 , n28093 , n27893 );
and ( n28095 , n28092 , n28094 );
xor ( n28096 , n27840 , n27845 );
xor ( n28097 , n28096 , n27882 );
xnor ( n28098 , n27944 , n27946 );
and ( n28099 , n28097 , n28098 );
and ( n28100 , n22824 , n27246 );
and ( n28101 , n22702 , n27558 );
and ( n28102 , n28100 , n28101 );
xor ( n28103 , n27820 , n27821 );
xor ( n28104 , n28103 , n27823 );
and ( n28105 , n28101 , n28104 );
and ( n28106 , n28100 , n28104 );
or ( n28107 , n28102 , n28105 , n28106 );
and ( n28108 , n24052 , n24064 );
and ( n28109 , n23903 , n24540 );
and ( n28110 , n28108 , n28109 );
and ( n28111 , n23620 , n25284 );
and ( n28112 , n28109 , n28111 );
and ( n28113 , n28108 , n28111 );
or ( n28114 , n28110 , n28112 , n28113 );
buf ( n28115 , n22589 );
buf ( n28116 , n762 );
buf ( n28117 , n28116 );
buf ( n28118 , n763 );
buf ( n28119 , n28118 );
buf ( n28120 , n764 );
buf ( n28121 , n28120 );
and ( n28122 , n28119 , n28121 );
not ( n28123 , n28122 );
and ( n28124 , n28117 , n28123 );
not ( n28125 , n28124 );
and ( n28126 , n28115 , n28125 );
and ( n28127 , n28114 , n28126 );
buf ( n28128 , n17316 );
buf ( n28129 , n28128 );
and ( n28130 , n28129 , n20877 );
and ( n28131 , n27863 , n20909 );
and ( n28132 , n28130 , n28131 );
and ( n28133 , n26678 , n21429 );
and ( n28134 , n28131 , n28133 );
and ( n28135 , n28130 , n28133 );
or ( n28136 , n28132 , n28134 , n28135 );
and ( n28137 , n28126 , n28136 );
and ( n28138 , n28114 , n28136 );
or ( n28139 , n28127 , n28137 , n28138 );
and ( n28140 , n28107 , n28139 );
and ( n28141 , n25742 , n21990 );
and ( n28142 , n23336 , n26229 );
and ( n28143 , n28141 , n28142 );
and ( n28144 , n23089 , n26876 );
and ( n28145 , n28142 , n28144 );
and ( n28146 , n28141 , n28144 );
or ( n28147 , n28143 , n28145 , n28146 );
xor ( n28148 , n28023 , n28024 );
xor ( n28149 , n28148 , n28026 );
and ( n28150 , n28147 , n28149 );
xor ( n28151 , n28031 , n28032 );
xor ( n28152 , n28151 , n28034 );
and ( n28153 , n28149 , n28152 );
and ( n28154 , n28147 , n28152 );
or ( n28155 , n28150 , n28153 , n28154 );
and ( n28156 , n28139 , n28155 );
and ( n28157 , n28107 , n28155 );
or ( n28158 , n28140 , n28156 , n28157 );
xor ( n28159 , n27848 , n27858 );
xor ( n28160 , n28159 , n27879 );
and ( n28161 , n28158 , n28160 );
xor ( n28162 , n27936 , n27938 );
xor ( n28163 , n28162 , n27941 );
and ( n28164 , n28160 , n28163 );
and ( n28165 , n28158 , n28163 );
or ( n28166 , n28161 , n28164 , n28165 );
and ( n28167 , n28098 , n28166 );
and ( n28168 , n28097 , n28166 );
or ( n28169 , n28099 , n28167 , n28168 );
xor ( n28170 , n27978 , n27980 );
xor ( n28171 , n27986 , n28007 );
and ( n28172 , n28170 , n28171 );
and ( n28173 , n25220 , n22562 );
and ( n28174 , n24731 , n22987 );
and ( n28175 , n28173 , n28174 );
and ( n28176 , n24546 , n23508 );
and ( n28177 , n28174 , n28176 );
and ( n28178 , n28173 , n28176 );
or ( n28179 , n28175 , n28177 , n28178 );
and ( n28180 , n23903 , n25026 );
and ( n28181 , n23336 , n26376 );
and ( n28182 , n28180 , n28181 );
and ( n28183 , n22936 , n27558 );
and ( n28184 , n28181 , n28183 );
and ( n28185 , n28180 , n28183 );
or ( n28186 , n28182 , n28184 , n28185 );
and ( n28187 , n24624 , n23322 );
and ( n28188 , n28186 , n28187 );
and ( n28189 , n24337 , n23758 );
and ( n28190 , n28187 , n28189 );
and ( n28191 , n28186 , n28189 );
or ( n28192 , n28188 , n28190 , n28191 );
and ( n28193 , n28179 , n28192 );
and ( n28194 , n26399 , n21429 );
and ( n28195 , n28192 , n28194 );
and ( n28196 , n28179 , n28194 );
or ( n28197 , n28193 , n28195 , n28196 );
and ( n28198 , n26782 , n21296 );
and ( n28199 , n25959 , n21827 );
and ( n28200 , n28198 , n28199 );
and ( n28201 , n25623 , n22172 );
and ( n28202 , n28199 , n28201 );
and ( n28203 , n28198 , n28201 );
or ( n28204 , n28200 , n28202 , n28203 );
and ( n28205 , n23215 , n26876 );
and ( n28206 , n23089 , n27246 );
and ( n28207 , n28205 , n28206 );
buf ( n28208 , n10921 );
buf ( n28209 , n28208 );
and ( n28210 , n22824 , n28209 );
not ( n28211 , n28210 );
and ( n28212 , n28206 , n28211 );
and ( n28213 , n28205 , n28211 );
or ( n28214 , n28207 , n28212 , n28213 );
and ( n28215 , n25451 , n22337 );
and ( n28216 , n28214 , n28215 );
and ( n28217 , n24993 , n22784 );
and ( n28218 , n28215 , n28217 );
and ( n28219 , n28214 , n28217 );
or ( n28220 , n28216 , n28218 , n28219 );
and ( n28221 , n28204 , n28220 );
xor ( n28222 , n27993 , n27994 );
xor ( n28223 , n28222 , n27996 );
and ( n28224 , n28220 , n28223 );
and ( n28225 , n28204 , n28223 );
or ( n28226 , n28221 , n28224 , n28225 );
and ( n28227 , n28197 , n28226 );
xor ( n28228 , n27930 , n27931 );
xor ( n28229 , n28228 , n27933 );
and ( n28230 , n28226 , n28229 );
and ( n28231 , n28197 , n28229 );
or ( n28232 , n28227 , n28230 , n28231 );
and ( n28233 , n28171 , n28232 );
and ( n28234 , n28170 , n28232 );
or ( n28235 , n28172 , n28233 , n28234 );
and ( n28236 , n27962 , n20890 );
and ( n28237 , n27591 , n20949 );
and ( n28238 , n28236 , n28237 );
xor ( n28239 , n27987 , n27988 );
xor ( n28240 , n28239 , n27990 );
and ( n28241 , n28237 , n28240 );
and ( n28242 , n28236 , n28240 );
or ( n28243 , n28238 , n28241 , n28242 );
and ( n28244 , n26980 , n21039 );
and ( n28245 , n28243 , n28244 );
xor ( n28246 , n27924 , n27925 );
xor ( n28247 , n28246 , n27927 );
and ( n28248 , n28244 , n28247 );
and ( n28249 , n28243 , n28247 );
or ( n28250 , n28245 , n28248 , n28249 );
xor ( n28251 , n27999 , n28001 );
xor ( n28252 , n28251 , n28004 );
or ( n28253 , n28250 , n28252 );
xor ( n28254 , n27861 , n27868 );
xor ( n28255 , n28254 , n27876 );
xor ( n28256 , n28022 , n28029 );
xor ( n28257 , n28256 , n28037 );
and ( n28258 , n28255 , n28257 );
xor ( n28259 , n27970 , n27972 );
xor ( n28260 , n28259 , n27975 );
and ( n28261 , n28257 , n28260 );
and ( n28262 , n28255 , n28260 );
or ( n28263 , n28258 , n28261 , n28262 );
and ( n28264 , n28253 , n28263 );
buf ( n28265 , n28210 );
and ( n28266 , n23483 , n25617 );
and ( n28267 , n28265 , n28266 );
and ( n28268 , n23215 , n26376 );
and ( n28269 , n28266 , n28268 );
and ( n28270 , n28265 , n28268 );
or ( n28271 , n28267 , n28269 , n28270 );
and ( n28272 , n25742 , n21827 );
and ( n28273 , n28271 , n28272 );
and ( n28274 , n25451 , n22172 );
and ( n28275 , n28272 , n28274 );
and ( n28276 , n28271 , n28274 );
or ( n28277 , n28273 , n28275 , n28276 );
xor ( n28278 , n27963 , n27964 );
xor ( n28279 , n28278 , n27967 );
and ( n28280 , n26980 , n21085 );
and ( n28281 , n26933 , n21178 );
and ( n28282 , n28280 , n28281 );
xor ( n28283 , n28108 , n28109 );
xor ( n28284 , n28283 , n28111 );
and ( n28285 , n28281 , n28284 );
and ( n28286 , n28280 , n28284 );
or ( n28287 , n28282 , n28285 , n28286 );
and ( n28288 , n28279 , n28287 );
and ( n28289 , n22702 , n28209 );
xor ( n28290 , n28198 , n28199 );
xor ( n28291 , n28290 , n28201 );
and ( n28292 , n28289 , n28291 );
xor ( n28293 , n28115 , n28125 );
and ( n28294 , n28291 , n28293 );
and ( n28295 , n28289 , n28293 );
or ( n28296 , n28292 , n28294 , n28295 );
and ( n28297 , n28287 , n28296 );
and ( n28298 , n28279 , n28296 );
or ( n28299 , n28288 , n28297 , n28298 );
and ( n28300 , n28277 , n28299 );
and ( n28301 , n23742 , n25284 );
and ( n28302 , n23620 , n25617 );
and ( n28303 , n28301 , n28302 );
and ( n28304 , n23483 , n26229 );
and ( n28305 , n28302 , n28304 );
and ( n28306 , n28301 , n28304 );
or ( n28307 , n28303 , n28305 , n28306 );
and ( n28308 , n27863 , n20949 );
and ( n28309 , n24731 , n23322 );
and ( n28310 , n28308 , n28309 );
and ( n28311 , n24546 , n23758 );
and ( n28312 , n28309 , n28311 );
and ( n28313 , n28308 , n28311 );
or ( n28314 , n28310 , n28312 , n28313 );
and ( n28315 , n28307 , n28314 );
and ( n28316 , n27591 , n21039 );
and ( n28317 , n26782 , n21429 );
and ( n28318 , n28316 , n28317 );
and ( n28319 , n25451 , n22562 );
and ( n28320 , n28317 , n28319 );
and ( n28321 , n28316 , n28319 );
or ( n28322 , n28318 , n28320 , n28321 );
and ( n28323 , n28314 , n28322 );
and ( n28324 , n28307 , n28322 );
or ( n28325 , n28315 , n28323 , n28324 );
and ( n28326 , n24624 , n23508 );
and ( n28327 , n24337 , n24064 );
and ( n28328 , n28326 , n28327 );
and ( n28329 , n24052 , n24540 );
and ( n28330 , n28327 , n28329 );
and ( n28331 , n28326 , n28329 );
or ( n28332 , n28328 , n28330 , n28331 );
xor ( n28333 , n28130 , n28131 );
xor ( n28334 , n28333 , n28133 );
and ( n28335 , n28332 , n28334 );
xor ( n28336 , n28141 , n28142 );
xor ( n28337 , n28336 , n28144 );
and ( n28338 , n28334 , n28337 );
and ( n28339 , n28332 , n28337 );
or ( n28340 , n28335 , n28338 , n28339 );
and ( n28341 , n28325 , n28340 );
xor ( n28342 , n28100 , n28101 );
xor ( n28343 , n28342 , n28104 );
and ( n28344 , n28340 , n28343 );
and ( n28345 , n28325 , n28343 );
or ( n28346 , n28341 , n28344 , n28345 );
and ( n28347 , n28299 , n28346 );
and ( n28348 , n28277 , n28346 );
or ( n28349 , n28300 , n28347 , n28348 );
and ( n28350 , n28263 , n28349 );
and ( n28351 , n28253 , n28349 );
or ( n28352 , n28264 , n28350 , n28351 );
and ( n28353 , n28235 , n28352 );
xor ( n28354 , n27949 , n27951 );
xor ( n28355 , n28354 , n27954 );
and ( n28356 , n28352 , n28355 );
and ( n28357 , n28235 , n28355 );
or ( n28358 , n28353 , n28356 , n28357 );
and ( n28359 , n28169 , n28358 );
xor ( n28360 , n27915 , n27917 );
xor ( n28361 , n28360 , n27920 );
and ( n28362 , n28358 , n28361 );
and ( n28363 , n28169 , n28361 );
or ( n28364 , n28359 , n28362 , n28363 );
and ( n28365 , n28094 , n28364 );
and ( n28366 , n28092 , n28364 );
or ( n28367 , n28095 , n28365 , n28366 );
xor ( n28368 , n27913 , n28081 );
xor ( n28369 , n28368 , n28084 );
and ( n28370 , n28367 , n28369 );
xor ( n28371 , n27923 , n28014 );
xor ( n28372 , n28371 , n28078 );
xor ( n28373 , n27947 , n27957 );
xor ( n28374 , n28373 , n28011 );
xor ( n28375 , n28070 , n28072 );
xor ( n28376 , n28375 , n28075 );
and ( n28377 , n28374 , n28376 );
xor ( n28378 , n27960 , n27981 );
xor ( n28379 , n28378 , n28008 );
xor ( n28380 , n28048 , n28064 );
xor ( n28381 , n28380 , n28067 );
and ( n28382 , n28379 , n28381 );
xor ( n28383 , n28040 , n28042 );
xor ( n28384 , n28383 , n28045 );
xor ( n28385 , n28050 , n28051 );
xor ( n28386 , n28385 , n28061 );
and ( n28387 , n28384 , n28386 );
xor ( n28388 , n28054 , n28056 );
xor ( n28389 , n28388 , n28058 );
xor ( n28390 , n28107 , n28139 );
xor ( n28391 , n28390 , n28155 );
and ( n28392 , n28389 , n28391 );
xor ( n28393 , n28197 , n28226 );
xor ( n28394 , n28393 , n28229 );
and ( n28395 , n28391 , n28394 );
and ( n28396 , n28389 , n28394 );
or ( n28397 , n28392 , n28395 , n28396 );
and ( n28398 , n28386 , n28397 );
and ( n28399 , n28384 , n28397 );
or ( n28400 , n28387 , n28398 , n28399 );
and ( n28401 , n28381 , n28400 );
and ( n28402 , n28379 , n28400 );
or ( n28403 , n28382 , n28401 , n28402 );
and ( n28404 , n28376 , n28403 );
and ( n28405 , n28374 , n28403 );
or ( n28406 , n28377 , n28404 , n28405 );
and ( n28407 , n28372 , n28406 );
xor ( n28408 , n28092 , n28094 );
xor ( n28409 , n28408 , n28364 );
and ( n28410 , n28406 , n28409 );
and ( n28411 , n28372 , n28409 );
or ( n28412 , n28407 , n28410 , n28411 );
and ( n28413 , n28369 , n28412 );
and ( n28414 , n28367 , n28412 );
or ( n28415 , n28370 , n28413 , n28414 );
and ( n28416 , n28089 , n28415 );
and ( n28417 , n28087 , n28415 );
or ( n28418 , n28090 , n28416 , n28417 );
and ( n28419 , n27910 , n28418 );
and ( n28420 , n27908 , n28418 );
or ( n28421 , n27911 , n28419 , n28420 );
and ( n28422 , n27656 , n28421 );
and ( n28423 , n27654 , n28421 );
or ( n28424 , n27657 , n28422 , n28423 );
or ( n28425 , n27652 , n28424 );
and ( n28426 , n27649 , n28425 );
and ( n28427 , n27647 , n28425 );
or ( n28428 , n27650 , n28426 , n28427 );
and ( n28429 , n27476 , n28428 );
xor ( n28430 , n27476 , n28428 );
xor ( n28431 , n27647 , n27649 );
xor ( n28432 , n28431 , n28425 );
xnor ( n28433 , n27652 , n28424 );
xor ( n28434 , n27654 , n27656 );
xor ( n28435 , n28434 , n28421 );
not ( n28436 , n28435 );
xor ( n28437 , n27908 , n27910 );
xor ( n28438 , n28437 , n28418 );
xor ( n28439 , n28087 , n28089 );
xor ( n28440 , n28439 , n28415 );
xor ( n28441 , n28367 , n28369 );
xor ( n28442 , n28441 , n28412 );
xnor ( n28443 , n28250 , n28252 );
and ( n28444 , n25220 , n22784 );
and ( n28445 , n24993 , n22987 );
and ( n28446 , n28444 , n28445 );
xor ( n28447 , n28180 , n28181 );
xor ( n28448 , n28447 , n28183 );
and ( n28449 , n28445 , n28448 );
and ( n28450 , n28444 , n28448 );
or ( n28451 , n28446 , n28449 , n28450 );
and ( n28452 , n27389 , n21039 );
and ( n28453 , n28451 , n28452 );
xor ( n28454 , n28186 , n28187 );
xor ( n28455 , n28454 , n28189 );
and ( n28456 , n28452 , n28455 );
and ( n28457 , n28451 , n28455 );
or ( n28458 , n28453 , n28456 , n28457 );
xor ( n28459 , n27849 , n27850 );
xor ( n28460 , n28459 , n27852 );
and ( n28461 , n28458 , n28460 );
xor ( n28462 , n28179 , n28192 );
xor ( n28463 , n28462 , n28194 );
and ( n28464 , n28460 , n28463 );
and ( n28465 , n28458 , n28463 );
or ( n28466 , n28461 , n28464 , n28465 );
and ( n28467 , n28443 , n28466 );
xor ( n28468 , n28016 , n28017 );
xor ( n28469 , n28468 , n28019 );
xor ( n28470 , n28271 , n28272 );
xor ( n28471 , n28470 , n28274 );
or ( n28472 , n28469 , n28471 );
and ( n28473 , n28466 , n28472 );
and ( n28474 , n28443 , n28472 );
or ( n28475 , n28467 , n28473 , n28474 );
xor ( n28476 , n28114 , n28126 );
xor ( n28477 , n28476 , n28136 );
xor ( n28478 , n28147 , n28149 );
xor ( n28479 , n28478 , n28152 );
and ( n28480 , n28477 , n28479 );
xor ( n28481 , n28243 , n28244 );
xor ( n28482 , n28481 , n28247 );
and ( n28483 , n28479 , n28482 );
and ( n28484 , n28477 , n28482 );
or ( n28485 , n28480 , n28483 , n28484 );
and ( n28486 , n26399 , n21527 );
and ( n28487 , n26148 , n21666 );
and ( n28488 , n28486 , n28487 );
xor ( n28489 , n28265 , n28266 );
xor ( n28490 , n28489 , n28268 );
and ( n28491 , n28487 , n28490 );
and ( n28492 , n28486 , n28490 );
or ( n28493 , n28488 , n28491 , n28492 );
xor ( n28494 , n28236 , n28237 );
xor ( n28495 , n28494 , n28240 );
xor ( n28496 , n28280 , n28281 );
xor ( n28497 , n28496 , n28284 );
and ( n28498 , n28495 , n28497 );
and ( n28499 , n26399 , n21666 );
and ( n28500 , n25959 , n21990 );
and ( n28501 , n28499 , n28500 );
xor ( n28502 , n28301 , n28302 );
xor ( n28503 , n28502 , n28304 );
and ( n28504 , n28500 , n28503 );
and ( n28505 , n28499 , n28503 );
or ( n28506 , n28501 , n28504 , n28505 );
and ( n28507 , n28497 , n28506 );
and ( n28508 , n28495 , n28506 );
or ( n28509 , n28498 , n28507 , n28508 );
and ( n28510 , n28493 , n28509 );
and ( n28511 , n27591 , n21085 );
and ( n28512 , n27389 , n21178 );
and ( n28513 , n28511 , n28512 );
and ( n28514 , n26782 , n21527 );
and ( n28515 , n28512 , n28514 );
and ( n28516 , n28511 , n28514 );
or ( n28517 , n28513 , n28515 , n28516 );
and ( n28518 , n28124 , n28517 );
and ( n28519 , n23089 , n27558 );
and ( n28520 , n22936 , n28209 );
or ( n28521 , n28519 , n28520 );
and ( n28522 , n28517 , n28521 );
and ( n28523 , n28124 , n28521 );
or ( n28524 , n28518 , n28522 , n28523 );
buf ( n28525 , n22702 );
buf ( n28526 , n765 );
buf ( n28527 , n28526 );
buf ( n28528 , n766 );
buf ( n28529 , n28528 );
and ( n28530 , n28527 , n28529 );
not ( n28531 , n28530 );
and ( n28532 , n28121 , n28531 );
not ( n28533 , n28532 );
and ( n28534 , n28525 , n28533 );
and ( n28535 , n26678 , n21666 );
and ( n28536 , n26148 , n21990 );
and ( n28537 , n28535 , n28536 );
buf ( n28538 , n778 );
buf ( n28539 , n28538 );
buf ( n28540 , n28539 );
buf ( n28541 , n779 );
buf ( n28542 , n28541 );
and ( n28543 , n28539 , n28542 );
buf ( n28544 , n779 );
buf ( n28545 , n28544 );
buf ( n28546 , n778 );
buf ( n28547 , n28546 );
and ( n28548 , n28545 , n28547 );
and ( n28549 , n28543 , n28548 );
and ( n28550 , n28540 , n28549 );
xor ( n28551 , n28543 , n28548 );
buf ( n28552 , n780 );
buf ( n28553 , n28552 );
and ( n28554 , n28539 , n28553 );
buf ( n28555 , n780 );
buf ( n28556 , n28555 );
and ( n28557 , n28556 , n28547 );
and ( n28558 , n28554 , n28557 );
and ( n28559 , n28551 , n28558 );
buf ( n28560 , n28545 );
xor ( n28561 , n28554 , n28557 );
and ( n28562 , n28560 , n28561 );
buf ( n28563 , n781 );
buf ( n28564 , n28563 );
and ( n28565 , n28539 , n28564 );
buf ( n28566 , n781 );
buf ( n28567 , n28566 );
and ( n28568 , n28567 , n28547 );
and ( n28569 , n28565 , n28568 );
and ( n28570 , n28561 , n28569 );
and ( n28571 , n28560 , n28569 );
or ( n28572 , n28562 , n28570 , n28571 );
and ( n28573 , n28558 , n28572 );
and ( n28574 , n28551 , n28572 );
or ( n28575 , n28559 , n28573 , n28574 );
and ( n28576 , n28549 , n28575 );
and ( n28577 , n28540 , n28575 );
or ( n28578 , n28550 , n28576 , n28577 );
xor ( n28579 , n28540 , n28549 );
xor ( n28580 , n28579 , n28575 );
buf ( n28581 , n782 );
buf ( n28582 , n28581 );
and ( n28583 , n28582 , n28547 );
and ( n28584 , n28567 , n28542 );
or ( n28585 , n28583 , n28584 );
buf ( n28586 , n782 );
buf ( n28587 , n28586 );
and ( n28588 , n28539 , n28587 );
and ( n28589 , n28545 , n28564 );
or ( n28590 , n28588 , n28589 );
and ( n28591 , n28585 , n28590 );
and ( n28592 , n28556 , n28542 );
and ( n28593 , n28545 , n28553 );
and ( n28594 , n28592 , n28593 );
xor ( n28595 , n28565 , n28568 );
and ( n28596 , n28593 , n28595 );
and ( n28597 , n28592 , n28595 );
or ( n28598 , n28594 , n28596 , n28597 );
and ( n28599 , n28591 , n28598 );
xor ( n28600 , n28560 , n28561 );
xor ( n28601 , n28600 , n28569 );
and ( n28602 , n28598 , n28601 );
and ( n28603 , n28591 , n28601 );
or ( n28604 , n28599 , n28602 , n28603 );
xor ( n28605 , n28551 , n28558 );
xor ( n28606 , n28605 , n28572 );
and ( n28607 , n28604 , n28606 );
xor ( n28608 , n28585 , n28590 );
xnor ( n28609 , n28583 , n28584 );
xnor ( n28610 , n28588 , n28589 );
and ( n28611 , n28609 , n28610 );
and ( n28612 , n28608 , n28611 );
buf ( n28613 , n28556 );
buf ( n28614 , n783 );
buf ( n28615 , n28614 );
and ( n28616 , n28539 , n28615 );
buf ( n28617 , n783 );
buf ( n28618 , n28617 );
and ( n28619 , n28618 , n28547 );
and ( n28620 , n28616 , n28619 );
and ( n28621 , n28613 , n28620 );
and ( n28622 , n28545 , n28587 );
and ( n28623 , n28582 , n28542 );
and ( n28624 , n28622 , n28623 );
and ( n28625 , n28620 , n28624 );
and ( n28626 , n28613 , n28624 );
or ( n28627 , n28621 , n28625 , n28626 );
and ( n28628 , n28611 , n28627 );
and ( n28629 , n28608 , n28627 );
or ( n28630 , n28612 , n28628 , n28629 );
xor ( n28631 , n28591 , n28598 );
xor ( n28632 , n28631 , n28601 );
and ( n28633 , n28630 , n28632 );
xor ( n28634 , n28592 , n28593 );
xor ( n28635 , n28634 , n28595 );
and ( n28636 , n28556 , n28564 );
and ( n28637 , n28567 , n28553 );
and ( n28638 , n28636 , n28637 );
xor ( n28639 , n28609 , n28610 );
and ( n28640 , n28638 , n28639 );
buf ( n28641 , n784 );
buf ( n28642 , n28641 );
and ( n28643 , n28642 , n28547 );
and ( n28644 , n28618 , n28542 );
and ( n28645 , n28643 , n28644 );
and ( n28646 , n28582 , n28553 );
and ( n28647 , n28644 , n28646 );
and ( n28648 , n28643 , n28646 );
or ( n28649 , n28645 , n28647 , n28648 );
buf ( n28650 , n784 );
buf ( n28651 , n28650 );
and ( n28652 , n28539 , n28651 );
and ( n28653 , n28545 , n28615 );
and ( n28654 , n28652 , n28653 );
and ( n28655 , n28556 , n28587 );
and ( n28656 , n28653 , n28655 );
and ( n28657 , n28652 , n28655 );
or ( n28658 , n28654 , n28656 , n28657 );
and ( n28659 , n28649 , n28658 );
and ( n28660 , n28639 , n28659 );
and ( n28661 , n28638 , n28659 );
or ( n28662 , n28640 , n28660 , n28661 );
and ( n28663 , n28635 , n28662 );
xor ( n28664 , n28608 , n28611 );
xor ( n28665 , n28664 , n28627 );
and ( n28666 , n28662 , n28665 );
and ( n28667 , n28635 , n28665 );
or ( n28668 , n28663 , n28666 , n28667 );
and ( n28669 , n28632 , n28668 );
and ( n28670 , n28630 , n28668 );
or ( n28671 , n28633 , n28669 , n28670 );
and ( n28672 , n28606 , n28671 );
and ( n28673 , n28604 , n28671 );
or ( n28674 , n28607 , n28672 , n28673 );
and ( n28675 , n28580 , n28674 );
xor ( n28676 , n28604 , n28606 );
xor ( n28677 , n28676 , n28671 );
xor ( n28678 , n28630 , n28632 );
xor ( n28679 , n28678 , n28668 );
xor ( n28680 , n28616 , n28619 );
xor ( n28681 , n28622 , n28623 );
and ( n28682 , n28680 , n28681 );
xor ( n28683 , n28636 , n28637 );
and ( n28684 , n28681 , n28683 );
and ( n28685 , n28680 , n28683 );
or ( n28686 , n28682 , n28684 , n28685 );
xor ( n28687 , n28613 , n28620 );
xor ( n28688 , n28687 , n28624 );
and ( n28689 , n28686 , n28688 );
xor ( n28690 , n28649 , n28658 );
xor ( n28691 , n28643 , n28644 );
xor ( n28692 , n28691 , n28646 );
xor ( n28693 , n28652 , n28653 );
xor ( n28694 , n28693 , n28655 );
and ( n28695 , n28692 , n28694 );
and ( n28696 , n28690 , n28695 );
xor ( n28697 , n28680 , n28681 );
xor ( n28698 , n28697 , n28683 );
and ( n28699 , n28695 , n28698 );
and ( n28700 , n28690 , n28698 );
or ( n28701 , n28696 , n28699 , n28700 );
and ( n28702 , n28688 , n28701 );
and ( n28703 , n28686 , n28701 );
or ( n28704 , n28689 , n28702 , n28703 );
xor ( n28705 , n28635 , n28662 );
xor ( n28706 , n28705 , n28665 );
and ( n28707 , n28704 , n28706 );
xor ( n28708 , n28638 , n28639 );
xor ( n28709 , n28708 , n28659 );
buf ( n28710 , n786 );
buf ( n28711 , n28710 );
and ( n28712 , n28539 , n28711 );
and ( n28713 , n28556 , n28651 );
and ( n28714 , n28712 , n28713 );
and ( n28715 , n28567 , n28615 );
and ( n28716 , n28713 , n28715 );
and ( n28717 , n28712 , n28715 );
or ( n28718 , n28714 , n28716 , n28717 );
buf ( n28719 , n785 );
buf ( n28720 , n28719 );
and ( n28721 , n28720 , n28547 );
and ( n28722 , n28718 , n28721 );
and ( n28723 , n28618 , n28553 );
and ( n28724 , n28721 , n28723 );
and ( n28725 , n28718 , n28723 );
or ( n28726 , n28722 , n28724 , n28725 );
buf ( n28727 , n786 );
buf ( n28728 , n28727 );
and ( n28729 , n28728 , n28547 );
and ( n28730 , n28642 , n28553 );
and ( n28731 , n28729 , n28730 );
and ( n28732 , n28618 , n28564 );
and ( n28733 , n28730 , n28732 );
and ( n28734 , n28729 , n28732 );
or ( n28735 , n28731 , n28733 , n28734 );
buf ( n28736 , n785 );
buf ( n28737 , n28736 );
and ( n28738 , n28539 , n28737 );
and ( n28739 , n28735 , n28738 );
and ( n28740 , n28556 , n28615 );
and ( n28741 , n28738 , n28740 );
and ( n28742 , n28735 , n28740 );
or ( n28743 , n28739 , n28741 , n28742 );
and ( n28744 , n28726 , n28743 );
buf ( n28745 , n28567 );
and ( n28746 , n28545 , n28651 );
and ( n28747 , n28642 , n28542 );
and ( n28748 , n28746 , n28747 );
and ( n28749 , n28745 , n28748 );
xor ( n28750 , n28692 , n28694 );
and ( n28751 , n28748 , n28750 );
and ( n28752 , n28745 , n28750 );
or ( n28753 , n28749 , n28751 , n28752 );
and ( n28754 , n28744 , n28753 );
xor ( n28755 , n28690 , n28695 );
xor ( n28756 , n28755 , n28698 );
and ( n28757 , n28753 , n28756 );
and ( n28758 , n28744 , n28756 );
or ( n28759 , n28754 , n28757 , n28758 );
and ( n28760 , n28709 , n28759 );
xor ( n28761 , n28686 , n28688 );
xor ( n28762 , n28761 , n28701 );
and ( n28763 , n28759 , n28762 );
and ( n28764 , n28709 , n28762 );
or ( n28765 , n28760 , n28763 , n28764 );
and ( n28766 , n28706 , n28765 );
and ( n28767 , n28704 , n28765 );
or ( n28768 , n28707 , n28766 , n28767 );
and ( n28769 , n28679 , n28768 );
xor ( n28770 , n28704 , n28706 );
xor ( n28771 , n28770 , n28765 );
xor ( n28772 , n28709 , n28759 );
xor ( n28773 , n28772 , n28762 );
and ( n28774 , n28582 , n28564 );
and ( n28775 , n28567 , n28587 );
and ( n28776 , n28774 , n28775 );
xor ( n28777 , n28746 , n28747 );
and ( n28778 , n28775 , n28777 );
and ( n28779 , n28774 , n28777 );
or ( n28780 , n28776 , n28778 , n28779 );
xor ( n28781 , n28726 , n28743 );
and ( n28782 , n28780 , n28781 );
xor ( n28783 , n28718 , n28721 );
xor ( n28784 , n28783 , n28723 );
xor ( n28785 , n28735 , n28738 );
xor ( n28786 , n28785 , n28740 );
and ( n28787 , n28784 , n28786 );
and ( n28788 , n28781 , n28787 );
and ( n28789 , n28780 , n28787 );
or ( n28790 , n28782 , n28788 , n28789 );
xor ( n28791 , n28744 , n28753 );
xor ( n28792 , n28791 , n28756 );
and ( n28793 , n28790 , n28792 );
and ( n28794 , n28545 , n28737 );
and ( n28795 , n28720 , n28542 );
and ( n28796 , n28794 , n28795 );
and ( n28797 , n28728 , n28542 );
and ( n28798 , n28642 , n28564 );
or ( n28799 , n28797 , n28798 );
and ( n28800 , n28545 , n28711 );
and ( n28801 , n28567 , n28651 );
or ( n28802 , n28800 , n28801 );
and ( n28803 , n28799 , n28802 );
and ( n28804 , n28796 , n28803 );
xor ( n28805 , n28729 , n28730 );
xor ( n28806 , n28805 , n28732 );
xor ( n28807 , n28712 , n28713 );
xor ( n28808 , n28807 , n28715 );
and ( n28809 , n28806 , n28808 );
and ( n28810 , n28803 , n28809 );
and ( n28811 , n28796 , n28809 );
or ( n28812 , n28804 , n28810 , n28811 );
xor ( n28813 , n28745 , n28748 );
xor ( n28814 , n28813 , n28750 );
and ( n28815 , n28812 , n28814 );
buf ( n28816 , n28582 );
xor ( n28817 , n28794 , n28795 );
and ( n28818 , n28816 , n28817 );
and ( n28819 , n28556 , n28737 );
and ( n28820 , n28720 , n28553 );
and ( n28821 , n28819 , n28820 );
and ( n28822 , n28817 , n28821 );
and ( n28823 , n28816 , n28821 );
or ( n28824 , n28818 , n28822 , n28823 );
xor ( n28825 , n28774 , n28775 );
xor ( n28826 , n28825 , n28777 );
and ( n28827 , n28824 , n28826 );
xor ( n28828 , n28784 , n28786 );
and ( n28829 , n28826 , n28828 );
and ( n28830 , n28824 , n28828 );
or ( n28831 , n28827 , n28829 , n28830 );
and ( n28832 , n28814 , n28831 );
and ( n28833 , n28812 , n28831 );
or ( n28834 , n28815 , n28832 , n28833 );
and ( n28835 , n28792 , n28834 );
and ( n28836 , n28790 , n28834 );
or ( n28837 , n28793 , n28835 , n28836 );
and ( n28838 , n28773 , n28837 );
buf ( n28839 , n787 );
buf ( n28840 , n28839 );
and ( n28841 , n28840 , n28547 );
not ( n28842 , n28841 );
xnor ( n28843 , n28800 , n28801 );
and ( n28844 , n28842 , n28843 );
buf ( n28845 , n787 );
buf ( n28846 , n28845 );
and ( n28847 , n28539 , n28846 );
not ( n28848 , n28847 );
xnor ( n28849 , n28797 , n28798 );
and ( n28850 , n28848 , n28849 );
and ( n28851 , n28844 , n28850 );
buf ( n28852 , n28841 );
buf ( n28853 , n28847 );
and ( n28854 , n28852 , n28853 );
and ( n28855 , n28851 , n28854 );
xor ( n28856 , n28799 , n28802 );
xor ( n28857 , n28806 , n28808 );
and ( n28858 , n28856 , n28857 );
and ( n28859 , n28840 , n28542 );
and ( n28860 , n28720 , n28564 );
and ( n28861 , n28859 , n28860 );
and ( n28862 , n28642 , n28587 );
and ( n28863 , n28860 , n28862 );
and ( n28864 , n28859 , n28862 );
or ( n28865 , n28861 , n28863 , n28864 );
and ( n28866 , n28545 , n28846 );
and ( n28867 , n28567 , n28737 );
and ( n28868 , n28866 , n28867 );
and ( n28869 , n28582 , n28651 );
and ( n28870 , n28867 , n28869 );
and ( n28871 , n28866 , n28869 );
or ( n28872 , n28868 , n28870 , n28871 );
and ( n28873 , n28865 , n28872 );
and ( n28874 , n28857 , n28873 );
and ( n28875 , n28856 , n28873 );
or ( n28876 , n28858 , n28874 , n28875 );
and ( n28877 , n28854 , n28876 );
and ( n28878 , n28851 , n28876 );
or ( n28879 , n28855 , n28877 , n28878 );
xor ( n28880 , n28780 , n28781 );
xor ( n28881 , n28880 , n28787 );
and ( n28882 , n28879 , n28881 );
xor ( n28883 , n28796 , n28803 );
xor ( n28884 , n28883 , n28809 );
and ( n28885 , n28618 , n28587 );
and ( n28886 , n28582 , n28615 );
and ( n28887 , n28885 , n28886 );
xor ( n28888 , n28819 , n28820 );
and ( n28889 , n28886 , n28888 );
and ( n28890 , n28885 , n28888 );
or ( n28891 , n28887 , n28889 , n28890 );
xor ( n28892 , n28816 , n28817 );
xor ( n28893 , n28892 , n28821 );
and ( n28894 , n28891 , n28893 );
xor ( n28895 , n28844 , n28850 );
and ( n28896 , n28893 , n28895 );
and ( n28897 , n28891 , n28895 );
or ( n28898 , n28894 , n28896 , n28897 );
and ( n28899 , n28884 , n28898 );
xor ( n28900 , n28852 , n28853 );
buf ( n28901 , n788 );
buf ( n28902 , n28901 );
and ( n28903 , n28545 , n28902 );
and ( n28904 , n28556 , n28846 );
and ( n28905 , n28903 , n28904 );
and ( n28906 , n28582 , n28737 );
and ( n28907 , n28904 , n28906 );
and ( n28908 , n28903 , n28906 );
or ( n28909 , n28905 , n28907 , n28908 );
buf ( n28910 , n788 );
buf ( n28911 , n28910 );
and ( n28912 , n28911 , n28547 );
and ( n28913 , n28909 , n28912 );
and ( n28914 , n28728 , n28553 );
and ( n28915 , n28912 , n28914 );
and ( n28916 , n28909 , n28914 );
or ( n28917 , n28913 , n28915 , n28916 );
and ( n28918 , n28911 , n28542 );
and ( n28919 , n28840 , n28553 );
and ( n28920 , n28918 , n28919 );
and ( n28921 , n28720 , n28587 );
and ( n28922 , n28919 , n28921 );
and ( n28923 , n28918 , n28921 );
or ( n28924 , n28920 , n28922 , n28923 );
and ( n28925 , n28539 , n28902 );
and ( n28926 , n28924 , n28925 );
and ( n28927 , n28556 , n28711 );
and ( n28928 , n28925 , n28927 );
and ( n28929 , n28924 , n28927 );
or ( n28930 , n28926 , n28928 , n28929 );
and ( n28931 , n28917 , n28930 );
and ( n28932 , n28900 , n28931 );
xor ( n28933 , n28842 , n28843 );
xor ( n28934 , n28848 , n28849 );
and ( n28935 , n28933 , n28934 );
and ( n28936 , n28931 , n28935 );
and ( n28937 , n28900 , n28935 );
or ( n28938 , n28932 , n28936 , n28937 );
and ( n28939 , n28898 , n28938 );
and ( n28940 , n28884 , n28938 );
or ( n28941 , n28899 , n28939 , n28940 );
and ( n28942 , n28881 , n28941 );
and ( n28943 , n28879 , n28941 );
or ( n28944 , n28882 , n28942 , n28943 );
xor ( n28945 , n28790 , n28792 );
xor ( n28946 , n28945 , n28834 );
and ( n28947 , n28944 , n28946 );
xor ( n28948 , n28812 , n28814 );
xor ( n28949 , n28948 , n28831 );
xor ( n28950 , n28824 , n28826 );
xor ( n28951 , n28950 , n28828 );
xor ( n28952 , n28851 , n28854 );
xor ( n28953 , n28952 , n28876 );
and ( n28954 , n28951 , n28953 );
xor ( n28955 , n28865 , n28872 );
xor ( n28956 , n28859 , n28860 );
xor ( n28957 , n28956 , n28862 );
xor ( n28958 , n28866 , n28867 );
xor ( n28959 , n28958 , n28869 );
and ( n28960 , n28957 , n28959 );
and ( n28961 , n28955 , n28960 );
buf ( n28962 , n28618 );
buf ( n28963 , n789 );
buf ( n28964 , n28963 );
and ( n28965 , n28539 , n28964 );
buf ( n28966 , n789 );
buf ( n28967 , n28966 );
and ( n28968 , n28967 , n28547 );
and ( n28969 , n28965 , n28968 );
and ( n28970 , n28962 , n28969 );
and ( n28971 , n28567 , n28711 );
and ( n28972 , n28728 , n28564 );
and ( n28973 , n28971 , n28972 );
and ( n28974 , n28969 , n28973 );
and ( n28975 , n28962 , n28973 );
or ( n28976 , n28970 , n28974 , n28975 );
and ( n28977 , n28960 , n28976 );
and ( n28978 , n28955 , n28976 );
or ( n28979 , n28961 , n28977 , n28978 );
xor ( n28980 , n28856 , n28857 );
xor ( n28981 , n28980 , n28873 );
and ( n28982 , n28979 , n28981 );
xor ( n28983 , n28885 , n28886 );
xor ( n28984 , n28983 , n28888 );
xor ( n28985 , n28917 , n28930 );
and ( n28986 , n28984 , n28985 );
xor ( n28987 , n28933 , n28934 );
and ( n28988 , n28985 , n28987 );
and ( n28989 , n28984 , n28987 );
or ( n28990 , n28986 , n28988 , n28989 );
and ( n28991 , n28981 , n28990 );
and ( n28992 , n28979 , n28990 );
or ( n28993 , n28982 , n28991 , n28992 );
and ( n28994 , n28953 , n28993 );
and ( n28995 , n28951 , n28993 );
or ( n28996 , n28954 , n28994 , n28995 );
and ( n28997 , n28949 , n28996 );
xor ( n28998 , n28879 , n28881 );
xor ( n28999 , n28998 , n28941 );
and ( n29000 , n28996 , n28999 );
and ( n29001 , n28949 , n28999 );
or ( n29002 , n28997 , n29000 , n29001 );
and ( n29003 , n28946 , n29002 );
and ( n29004 , n28944 , n29002 );
or ( n29005 , n28947 , n29003 , n29004 );
and ( n29006 , n28837 , n29005 );
and ( n29007 , n28773 , n29005 );
or ( n29008 , n28838 , n29006 , n29007 );
and ( n29009 , n28771 , n29008 );
xor ( n29010 , n28773 , n28837 );
xor ( n29011 , n29010 , n29005 );
xor ( n29012 , n28944 , n28946 );
xor ( n29013 , n29012 , n29002 );
xor ( n29014 , n28909 , n28912 );
xor ( n29015 , n29014 , n28914 );
xor ( n29016 , n28924 , n28925 );
xor ( n29017 , n29016 , n28927 );
and ( n29018 , n29015 , n29017 );
and ( n29019 , n28618 , n28651 );
and ( n29020 , n28642 , n28615 );
and ( n29021 , n29019 , n29020 );
xor ( n29022 , n28957 , n28959 );
and ( n29023 , n29021 , n29022 );
and ( n29024 , n28911 , n28553 );
and ( n29025 , n28728 , n28587 );
or ( n29026 , n29024 , n29025 );
and ( n29027 , n28556 , n28902 );
and ( n29028 , n28582 , n28711 );
or ( n29029 , n29027 , n29028 );
and ( n29030 , n29026 , n29029 );
and ( n29031 , n29022 , n29030 );
and ( n29032 , n29021 , n29030 );
or ( n29033 , n29023 , n29031 , n29032 );
and ( n29034 , n29018 , n29033 );
and ( n29035 , n28967 , n28542 );
and ( n29036 , n28840 , n28564 );
or ( n29037 , n29035 , n29036 );
and ( n29038 , n28545 , n28964 );
and ( n29039 , n28567 , n28846 );
or ( n29040 , n29038 , n29039 );
and ( n29041 , n29037 , n29040 );
xor ( n29042 , n28918 , n28919 );
xor ( n29043 , n29042 , n28921 );
xor ( n29044 , n28903 , n28904 );
xor ( n29045 , n29044 , n28906 );
and ( n29046 , n29043 , n29045 );
and ( n29047 , n29041 , n29046 );
xor ( n29048 , n28965 , n28968 );
xor ( n29049 , n28971 , n28972 );
and ( n29050 , n29048 , n29049 );
xor ( n29051 , n29019 , n29020 );
and ( n29052 , n29049 , n29051 );
and ( n29053 , n29048 , n29051 );
or ( n29054 , n29050 , n29052 , n29053 );
and ( n29055 , n29046 , n29054 );
and ( n29056 , n29041 , n29054 );
or ( n29057 , n29047 , n29055 , n29056 );
and ( n29058 , n29033 , n29057 );
and ( n29059 , n29018 , n29057 );
or ( n29060 , n29034 , n29058 , n29059 );
xor ( n29061 , n28891 , n28893 );
xor ( n29062 , n29061 , n28895 );
and ( n29063 , n29060 , n29062 );
xor ( n29064 , n28900 , n28931 );
xor ( n29065 , n29064 , n28935 );
and ( n29066 , n29062 , n29065 );
and ( n29067 , n29060 , n29065 );
or ( n29068 , n29063 , n29066 , n29067 );
xor ( n29069 , n28884 , n28898 );
xor ( n29070 , n29069 , n28938 );
and ( n29071 , n29068 , n29070 );
xor ( n29072 , n28955 , n28960 );
xor ( n29073 , n29072 , n28976 );
xor ( n29074 , n28962 , n28969 );
xor ( n29075 , n29074 , n28973 );
xor ( n29076 , n29015 , n29017 );
and ( n29077 , n29075 , n29076 );
and ( n29078 , n28720 , n28615 );
xnor ( n29079 , n29027 , n29028 );
or ( n29080 , n29078 , n29079 );
and ( n29081 , n28618 , n28737 );
xnor ( n29082 , n29024 , n29025 );
or ( n29083 , n29081 , n29082 );
and ( n29084 , n29080 , n29083 );
and ( n29085 , n29076 , n29084 );
and ( n29086 , n29075 , n29084 );
or ( n29087 , n29077 , n29085 , n29086 );
and ( n29088 , n29073 , n29087 );
buf ( n29089 , n790 );
buf ( n29090 , n29089 );
and ( n29091 , n29090 , n28547 );
xnor ( n29092 , n29038 , n29039 );
or ( n29093 , n29091 , n29092 );
buf ( n29094 , n790 );
buf ( n29095 , n29094 );
and ( n29096 , n28539 , n29095 );
xnor ( n29097 , n29035 , n29036 );
or ( n29098 , n29096 , n29097 );
and ( n29099 , n29093 , n29098 );
xor ( n29100 , n29026 , n29029 );
xor ( n29101 , n29037 , n29040 );
and ( n29102 , n29100 , n29101 );
xor ( n29103 , n29043 , n29045 );
and ( n29104 , n29101 , n29103 );
and ( n29105 , n29100 , n29103 );
or ( n29106 , n29102 , n29104 , n29105 );
and ( n29107 , n29099 , n29106 );
buf ( n29108 , n791 );
buf ( n29109 , n29108 );
and ( n29110 , n29109 , n28547 );
and ( n29111 , n28911 , n28564 );
and ( n29112 , n29110 , n29111 );
and ( n29113 , n28728 , n28615 );
and ( n29114 , n29111 , n29113 );
and ( n29115 , n29110 , n29113 );
or ( n29116 , n29112 , n29114 , n29115 );
buf ( n29117 , n791 );
buf ( n29118 , n29117 );
and ( n29119 , n28539 , n29118 );
and ( n29120 , n28567 , n28902 );
and ( n29121 , n29119 , n29120 );
and ( n29122 , n28618 , n28711 );
and ( n29123 , n29120 , n29122 );
and ( n29124 , n29119 , n29122 );
or ( n29125 , n29121 , n29123 , n29124 );
and ( n29126 , n29116 , n29125 );
and ( n29127 , n29090 , n28542 );
and ( n29128 , n28967 , n28553 );
or ( n29129 , n29127 , n29128 );
and ( n29130 , n28545 , n29095 );
and ( n29131 , n28556 , n28964 );
or ( n29132 , n29130 , n29131 );
and ( n29133 , n29129 , n29132 );
and ( n29134 , n29126 , n29133 );
xor ( n29135 , n29048 , n29049 );
xor ( n29136 , n29135 , n29051 );
and ( n29137 , n29133 , n29136 );
and ( n29138 , n29126 , n29136 );
or ( n29139 , n29134 , n29137 , n29138 );
and ( n29140 , n29106 , n29139 );
and ( n29141 , n29099 , n29139 );
or ( n29142 , n29107 , n29140 , n29141 );
and ( n29143 , n29087 , n29142 );
and ( n29144 , n29073 , n29142 );
or ( n29145 , n29088 , n29143 , n29144 );
xor ( n29146 , n28979 , n28981 );
xor ( n29147 , n29146 , n28990 );
and ( n29148 , n29145 , n29147 );
xor ( n29149 , n29060 , n29062 );
xor ( n29150 , n29149 , n29065 );
and ( n29151 , n29147 , n29150 );
and ( n29152 , n29145 , n29150 );
or ( n29153 , n29148 , n29151 , n29152 );
and ( n29154 , n29070 , n29153 );
and ( n29155 , n29068 , n29153 );
or ( n29156 , n29071 , n29154 , n29155 );
xor ( n29157 , n28949 , n28996 );
xor ( n29158 , n29157 , n28999 );
and ( n29159 , n29156 , n29158 );
xor ( n29160 , n28951 , n28953 );
xor ( n29161 , n29160 , n28993 );
xor ( n29162 , n29068 , n29070 );
xor ( n29163 , n29162 , n29153 );
and ( n29164 , n29161 , n29163 );
xor ( n29165 , n28984 , n28985 );
xor ( n29166 , n29165 , n28987 );
xor ( n29167 , n29018 , n29033 );
xor ( n29168 , n29167 , n29057 );
and ( n29169 , n29166 , n29168 );
xor ( n29170 , n29021 , n29022 );
xor ( n29171 , n29170 , n29030 );
xor ( n29172 , n29041 , n29046 );
xor ( n29173 , n29172 , n29054 );
and ( n29174 , n29171 , n29173 );
xor ( n29175 , n29080 , n29083 );
xor ( n29176 , n29093 , n29098 );
and ( n29177 , n29175 , n29176 );
xnor ( n29178 , n29078 , n29079 );
xnor ( n29179 , n29081 , n29082 );
and ( n29180 , n29178 , n29179 );
and ( n29181 , n29176 , n29180 );
and ( n29182 , n29175 , n29180 );
or ( n29183 , n29177 , n29181 , n29182 );
and ( n29184 , n29173 , n29183 );
and ( n29185 , n29171 , n29183 );
or ( n29186 , n29174 , n29184 , n29185 );
and ( n29187 , n29168 , n29186 );
and ( n29188 , n29166 , n29186 );
or ( n29189 , n29169 , n29187 , n29188 );
xor ( n29190 , n29145 , n29147 );
xor ( n29191 , n29190 , n29150 );
and ( n29192 , n29189 , n29191 );
xnor ( n29193 , n29091 , n29092 );
xnor ( n29194 , n29096 , n29097 );
and ( n29195 , n29193 , n29194 );
buf ( n29196 , n28642 );
and ( n29197 , n28582 , n28846 );
and ( n29198 , n28840 , n28587 );
and ( n29199 , n29197 , n29198 );
and ( n29200 , n29196 , n29199 );
xor ( n29201 , n29116 , n29125 );
and ( n29202 , n29199 , n29201 );
and ( n29203 , n29196 , n29201 );
or ( n29204 , n29200 , n29202 , n29203 );
and ( n29205 , n29195 , n29204 );
xor ( n29206 , n29129 , n29132 );
and ( n29207 , n28840 , n28615 );
and ( n29208 , n28728 , n28651 );
or ( n29209 , n29207 , n29208 );
and ( n29210 , n28618 , n28846 );
and ( n29211 , n28642 , n28711 );
or ( n29212 , n29210 , n29211 );
and ( n29213 , n29209 , n29212 );
and ( n29214 , n29206 , n29213 );
xor ( n29215 , n29110 , n29111 );
xor ( n29216 , n29215 , n29113 );
xor ( n29217 , n29119 , n29120 );
xor ( n29218 , n29217 , n29122 );
and ( n29219 , n29216 , n29218 );
and ( n29220 , n29213 , n29219 );
and ( n29221 , n29206 , n29219 );
or ( n29222 , n29214 , n29220 , n29221 );
and ( n29223 , n29204 , n29222 );
and ( n29224 , n29195 , n29222 );
or ( n29225 , n29205 , n29223 , n29224 );
xnor ( n29226 , n29127 , n29128 );
xnor ( n29227 , n29130 , n29131 );
and ( n29228 , n29226 , n29227 );
and ( n29229 , n28720 , n28651 );
and ( n29230 , n28642 , n28737 );
and ( n29231 , n29229 , n29230 );
xor ( n29232 , n29197 , n29198 );
and ( n29233 , n29230 , n29232 );
and ( n29234 , n29229 , n29232 );
or ( n29235 , n29231 , n29233 , n29234 );
and ( n29236 , n29228 , n29235 );
and ( n29237 , n28545 , n29118 );
and ( n29238 , n29109 , n28542 );
and ( n29239 , n29237 , n29238 );
and ( n29240 , n28556 , n29095 );
and ( n29241 , n29090 , n28553 );
and ( n29242 , n29240 , n29241 );
and ( n29243 , n29239 , n29242 );
and ( n29244 , n28567 , n28964 );
and ( n29245 , n28967 , n28564 );
and ( n29246 , n29244 , n29245 );
and ( n29247 , n29242 , n29246 );
and ( n29248 , n29239 , n29246 );
or ( n29249 , n29243 , n29247 , n29248 );
and ( n29250 , n29235 , n29249 );
and ( n29251 , n29228 , n29249 );
or ( n29252 , n29236 , n29250 , n29251 );
xor ( n29253 , n29100 , n29101 );
xor ( n29254 , n29253 , n29103 );
and ( n29255 , n29252 , n29254 );
xor ( n29256 , n29126 , n29133 );
xor ( n29257 , n29256 , n29136 );
and ( n29258 , n29254 , n29257 );
and ( n29259 , n29252 , n29257 );
or ( n29260 , n29255 , n29258 , n29259 );
and ( n29261 , n29225 , n29260 );
xor ( n29262 , n29075 , n29076 );
xor ( n29263 , n29262 , n29084 );
and ( n29264 , n29260 , n29263 );
and ( n29265 , n29225 , n29263 );
or ( n29266 , n29261 , n29264 , n29265 );
xor ( n29267 , n29073 , n29087 );
xor ( n29268 , n29267 , n29142 );
and ( n29269 , n29266 , n29268 );
xor ( n29270 , n29099 , n29106 );
xor ( n29271 , n29270 , n29139 );
xor ( n29272 , n29178 , n29179 );
xor ( n29273 , n29193 , n29194 );
and ( n29274 , n29272 , n29273 );
and ( n29275 , n28582 , n28902 );
and ( n29276 , n28911 , n28587 );
and ( n29277 , n29275 , n29276 );
xor ( n29278 , n29209 , n29212 );
and ( n29279 , n29277 , n29278 );
xor ( n29280 , n29216 , n29218 );
and ( n29281 , n29278 , n29280 );
and ( n29282 , n29277 , n29280 );
or ( n29283 , n29279 , n29281 , n29282 );
and ( n29284 , n29273 , n29283 );
and ( n29285 , n29272 , n29283 );
or ( n29286 , n29274 , n29284 , n29285 );
xor ( n29287 , n29226 , n29227 );
buf ( n29288 , n793 );
buf ( n29289 , n29288 );
and ( n29290 , n29289 , n28547 );
buf ( n29291 , n792 );
buf ( n29292 , n29291 );
and ( n29293 , n29292 , n28542 );
and ( n29294 , n29290 , n29293 );
and ( n29295 , n28911 , n28615 );
and ( n29296 , n29293 , n29295 );
and ( n29297 , n29290 , n29295 );
or ( n29298 , n29294 , n29296 , n29297 );
and ( n29299 , n28720 , n28711 );
and ( n29300 , n28728 , n28737 );
and ( n29301 , n29299 , n29300 );
and ( n29302 , n29298 , n29301 );
buf ( n29303 , n792 );
buf ( n29304 , n29303 );
and ( n29305 , n28539 , n29304 );
and ( n29306 , n29301 , n29305 );
and ( n29307 , n29298 , n29305 );
or ( n29308 , n29302 , n29306 , n29307 );
and ( n29309 , n29287 , n29308 );
xnor ( n29310 , n29207 , n29208 );
xnor ( n29311 , n29210 , n29211 );
and ( n29312 , n29310 , n29311 );
and ( n29313 , n29308 , n29312 );
and ( n29314 , n29287 , n29312 );
or ( n29315 , n29309 , n29313 , n29314 );
and ( n29316 , n29292 , n28547 );
buf ( n29317 , n28720 );
and ( n29318 , n29316 , n29317 );
xor ( n29319 , n29237 , n29238 );
and ( n29320 , n29317 , n29319 );
and ( n29321 , n29316 , n29319 );
or ( n29322 , n29318 , n29320 , n29321 );
xor ( n29323 , n29240 , n29241 );
xor ( n29324 , n29244 , n29245 );
and ( n29325 , n29323 , n29324 );
xor ( n29326 , n29275 , n29276 );
and ( n29327 , n29324 , n29326 );
and ( n29328 , n29323 , n29326 );
or ( n29329 , n29325 , n29327 , n29328 );
and ( n29330 , n29322 , n29329 );
buf ( n29331 , n793 );
buf ( n29332 , n29331 );
and ( n29333 , n28539 , n29332 );
and ( n29334 , n28545 , n29304 );
and ( n29335 , n29333 , n29334 );
and ( n29336 , n28618 , n28902 );
and ( n29337 , n29334 , n29336 );
and ( n29338 , n29333 , n29336 );
or ( n29339 , n29335 , n29337 , n29338 );
and ( n29340 , n28556 , n29118 );
and ( n29341 , n29109 , n28553 );
and ( n29342 , n29340 , n29341 );
and ( n29343 , n29339 , n29342 );
and ( n29344 , n28567 , n29095 );
and ( n29345 , n29090 , n28564 );
and ( n29346 , n29344 , n29345 );
and ( n29347 , n29342 , n29346 );
and ( n29348 , n29339 , n29346 );
or ( n29349 , n29343 , n29347 , n29348 );
and ( n29350 , n29329 , n29349 );
and ( n29351 , n29322 , n29349 );
or ( n29352 , n29330 , n29350 , n29351 );
and ( n29353 , n29315 , n29352 );
xor ( n29354 , n29196 , n29199 );
xor ( n29355 , n29354 , n29201 );
and ( n29356 , n29352 , n29355 );
and ( n29357 , n29315 , n29355 );
or ( n29358 , n29353 , n29356 , n29357 );
and ( n29359 , n29286 , n29358 );
xor ( n29360 , n29175 , n29176 );
xor ( n29361 , n29360 , n29180 );
and ( n29362 , n29358 , n29361 );
and ( n29363 , n29286 , n29361 );
or ( n29364 , n29359 , n29362 , n29363 );
and ( n29365 , n29271 , n29364 );
xor ( n29366 , n29171 , n29173 );
xor ( n29367 , n29366 , n29183 );
and ( n29368 , n29364 , n29367 );
and ( n29369 , n29271 , n29367 );
or ( n29370 , n29365 , n29368 , n29369 );
and ( n29371 , n29268 , n29370 );
and ( n29372 , n29266 , n29370 );
or ( n29373 , n29269 , n29371 , n29372 );
and ( n29374 , n29191 , n29373 );
and ( n29375 , n29189 , n29373 );
or ( n29376 , n29192 , n29374 , n29375 );
and ( n29377 , n29163 , n29376 );
and ( n29378 , n29161 , n29376 );
or ( n29379 , n29164 , n29377 , n29378 );
and ( n29380 , n29158 , n29379 );
and ( n29381 , n29156 , n29379 );
or ( n29382 , n29159 , n29380 , n29381 );
or ( n29383 , n29013 , n29382 );
or ( n29384 , n29011 , n29383 );
and ( n29385 , n29008 , n29384 );
and ( n29386 , n28771 , n29384 );
or ( n29387 , n29009 , n29385 , n29386 );
and ( n29388 , n28768 , n29387 );
and ( n29389 , n28679 , n29387 );
or ( n29390 , n28769 , n29388 , n29389 );
or ( n29391 , n28677 , n29390 );
and ( n29392 , n28674 , n29391 );
and ( n29393 , n28580 , n29391 );
or ( n29394 , n28675 , n29392 , n29393 );
xnor ( n29395 , n28578 , n29394 );
xor ( n29396 , n28580 , n28674 );
xor ( n29397 , n29396 , n29391 );
not ( n29398 , n29397 );
xnor ( n29399 , n28677 , n29390 );
xor ( n29400 , n28679 , n28768 );
xor ( n29401 , n29400 , n29387 );
not ( n29402 , n29401 );
xor ( n29403 , n28771 , n29008 );
xor ( n29404 , n29403 , n29384 );
xnor ( n29405 , n29011 , n29383 );
xnor ( n29406 , n29013 , n29382 );
xor ( n29407 , n29156 , n29158 );
xor ( n29408 , n29407 , n29379 );
not ( n29409 , n29408 );
xor ( n29410 , n29161 , n29163 );
xor ( n29411 , n29410 , n29376 );
xor ( n29412 , n29166 , n29168 );
xor ( n29413 , n29412 , n29186 );
xor ( n29414 , n29225 , n29260 );
xor ( n29415 , n29414 , n29263 );
xor ( n29416 , n29195 , n29204 );
xor ( n29417 , n29416 , n29222 );
xor ( n29418 , n29252 , n29254 );
xor ( n29419 , n29418 , n29257 );
and ( n29420 , n29417 , n29419 );
xor ( n29421 , n29206 , n29213 );
xor ( n29422 , n29421 , n29219 );
xor ( n29423 , n29228 , n29235 );
xor ( n29424 , n29423 , n29249 );
and ( n29425 , n29422 , n29424 );
xor ( n29426 , n29229 , n29230 );
xor ( n29427 , n29426 , n29232 );
xor ( n29428 , n29239 , n29242 );
xor ( n29429 , n29428 , n29246 );
and ( n29430 , n29427 , n29429 );
and ( n29431 , n28582 , n28964 );
and ( n29432 , n28967 , n28587 );
and ( n29433 , n29431 , n29432 );
and ( n29434 , n28642 , n28846 );
and ( n29435 , n28840 , n28651 );
and ( n29436 , n29434 , n29435 );
and ( n29437 , n29433 , n29436 );
xor ( n29438 , n29298 , n29301 );
xor ( n29439 , n29438 , n29305 );
and ( n29440 , n29436 , n29439 );
and ( n29441 , n29433 , n29439 );
or ( n29442 , n29437 , n29440 , n29441 );
and ( n29443 , n29429 , n29442 );
and ( n29444 , n29427 , n29442 );
or ( n29445 , n29430 , n29443 , n29444 );
and ( n29446 , n29424 , n29445 );
and ( n29447 , n29422 , n29445 );
or ( n29448 , n29425 , n29446 , n29447 );
and ( n29449 , n29419 , n29448 );
and ( n29450 , n29417 , n29448 );
or ( n29451 , n29420 , n29449 , n29450 );
and ( n29452 , n29415 , n29451 );
xor ( n29453 , n29271 , n29364 );
xor ( n29454 , n29453 , n29367 );
and ( n29455 , n29451 , n29454 );
and ( n29456 , n29415 , n29454 );
or ( n29457 , n29452 , n29455 , n29456 );
and ( n29458 , n29413 , n29457 );
xor ( n29459 , n29266 , n29268 );
xor ( n29460 , n29459 , n29370 );
and ( n29461 , n29457 , n29460 );
and ( n29462 , n29413 , n29460 );
or ( n29463 , n29458 , n29461 , n29462 );
xor ( n29464 , n29189 , n29191 );
xor ( n29465 , n29464 , n29373 );
and ( n29466 , n29463 , n29465 );
xor ( n29467 , n29413 , n29457 );
xor ( n29468 , n29467 , n29460 );
xor ( n29469 , n29310 , n29311 );
and ( n29470 , n29109 , n28564 );
and ( n29471 , n29090 , n28587 );
and ( n29472 , n29470 , n29471 );
and ( n29473 , n28967 , n28615 );
and ( n29474 , n29471 , n29473 );
and ( n29475 , n29470 , n29473 );
or ( n29476 , n29472 , n29474 , n29475 );
and ( n29477 , n28567 , n29118 );
and ( n29478 , n28582 , n29095 );
and ( n29479 , n29477 , n29478 );
and ( n29480 , n28618 , n28964 );
and ( n29481 , n29478 , n29480 );
and ( n29482 , n29477 , n29480 );
or ( n29483 , n29479 , n29481 , n29482 );
and ( n29484 , n29476 , n29483 );
and ( n29485 , n29469 , n29484 );
and ( n29486 , n29289 , n28542 );
and ( n29487 , n29292 , n28553 );
or ( n29488 , n29486 , n29487 );
and ( n29489 , n28545 , n29332 );
and ( n29490 , n28556 , n29304 );
or ( n29491 , n29489 , n29490 );
and ( n29492 , n29488 , n29491 );
and ( n29493 , n29484 , n29492 );
and ( n29494 , n29469 , n29492 );
or ( n29495 , n29485 , n29493 , n29494 );
and ( n29496 , n28911 , n28651 );
not ( n29497 , n29496 );
and ( n29498 , n28840 , n28737 );
and ( n29499 , n29497 , n29498 );
and ( n29500 , n28642 , n28902 );
not ( n29501 , n29500 );
and ( n29502 , n28720 , n28846 );
and ( n29503 , n29501 , n29502 );
and ( n29504 , n29499 , n29503 );
buf ( n29505 , n29496 );
buf ( n29506 , n29500 );
and ( n29507 , n29505 , n29506 );
and ( n29508 , n29504 , n29507 );
xor ( n29509 , n29290 , n29293 );
xor ( n29510 , n29509 , n29295 );
xor ( n29511 , n29333 , n29334 );
xor ( n29512 , n29511 , n29336 );
and ( n29513 , n29510 , n29512 );
and ( n29514 , n29507 , n29513 );
and ( n29515 , n29504 , n29513 );
or ( n29516 , n29508 , n29514 , n29515 );
and ( n29517 , n29495 , n29516 );
xor ( n29518 , n29340 , n29341 );
xor ( n29519 , n29344 , n29345 );
and ( n29520 , n29518 , n29519 );
xor ( n29521 , n29431 , n29432 );
and ( n29522 , n29519 , n29521 );
and ( n29523 , n29518 , n29521 );
or ( n29524 , n29520 , n29522 , n29523 );
xor ( n29525 , n29316 , n29317 );
xor ( n29526 , n29525 , n29319 );
and ( n29527 , n29524 , n29526 );
xor ( n29528 , n29323 , n29324 );
xor ( n29529 , n29528 , n29326 );
and ( n29530 , n29526 , n29529 );
and ( n29531 , n29524 , n29529 );
or ( n29532 , n29527 , n29530 , n29531 );
and ( n29533 , n29516 , n29532 );
and ( n29534 , n29495 , n29532 );
or ( n29535 , n29517 , n29533 , n29534 );
xor ( n29536 , n29277 , n29278 );
xor ( n29537 , n29536 , n29280 );
xor ( n29538 , n29287 , n29308 );
xor ( n29539 , n29538 , n29312 );
and ( n29540 , n29537 , n29539 );
xor ( n29541 , n29322 , n29329 );
xor ( n29542 , n29541 , n29349 );
and ( n29543 , n29539 , n29542 );
and ( n29544 , n29537 , n29542 );
or ( n29545 , n29540 , n29543 , n29544 );
and ( n29546 , n29535 , n29545 );
xor ( n29547 , n29272 , n29273 );
xor ( n29548 , n29547 , n29283 );
and ( n29549 , n29545 , n29548 );
and ( n29550 , n29535 , n29548 );
or ( n29551 , n29546 , n29549 , n29550 );
xor ( n29552 , n29286 , n29358 );
xor ( n29553 , n29552 , n29361 );
and ( n29554 , n29551 , n29553 );
xor ( n29555 , n29315 , n29352 );
xor ( n29556 , n29555 , n29355 );
xor ( n29557 , n29339 , n29342 );
xor ( n29558 , n29557 , n29346 );
xnor ( n29559 , n29489 , n29490 );
not ( n29560 , n29559 );
xor ( n29561 , n29501 , n29502 );
and ( n29562 , n29560 , n29561 );
xnor ( n29563 , n29486 , n29487 );
not ( n29564 , n29563 );
xor ( n29565 , n29497 , n29498 );
and ( n29566 , n29564 , n29565 );
and ( n29567 , n29562 , n29566 );
and ( n29568 , n29558 , n29567 );
buf ( n29569 , n29559 );
buf ( n29570 , n29563 );
and ( n29571 , n29569 , n29570 );
and ( n29572 , n29567 , n29571 );
and ( n29573 , n29558 , n29571 );
or ( n29574 , n29568 , n29572 , n29573 );
xor ( n29575 , n29434 , n29435 );
xor ( n29576 , n29299 , n29300 );
and ( n29577 , n29575 , n29576 );
xor ( n29578 , n29476 , n29483 );
and ( n29579 , n29576 , n29578 );
and ( n29580 , n29575 , n29578 );
or ( n29581 , n29577 , n29579 , n29580 );
xor ( n29582 , n29488 , n29491 );
xor ( n29583 , n29499 , n29503 );
and ( n29584 , n29582 , n29583 );
xor ( n29585 , n29505 , n29506 );
and ( n29586 , n29583 , n29585 );
and ( n29587 , n29582 , n29585 );
or ( n29588 , n29584 , n29586 , n29587 );
and ( n29589 , n29581 , n29588 );
xor ( n29590 , n29510 , n29512 );
and ( n29591 , n29292 , n28564 );
and ( n29592 , n29109 , n28587 );
and ( n29593 , n29591 , n29592 );
and ( n29594 , n28911 , n28737 );
and ( n29595 , n29592 , n29594 );
and ( n29596 , n29591 , n29594 );
or ( n29597 , n29593 , n29595 , n29596 );
and ( n29598 , n29289 , n28553 );
and ( n29599 , n29090 , n28615 );
and ( n29600 , n29598 , n29599 );
and ( n29601 , n28967 , n28651 );
and ( n29602 , n29599 , n29601 );
and ( n29603 , n29598 , n29601 );
or ( n29604 , n29600 , n29602 , n29603 );
and ( n29605 , n29597 , n29604 );
and ( n29606 , n28728 , n28846 );
and ( n29607 , n28840 , n28711 );
and ( n29608 , n29606 , n29607 );
and ( n29609 , n29604 , n29608 );
and ( n29610 , n29597 , n29608 );
or ( n29611 , n29605 , n29609 , n29610 );
and ( n29612 , n29590 , n29611 );
buf ( n29613 , n28728 );
and ( n29614 , n28567 , n29304 );
and ( n29615 , n28582 , n29118 );
and ( n29616 , n29614 , n29615 );
and ( n29617 , n28720 , n28902 );
and ( n29618 , n29615 , n29617 );
and ( n29619 , n29614 , n29617 );
or ( n29620 , n29616 , n29618 , n29619 );
and ( n29621 , n29613 , n29620 );
and ( n29622 , n28556 , n29332 );
and ( n29623 , n28618 , n29095 );
and ( n29624 , n29622 , n29623 );
and ( n29625 , n28642 , n28964 );
and ( n29626 , n29623 , n29625 );
and ( n29627 , n29622 , n29625 );
or ( n29628 , n29624 , n29626 , n29627 );
and ( n29629 , n29620 , n29628 );
and ( n29630 , n29613 , n29628 );
or ( n29631 , n29621 , n29629 , n29630 );
and ( n29632 , n29611 , n29631 );
and ( n29633 , n29590 , n29631 );
or ( n29634 , n29612 , n29632 , n29633 );
and ( n29635 , n29588 , n29634 );
and ( n29636 , n29581 , n29634 );
or ( n29637 , n29589 , n29635 , n29636 );
and ( n29638 , n29574 , n29637 );
xor ( n29639 , n29433 , n29436 );
xor ( n29640 , n29639 , n29439 );
xor ( n29641 , n29469 , n29484 );
xor ( n29642 , n29641 , n29492 );
and ( n29643 , n29640 , n29642 );
xor ( n29644 , n29504 , n29507 );
xor ( n29645 , n29644 , n29513 );
and ( n29646 , n29642 , n29645 );
and ( n29647 , n29640 , n29645 );
or ( n29648 , n29643 , n29646 , n29647 );
and ( n29649 , n29637 , n29648 );
and ( n29650 , n29574 , n29648 );
or ( n29651 , n29638 , n29649 , n29650 );
and ( n29652 , n29556 , n29651 );
xor ( n29653 , n29427 , n29429 );
xor ( n29654 , n29653 , n29442 );
xor ( n29655 , n29495 , n29516 );
xor ( n29656 , n29655 , n29532 );
and ( n29657 , n29654 , n29656 );
xor ( n29658 , n29537 , n29539 );
xor ( n29659 , n29658 , n29542 );
and ( n29660 , n29656 , n29659 );
and ( n29661 , n29654 , n29659 );
or ( n29662 , n29657 , n29660 , n29661 );
and ( n29663 , n29651 , n29662 );
and ( n29664 , n29556 , n29662 );
or ( n29665 , n29652 , n29663 , n29664 );
and ( n29666 , n29553 , n29665 );
and ( n29667 , n29551 , n29665 );
or ( n29668 , n29554 , n29666 , n29667 );
xor ( n29669 , n29415 , n29451 );
xor ( n29670 , n29669 , n29454 );
and ( n29671 , n29668 , n29670 );
xor ( n29672 , n29417 , n29419 );
xor ( n29673 , n29672 , n29448 );
xor ( n29674 , n29422 , n29424 );
xor ( n29675 , n29674 , n29445 );
xor ( n29676 , n29535 , n29545 );
xor ( n29677 , n29676 , n29548 );
and ( n29678 , n29675 , n29677 );
xor ( n29679 , n29524 , n29526 );
xor ( n29680 , n29679 , n29529 );
xor ( n29681 , n29477 , n29478 );
xor ( n29682 , n29681 , n29480 );
not ( n29683 , n29682 );
xor ( n29684 , n29564 , n29565 );
and ( n29685 , n29683 , n29684 );
xor ( n29686 , n29470 , n29471 );
xor ( n29687 , n29686 , n29473 );
not ( n29688 , n29687 );
xor ( n29689 , n29560 , n29561 );
and ( n29690 , n29688 , n29689 );
and ( n29691 , n29685 , n29690 );
and ( n29692 , n29680 , n29691 );
buf ( n29693 , n29682 );
buf ( n29694 , n29687 );
and ( n29695 , n29693 , n29694 );
and ( n29696 , n29691 , n29695 );
and ( n29697 , n29680 , n29695 );
or ( n29698 , n29692 , n29696 , n29697 );
xor ( n29699 , n29518 , n29519 );
xor ( n29700 , n29699 , n29521 );
xor ( n29701 , n29562 , n29566 );
and ( n29702 , n29700 , n29701 );
xor ( n29703 , n29569 , n29570 );
and ( n29704 , n29701 , n29703 );
and ( n29705 , n29700 , n29703 );
or ( n29706 , n29702 , n29704 , n29705 );
xor ( n29707 , n29591 , n29592 );
xor ( n29708 , n29707 , n29594 );
xor ( n29709 , n29598 , n29599 );
xor ( n29710 , n29709 , n29601 );
or ( n29711 , n29708 , n29710 );
and ( n29712 , n29292 , n28587 );
and ( n29713 , n29109 , n28615 );
and ( n29714 , n29712 , n29713 );
and ( n29715 , n29090 , n28651 );
and ( n29716 , n29713 , n29715 );
and ( n29717 , n29712 , n29715 );
or ( n29718 , n29714 , n29716 , n29717 );
and ( n29719 , n28582 , n29304 );
and ( n29720 , n28618 , n29118 );
and ( n29721 , n29719 , n29720 );
and ( n29722 , n28642 , n29095 );
and ( n29723 , n29720 , n29722 );
and ( n29724 , n29719 , n29722 );
or ( n29725 , n29721 , n29723 , n29724 );
and ( n29726 , n29718 , n29725 );
and ( n29727 , n29711 , n29726 );
and ( n29728 , n28967 , n28737 );
and ( n29729 , n28911 , n28711 );
and ( n29730 , n29728 , n29729 );
and ( n29731 , n28720 , n28964 );
and ( n29732 , n28728 , n28902 );
and ( n29733 , n29731 , n29732 );
and ( n29734 , n29730 , n29733 );
and ( n29735 , n29726 , n29734 );
and ( n29736 , n29711 , n29734 );
or ( n29737 , n29727 , n29735 , n29736 );
xor ( n29738 , n29575 , n29576 );
xor ( n29739 , n29738 , n29578 );
and ( n29740 , n29737 , n29739 );
xor ( n29741 , n29582 , n29583 );
xor ( n29742 , n29741 , n29585 );
and ( n29743 , n29739 , n29742 );
and ( n29744 , n29737 , n29742 );
or ( n29745 , n29740 , n29743 , n29744 );
and ( n29746 , n29706 , n29745 );
xor ( n29747 , n29558 , n29567 );
xor ( n29748 , n29747 , n29571 );
and ( n29749 , n29745 , n29748 );
and ( n29750 , n29706 , n29748 );
or ( n29751 , n29746 , n29749 , n29750 );
and ( n29752 , n29698 , n29751 );
xor ( n29753 , n29574 , n29637 );
xor ( n29754 , n29753 , n29648 );
and ( n29755 , n29751 , n29754 );
and ( n29756 , n29698 , n29754 );
or ( n29757 , n29752 , n29755 , n29756 );
and ( n29758 , n29677 , n29757 );
and ( n29759 , n29675 , n29757 );
or ( n29760 , n29678 , n29758 , n29759 );
and ( n29761 , n29673 , n29760 );
xor ( n29762 , n29551 , n29553 );
xor ( n29763 , n29762 , n29665 );
and ( n29764 , n29760 , n29763 );
and ( n29765 , n29673 , n29763 );
or ( n29766 , n29761 , n29764 , n29765 );
and ( n29767 , n29670 , n29766 );
and ( n29768 , n29668 , n29766 );
or ( n29769 , n29671 , n29767 , n29768 );
and ( n29770 , n29468 , n29769 );
xor ( n29771 , n29668 , n29670 );
xor ( n29772 , n29771 , n29766 );
xor ( n29773 , n29556 , n29651 );
xor ( n29774 , n29773 , n29662 );
xor ( n29775 , n29654 , n29656 );
xor ( n29776 , n29775 , n29659 );
xor ( n29777 , n29581 , n29588 );
xor ( n29778 , n29777 , n29634 );
xor ( n29779 , n29640 , n29642 );
xor ( n29780 , n29779 , n29645 );
and ( n29781 , n29778 , n29780 );
xor ( n29782 , n29590 , n29611 );
xor ( n29783 , n29782 , n29631 );
xor ( n29784 , n29685 , n29690 );
and ( n29785 , n29783 , n29784 );
xor ( n29786 , n29693 , n29694 );
and ( n29787 , n29784 , n29786 );
and ( n29788 , n29783 , n29786 );
or ( n29789 , n29785 , n29787 , n29788 );
and ( n29790 , n29780 , n29789 );
and ( n29791 , n29778 , n29789 );
or ( n29792 , n29781 , n29790 , n29791 );
and ( n29793 , n29776 , n29792 );
xor ( n29794 , n29731 , n29732 );
and ( n29795 , n28840 , n28902 );
and ( n29796 , n28911 , n28846 );
and ( n29797 , n29795 , n29796 );
and ( n29798 , n29794 , n29797 );
and ( n29799 , n28567 , n29332 );
and ( n29800 , n29797 , n29799 );
and ( n29801 , n29794 , n29799 );
or ( n29802 , n29798 , n29800 , n29801 );
xor ( n29803 , n29614 , n29615 );
xor ( n29804 , n29803 , n29617 );
and ( n29805 , n29802 , n29804 );
xor ( n29806 , n29622 , n29623 );
xor ( n29807 , n29806 , n29625 );
and ( n29808 , n29804 , n29807 );
and ( n29809 , n29802 , n29807 );
or ( n29810 , n29805 , n29808 , n29809 );
xor ( n29811 , n29597 , n29604 );
xor ( n29812 , n29811 , n29608 );
and ( n29813 , n29810 , n29812 );
xor ( n29814 , n29683 , n29684 );
xor ( n29815 , n29688 , n29689 );
and ( n29816 , n29814 , n29815 );
and ( n29817 , n29813 , n29816 );
xor ( n29818 , n29613 , n29620 );
xor ( n29819 , n29818 , n29628 );
xor ( n29820 , n29606 , n29607 );
xnor ( n29821 , n29708 , n29710 );
and ( n29822 , n29820 , n29821 );
xor ( n29823 , n29718 , n29725 );
and ( n29824 , n29821 , n29823 );
and ( n29825 , n29820 , n29823 );
or ( n29826 , n29822 , n29824 , n29825 );
and ( n29827 , n29819 , n29826 );
xor ( n29828 , n29711 , n29726 );
xor ( n29829 , n29828 , n29734 );
and ( n29830 , n29826 , n29829 );
and ( n29831 , n29819 , n29829 );
or ( n29832 , n29827 , n29830 , n29831 );
and ( n29833 , n29816 , n29832 );
and ( n29834 , n29813 , n29832 );
or ( n29835 , n29817 , n29833 , n29834 );
xor ( n29836 , n29680 , n29691 );
xor ( n29837 , n29836 , n29695 );
and ( n29838 , n29835 , n29837 );
xor ( n29839 , n29706 , n29745 );
xor ( n29840 , n29839 , n29748 );
and ( n29841 , n29837 , n29840 );
and ( n29842 , n29835 , n29840 );
or ( n29843 , n29838 , n29841 , n29842 );
and ( n29844 , n29792 , n29843 );
and ( n29845 , n29776 , n29843 );
or ( n29846 , n29793 , n29844 , n29845 );
and ( n29847 , n29774 , n29846 );
xor ( n29848 , n29675 , n29677 );
xor ( n29849 , n29848 , n29757 );
and ( n29850 , n29846 , n29849 );
and ( n29851 , n29774 , n29849 );
or ( n29852 , n29847 , n29850 , n29851 );
xor ( n29853 , n29673 , n29760 );
xor ( n29854 , n29853 , n29763 );
and ( n29855 , n29852 , n29854 );
xor ( n29856 , n29698 , n29751 );
xor ( n29857 , n29856 , n29754 );
xor ( n29858 , n29700 , n29701 );
xor ( n29859 , n29858 , n29703 );
xor ( n29860 , n29737 , n29739 );
xor ( n29861 , n29860 , n29742 );
and ( n29862 , n29859 , n29861 );
xor ( n29863 , n29810 , n29812 );
xor ( n29864 , n29814 , n29815 );
and ( n29865 , n29863 , n29864 );
and ( n29866 , n28642 , n29118 );
and ( n29867 , n28720 , n29095 );
and ( n29868 , n29866 , n29867 );
and ( n29869 , n28728 , n28964 );
and ( n29870 , n29867 , n29869 );
and ( n29871 , n29866 , n29869 );
or ( n29872 , n29868 , n29870 , n29871 );
and ( n29873 , n29090 , n28711 );
and ( n29874 , n28967 , n28846 );
and ( n29875 , n29873 , n29874 );
and ( n29876 , n28582 , n29332 );
and ( n29877 , n29875 , n29876 );
and ( n29878 , n28618 , n29304 );
and ( n29879 , n29876 , n29878 );
and ( n29880 , n29875 , n29878 );
or ( n29881 , n29877 , n29879 , n29880 );
and ( n29882 , n29872 , n29881 );
xor ( n29883 , n29712 , n29713 );
xor ( n29884 , n29883 , n29715 );
and ( n29885 , n29881 , n29884 );
and ( n29886 , n29872 , n29884 );
or ( n29887 , n29882 , n29885 , n29886 );
and ( n29888 , n29109 , n28651 );
and ( n29889 , n29090 , n28737 );
and ( n29890 , n29888 , n29889 );
and ( n29891 , n28967 , n28711 );
and ( n29892 , n29889 , n29891 );
and ( n29893 , n29888 , n29891 );
or ( n29894 , n29890 , n29892 , n29893 );
and ( n29895 , n28728 , n29095 );
and ( n29896 , n28840 , n28964 );
and ( n29897 , n29895 , n29896 );
and ( n29898 , n29289 , n28587 );
and ( n29899 , n29897 , n29898 );
and ( n29900 , n29292 , n28615 );
and ( n29901 , n29898 , n29900 );
and ( n29902 , n29897 , n29900 );
or ( n29903 , n29899 , n29901 , n29902 );
and ( n29904 , n29894 , n29903 );
xor ( n29905 , n29719 , n29720 );
xor ( n29906 , n29905 , n29722 );
and ( n29907 , n29903 , n29906 );
and ( n29908 , n29894 , n29906 );
or ( n29909 , n29904 , n29907 , n29908 );
and ( n29910 , n29887 , n29909 );
and ( n29911 , n29864 , n29910 );
and ( n29912 , n29863 , n29910 );
or ( n29913 , n29865 , n29911 , n29912 );
and ( n29914 , n29861 , n29913 );
and ( n29915 , n29859 , n29913 );
or ( n29916 , n29862 , n29914 , n29915 );
xor ( n29917 , n29778 , n29780 );
xor ( n29918 , n29917 , n29789 );
and ( n29919 , n29916 , n29918 );
xor ( n29920 , n29835 , n29837 );
xor ( n29921 , n29920 , n29840 );
and ( n29922 , n29918 , n29921 );
and ( n29923 , n29916 , n29921 );
or ( n29924 , n29919 , n29922 , n29923 );
and ( n29925 , n29857 , n29924 );
xor ( n29926 , n29776 , n29792 );
xor ( n29927 , n29926 , n29843 );
and ( n29928 , n29924 , n29927 );
and ( n29929 , n29857 , n29927 );
or ( n29930 , n29925 , n29928 , n29929 );
xor ( n29931 , n29774 , n29846 );
xor ( n29932 , n29931 , n29849 );
and ( n29933 , n29930 , n29932 );
xor ( n29934 , n29857 , n29924 );
xor ( n29935 , n29934 , n29927 );
xor ( n29936 , n29783 , n29784 );
xor ( n29937 , n29936 , n29786 );
xor ( n29938 , n29813 , n29816 );
xor ( n29939 , n29938 , n29832 );
and ( n29940 , n29937 , n29939 );
xor ( n29941 , n29730 , n29733 );
and ( n29942 , n29289 , n28564 );
buf ( n29943 , n28840 );
and ( n29944 , n29942 , n29943 );
xor ( n29945 , n29728 , n29729 );
and ( n29946 , n29943 , n29945 );
and ( n29947 , n29942 , n29945 );
or ( n29948 , n29944 , n29946 , n29947 );
and ( n29949 , n29941 , n29948 );
xor ( n29950 , n29802 , n29804 );
xor ( n29951 , n29950 , n29807 );
and ( n29952 , n29948 , n29951 );
and ( n29953 , n29941 , n29951 );
or ( n29954 , n29949 , n29952 , n29953 );
xor ( n29955 , n29819 , n29826 );
xor ( n29956 , n29955 , n29829 );
and ( n29957 , n29954 , n29956 );
xor ( n29958 , n29794 , n29797 );
xor ( n29959 , n29958 , n29799 );
and ( n29960 , n29289 , n28615 );
and ( n29961 , n29292 , n28651 );
and ( n29962 , n29960 , n29961 );
and ( n29963 , n29109 , n28737 );
and ( n29964 , n29961 , n29963 );
and ( n29965 , n29960 , n29963 );
or ( n29966 , n29962 , n29964 , n29965 );
and ( n29967 , n28618 , n29332 );
and ( n29968 , n28642 , n29304 );
and ( n29969 , n29967 , n29968 );
and ( n29970 , n28720 , n29118 );
and ( n29971 , n29968 , n29970 );
and ( n29972 , n29967 , n29970 );
or ( n29973 , n29969 , n29971 , n29972 );
and ( n29974 , n29966 , n29973 );
and ( n29975 , n29959 , n29974 );
xor ( n29976 , n29888 , n29889 );
xor ( n29977 , n29976 , n29891 );
xor ( n29978 , n29866 , n29867 );
xor ( n29979 , n29978 , n29869 );
and ( n29980 , n29977 , n29979 );
and ( n29981 , n29974 , n29980 );
and ( n29982 , n29959 , n29980 );
or ( n29983 , n29975 , n29981 , n29982 );
xor ( n29984 , n29820 , n29821 );
xor ( n29985 , n29984 , n29823 );
and ( n29986 , n29983 , n29985 );
xor ( n29987 , n29887 , n29909 );
and ( n29988 , n29985 , n29987 );
and ( n29989 , n29983 , n29987 );
or ( n29990 , n29986 , n29988 , n29989 );
and ( n29991 , n29956 , n29990 );
and ( n29992 , n29954 , n29990 );
or ( n29993 , n29957 , n29991 , n29992 );
and ( n29994 , n29939 , n29993 );
and ( n29995 , n29937 , n29993 );
or ( n29996 , n29940 , n29994 , n29995 );
xor ( n29997 , n29916 , n29918 );
xor ( n29998 , n29997 , n29921 );
and ( n29999 , n29996 , n29998 );
xor ( n30000 , n29859 , n29861 );
xor ( n30001 , n30000 , n29913 );
xor ( n30002 , n29872 , n29881 );
xor ( n30003 , n30002 , n29884 );
xor ( n30004 , n29894 , n29903 );
xor ( n30005 , n30004 , n29906 );
and ( n30006 , n30003 , n30005 );
xor ( n30007 , n29942 , n29943 );
xor ( n30008 , n30007 , n29945 );
xor ( n30009 , n29895 , n29896 );
and ( n30010 , n29292 , n28737 );
and ( n30011 , n29109 , n28711 );
and ( n30012 , n30010 , n30011 );
and ( n30013 , n29090 , n28846 );
and ( n30014 , n30011 , n30013 );
and ( n30015 , n30010 , n30013 );
or ( n30016 , n30012 , n30014 , n30015 );
and ( n30017 , n30009 , n30016 );
and ( n30018 , n28911 , n28964 );
and ( n30019 , n28967 , n28902 );
and ( n30020 , n30018 , n30019 );
and ( n30021 , n30016 , n30020 );
and ( n30022 , n30009 , n30020 );
or ( n30023 , n30017 , n30021 , n30022 );
xor ( n30024 , n29897 , n29898 );
xor ( n30025 , n30024 , n29900 );
and ( n30026 , n30023 , n30025 );
and ( n30027 , n30008 , n30026 );
xor ( n30028 , n29795 , n29796 );
xor ( n30029 , n29875 , n29876 );
xor ( n30030 , n30029 , n29878 );
and ( n30031 , n30028 , n30030 );
xor ( n30032 , n29966 , n29973 );
and ( n30033 , n30030 , n30032 );
and ( n30034 , n30028 , n30032 );
or ( n30035 , n30031 , n30033 , n30034 );
and ( n30036 , n30026 , n30035 );
and ( n30037 , n30008 , n30035 );
or ( n30038 , n30027 , n30036 , n30037 );
and ( n30039 , n30006 , n30038 );
xor ( n30040 , n29941 , n29948 );
xor ( n30041 , n30040 , n29951 );
and ( n30042 , n30038 , n30041 );
and ( n30043 , n30006 , n30041 );
or ( n30044 , n30039 , n30042 , n30043 );
xor ( n30045 , n29863 , n29864 );
xor ( n30046 , n30045 , n29910 );
and ( n30047 , n30044 , n30046 );
xor ( n30048 , n29977 , n29979 );
xor ( n30049 , n29960 , n29961 );
xor ( n30050 , n30049 , n29963 );
xor ( n30051 , n29967 , n29968 );
xor ( n30052 , n30051 , n29970 );
and ( n30053 , n30050 , n30052 );
and ( n30054 , n30048 , n30053 );
buf ( n30055 , n28911 );
xor ( n30056 , n29873 , n29874 );
and ( n30057 , n30055 , n30056 );
and ( n30058 , n28720 , n29304 );
and ( n30059 , n28728 , n29118 );
and ( n30060 , n30058 , n30059 );
and ( n30061 , n28840 , n29095 );
and ( n30062 , n30059 , n30061 );
and ( n30063 , n30058 , n30061 );
or ( n30064 , n30060 , n30062 , n30063 );
and ( n30065 , n30056 , n30064 );
and ( n30066 , n30055 , n30064 );
or ( n30067 , n30057 , n30065 , n30066 );
and ( n30068 , n30053 , n30067 );
and ( n30069 , n30048 , n30067 );
or ( n30070 , n30054 , n30068 , n30069 );
xor ( n30071 , n29959 , n29974 );
xor ( n30072 , n30071 , n29980 );
and ( n30073 , n30070 , n30072 );
xor ( n30074 , n30003 , n30005 );
and ( n30075 , n30072 , n30074 );
and ( n30076 , n30070 , n30074 );
or ( n30077 , n30073 , n30075 , n30076 );
xor ( n30078 , n29983 , n29985 );
xor ( n30079 , n30078 , n29987 );
and ( n30080 , n30077 , n30079 );
xor ( n30081 , n30006 , n30038 );
xor ( n30082 , n30081 , n30041 );
and ( n30083 , n30079 , n30082 );
and ( n30084 , n30077 , n30082 );
or ( n30085 , n30080 , n30083 , n30084 );
and ( n30086 , n30046 , n30085 );
and ( n30087 , n30044 , n30085 );
or ( n30088 , n30047 , n30086 , n30087 );
and ( n30089 , n30001 , n30088 );
xor ( n30090 , n29937 , n29939 );
xor ( n30091 , n30090 , n29993 );
and ( n30092 , n30088 , n30091 );
and ( n30093 , n30001 , n30091 );
or ( n30094 , n30089 , n30092 , n30093 );
and ( n30095 , n29998 , n30094 );
and ( n30096 , n29996 , n30094 );
or ( n30097 , n29999 , n30095 , n30096 );
and ( n30098 , n29935 , n30097 );
xor ( n30099 , n29996 , n29998 );
xor ( n30100 , n30099 , n30094 );
xor ( n30101 , n30001 , n30088 );
xor ( n30102 , n30101 , n30091 );
xor ( n30103 , n29954 , n29956 );
xor ( n30104 , n30103 , n29990 );
xor ( n30105 , n30044 , n30046 );
xor ( n30106 , n30105 , n30085 );
and ( n30107 , n30104 , n30106 );
xor ( n30108 , n30023 , n30025 );
and ( n30109 , n28840 , n29118 );
and ( n30110 , n28911 , n29095 );
and ( n30111 , n30109 , n30110 );
and ( n30112 , n29289 , n28651 );
and ( n30113 , n30111 , n30112 );
and ( n30114 , n29109 , n28846 );
and ( n30115 , n29090 , n28902 );
and ( n30116 , n30114 , n30115 );
and ( n30117 , n28642 , n29332 );
and ( n30118 , n30116 , n30117 );
and ( n30119 , n30113 , n30118 );
and ( n30120 , n30108 , n30119 );
xor ( n30121 , n30009 , n30016 );
xor ( n30122 , n30121 , n30020 );
xor ( n30123 , n30050 , n30052 );
and ( n30124 , n30122 , n30123 );
xor ( n30125 , n30058 , n30059 );
xor ( n30126 , n30125 , n30061 );
xor ( n30127 , n30018 , n30019 );
and ( n30128 , n30126 , n30127 );
and ( n30129 , n29289 , n28737 );
and ( n30130 , n29292 , n28711 );
and ( n30131 , n30129 , n30130 );
and ( n30132 , n30127 , n30131 );
and ( n30133 , n30126 , n30131 );
or ( n30134 , n30128 , n30132 , n30133 );
and ( n30135 , n30123 , n30134 );
and ( n30136 , n30122 , n30134 );
or ( n30137 , n30124 , n30135 , n30136 );
and ( n30138 , n30119 , n30137 );
and ( n30139 , n30108 , n30137 );
or ( n30140 , n30120 , n30138 , n30139 );
xor ( n30141 , n30008 , n30026 );
xor ( n30142 , n30141 , n30035 );
and ( n30143 , n30140 , n30142 );
xor ( n30144 , n30028 , n30030 );
xor ( n30145 , n30144 , n30032 );
xor ( n30146 , n30048 , n30053 );
xor ( n30147 , n30146 , n30067 );
and ( n30148 , n30145 , n30147 );
xor ( n30149 , n30055 , n30056 );
xor ( n30150 , n30149 , n30064 );
xor ( n30151 , n30113 , n30118 );
and ( n30152 , n30150 , n30151 );
and ( n30153 , n28967 , n29095 );
and ( n30154 , n29090 , n28964 );
and ( n30155 , n30153 , n30154 );
and ( n30156 , n28720 , n29332 );
and ( n30157 , n30155 , n30156 );
and ( n30158 , n28728 , n29304 );
and ( n30159 , n30156 , n30158 );
and ( n30160 , n30155 , n30158 );
or ( n30161 , n30157 , n30159 , n30160 );
xor ( n30162 , n30010 , n30011 );
xor ( n30163 , n30162 , n30013 );
and ( n30164 , n30161 , n30163 );
and ( n30165 , n30151 , n30164 );
and ( n30166 , n30150 , n30164 );
or ( n30167 , n30152 , n30165 , n30166 );
and ( n30168 , n30147 , n30167 );
and ( n30169 , n30145 , n30167 );
or ( n30170 , n30148 , n30168 , n30169 );
and ( n30171 , n30142 , n30170 );
and ( n30172 , n30140 , n30170 );
or ( n30173 , n30143 , n30171 , n30172 );
xor ( n30174 , n30077 , n30079 );
xor ( n30175 , n30174 , n30082 );
and ( n30176 , n30173 , n30175 );
xor ( n30177 , n30070 , n30072 );
xor ( n30178 , n30177 , n30074 );
xor ( n30179 , n30108 , n30119 );
xor ( n30180 , n30179 , n30137 );
xor ( n30181 , n30111 , n30112 );
xor ( n30182 , n30116 , n30117 );
and ( n30183 , n30181 , n30182 );
xor ( n30184 , n30122 , n30123 );
xor ( n30185 , n30184 , n30134 );
and ( n30186 , n30183 , n30185 );
and ( n30187 , n28728 , n29332 );
and ( n30188 , n28840 , n29304 );
and ( n30189 , n30187 , n30188 );
and ( n30190 , n28911 , n29118 );
and ( n30191 , n30188 , n30190 );
and ( n30192 , n30187 , n30190 );
or ( n30193 , n30189 , n30191 , n30192 );
xor ( n30194 , n30114 , n30115 );
and ( n30195 , n30193 , n30194 );
xor ( n30196 , n30126 , n30127 );
xor ( n30197 , n30196 , n30131 );
and ( n30198 , n30195 , n30197 );
xor ( n30199 , n30161 , n30163 );
and ( n30200 , n30197 , n30199 );
and ( n30201 , n30195 , n30199 );
or ( n30202 , n30198 , n30200 , n30201 );
and ( n30203 , n30185 , n30202 );
and ( n30204 , n30183 , n30202 );
or ( n30205 , n30186 , n30203 , n30204 );
and ( n30206 , n30180 , n30205 );
xor ( n30207 , n30145 , n30147 );
xor ( n30208 , n30207 , n30167 );
and ( n30209 , n30205 , n30208 );
and ( n30210 , n30180 , n30208 );
or ( n30211 , n30206 , n30209 , n30210 );
and ( n30212 , n30178 , n30211 );
xor ( n30213 , n30140 , n30142 );
xor ( n30214 , n30213 , n30170 );
and ( n30215 , n30211 , n30214 );
and ( n30216 , n30178 , n30214 );
or ( n30217 , n30212 , n30215 , n30216 );
and ( n30218 , n30175 , n30217 );
and ( n30219 , n30173 , n30217 );
or ( n30220 , n30176 , n30218 , n30219 );
and ( n30221 , n30106 , n30220 );
and ( n30222 , n30104 , n30220 );
or ( n30223 , n30107 , n30221 , n30222 );
or ( n30224 , n30102 , n30223 );
or ( n30225 , n30100 , n30224 );
and ( n30226 , n30097 , n30225 );
and ( n30227 , n29935 , n30225 );
or ( n30228 , n30098 , n30226 , n30227 );
and ( n30229 , n29932 , n30228 );
and ( n30230 , n29930 , n30228 );
or ( n30231 , n29933 , n30229 , n30230 );
and ( n30232 , n29854 , n30231 );
and ( n30233 , n29852 , n30231 );
or ( n30234 , n29855 , n30232 , n30233 );
or ( n30235 , n29772 , n30234 );
and ( n30236 , n29769 , n30235 );
and ( n30237 , n29468 , n30235 );
or ( n30238 , n29770 , n30236 , n30237 );
and ( n30239 , n29465 , n30238 );
and ( n30240 , n29463 , n30238 );
or ( n30241 , n29466 , n30239 , n30240 );
and ( n30242 , n29411 , n30241 );
xor ( n30243 , n29411 , n30241 );
xor ( n30244 , n29463 , n29465 );
xor ( n30245 , n30244 , n30238 );
not ( n30246 , n30245 );
xor ( n30247 , n29468 , n29769 );
xor ( n30248 , n30247 , n30235 );
xnor ( n30249 , n29772 , n30234 );
xor ( n30250 , n29852 , n29854 );
xor ( n30251 , n30250 , n30231 );
xor ( n30252 , n29930 , n29932 );
xor ( n30253 , n30252 , n30228 );
not ( n30254 , n30253 );
xor ( n30255 , n29935 , n30097 );
xor ( n30256 , n30255 , n30225 );
not ( n30257 , n30256 );
xnor ( n30258 , n30100 , n30224 );
xnor ( n30259 , n30102 , n30223 );
xor ( n30260 , n30104 , n30106 );
xor ( n30261 , n30260 , n30220 );
not ( n30262 , n30261 );
xor ( n30263 , n30173 , n30175 );
xor ( n30264 , n30263 , n30217 );
xor ( n30265 , n30178 , n30211 );
xor ( n30266 , n30265 , n30214 );
xor ( n30267 , n30181 , n30182 );
xor ( n30268 , n30109 , n30110 );
and ( n30269 , n29289 , n28711 );
and ( n30270 , n29292 , n28846 );
and ( n30271 , n30269 , n30270 );
and ( n30272 , n29109 , n28902 );
and ( n30273 , n30270 , n30272 );
and ( n30274 , n30269 , n30272 );
or ( n30275 , n30271 , n30273 , n30274 );
and ( n30276 , n30268 , n30275 );
xor ( n30277 , n30155 , n30156 );
xor ( n30278 , n30277 , n30158 );
and ( n30279 , n30275 , n30278 );
and ( n30280 , n30268 , n30278 );
or ( n30281 , n30276 , n30279 , n30280 );
and ( n30282 , n30267 , n30281 );
buf ( n30283 , n28967 );
xor ( n30284 , n30129 , n30130 );
and ( n30285 , n30283 , n30284 );
xor ( n30286 , n30193 , n30194 );
and ( n30287 , n30284 , n30286 );
and ( n30288 , n30283 , n30286 );
or ( n30289 , n30285 , n30287 , n30288 );
and ( n30290 , n30281 , n30289 );
and ( n30291 , n30267 , n30289 );
or ( n30292 , n30282 , n30290 , n30291 );
xor ( n30293 , n30150 , n30151 );
xor ( n30294 , n30293 , n30164 );
and ( n30295 , n30292 , n30294 );
and ( n30296 , n29292 , n28902 );
and ( n30297 , n29109 , n28964 );
and ( n30298 , n30296 , n30297 );
and ( n30299 , n28911 , n29304 );
and ( n30300 , n28967 , n29118 );
and ( n30301 , n30299 , n30300 );
and ( n30302 , n30298 , n30301 );
xor ( n30303 , n30269 , n30270 );
xor ( n30304 , n30303 , n30272 );
xor ( n30305 , n30187 , n30188 );
xor ( n30306 , n30305 , n30190 );
and ( n30307 , n30304 , n30306 );
and ( n30308 , n30302 , n30307 );
xor ( n30309 , n30268 , n30275 );
xor ( n30310 , n30309 , n30278 );
and ( n30311 , n30307 , n30310 );
and ( n30312 , n30302 , n30310 );
or ( n30313 , n30308 , n30311 , n30312 );
xor ( n30314 , n30153 , n30154 );
xor ( n30315 , n30298 , n30301 );
and ( n30316 , n30314 , n30315 );
xor ( n30317 , n30304 , n30306 );
and ( n30318 , n30315 , n30317 );
and ( n30319 , n30314 , n30317 );
or ( n30320 , n30316 , n30318 , n30319 );
xor ( n30321 , n30299 , n30300 );
and ( n30322 , n29090 , n29118 );
and ( n30323 , n29109 , n29095 );
and ( n30324 , n30322 , n30323 );
and ( n30325 , n30321 , n30324 );
and ( n30326 , n28840 , n29332 );
and ( n30327 , n30324 , n30326 );
and ( n30328 , n30321 , n30326 );
or ( n30329 , n30325 , n30327 , n30328 );
and ( n30330 , n29289 , n28902 );
and ( n30331 , n29292 , n28964 );
and ( n30332 , n30330 , n30331 );
and ( n30333 , n28911 , n29332 );
and ( n30334 , n28967 , n29304 );
and ( n30335 , n30333 , n30334 );
and ( n30336 , n30332 , n30335 );
and ( n30337 , n30329 , n30336 );
and ( n30338 , n29289 , n28846 );
buf ( n30339 , n29090 );
and ( n30340 , n30338 , n30339 );
xor ( n30341 , n30296 , n30297 );
and ( n30342 , n30339 , n30341 );
and ( n30343 , n30338 , n30341 );
or ( n30344 , n30340 , n30342 , n30343 );
and ( n30345 , n30336 , n30344 );
and ( n30346 , n30329 , n30344 );
or ( n30347 , n30337 , n30345 , n30346 );
and ( n30348 , n30320 , n30347 );
xor ( n30349 , n30283 , n30284 );
xor ( n30350 , n30349 , n30286 );
and ( n30351 , n30347 , n30350 );
and ( n30352 , n30320 , n30350 );
or ( n30353 , n30348 , n30351 , n30352 );
and ( n30354 , n30313 , n30353 );
xor ( n30355 , n30195 , n30197 );
xor ( n30356 , n30355 , n30199 );
and ( n30357 , n30353 , n30356 );
and ( n30358 , n30313 , n30356 );
or ( n30359 , n30354 , n30357 , n30358 );
and ( n30360 , n30294 , n30359 );
and ( n30361 , n30292 , n30359 );
or ( n30362 , n30295 , n30360 , n30361 );
xor ( n30363 , n30180 , n30205 );
xor ( n30364 , n30363 , n30208 );
and ( n30365 , n30362 , n30364 );
xor ( n30366 , n30183 , n30185 );
xor ( n30367 , n30366 , n30202 );
xor ( n30368 , n30267 , n30281 );
xor ( n30369 , n30368 , n30289 );
xor ( n30370 , n30321 , n30324 );
xor ( n30371 , n30370 , n30326 );
xor ( n30372 , n30332 , n30335 );
and ( n30373 , n30371 , n30372 );
and ( n30374 , n29289 , n28964 );
and ( n30375 , n29292 , n29095 );
and ( n30376 , n30374 , n30375 );
and ( n30377 , n28967 , n29332 );
and ( n30378 , n29090 , n29304 );
and ( n30379 , n30377 , n30378 );
and ( n30380 , n30376 , n30379 );
and ( n30381 , n30372 , n30380 );
and ( n30382 , n30371 , n30380 );
or ( n30383 , n30373 , n30381 , n30382 );
xor ( n30384 , n30314 , n30315 );
xor ( n30385 , n30384 , n30317 );
and ( n30386 , n30383 , n30385 );
xor ( n30387 , n30329 , n30336 );
xor ( n30388 , n30387 , n30344 );
and ( n30389 , n30385 , n30388 );
and ( n30390 , n30383 , n30388 );
or ( n30391 , n30386 , n30389 , n30390 );
xor ( n30392 , n30302 , n30307 );
xor ( n30393 , n30392 , n30310 );
and ( n30394 , n30391 , n30393 );
xor ( n30395 , n30320 , n30347 );
xor ( n30396 , n30395 , n30350 );
and ( n30397 , n30393 , n30396 );
and ( n30398 , n30391 , n30396 );
or ( n30399 , n30394 , n30397 , n30398 );
and ( n30400 , n30369 , n30399 );
xor ( n30401 , n30313 , n30353 );
xor ( n30402 , n30401 , n30356 );
and ( n30403 , n30399 , n30402 );
and ( n30404 , n30369 , n30402 );
or ( n30405 , n30400 , n30403 , n30404 );
and ( n30406 , n30367 , n30405 );
xor ( n30407 , n30292 , n30294 );
xor ( n30408 , n30407 , n30359 );
and ( n30409 , n30405 , n30408 );
and ( n30410 , n30367 , n30408 );
or ( n30411 , n30406 , n30409 , n30410 );
and ( n30412 , n30364 , n30411 );
and ( n30413 , n30362 , n30411 );
or ( n30414 , n30365 , n30412 , n30413 );
and ( n30415 , n30266 , n30414 );
xor ( n30416 , n30362 , n30364 );
xor ( n30417 , n30416 , n30411 );
xor ( n30418 , n30367 , n30405 );
xor ( n30419 , n30418 , n30408 );
xor ( n30420 , n30369 , n30399 );
xor ( n30421 , n30420 , n30402 );
xor ( n30422 , n30391 , n30393 );
xor ( n30423 , n30422 , n30396 );
xor ( n30424 , n30330 , n30331 );
xor ( n30425 , n30333 , n30334 );
and ( n30426 , n30424 , n30425 );
xor ( n30427 , n30338 , n30339 );
xor ( n30428 , n30427 , n30341 );
and ( n30429 , n30426 , n30428 );
xor ( n30430 , n30322 , n30323 );
xor ( n30431 , n30376 , n30379 );
and ( n30432 , n30430 , n30431 );
xor ( n30433 , n30424 , n30425 );
and ( n30434 , n30431 , n30433 );
and ( n30435 , n30430 , n30433 );
or ( n30436 , n30432 , n30434 , n30435 );
and ( n30437 , n30428 , n30436 );
and ( n30438 , n30426 , n30436 );
or ( n30439 , n30429 , n30437 , n30438 );
xor ( n30440 , n30383 , n30385 );
xor ( n30441 , n30440 , n30388 );
and ( n30442 , n30439 , n30441 );
xor ( n30443 , n30371 , n30372 );
xor ( n30444 , n30443 , n30380 );
and ( n30445 , n29090 , n29332 );
and ( n30446 , n29289 , n29095 );
and ( n30447 , n30445 , n30446 );
buf ( n30448 , n29109 );
or ( n30449 , n30447 , n30448 );
xor ( n30450 , n30374 , n30375 );
xor ( n30451 , n30377 , n30378 );
and ( n30452 , n30450 , n30451 );
and ( n30453 , n30449 , n30452 );
and ( n30454 , n29109 , n29304 );
and ( n30455 , n29292 , n29118 );
and ( n30456 , n30454 , n30455 );
xnor ( n30457 , n30447 , n30448 );
or ( n30458 , n30456 , n30457 );
and ( n30459 , n30452 , n30458 );
and ( n30460 , n30449 , n30458 );
or ( n30461 , n30453 , n30459 , n30460 );
and ( n30462 , n30444 , n30461 );
xor ( n30463 , n30426 , n30428 );
xor ( n30464 , n30463 , n30436 );
and ( n30465 , n30461 , n30464 );
and ( n30466 , n30444 , n30464 );
or ( n30467 , n30462 , n30465 , n30466 );
and ( n30468 , n30441 , n30467 );
and ( n30469 , n30439 , n30467 );
or ( n30470 , n30442 , n30468 , n30469 );
and ( n30471 , n30423 , n30470 );
xor ( n30472 , n30430 , n30431 );
xor ( n30473 , n30472 , n30433 );
xor ( n30474 , n30450 , n30451 );
xnor ( n30475 , n30456 , n30457 );
and ( n30476 , n30474 , n30475 );
xor ( n30477 , n30445 , n30446 );
xor ( n30478 , n30454 , n30455 );
and ( n30479 , n30477 , n30478 );
and ( n30480 , n29292 , n29332 );
and ( n30481 , n29289 , n29304 );
and ( n30482 , n30480 , n30481 );
and ( n30483 , n29109 , n29332 );
and ( n30484 , n30482 , n30483 );
and ( n30485 , n30478 , n30484 );
and ( n30486 , n30477 , n30484 );
or ( n30487 , n30479 , n30485 , n30486 );
and ( n30488 , n30475 , n30487 );
and ( n30489 , n30474 , n30487 );
or ( n30490 , n30476 , n30488 , n30489 );
and ( n30491 , n30473 , n30490 );
xor ( n30492 , n30449 , n30452 );
xor ( n30493 , n30492 , n30458 );
and ( n30494 , n30490 , n30493 );
and ( n30495 , n30473 , n30493 );
or ( n30496 , n30491 , n30494 , n30495 );
xor ( n30497 , n30444 , n30461 );
xor ( n30498 , n30497 , n30464 );
or ( n30499 , n30496 , n30498 );
xor ( n30500 , n30439 , n30441 );
xor ( n30501 , n30500 , n30467 );
or ( n30502 , n30499 , n30501 );
and ( n30503 , n30470 , n30502 );
and ( n30504 , n30423 , n30502 );
or ( n30505 , n30471 , n30503 , n30504 );
or ( n30506 , n30421 , n30505 );
or ( n30507 , n30419 , n30506 );
or ( n30508 , n30417 , n30507 );
and ( n30509 , n30414 , n30508 );
and ( n30510 , n30266 , n30508 );
or ( n30511 , n30415 , n30509 , n30510 );
and ( n30512 , n30264 , n30511 );
xor ( n30513 , n30264 , n30511 );
xor ( n30514 , n30266 , n30414 );
xor ( n30515 , n30514 , n30508 );
not ( n30516 , n30515 );
xnor ( n30517 , n30417 , n30507 );
xnor ( n30518 , n30419 , n30506 );
xnor ( n30519 , n30421 , n30505 );
xor ( n30520 , n30423 , n30470 );
xor ( n30521 , n30520 , n30502 );
not ( n30522 , n30521 );
xnor ( n30523 , n30499 , n30501 );
xnor ( n30524 , n30496 , n30498 );
xor ( n30525 , n30473 , n30490 );
xor ( n30526 , n30525 , n30493 );
buf ( n30527 , n29292 );
not ( n30528 , n30527 );
xor ( n30529 , n30482 , n30483 );
and ( n30530 , n30528 , n30529 );
buf ( n30531 , n30527 );
and ( n30532 , n30530 , n30531 );
xor ( n30533 , n30477 , n30478 );
xor ( n30534 , n30533 , n30484 );
and ( n30535 , n30531 , n30534 );
and ( n30536 , n30530 , n30534 );
or ( n30537 , n30532 , n30535 , n30536 );
xor ( n30538 , n30474 , n30475 );
xor ( n30539 , n30538 , n30487 );
and ( n30540 , n30537 , n30539 );
and ( n30541 , n29289 , n29118 );
xor ( n30542 , n30528 , n30529 );
or ( n30543 , n30541 , n30542 );
xor ( n30544 , n30530 , n30531 );
xor ( n30545 , n30544 , n30534 );
or ( n30546 , n30543 , n30545 );
and ( n30547 , n30539 , n30546 );
and ( n30548 , n30537 , n30546 );
or ( n30549 , n30540 , n30547 , n30548 );
and ( n30550 , n30526 , n30549 );
xor ( n30551 , n30526 , n30549 );
xor ( n30552 , n30537 , n30539 );
xor ( n30553 , n30552 , n30546 );
and ( n30554 , n30551 , n30553 );
or ( n30555 , n30550 , n30554 );
and ( n30556 , n30524 , n30555 );
and ( n30557 , n30523 , n30556 );
and ( n30558 , n30522 , n30557 );
or ( n30559 , n30521 , n30558 );
and ( n30560 , n30519 , n30559 );
and ( n30561 , n30518 , n30560 );
and ( n30562 , n30517 , n30561 );
and ( n30563 , n30516 , n30562 );
or ( n30564 , n30515 , n30563 );
and ( n30565 , n30513 , n30564 );
or ( n30566 , n30512 , n30565 );
and ( n30567 , n30262 , n30566 );
or ( n30568 , n30261 , n30567 );
and ( n30569 , n30259 , n30568 );
and ( n30570 , n30258 , n30569 );
and ( n30571 , n30257 , n30570 );
or ( n30572 , n30256 , n30571 );
and ( n30573 , n30254 , n30572 );
or ( n30574 , n30253 , n30573 );
and ( n30575 , n30251 , n30574 );
and ( n30576 , n30249 , n30575 );
and ( n30577 , n30248 , n30576 );
and ( n30578 , n30246 , n30577 );
or ( n30579 , n30245 , n30578 );
and ( n30580 , n30243 , n30579 );
or ( n30581 , n30242 , n30580 );
and ( n30582 , n29409 , n30581 );
or ( n30583 , n29408 , n30582 );
and ( n30584 , n29406 , n30583 );
and ( n30585 , n29405 , n30584 );
and ( n30586 , n29404 , n30585 );
and ( n30587 , n29402 , n30586 );
or ( n30588 , n29401 , n30587 );
and ( n30589 , n29399 , n30588 );
and ( n30590 , n29398 , n30589 );
or ( n30591 , n29397 , n30590 );
xor ( n30592 , n29395 , n30591 );
buf ( n30593 , n30592 );
buf ( n30594 , n30593 );
buf ( n30595 , n30594 );
buf ( n30596 , n778 );
buf ( n30597 , n30596 );
buf ( n30598 , n779 );
buf ( n30599 , n30598 );
xor ( n30600 , n30597 , n30599 );
buf ( n30601 , n780 );
buf ( n30602 , n30601 );
xor ( n30603 , n30599 , n30602 );
not ( n30604 , n30603 );
and ( n30605 , n30600 , n30604 );
and ( n30606 , n30595 , n30605 );
not ( n30607 , n30606 );
and ( n30608 , n30599 , n30602 );
not ( n30609 , n30608 );
and ( n30610 , n30597 , n30609 );
xnor ( n30611 , n30607 , n30610 );
buf ( n30612 , n30611 );
buf ( n30613 , n781 );
buf ( n30614 , n30613 );
buf ( n30615 , n782 );
buf ( n30616 , n30615 );
and ( n30617 , n30614 , n30616 );
not ( n30618 , n30617 );
and ( n30619 , n30602 , n30618 );
not ( n30620 , n30619 );
xor ( n30621 , n29398 , n30589 );
buf ( n30622 , n30621 );
buf ( n30623 , n30622 );
buf ( n30624 , n30623 );
and ( n30625 , n30624 , n30605 );
and ( n30626 , n30595 , n30603 );
nor ( n30627 , n30625 , n30626 );
xnor ( n30628 , n30627 , n30610 );
and ( n30629 , n30620 , n30628 );
xor ( n30630 , n29399 , n30588 );
buf ( n30631 , n30630 );
buf ( n30632 , n30631 );
buf ( n30633 , n30632 );
and ( n30634 , n30633 , n30597 );
and ( n30635 , n30628 , n30634 );
and ( n30636 , n30620 , n30634 );
or ( n30637 , n30629 , n30635 , n30636 );
not ( n30638 , n30611 );
xor ( n30639 , n30637 , n30638 );
and ( n30640 , n30624 , n30597 );
xor ( n30641 , n30639 , n30640 );
xor ( n30642 , n30602 , n30614 );
xor ( n30643 , n30614 , n30616 );
not ( n30644 , n30643 );
and ( n30645 , n30642 , n30644 );
and ( n30646 , n30595 , n30645 );
not ( n30647 , n30646 );
xnor ( n30648 , n30647 , n30619 );
not ( n30649 , n30648 );
and ( n30650 , n30633 , n30605 );
and ( n30651 , n30624 , n30603 );
nor ( n30652 , n30650 , n30651 );
xnor ( n30653 , n30652 , n30610 );
and ( n30654 , n30649 , n30653 );
xor ( n30655 , n29402 , n30586 );
buf ( n30656 , n30655 );
buf ( n30657 , n30656 );
buf ( n30658 , n30657 );
and ( n30659 , n30658 , n30597 );
and ( n30660 , n30653 , n30659 );
and ( n30661 , n30649 , n30659 );
or ( n30662 , n30654 , n30660 , n30661 );
buf ( n30663 , n30648 );
and ( n30664 , n30662 , n30663 );
xor ( n30665 , n30620 , n30628 );
xor ( n30666 , n30665 , n30634 );
and ( n30667 , n30663 , n30666 );
and ( n30668 , n30662 , n30666 );
or ( n30669 , n30664 , n30667 , n30668 );
and ( n30670 , n30641 , n30669 );
xor ( n30671 , n30612 , n30670 );
not ( n30672 , n30610 );
and ( n30673 , n30595 , n30597 );
xor ( n30674 , n30672 , n30673 );
and ( n30675 , n30637 , n30638 );
and ( n30676 , n30638 , n30640 );
and ( n30677 , n30637 , n30640 );
or ( n30678 , n30675 , n30676 , n30677 );
xor ( n30679 , n30674 , n30678 );
xor ( n30680 , n30671 , n30679 );
xor ( n30681 , n30641 , n30669 );
xor ( n30682 , n30662 , n30663 );
xor ( n30683 , n30682 , n30666 );
buf ( n30684 , n783 );
buf ( n30685 , n30684 );
xor ( n30686 , n30616 , n30685 );
buf ( n30687 , n784 );
buf ( n30688 , n30687 );
xor ( n30689 , n30685 , n30688 );
not ( n30690 , n30689 );
and ( n30691 , n30686 , n30690 );
and ( n30692 , n30595 , n30691 );
not ( n30693 , n30692 );
and ( n30694 , n30685 , n30688 );
not ( n30695 , n30694 );
and ( n30696 , n30616 , n30695 );
xnor ( n30697 , n30693 , n30696 );
buf ( n30698 , n30697 );
not ( n30699 , n30696 );
and ( n30700 , n30698 , n30699 );
xor ( n30701 , n29404 , n30585 );
buf ( n30702 , n30701 );
buf ( n30703 , n30702 );
buf ( n30704 , n30703 );
and ( n30705 , n30704 , n30597 );
and ( n30706 , n30699 , n30705 );
and ( n30707 , n30698 , n30705 );
or ( n30708 , n30700 , n30706 , n30707 );
not ( n30709 , n30697 );
and ( n30710 , n30704 , n30605 );
and ( n30711 , n30658 , n30603 );
nor ( n30712 , n30710 , n30711 );
xnor ( n30713 , n30712 , n30610 );
and ( n30714 , n30709 , n30713 );
xor ( n30715 , n29405 , n30584 );
buf ( n30716 , n30715 );
buf ( n30717 , n30716 );
buf ( n30718 , n30717 );
and ( n30719 , n30718 , n30597 );
and ( n30720 , n30713 , n30719 );
and ( n30721 , n30709 , n30719 );
or ( n30722 , n30714 , n30720 , n30721 );
and ( n30723 , n30624 , n30645 );
and ( n30724 , n30595 , n30643 );
nor ( n30725 , n30723 , n30724 );
xnor ( n30726 , n30725 , n30619 );
and ( n30727 , n30722 , n30726 );
and ( n30728 , n30658 , n30605 );
and ( n30729 , n30633 , n30603 );
nor ( n30730 , n30728 , n30729 );
xnor ( n30731 , n30730 , n30610 );
and ( n30732 , n30726 , n30731 );
and ( n30733 , n30722 , n30731 );
or ( n30734 , n30727 , n30732 , n30733 );
and ( n30735 , n30708 , n30734 );
xor ( n30736 , n30649 , n30653 );
xor ( n30737 , n30736 , n30659 );
and ( n30738 , n30734 , n30737 );
and ( n30739 , n30708 , n30737 );
or ( n30740 , n30735 , n30738 , n30739 );
and ( n30741 , n30683 , n30740 );
and ( n30742 , n30681 , n30741 );
xor ( n30743 , n30683 , n30740 );
xor ( n30744 , n30708 , n30734 );
xor ( n30745 , n30744 , n30737 );
buf ( n30746 , n785 );
buf ( n30747 , n30746 );
buf ( n30748 , n786 );
buf ( n30749 , n30748 );
and ( n30750 , n30747 , n30749 );
not ( n30751 , n30750 );
and ( n30752 , n30688 , n30751 );
not ( n30753 , n30752 );
and ( n30754 , n30624 , n30691 );
and ( n30755 , n30595 , n30689 );
nor ( n30756 , n30754 , n30755 );
xnor ( n30757 , n30756 , n30696 );
and ( n30758 , n30753 , n30757 );
xor ( n30759 , n29406 , n30583 );
buf ( n30760 , n30759 );
buf ( n30761 , n30760 );
buf ( n30762 , n30761 );
and ( n30763 , n30762 , n30597 );
and ( n30764 , n30757 , n30763 );
and ( n30765 , n30753 , n30763 );
or ( n30766 , n30758 , n30764 , n30765 );
xor ( n30767 , n30688 , n30747 );
xor ( n30768 , n30747 , n30749 );
not ( n30769 , n30768 );
and ( n30770 , n30767 , n30769 );
and ( n30771 , n30595 , n30770 );
not ( n30772 , n30771 );
xnor ( n30773 , n30772 , n30752 );
buf ( n30774 , n30773 );
and ( n30775 , n30658 , n30645 );
and ( n30776 , n30633 , n30643 );
nor ( n30777 , n30775 , n30776 );
xnor ( n30778 , n30777 , n30619 );
and ( n30779 , n30774 , n30778 );
and ( n30780 , n30718 , n30605 );
and ( n30781 , n30704 , n30603 );
nor ( n30782 , n30780 , n30781 );
xnor ( n30783 , n30782 , n30610 );
and ( n30784 , n30778 , n30783 );
and ( n30785 , n30774 , n30783 );
or ( n30786 , n30779 , n30784 , n30785 );
and ( n30787 , n30766 , n30786 );
and ( n30788 , n30633 , n30645 );
and ( n30789 , n30624 , n30643 );
nor ( n30790 , n30788 , n30789 );
xnor ( n30791 , n30790 , n30619 );
and ( n30792 , n30786 , n30791 );
and ( n30793 , n30766 , n30791 );
or ( n30794 , n30787 , n30792 , n30793 );
xor ( n30795 , n30698 , n30699 );
xor ( n30796 , n30795 , n30705 );
and ( n30797 , n30794 , n30796 );
xor ( n30798 , n30722 , n30726 );
xor ( n30799 , n30798 , n30731 );
and ( n30800 , n30796 , n30799 );
and ( n30801 , n30794 , n30799 );
or ( n30802 , n30797 , n30800 , n30801 );
and ( n30803 , n30745 , n30802 );
and ( n30804 , n30743 , n30803 );
xor ( n30805 , n30794 , n30796 );
xor ( n30806 , n30805 , n30799 );
not ( n30807 , n30773 );
and ( n30808 , n30704 , n30645 );
and ( n30809 , n30658 , n30643 );
nor ( n30810 , n30808 , n30809 );
xnor ( n30811 , n30810 , n30619 );
and ( n30812 , n30807 , n30811 );
xor ( n30813 , n29409 , n30581 );
buf ( n30814 , n30813 );
buf ( n30815 , n30814 );
buf ( n30816 , n30815 );
and ( n30817 , n30816 , n30597 );
and ( n30818 , n30811 , n30817 );
and ( n30819 , n30807 , n30817 );
or ( n30820 , n30812 , n30818 , n30819 );
xor ( n30821 , n30753 , n30757 );
xor ( n30822 , n30821 , n30763 );
and ( n30823 , n30820 , n30822 );
xor ( n30824 , n30774 , n30778 );
xor ( n30825 , n30824 , n30783 );
and ( n30826 , n30822 , n30825 );
and ( n30827 , n30820 , n30825 );
or ( n30828 , n30823 , n30826 , n30827 );
xor ( n30829 , n30766 , n30786 );
xor ( n30830 , n30829 , n30791 );
and ( n30831 , n30828 , n30830 );
xor ( n30832 , n30709 , n30713 );
xor ( n30833 , n30832 , n30719 );
and ( n30834 , n30830 , n30833 );
and ( n30835 , n30828 , n30833 );
or ( n30836 , n30831 , n30834 , n30835 );
and ( n30837 , n30806 , n30836 );
xor ( n30838 , n30745 , n30802 );
and ( n30839 , n30837 , n30838 );
xor ( n30840 , n30828 , n30830 );
xor ( n30841 , n30840 , n30833 );
buf ( n30842 , n787 );
buf ( n30843 , n30842 );
buf ( n30844 , n788 );
buf ( n30845 , n30844 );
and ( n30846 , n30843 , n30845 );
not ( n30847 , n30846 );
and ( n30848 , n30749 , n30847 );
not ( n30849 , n30848 );
and ( n30850 , n30658 , n30691 );
and ( n30851 , n30633 , n30689 );
nor ( n30852 , n30850 , n30851 );
xnor ( n30853 , n30852 , n30696 );
and ( n30854 , n30849 , n30853 );
xor ( n30855 , n30243 , n30579 );
buf ( n30856 , n30855 );
buf ( n30857 , n30856 );
buf ( n30858 , n30857 );
and ( n30859 , n30858 , n30597 );
and ( n30860 , n30853 , n30859 );
and ( n30861 , n30849 , n30859 );
or ( n30862 , n30854 , n30860 , n30861 );
and ( n30863 , n30633 , n30691 );
and ( n30864 , n30624 , n30689 );
nor ( n30865 , n30863 , n30864 );
xnor ( n30866 , n30865 , n30696 );
and ( n30867 , n30862 , n30866 );
and ( n30868 , n30762 , n30605 );
and ( n30869 , n30718 , n30603 );
nor ( n30870 , n30868 , n30869 );
xnor ( n30871 , n30870 , n30610 );
and ( n30872 , n30866 , n30871 );
and ( n30873 , n30862 , n30871 );
or ( n30874 , n30867 , n30872 , n30873 );
and ( n30875 , n30624 , n30770 );
and ( n30876 , n30595 , n30768 );
nor ( n30877 , n30875 , n30876 );
xnor ( n30878 , n30877 , n30752 );
and ( n30879 , n30718 , n30645 );
and ( n30880 , n30704 , n30643 );
nor ( n30881 , n30879 , n30880 );
xnor ( n30882 , n30881 , n30619 );
and ( n30883 , n30878 , n30882 );
and ( n30884 , n30816 , n30605 );
and ( n30885 , n30762 , n30603 );
nor ( n30886 , n30884 , n30885 );
xnor ( n30887 , n30886 , n30610 );
and ( n30888 , n30882 , n30887 );
and ( n30889 , n30878 , n30887 );
or ( n30890 , n30883 , n30888 , n30889 );
and ( n30891 , n30762 , n30645 );
and ( n30892 , n30718 , n30643 );
nor ( n30893 , n30891 , n30892 );
xnor ( n30894 , n30893 , n30619 );
and ( n30895 , n30858 , n30605 );
and ( n30896 , n30816 , n30603 );
nor ( n30897 , n30895 , n30896 );
xnor ( n30898 , n30897 , n30610 );
and ( n30899 , n30894 , n30898 );
xor ( n30900 , n30246 , n30577 );
buf ( n30901 , n30900 );
buf ( n30902 , n30901 );
buf ( n30903 , n30902 );
and ( n30904 , n30903 , n30597 );
and ( n30905 , n30898 , n30904 );
and ( n30906 , n30894 , n30904 );
or ( n30907 , n30899 , n30905 , n30906 );
xor ( n30908 , n30749 , n30843 );
xor ( n30909 , n30843 , n30845 );
not ( n30910 , n30909 );
and ( n30911 , n30908 , n30910 );
and ( n30912 , n30595 , n30911 );
not ( n30913 , n30912 );
xnor ( n30914 , n30913 , n30848 );
not ( n30915 , n30914 );
and ( n30916 , n30633 , n30770 );
and ( n30917 , n30624 , n30768 );
nor ( n30918 , n30916 , n30917 );
xnor ( n30919 , n30918 , n30752 );
and ( n30920 , n30915 , n30919 );
and ( n30921 , n30704 , n30691 );
and ( n30922 , n30658 , n30689 );
nor ( n30923 , n30921 , n30922 );
xnor ( n30924 , n30923 , n30696 );
and ( n30925 , n30919 , n30924 );
and ( n30926 , n30915 , n30924 );
or ( n30927 , n30920 , n30925 , n30926 );
and ( n30928 , n30907 , n30927 );
buf ( n30929 , n30914 );
and ( n30930 , n30927 , n30929 );
and ( n30931 , n30907 , n30929 );
or ( n30932 , n30928 , n30930 , n30931 );
and ( n30933 , n30890 , n30932 );
xor ( n30934 , n30807 , n30811 );
xor ( n30935 , n30934 , n30817 );
and ( n30936 , n30932 , n30935 );
and ( n30937 , n30890 , n30935 );
or ( n30938 , n30933 , n30936 , n30937 );
and ( n30939 , n30874 , n30938 );
xor ( n30940 , n30820 , n30822 );
xor ( n30941 , n30940 , n30825 );
and ( n30942 , n30938 , n30941 );
and ( n30943 , n30874 , n30941 );
or ( n30944 , n30939 , n30942 , n30943 );
and ( n30945 , n30841 , n30944 );
xor ( n30946 , n30806 , n30836 );
and ( n30947 , n30945 , n30946 );
xor ( n30948 , n30841 , n30944 );
xor ( n30949 , n30874 , n30938 );
xor ( n30950 , n30949 , n30941 );
buf ( n30951 , n789 );
buf ( n30952 , n30951 );
buf ( n30953 , n790 );
buf ( n30954 , n30953 );
and ( n30955 , n30952 , n30954 );
not ( n30956 , n30955 );
and ( n30957 , n30845 , n30956 );
not ( n30958 , n30957 );
and ( n30959 , n30903 , n30605 );
and ( n30960 , n30858 , n30603 );
nor ( n30961 , n30959 , n30960 );
xnor ( n30962 , n30961 , n30610 );
and ( n30963 , n30958 , n30962 );
xor ( n30964 , n30248 , n30576 );
buf ( n30965 , n30964 );
buf ( n30966 , n30965 );
buf ( n30967 , n30966 );
and ( n30968 , n30967 , n30597 );
and ( n30969 , n30962 , n30968 );
and ( n30970 , n30958 , n30968 );
or ( n30971 , n30963 , n30969 , n30970 );
xor ( n30972 , n30845 , n30952 );
xor ( n30973 , n30952 , n30954 );
not ( n30974 , n30973 );
and ( n30975 , n30972 , n30974 );
and ( n30976 , n30595 , n30975 );
not ( n30977 , n30976 );
xnor ( n30978 , n30977 , n30957 );
buf ( n30979 , n30978 );
and ( n30980 , n30624 , n30911 );
and ( n30981 , n30595 , n30909 );
nor ( n30982 , n30980 , n30981 );
xnor ( n30983 , n30982 , n30848 );
and ( n30984 , n30979 , n30983 );
and ( n30985 , n30816 , n30645 );
and ( n30986 , n30762 , n30643 );
nor ( n30987 , n30985 , n30986 );
xnor ( n30988 , n30987 , n30619 );
and ( n30989 , n30983 , n30988 );
and ( n30990 , n30979 , n30988 );
or ( n30991 , n30984 , n30989 , n30990 );
and ( n30992 , n30971 , n30991 );
xor ( n30993 , n30894 , n30898 );
xor ( n30994 , n30993 , n30904 );
and ( n30995 , n30991 , n30994 );
and ( n30996 , n30971 , n30994 );
or ( n30997 , n30992 , n30995 , n30996 );
xor ( n30998 , n30849 , n30853 );
xor ( n30999 , n30998 , n30859 );
and ( n31000 , n30997 , n30999 );
xor ( n31001 , n30878 , n30882 );
xor ( n31002 , n31001 , n30887 );
and ( n31003 , n30999 , n31002 );
and ( n31004 , n30997 , n31002 );
or ( n31005 , n31000 , n31003 , n31004 );
xor ( n31006 , n30862 , n30866 );
xor ( n31007 , n31006 , n30871 );
and ( n31008 , n31005 , n31007 );
xor ( n31009 , n30890 , n30932 );
xor ( n31010 , n31009 , n30935 );
and ( n31011 , n31007 , n31010 );
and ( n31012 , n31005 , n31010 );
or ( n31013 , n31008 , n31011 , n31012 );
and ( n31014 , n30950 , n31013 );
and ( n31015 , n30948 , n31014 );
xor ( n31016 , n30907 , n30927 );
xor ( n31017 , n31016 , n30929 );
xor ( n31018 , n30915 , n30919 );
xor ( n31019 , n31018 , n30924 );
and ( n31020 , n30658 , n30770 );
and ( n31021 , n30633 , n30768 );
nor ( n31022 , n31020 , n31021 );
xnor ( n31023 , n31022 , n30752 );
and ( n31024 , n30718 , n30691 );
and ( n31025 , n30704 , n30689 );
nor ( n31026 , n31024 , n31025 );
xnor ( n31027 , n31026 , n30696 );
and ( n31028 , n31023 , n31027 );
and ( n31029 , n31019 , n31028 );
and ( n31030 , n31017 , n31029 );
xor ( n31031 , n31005 , n31007 );
xor ( n31032 , n31031 , n31010 );
and ( n31033 , n31030 , n31032 );
xor ( n31034 , n30950 , n31013 );
and ( n31035 , n31033 , n31034 );
xor ( n31036 , n31017 , n31029 );
xor ( n31037 , n30997 , n30999 );
xor ( n31038 , n31037 , n31002 );
and ( n31039 , n31036 , n31038 );
xor ( n31040 , n31023 , n31027 );
and ( n31041 , n30858 , n30645 );
and ( n31042 , n30816 , n30643 );
nor ( n31043 , n31041 , n31042 );
xnor ( n31044 , n31043 , n30619 );
and ( n31045 , n30967 , n30605 );
and ( n31046 , n30903 , n30603 );
nor ( n31047 , n31045 , n31046 );
xnor ( n31048 , n31047 , n30610 );
and ( n31049 , n31044 , n31048 );
xor ( n31050 , n30249 , n30575 );
buf ( n31051 , n31050 );
buf ( n31052 , n31051 );
buf ( n31053 , n31052 );
and ( n31054 , n31053 , n30597 );
and ( n31055 , n31048 , n31054 );
and ( n31056 , n31044 , n31054 );
or ( n31057 , n31049 , n31055 , n31056 );
and ( n31058 , n31040 , n31057 );
xor ( n31059 , n31019 , n31028 );
and ( n31060 , n31058 , n31059 );
xor ( n31061 , n30971 , n30991 );
xor ( n31062 , n31061 , n30994 );
and ( n31063 , n31059 , n31062 );
and ( n31064 , n31058 , n31062 );
or ( n31065 , n31060 , n31063 , n31064 );
and ( n31066 , n31038 , n31065 );
and ( n31067 , n31036 , n31065 );
or ( n31068 , n31039 , n31066 , n31067 );
xor ( n31069 , n31030 , n31032 );
and ( n31070 , n31068 , n31069 );
not ( n31071 , n30978 );
and ( n31072 , n30704 , n30770 );
and ( n31073 , n30658 , n30768 );
nor ( n31074 , n31072 , n31073 );
xnor ( n31075 , n31074 , n30752 );
and ( n31076 , n31071 , n31075 );
and ( n31077 , n30762 , n30691 );
and ( n31078 , n30718 , n30689 );
nor ( n31079 , n31077 , n31078 );
xnor ( n31080 , n31079 , n30696 );
and ( n31081 , n31075 , n31080 );
and ( n31082 , n31071 , n31080 );
or ( n31083 , n31076 , n31081 , n31082 );
xor ( n31084 , n30958 , n30962 );
xor ( n31085 , n31084 , n30968 );
and ( n31086 , n31083 , n31085 );
xor ( n31087 , n30979 , n30983 );
xor ( n31088 , n31087 , n30988 );
and ( n31089 , n31085 , n31088 );
and ( n31090 , n31083 , n31088 );
or ( n31091 , n31086 , n31089 , n31090 );
xor ( n31092 , n31071 , n31075 );
xor ( n31093 , n31092 , n31080 );
and ( n31094 , n30624 , n30975 );
and ( n31095 , n30595 , n30973 );
nor ( n31096 , n31094 , n31095 );
xnor ( n31097 , n31096 , n30957 );
and ( n31098 , n30903 , n30645 );
and ( n31099 , n30858 , n30643 );
nor ( n31100 , n31098 , n31099 );
xnor ( n31101 , n31100 , n30619 );
and ( n31102 , n31097 , n31101 );
and ( n31103 , n31053 , n30605 );
and ( n31104 , n30967 , n30603 );
nor ( n31105 , n31103 , n31104 );
xnor ( n31106 , n31105 , n30610 );
and ( n31107 , n31101 , n31106 );
and ( n31108 , n31097 , n31106 );
or ( n31109 , n31102 , n31107 , n31108 );
and ( n31110 , n31093 , n31109 );
xor ( n31111 , n31040 , n31057 );
and ( n31112 , n31110 , n31111 );
xor ( n31113 , n31083 , n31085 );
xor ( n31114 , n31113 , n31088 );
and ( n31115 , n31111 , n31114 );
and ( n31116 , n31110 , n31114 );
or ( n31117 , n31112 , n31115 , n31116 );
and ( n31118 , n31091 , n31117 );
xor ( n31119 , n31058 , n31059 );
xor ( n31120 , n31119 , n31062 );
and ( n31121 , n31117 , n31120 );
and ( n31122 , n31091 , n31120 );
or ( n31123 , n31118 , n31121 , n31122 );
xor ( n31124 , n31036 , n31038 );
xor ( n31125 , n31124 , n31065 );
and ( n31126 , n31123 , n31125 );
xor ( n31127 , n31091 , n31117 );
xor ( n31128 , n31127 , n31120 );
and ( n31129 , n30658 , n30911 );
and ( n31130 , n30633 , n30909 );
nor ( n31131 , n31129 , n31130 );
xnor ( n31132 , n31131 , n30848 );
and ( n31133 , n30718 , n30770 );
and ( n31134 , n30704 , n30768 );
nor ( n31135 , n31133 , n31134 );
xnor ( n31136 , n31135 , n30752 );
and ( n31137 , n31132 , n31136 );
and ( n31138 , n30816 , n30691 );
and ( n31139 , n30762 , n30689 );
nor ( n31140 , n31138 , n31139 );
xnor ( n31141 , n31140 , n30696 );
and ( n31142 , n31136 , n31141 );
and ( n31143 , n31132 , n31141 );
or ( n31144 , n31137 , n31142 , n31143 );
buf ( n31145 , n792 );
buf ( n31146 , n31145 );
not ( n31147 , n31146 );
buf ( n31148 , n31147 );
buf ( n31149 , n31148 );
buf ( n31150 , n791 );
buf ( n31151 , n31150 );
and ( n31152 , n31151 , n31146 );
not ( n31153 , n31152 );
and ( n31154 , n30954 , n31153 );
not ( n31155 , n31154 );
and ( n31156 , n31149 , n31155 );
xor ( n31157 , n30251 , n30574 );
buf ( n31158 , n31157 );
buf ( n31159 , n31158 );
buf ( n31160 , n31159 );
and ( n31161 , n31160 , n30597 );
and ( n31162 , n31155 , n31161 );
and ( n31163 , n31149 , n31161 );
or ( n31164 , n31156 , n31162 , n31163 );
and ( n31165 , n31144 , n31164 );
and ( n31166 , n30633 , n30911 );
and ( n31167 , n30624 , n30909 );
nor ( n31168 , n31166 , n31167 );
xnor ( n31169 , n31168 , n30848 );
and ( n31170 , n31164 , n31169 );
and ( n31171 , n31144 , n31169 );
or ( n31172 , n31165 , n31170 , n31171 );
xor ( n31173 , n31110 , n31111 );
xor ( n31174 , n31173 , n31114 );
and ( n31175 , n31172 , n31174 );
and ( n31176 , n30633 , n30975 );
and ( n31177 , n30624 , n30973 );
nor ( n31178 , n31176 , n31177 );
xnor ( n31179 , n31178 , n30957 );
and ( n31180 , n30704 , n30911 );
and ( n31181 , n30658 , n30909 );
nor ( n31182 , n31180 , n31181 );
xnor ( n31183 , n31182 , n30848 );
and ( n31184 , n31179 , n31183 );
and ( n31185 , n30762 , n30770 );
and ( n31186 , n30718 , n30768 );
nor ( n31187 , n31185 , n31186 );
xnor ( n31188 , n31187 , n30752 );
and ( n31189 , n31183 , n31188 );
and ( n31190 , n31179 , n31188 );
or ( n31191 , n31184 , n31189 , n31190 );
xor ( n31192 , n31097 , n31101 );
xor ( n31193 , n31192 , n31106 );
and ( n31194 , n31191 , n31193 );
xor ( n31195 , n31132 , n31136 );
xor ( n31196 , n31195 , n31141 );
and ( n31197 , n31193 , n31196 );
and ( n31198 , n31191 , n31196 );
or ( n31199 , n31194 , n31197 , n31198 );
and ( n31200 , n30858 , n30691 );
and ( n31201 , n30816 , n30689 );
nor ( n31202 , n31200 , n31201 );
xnor ( n31203 , n31202 , n30696 );
and ( n31204 , n30967 , n30645 );
and ( n31205 , n30903 , n30643 );
nor ( n31206 , n31204 , n31205 );
xnor ( n31207 , n31206 , n30619 );
and ( n31208 , n31203 , n31207 );
and ( n31209 , n31160 , n30605 );
and ( n31210 , n31053 , n30603 );
nor ( n31211 , n31209 , n31210 );
xnor ( n31212 , n31211 , n30610 );
and ( n31213 , n31207 , n31212 );
and ( n31214 , n31203 , n31212 );
or ( n31215 , n31208 , n31213 , n31214 );
not ( n31216 , n31148 );
xor ( n31217 , n30954 , n31151 );
xor ( n31218 , n31151 , n31146 );
not ( n31219 , n31218 );
and ( n31220 , n31217 , n31219 );
and ( n31221 , n30595 , n31220 );
not ( n31222 , n31221 );
xnor ( n31223 , n31222 , n31154 );
and ( n31224 , n31216 , n31223 );
xor ( n31225 , n30254 , n30572 );
buf ( n31226 , n31225 );
buf ( n31227 , n31226 );
buf ( n31228 , n31227 );
and ( n31229 , n31228 , n30597 );
and ( n31230 , n31223 , n31229 );
and ( n31231 , n31216 , n31229 );
or ( n31232 , n31224 , n31230 , n31231 );
and ( n31233 , n31215 , n31232 );
xor ( n31234 , n31149 , n31155 );
xor ( n31235 , n31234 , n31161 );
and ( n31236 , n31232 , n31235 );
and ( n31237 , n31215 , n31235 );
or ( n31238 , n31233 , n31236 , n31237 );
and ( n31239 , n31199 , n31238 );
xor ( n31240 , n31144 , n31164 );
xor ( n31241 , n31240 , n31169 );
and ( n31242 , n31238 , n31241 );
and ( n31243 , n31199 , n31241 );
or ( n31244 , n31239 , n31242 , n31243 );
and ( n31245 , n31174 , n31244 );
and ( n31246 , n31172 , n31244 );
or ( n31247 , n31175 , n31245 , n31246 );
and ( n31248 , n31128 , n31247 );
xor ( n31249 , n31044 , n31048 );
xor ( n31250 , n31249 , n31054 );
xor ( n31251 , n31093 , n31109 );
and ( n31252 , n31250 , n31251 );
xor ( n31253 , n31199 , n31238 );
xor ( n31254 , n31253 , n31241 );
and ( n31255 , n31251 , n31254 );
and ( n31256 , n31250 , n31254 );
or ( n31257 , n31252 , n31255 , n31256 );
xor ( n31258 , n31172 , n31174 );
xor ( n31259 , n31258 , n31244 );
and ( n31260 , n31257 , n31259 );
and ( n31261 , n30718 , n30911 );
and ( n31262 , n30704 , n30909 );
nor ( n31263 , n31261 , n31262 );
xnor ( n31264 , n31263 , n30848 );
and ( n31265 , n30903 , n30691 );
and ( n31266 , n30858 , n30689 );
nor ( n31267 , n31265 , n31266 );
xnor ( n31268 , n31267 , n30696 );
and ( n31269 , n31264 , n31268 );
and ( n31270 , n31053 , n30645 );
and ( n31271 , n30967 , n30643 );
nor ( n31272 , n31270 , n31271 );
xnor ( n31273 , n31272 , n30619 );
and ( n31274 , n31268 , n31273 );
and ( n31275 , n31264 , n31273 );
or ( n31276 , n31269 , n31274 , n31275 );
and ( n31277 , n30624 , n31220 );
and ( n31278 , n30595 , n31218 );
nor ( n31279 , n31277 , n31278 );
xnor ( n31280 , n31279 , n31154 );
and ( n31281 , n30658 , n30975 );
and ( n31282 , n30633 , n30973 );
nor ( n31283 , n31281 , n31282 );
xnor ( n31284 , n31283 , n30957 );
and ( n31285 , n31280 , n31284 );
and ( n31286 , n30816 , n30770 );
and ( n31287 , n30762 , n30768 );
nor ( n31288 , n31286 , n31287 );
xnor ( n31289 , n31288 , n30752 );
and ( n31290 , n31284 , n31289 );
and ( n31291 , n31280 , n31289 );
or ( n31292 , n31285 , n31290 , n31291 );
and ( n31293 , n31276 , n31292 );
xor ( n31294 , n31179 , n31183 );
xor ( n31295 , n31294 , n31188 );
and ( n31296 , n31292 , n31295 );
and ( n31297 , n31276 , n31295 );
or ( n31298 , n31293 , n31296 , n31297 );
and ( n31299 , n31228 , n30605 );
and ( n31300 , n31160 , n30603 );
nor ( n31301 , n31299 , n31300 );
xnor ( n31302 , n31301 , n30610 );
and ( n31303 , n31146 , n31302 );
xor ( n31304 , n30257 , n30570 );
buf ( n31305 , n31304 );
buf ( n31306 , n31305 );
buf ( n31307 , n31306 );
and ( n31308 , n31307 , n30597 );
and ( n31309 , n31302 , n31308 );
and ( n31310 , n31146 , n31308 );
or ( n31311 , n31303 , n31309 , n31310 );
xor ( n31312 , n31203 , n31207 );
xor ( n31313 , n31312 , n31212 );
and ( n31314 , n31311 , n31313 );
xor ( n31315 , n31216 , n31223 );
xor ( n31316 , n31315 , n31229 );
and ( n31317 , n31313 , n31316 );
and ( n31318 , n31311 , n31316 );
or ( n31319 , n31314 , n31317 , n31318 );
and ( n31320 , n31298 , n31319 );
xor ( n31321 , n31215 , n31232 );
xor ( n31322 , n31321 , n31235 );
and ( n31323 , n31319 , n31322 );
and ( n31324 , n31298 , n31322 );
or ( n31325 , n31320 , n31323 , n31324 );
and ( n31326 , n30633 , n31220 );
and ( n31327 , n30624 , n31218 );
nor ( n31328 , n31326 , n31327 );
xnor ( n31329 , n31328 , n31154 );
and ( n31330 , n30704 , n30975 );
and ( n31331 , n30658 , n30973 );
nor ( n31332 , n31330 , n31331 );
xnor ( n31333 , n31332 , n30957 );
and ( n31334 , n31329 , n31333 );
and ( n31335 , n30762 , n30911 );
and ( n31336 , n30718 , n30909 );
nor ( n31337 , n31335 , n31336 );
xnor ( n31338 , n31337 , n30848 );
and ( n31339 , n31333 , n31338 );
and ( n31340 , n31329 , n31338 );
or ( n31341 , n31334 , n31339 , n31340 );
xor ( n31342 , n31264 , n31268 );
xor ( n31343 , n31342 , n31273 );
and ( n31344 , n31341 , n31343 );
xor ( n31345 , n31280 , n31284 );
xor ( n31346 , n31345 , n31289 );
and ( n31347 , n31343 , n31346 );
and ( n31348 , n31341 , n31346 );
or ( n31349 , n31344 , n31347 , n31348 );
buf ( n31350 , n793 );
buf ( n31351 , n31350 );
xor ( n31352 , n31146 , n31351 );
not ( n31353 , n31351 );
and ( n31354 , n31352 , n31353 );
and ( n31355 , n30595 , n31354 );
not ( n31356 , n31355 );
xnor ( n31357 , n31356 , n31146 );
and ( n31358 , n31307 , n30605 );
and ( n31359 , n31228 , n30603 );
nor ( n31360 , n31358 , n31359 );
xnor ( n31361 , n31360 , n30610 );
and ( n31362 , n31357 , n31361 );
xor ( n31363 , n30258 , n30569 );
buf ( n31364 , n31363 );
buf ( n31365 , n31364 );
buf ( n31366 , n31365 );
and ( n31367 , n31366 , n30597 );
and ( n31368 , n31361 , n31367 );
and ( n31369 , n31357 , n31367 );
or ( n31370 , n31362 , n31368 , n31369 );
and ( n31371 , n30858 , n30770 );
and ( n31372 , n30816 , n30768 );
nor ( n31373 , n31371 , n31372 );
xnor ( n31374 , n31373 , n30752 );
and ( n31375 , n30967 , n30691 );
and ( n31376 , n30903 , n30689 );
nor ( n31377 , n31375 , n31376 );
xnor ( n31378 , n31377 , n30696 );
and ( n31379 , n31374 , n31378 );
and ( n31380 , n31160 , n30645 );
and ( n31381 , n31053 , n30643 );
nor ( n31382 , n31380 , n31381 );
xnor ( n31383 , n31382 , n30619 );
and ( n31384 , n31378 , n31383 );
and ( n31385 , n31374 , n31383 );
or ( n31386 , n31379 , n31384 , n31385 );
and ( n31387 , n31370 , n31386 );
xor ( n31388 , n31146 , n31302 );
xor ( n31389 , n31388 , n31308 );
and ( n31390 , n31386 , n31389 );
and ( n31391 , n31370 , n31389 );
or ( n31392 , n31387 , n31390 , n31391 );
and ( n31393 , n31349 , n31392 );
xor ( n31394 , n31311 , n31313 );
xor ( n31395 , n31394 , n31316 );
and ( n31396 , n31392 , n31395 );
and ( n31397 , n31349 , n31395 );
or ( n31398 , n31393 , n31396 , n31397 );
xor ( n31399 , n31191 , n31193 );
xor ( n31400 , n31399 , n31196 );
and ( n31401 , n31398 , n31400 );
xor ( n31402 , n31298 , n31319 );
xor ( n31403 , n31402 , n31322 );
and ( n31404 , n31400 , n31403 );
and ( n31405 , n31398 , n31403 );
or ( n31406 , n31401 , n31404 , n31405 );
and ( n31407 , n31325 , n31406 );
xor ( n31408 , n31250 , n31251 );
xor ( n31409 , n31408 , n31254 );
and ( n31410 , n31406 , n31409 );
and ( n31411 , n31325 , n31409 );
or ( n31412 , n31407 , n31410 , n31411 );
and ( n31413 , n31259 , n31412 );
and ( n31414 , n31257 , n31412 );
or ( n31415 , n31260 , n31413 , n31414 );
and ( n31416 , n31247 , n31415 );
and ( n31417 , n31128 , n31415 );
or ( n31418 , n31248 , n31416 , n31417 );
and ( n31419 , n31125 , n31418 );
and ( n31420 , n31123 , n31418 );
or ( n31421 , n31126 , n31419 , n31420 );
and ( n31422 , n31069 , n31421 );
and ( n31423 , n31068 , n31421 );
or ( n31424 , n31070 , n31422 , n31423 );
and ( n31425 , n31034 , n31424 );
and ( n31426 , n31033 , n31424 );
or ( n31427 , n31035 , n31425 , n31426 );
and ( n31428 , n31014 , n31427 );
and ( n31429 , n30948 , n31427 );
or ( n31430 , n31015 , n31428 , n31429 );
and ( n31431 , n30946 , n31430 );
and ( n31432 , n30945 , n31430 );
or ( n31433 , n30947 , n31431 , n31432 );
and ( n31434 , n30838 , n31433 );
and ( n31435 , n30837 , n31433 );
or ( n31436 , n30839 , n31434 , n31435 );
and ( n31437 , n30803 , n31436 );
and ( n31438 , n30743 , n31436 );
or ( n31439 , n30804 , n31437 , n31438 );
and ( n31440 , n30741 , n31439 );
and ( n31441 , n30681 , n31439 );
or ( n31442 , n30742 , n31440 , n31441 );
xor ( n31443 , n30680 , n31442 );
xor ( n31444 , n30681 , n30741 );
xor ( n31445 , n31444 , n31439 );
xor ( n31446 , n30743 , n30803 );
xor ( n31447 , n31446 , n31436 );
xor ( n31448 , n30837 , n30838 );
xor ( n31449 , n31448 , n31433 );
xor ( n31450 , n30945 , n30946 );
xor ( n31451 , n31450 , n31430 );
xor ( n31452 , n30948 , n31014 );
xor ( n31453 , n31452 , n31427 );
xor ( n31454 , n31033 , n31034 );
xor ( n31455 , n31454 , n31424 );
xor ( n31456 , n31068 , n31069 );
xor ( n31457 , n31456 , n31421 );
xor ( n31458 , n31123 , n31125 );
xor ( n31459 , n31458 , n31418 );
xor ( n31460 , n31128 , n31247 );
xor ( n31461 , n31460 , n31415 );
xor ( n31462 , n31257 , n31259 );
xor ( n31463 , n31462 , n31412 );
and ( n31464 , n31228 , n30645 );
and ( n31465 , n31160 , n30643 );
nor ( n31466 , n31464 , n31465 );
xnor ( n31467 , n31466 , n30619 );
and ( n31468 , n31366 , n30605 );
and ( n31469 , n31307 , n30603 );
nor ( n31470 , n31468 , n31469 );
xnor ( n31471 , n31470 , n30610 );
and ( n31472 , n31467 , n31471 );
xor ( n31473 , n30259 , n30568 );
buf ( n31474 , n31473 );
buf ( n31475 , n31474 );
buf ( n31476 , n31475 );
and ( n31477 , n31476 , n30597 );
and ( n31478 , n31471 , n31477 );
and ( n31479 , n31467 , n31477 );
or ( n31480 , n31472 , n31478 , n31479 );
xor ( n31481 , n31357 , n31361 );
xor ( n31482 , n31481 , n31367 );
and ( n31483 , n31480 , n31482 );
xor ( n31484 , n31374 , n31378 );
xor ( n31485 , n31484 , n31383 );
and ( n31486 , n31482 , n31485 );
and ( n31487 , n31480 , n31485 );
or ( n31488 , n31483 , n31486 , n31487 );
and ( n31489 , n30658 , n31220 );
and ( n31490 , n30633 , n31218 );
nor ( n31491 , n31489 , n31490 );
xnor ( n31492 , n31491 , n31154 );
and ( n31493 , n30903 , n30770 );
and ( n31494 , n30858 , n30768 );
nor ( n31495 , n31493 , n31494 );
xnor ( n31496 , n31495 , n30752 );
and ( n31497 , n31492 , n31496 );
and ( n31498 , n31053 , n30691 );
and ( n31499 , n30967 , n30689 );
nor ( n31500 , n31498 , n31499 );
xnor ( n31501 , n31500 , n30696 );
and ( n31502 , n31496 , n31501 );
and ( n31503 , n31492 , n31501 );
or ( n31504 , n31497 , n31502 , n31503 );
and ( n31505 , n30624 , n31354 );
and ( n31506 , n30595 , n31351 );
nor ( n31507 , n31505 , n31506 );
xnor ( n31508 , n31507 , n31146 );
and ( n31509 , n30718 , n30975 );
and ( n31510 , n30704 , n30973 );
nor ( n31511 , n31509 , n31510 );
xnor ( n31512 , n31511 , n30957 );
and ( n31513 , n31508 , n31512 );
and ( n31514 , n30816 , n30911 );
and ( n31515 , n30762 , n30909 );
nor ( n31516 , n31514 , n31515 );
xnor ( n31517 , n31516 , n30848 );
and ( n31518 , n31512 , n31517 );
and ( n31519 , n31508 , n31517 );
or ( n31520 , n31513 , n31518 , n31519 );
and ( n31521 , n31504 , n31520 );
xor ( n31522 , n31329 , n31333 );
xor ( n31523 , n31522 , n31338 );
and ( n31524 , n31520 , n31523 );
and ( n31525 , n31504 , n31523 );
or ( n31526 , n31521 , n31524 , n31525 );
and ( n31527 , n31488 , n31526 );
xor ( n31528 , n31370 , n31386 );
xor ( n31529 , n31528 , n31389 );
and ( n31530 , n31526 , n31529 );
and ( n31531 , n31488 , n31529 );
or ( n31532 , n31527 , n31530 , n31531 );
xor ( n31533 , n31276 , n31292 );
xor ( n31534 , n31533 , n31295 );
and ( n31535 , n31532 , n31534 );
xor ( n31536 , n31349 , n31392 );
xor ( n31537 , n31536 , n31395 );
and ( n31538 , n31534 , n31537 );
and ( n31539 , n31532 , n31537 );
or ( n31540 , n31535 , n31538 , n31539 );
xor ( n31541 , n31398 , n31400 );
xor ( n31542 , n31541 , n31403 );
and ( n31543 , n31540 , n31542 );
xor ( n31544 , n31325 , n31406 );
xor ( n31545 , n31544 , n31409 );
and ( n31546 , n31543 , n31545 );
xor ( n31547 , n31543 , n31545 );
and ( n31548 , n31307 , n30645 );
and ( n31549 , n31228 , n30643 );
nor ( n31550 , n31548 , n31549 );
xnor ( n31551 , n31550 , n30619 );
and ( n31552 , n31476 , n30605 );
and ( n31553 , n31366 , n30603 );
nor ( n31554 , n31552 , n31553 );
xnor ( n31555 , n31554 , n30610 );
and ( n31556 , n31551 , n31555 );
xor ( n31557 , n30262 , n30566 );
buf ( n31558 , n31557 );
buf ( n31559 , n31558 );
buf ( n31560 , n31559 );
and ( n31561 , n31560 , n30597 );
and ( n31562 , n31555 , n31561 );
and ( n31563 , n31551 , n31561 );
or ( n31564 , n31556 , n31562 , n31563 );
and ( n31565 , n30858 , n30911 );
and ( n31566 , n30816 , n30909 );
nor ( n31567 , n31565 , n31566 );
xnor ( n31568 , n31567 , n30848 );
and ( n31569 , n30967 , n30770 );
and ( n31570 , n30903 , n30768 );
nor ( n31571 , n31569 , n31570 );
xnor ( n31572 , n31571 , n30752 );
and ( n31573 , n31568 , n31572 );
and ( n31574 , n31160 , n30691 );
and ( n31575 , n31053 , n30689 );
nor ( n31576 , n31574 , n31575 );
xnor ( n31577 , n31576 , n30696 );
and ( n31578 , n31572 , n31577 );
and ( n31579 , n31568 , n31577 );
or ( n31580 , n31573 , n31578 , n31579 );
and ( n31581 , n31564 , n31580 );
xor ( n31582 , n31467 , n31471 );
xor ( n31583 , n31582 , n31477 );
and ( n31584 , n31580 , n31583 );
and ( n31585 , n31564 , n31583 );
or ( n31586 , n31581 , n31584 , n31585 );
and ( n31587 , n30633 , n31354 );
and ( n31588 , n30624 , n31351 );
nor ( n31589 , n31587 , n31588 );
xnor ( n31590 , n31589 , n31146 );
and ( n31591 , n30704 , n31220 );
and ( n31592 , n30658 , n31218 );
nor ( n31593 , n31591 , n31592 );
xnor ( n31594 , n31593 , n31154 );
and ( n31595 , n31590 , n31594 );
and ( n31596 , n30762 , n30975 );
and ( n31597 , n30718 , n30973 );
nor ( n31598 , n31596 , n31597 );
xnor ( n31599 , n31598 , n30957 );
and ( n31600 , n31594 , n31599 );
and ( n31601 , n31590 , n31599 );
or ( n31602 , n31595 , n31600 , n31601 );
xor ( n31603 , n31492 , n31496 );
xor ( n31604 , n31603 , n31501 );
and ( n31605 , n31602 , n31604 );
xor ( n31606 , n31508 , n31512 );
xor ( n31607 , n31606 , n31517 );
and ( n31608 , n31604 , n31607 );
and ( n31609 , n31602 , n31607 );
or ( n31610 , n31605 , n31608 , n31609 );
and ( n31611 , n31586 , n31610 );
xor ( n31612 , n31480 , n31482 );
xor ( n31613 , n31612 , n31485 );
and ( n31614 , n31610 , n31613 );
and ( n31615 , n31586 , n31613 );
or ( n31616 , n31611 , n31614 , n31615 );
xor ( n31617 , n31341 , n31343 );
xor ( n31618 , n31617 , n31346 );
and ( n31619 , n31616 , n31618 );
xor ( n31620 , n31488 , n31526 );
xor ( n31621 , n31620 , n31529 );
and ( n31622 , n31618 , n31621 );
and ( n31623 , n31616 , n31621 );
or ( n31624 , n31619 , n31622 , n31623 );
xor ( n31625 , n31532 , n31534 );
xor ( n31626 , n31625 , n31537 );
and ( n31627 , n31624 , n31626 );
xor ( n31628 , n31540 , n31542 );
and ( n31629 , n31627 , n31628 );
xor ( n31630 , n31627 , n31628 );
xor ( n31631 , n31616 , n31618 );
xor ( n31632 , n31631 , n31621 );
and ( n31633 , n31228 , n30691 );
and ( n31634 , n31160 , n30689 );
nor ( n31635 , n31633 , n31634 );
xnor ( n31636 , n31635 , n30696 );
and ( n31637 , n31560 , n30605 );
and ( n31638 , n31476 , n30603 );
nor ( n31639 , n31637 , n31638 );
xnor ( n31640 , n31639 , n30610 );
and ( n31641 , n31636 , n31640 );
xor ( n31642 , n30513 , n30564 );
buf ( n31643 , n31642 );
buf ( n31644 , n31643 );
buf ( n31645 , n31644 );
and ( n31646 , n31645 , n30597 );
and ( n31647 , n31640 , n31646 );
and ( n31648 , n31636 , n31646 );
or ( n31649 , n31641 , n31647 , n31648 );
and ( n31650 , n30903 , n30911 );
and ( n31651 , n30858 , n30909 );
nor ( n31652 , n31650 , n31651 );
xnor ( n31653 , n31652 , n30848 );
and ( n31654 , n31053 , n30770 );
and ( n31655 , n30967 , n30768 );
nor ( n31656 , n31654 , n31655 );
xnor ( n31657 , n31656 , n30752 );
and ( n31658 , n31653 , n31657 );
and ( n31659 , n31366 , n30645 );
and ( n31660 , n31307 , n30643 );
nor ( n31661 , n31659 , n31660 );
xnor ( n31662 , n31661 , n30619 );
and ( n31663 , n31657 , n31662 );
and ( n31664 , n31653 , n31662 );
or ( n31665 , n31658 , n31663 , n31664 );
and ( n31666 , n31649 , n31665 );
xor ( n31667 , n31551 , n31555 );
xor ( n31668 , n31667 , n31561 );
and ( n31669 , n31665 , n31668 );
and ( n31670 , n31649 , n31668 );
or ( n31671 , n31666 , n31669 , n31670 );
and ( n31672 , n31476 , n30645 );
and ( n31673 , n31366 , n30643 );
nor ( n31674 , n31672 , n31673 );
xnor ( n31675 , n31674 , n30619 );
and ( n31676 , n31645 , n30605 );
and ( n31677 , n31560 , n30603 );
nor ( n31678 , n31676 , n31677 );
xnor ( n31679 , n31678 , n30610 );
and ( n31680 , n31675 , n31679 );
xor ( n31681 , n30516 , n30562 );
buf ( n31682 , n31681 );
buf ( n31683 , n31682 );
buf ( n31684 , n31683 );
and ( n31685 , n31684 , n30597 );
and ( n31686 , n31679 , n31685 );
and ( n31687 , n31675 , n31685 );
or ( n31688 , n31680 , n31686 , n31687 );
and ( n31689 , n30718 , n31220 );
and ( n31690 , n30704 , n31218 );
nor ( n31691 , n31689 , n31690 );
xnor ( n31692 , n31691 , n31154 );
and ( n31693 , n31688 , n31692 );
and ( n31694 , n30816 , n30975 );
and ( n31695 , n30762 , n30973 );
nor ( n31696 , n31694 , n31695 );
xnor ( n31697 , n31696 , n30957 );
and ( n31698 , n31692 , n31697 );
and ( n31699 , n31688 , n31697 );
or ( n31700 , n31693 , n31698 , n31699 );
xor ( n31701 , n31568 , n31572 );
xor ( n31702 , n31701 , n31577 );
and ( n31703 , n31700 , n31702 );
xor ( n31704 , n31590 , n31594 );
xor ( n31705 , n31704 , n31599 );
and ( n31706 , n31702 , n31705 );
and ( n31707 , n31700 , n31705 );
or ( n31708 , n31703 , n31706 , n31707 );
and ( n31709 , n31671 , n31708 );
xor ( n31710 , n31564 , n31580 );
xor ( n31711 , n31710 , n31583 );
and ( n31712 , n31708 , n31711 );
and ( n31713 , n31671 , n31711 );
or ( n31714 , n31709 , n31712 , n31713 );
xor ( n31715 , n31504 , n31520 );
xor ( n31716 , n31715 , n31523 );
and ( n31717 , n31714 , n31716 );
xor ( n31718 , n31586 , n31610 );
xor ( n31719 , n31718 , n31613 );
and ( n31720 , n31716 , n31719 );
and ( n31721 , n31714 , n31719 );
or ( n31722 , n31717 , n31720 , n31721 );
and ( n31723 , n31632 , n31722 );
xor ( n31724 , n31624 , n31626 );
and ( n31725 , n31723 , n31724 );
xor ( n31726 , n31723 , n31724 );
xor ( n31727 , n31714 , n31716 );
xor ( n31728 , n31727 , n31719 );
and ( n31729 , n31560 , n30645 );
and ( n31730 , n31476 , n30643 );
nor ( n31731 , n31729 , n31730 );
xnor ( n31732 , n31731 , n30619 );
and ( n31733 , n31684 , n30605 );
and ( n31734 , n31645 , n30603 );
nor ( n31735 , n31733 , n31734 );
xnor ( n31736 , n31735 , n30610 );
and ( n31737 , n31732 , n31736 );
xor ( n31738 , n30517 , n30561 );
buf ( n31739 , n31738 );
buf ( n31740 , n31739 );
buf ( n31741 , n31740 );
and ( n31742 , n31741 , n30597 );
and ( n31743 , n31736 , n31742 );
and ( n31744 , n31732 , n31742 );
or ( n31745 , n31737 , n31743 , n31744 );
and ( n31746 , n30858 , n30975 );
and ( n31747 , n30816 , n30973 );
nor ( n31748 , n31746 , n31747 );
xnor ( n31749 , n31748 , n30957 );
and ( n31750 , n31745 , n31749 );
and ( n31751 , n31307 , n30691 );
and ( n31752 , n31228 , n30689 );
nor ( n31753 , n31751 , n31752 );
xnor ( n31754 , n31753 , n30696 );
and ( n31755 , n31749 , n31754 );
and ( n31756 , n31745 , n31754 );
or ( n31757 , n31750 , n31755 , n31756 );
and ( n31758 , n30658 , n31354 );
and ( n31759 , n30633 , n31351 );
nor ( n31760 , n31758 , n31759 );
xnor ( n31761 , n31760 , n31146 );
and ( n31762 , n31757 , n31761 );
xor ( n31763 , n31636 , n31640 );
xor ( n31764 , n31763 , n31646 );
and ( n31765 , n31761 , n31764 );
and ( n31766 , n31757 , n31764 );
or ( n31767 , n31762 , n31765 , n31766 );
and ( n31768 , n30967 , n30911 );
and ( n31769 , n30903 , n30909 );
nor ( n31770 , n31768 , n31769 );
xnor ( n31771 , n31770 , n30848 );
and ( n31772 , n31160 , n30770 );
and ( n31773 , n31053 , n30768 );
nor ( n31774 , n31772 , n31773 );
xnor ( n31775 , n31774 , n30752 );
and ( n31776 , n31771 , n31775 );
xor ( n31777 , n31675 , n31679 );
xor ( n31778 , n31777 , n31685 );
and ( n31779 , n31775 , n31778 );
and ( n31780 , n31771 , n31778 );
or ( n31781 , n31776 , n31779 , n31780 );
xor ( n31782 , n31653 , n31657 );
xor ( n31783 , n31782 , n31662 );
and ( n31784 , n31781 , n31783 );
xor ( n31785 , n31688 , n31692 );
xor ( n31786 , n31785 , n31697 );
and ( n31787 , n31783 , n31786 );
and ( n31788 , n31781 , n31786 );
or ( n31789 , n31784 , n31787 , n31788 );
and ( n31790 , n31767 , n31789 );
xor ( n31791 , n31649 , n31665 );
xor ( n31792 , n31791 , n31668 );
and ( n31793 , n31789 , n31792 );
and ( n31794 , n31767 , n31792 );
or ( n31795 , n31790 , n31793 , n31794 );
xor ( n31796 , n31602 , n31604 );
xor ( n31797 , n31796 , n31607 );
and ( n31798 , n31795 , n31797 );
xor ( n31799 , n31671 , n31708 );
xor ( n31800 , n31799 , n31711 );
and ( n31801 , n31797 , n31800 );
and ( n31802 , n31795 , n31800 );
or ( n31803 , n31798 , n31801 , n31802 );
and ( n31804 , n31728 , n31803 );
xor ( n31805 , n31632 , n31722 );
and ( n31806 , n31804 , n31805 );
xor ( n31807 , n31804 , n31805 );
xor ( n31808 , n31728 , n31803 );
xor ( n31809 , n31795 , n31797 );
xor ( n31810 , n31809 , n31800 );
and ( n31811 , n31645 , n30645 );
and ( n31812 , n31560 , n30643 );
nor ( n31813 , n31811 , n31812 );
xnor ( n31814 , n31813 , n30619 );
and ( n31815 , n31741 , n30605 );
and ( n31816 , n31684 , n30603 );
nor ( n31817 , n31815 , n31816 );
xnor ( n31818 , n31817 , n30610 );
and ( n31819 , n31814 , n31818 );
xor ( n31820 , n30518 , n30560 );
buf ( n31821 , n31820 );
buf ( n31822 , n31821 );
buf ( n31823 , n31822 );
and ( n31824 , n31823 , n30597 );
and ( n31825 , n31818 , n31824 );
and ( n31826 , n31814 , n31824 );
or ( n31827 , n31819 , n31825 , n31826 );
and ( n31828 , n31228 , n30770 );
and ( n31829 , n31160 , n30768 );
nor ( n31830 , n31828 , n31829 );
xnor ( n31831 , n31830 , n30752 );
and ( n31832 , n31827 , n31831 );
and ( n31833 , n31366 , n30691 );
and ( n31834 , n31307 , n30689 );
nor ( n31835 , n31833 , n31834 );
xnor ( n31836 , n31835 , n30696 );
and ( n31837 , n31831 , n31836 );
and ( n31838 , n31827 , n31836 );
or ( n31839 , n31832 , n31837 , n31838 );
and ( n31840 , n30704 , n31354 );
and ( n31841 , n30658 , n31351 );
nor ( n31842 , n31840 , n31841 );
xnor ( n31843 , n31842 , n31146 );
and ( n31844 , n31839 , n31843 );
and ( n31845 , n30762 , n31220 );
and ( n31846 , n30718 , n31218 );
nor ( n31847 , n31845 , n31846 );
xnor ( n31848 , n31847 , n31154 );
and ( n31849 , n31843 , n31848 );
and ( n31850 , n31839 , n31848 );
or ( n31851 , n31844 , n31849 , n31850 );
and ( n31852 , n31684 , n30645 );
and ( n31853 , n31645 , n30643 );
nor ( n31854 , n31852 , n31853 );
xnor ( n31855 , n31854 , n30619 );
and ( n31856 , n31823 , n30605 );
and ( n31857 , n31741 , n30603 );
nor ( n31858 , n31856 , n31857 );
xnor ( n31859 , n31858 , n30610 );
and ( n31860 , n31855 , n31859 );
xor ( n31861 , n30519 , n30559 );
buf ( n31862 , n31861 );
buf ( n31863 , n31862 );
buf ( n31864 , n31863 );
and ( n31865 , n31864 , n30597 );
and ( n31866 , n31859 , n31865 );
and ( n31867 , n31855 , n31865 );
or ( n31868 , n31860 , n31866 , n31867 );
and ( n31869 , n31476 , n30691 );
and ( n31870 , n31366 , n30689 );
nor ( n31871 , n31869 , n31870 );
xnor ( n31872 , n31871 , n30696 );
and ( n31873 , n31868 , n31872 );
xor ( n31874 , n31814 , n31818 );
xor ( n31875 , n31874 , n31824 );
and ( n31876 , n31872 , n31875 );
and ( n31877 , n31868 , n31875 );
or ( n31878 , n31873 , n31876 , n31877 );
and ( n31879 , n30718 , n31354 );
and ( n31880 , n30704 , n31351 );
nor ( n31881 , n31879 , n31880 );
xnor ( n31882 , n31881 , n31146 );
and ( n31883 , n31878 , n31882 );
and ( n31884 , n30816 , n31220 );
and ( n31885 , n30762 , n31218 );
nor ( n31886 , n31884 , n31885 );
xnor ( n31887 , n31886 , n31154 );
and ( n31888 , n31882 , n31887 );
and ( n31889 , n31878 , n31887 );
or ( n31890 , n31883 , n31888 , n31889 );
and ( n31891 , n30903 , n30975 );
and ( n31892 , n30858 , n30973 );
nor ( n31893 , n31891 , n31892 );
xnor ( n31894 , n31893 , n30957 );
and ( n31895 , n31053 , n30911 );
and ( n31896 , n30967 , n30909 );
nor ( n31897 , n31895 , n31896 );
xnor ( n31898 , n31897 , n30848 );
and ( n31899 , n31894 , n31898 );
xor ( n31900 , n31732 , n31736 );
xor ( n31901 , n31900 , n31742 );
and ( n31902 , n31898 , n31901 );
and ( n31903 , n31894 , n31901 );
or ( n31904 , n31899 , n31902 , n31903 );
and ( n31905 , n31890 , n31904 );
xor ( n31906 , n31745 , n31749 );
xor ( n31907 , n31906 , n31754 );
and ( n31908 , n31904 , n31907 );
and ( n31909 , n31890 , n31907 );
or ( n31910 , n31905 , n31908 , n31909 );
and ( n31911 , n31851 , n31910 );
xor ( n31912 , n31757 , n31761 );
xor ( n31913 , n31912 , n31764 );
and ( n31914 , n31910 , n31913 );
and ( n31915 , n31851 , n31913 );
or ( n31916 , n31911 , n31914 , n31915 );
xor ( n31917 , n31700 , n31702 );
xor ( n31918 , n31917 , n31705 );
and ( n31919 , n31916 , n31918 );
xor ( n31920 , n31767 , n31789 );
xor ( n31921 , n31920 , n31792 );
and ( n31922 , n31918 , n31921 );
and ( n31923 , n31916 , n31921 );
or ( n31924 , n31919 , n31922 , n31923 );
and ( n31925 , n31810 , n31924 );
and ( n31926 , n31808 , n31925 );
xor ( n31927 , n31808 , n31925 );
xor ( n31928 , n31916 , n31918 );
xor ( n31929 , n31928 , n31921 );
xor ( n31930 , n31839 , n31843 );
xor ( n31931 , n31930 , n31848 );
xor ( n31932 , n31771 , n31775 );
xor ( n31933 , n31932 , n31778 );
and ( n31934 , n31931 , n31933 );
xor ( n31935 , n31890 , n31904 );
xor ( n31936 , n31935 , n31907 );
and ( n31937 , n31933 , n31936 );
and ( n31938 , n31931 , n31936 );
or ( n31939 , n31934 , n31937 , n31938 );
xor ( n31940 , n31781 , n31783 );
xor ( n31941 , n31940 , n31786 );
and ( n31942 , n31939 , n31941 );
xor ( n31943 , n31851 , n31910 );
xor ( n31944 , n31943 , n31913 );
and ( n31945 , n31941 , n31944 );
and ( n31946 , n31939 , n31944 );
or ( n31947 , n31942 , n31945 , n31946 );
and ( n31948 , n31929 , n31947 );
xor ( n31949 , n31810 , n31924 );
and ( n31950 , n31948 , n31949 );
xor ( n31951 , n31948 , n31949 );
xor ( n31952 , n31939 , n31941 );
xor ( n31953 , n31952 , n31944 );
and ( n31954 , n31741 , n30645 );
and ( n31955 , n31684 , n30643 );
nor ( n31956 , n31954 , n31955 );
xnor ( n31957 , n31956 , n30619 );
and ( n31958 , n31864 , n30605 );
and ( n31959 , n31823 , n30603 );
nor ( n31960 , n31958 , n31959 );
xnor ( n31961 , n31960 , n30610 );
and ( n31962 , n31957 , n31961 );
xor ( n31963 , n30522 , n30557 );
buf ( n31964 , n31963 );
buf ( n31965 , n31964 );
buf ( n31966 , n31965 );
and ( n31967 , n31966 , n30597 );
and ( n31968 , n31961 , n31967 );
and ( n31969 , n31957 , n31967 );
or ( n31970 , n31962 , n31968 , n31969 );
and ( n31971 , n31560 , n30691 );
and ( n31972 , n31476 , n30689 );
nor ( n31973 , n31971 , n31972 );
xnor ( n31974 , n31973 , n30696 );
and ( n31975 , n31970 , n31974 );
xor ( n31976 , n31855 , n31859 );
xor ( n31977 , n31976 , n31865 );
and ( n31978 , n31974 , n31977 );
and ( n31979 , n31970 , n31977 );
or ( n31980 , n31975 , n31978 , n31979 );
and ( n31981 , n30762 , n31354 );
and ( n31982 , n30718 , n31351 );
nor ( n31983 , n31981 , n31982 );
xnor ( n31984 , n31983 , n31146 );
and ( n31985 , n31980 , n31984 );
and ( n31986 , n30858 , n31220 );
and ( n31987 , n30816 , n31218 );
nor ( n31988 , n31986 , n31987 );
xnor ( n31989 , n31988 , n31154 );
and ( n31990 , n31984 , n31989 );
and ( n31991 , n31980 , n31989 );
or ( n31992 , n31985 , n31990 , n31991 );
and ( n31993 , n30903 , n31220 );
and ( n31994 , n30858 , n31218 );
nor ( n31995 , n31993 , n31994 );
xnor ( n31996 , n31995 , n31154 );
and ( n31997 , n31228 , n30911 );
and ( n31998 , n31160 , n30909 );
nor ( n31999 , n31997 , n31998 );
xnor ( n32000 , n31999 , n30848 );
and ( n32001 , n31996 , n32000 );
and ( n32002 , n31366 , n30770 );
and ( n32003 , n31307 , n30768 );
nor ( n32004 , n32002 , n32003 );
xnor ( n32005 , n32004 , n30752 );
and ( n32006 , n32000 , n32005 );
and ( n32007 , n31996 , n32005 );
or ( n32008 , n32001 , n32006 , n32007 );
and ( n32009 , n30967 , n30975 );
and ( n32010 , n30903 , n30973 );
nor ( n32011 , n32009 , n32010 );
xnor ( n32012 , n32011 , n30957 );
and ( n32013 , n31160 , n30911 );
and ( n32014 , n31053 , n30909 );
nor ( n32015 , n32013 , n32014 );
xnor ( n32016 , n32015 , n30848 );
xor ( n32017 , n32012 , n32016 );
and ( n32018 , n31307 , n30770 );
and ( n32019 , n31228 , n30768 );
nor ( n32020 , n32018 , n32019 );
xnor ( n32021 , n32020 , n30752 );
xor ( n32022 , n32017 , n32021 );
and ( n32023 , n32008 , n32022 );
xor ( n32024 , n31868 , n31872 );
xor ( n32025 , n32024 , n31875 );
and ( n32026 , n32022 , n32025 );
and ( n32027 , n32008 , n32025 );
or ( n32028 , n32023 , n32026 , n32027 );
and ( n32029 , n31992 , n32028 );
xor ( n32030 , n31878 , n31882 );
xor ( n32031 , n32030 , n31887 );
and ( n32032 , n32028 , n32031 );
and ( n32033 , n31992 , n32031 );
or ( n32034 , n32029 , n32032 , n32033 );
and ( n32035 , n32012 , n32016 );
and ( n32036 , n32016 , n32021 );
and ( n32037 , n32012 , n32021 );
or ( n32038 , n32035 , n32036 , n32037 );
xor ( n32039 , n31827 , n31831 );
xor ( n32040 , n32039 , n31836 );
and ( n32041 , n32038 , n32040 );
xor ( n32042 , n31894 , n31898 );
xor ( n32043 , n32042 , n31901 );
and ( n32044 , n32040 , n32043 );
and ( n32045 , n32038 , n32043 );
or ( n32046 , n32041 , n32044 , n32045 );
and ( n32047 , n32034 , n32046 );
xor ( n32048 , n31931 , n31933 );
xor ( n32049 , n32048 , n31936 );
and ( n32050 , n32046 , n32049 );
and ( n32051 , n32034 , n32049 );
or ( n32052 , n32047 , n32050 , n32051 );
and ( n32053 , n31953 , n32052 );
xor ( n32054 , n31929 , n31947 );
and ( n32055 , n32053 , n32054 );
xor ( n32056 , n32053 , n32054 );
xor ( n32057 , n32034 , n32046 );
xor ( n32058 , n32057 , n32049 );
and ( n32059 , n31823 , n30645 );
and ( n32060 , n31741 , n30643 );
nor ( n32061 , n32059 , n32060 );
xnor ( n32062 , n32061 , n30619 );
and ( n32063 , n31966 , n30605 );
and ( n32064 , n31864 , n30603 );
nor ( n32065 , n32063 , n32064 );
xnor ( n32066 , n32065 , n30610 );
and ( n32067 , n32062 , n32066 );
xor ( n32068 , n30523 , n30556 );
buf ( n32069 , n32068 );
buf ( n32070 , n32069 );
buf ( n32071 , n32070 );
and ( n32072 , n32071 , n30597 );
and ( n32073 , n32066 , n32072 );
and ( n32074 , n32062 , n32072 );
or ( n32075 , n32067 , n32073 , n32074 );
and ( n32076 , n31645 , n30691 );
and ( n32077 , n31560 , n30689 );
nor ( n32078 , n32076 , n32077 );
xnor ( n32079 , n32078 , n30696 );
and ( n32080 , n32075 , n32079 );
xor ( n32081 , n31957 , n31961 );
xor ( n32082 , n32081 , n31967 );
and ( n32083 , n32079 , n32082 );
and ( n32084 , n32075 , n32082 );
or ( n32085 , n32080 , n32083 , n32084 );
and ( n32086 , n30816 , n31354 );
and ( n32087 , n30762 , n31351 );
nor ( n32088 , n32086 , n32087 );
xnor ( n32089 , n32088 , n31146 );
and ( n32090 , n32085 , n32089 );
and ( n32091 , n31053 , n30975 );
and ( n32092 , n30967 , n30973 );
nor ( n32093 , n32091 , n32092 );
xnor ( n32094 , n32093 , n30957 );
and ( n32095 , n32089 , n32094 );
and ( n32096 , n32085 , n32094 );
or ( n32097 , n32090 , n32095 , n32096 );
and ( n32098 , n31864 , n30645 );
and ( n32099 , n31823 , n30643 );
nor ( n32100 , n32098 , n32099 );
xnor ( n32101 , n32100 , n30619 );
and ( n32102 , n32071 , n30605 );
and ( n32103 , n31966 , n30603 );
nor ( n32104 , n32102 , n32103 );
xnor ( n32105 , n32104 , n30610 );
and ( n32106 , n32101 , n32105 );
xor ( n32107 , n30524 , n30555 );
buf ( n32108 , n32107 );
buf ( n32109 , n32108 );
buf ( n32110 , n32109 );
and ( n32111 , n32110 , n30597 );
and ( n32112 , n32105 , n32111 );
and ( n32113 , n32101 , n32111 );
or ( n32114 , n32106 , n32112 , n32113 );
and ( n32115 , n31560 , n30770 );
and ( n32116 , n31476 , n30768 );
nor ( n32117 , n32115 , n32116 );
xnor ( n32118 , n32117 , n30752 );
and ( n32119 , n32114 , n32118 );
and ( n32120 , n31684 , n30691 );
and ( n32121 , n31645 , n30689 );
nor ( n32122 , n32120 , n32121 );
xnor ( n32123 , n32122 , n30696 );
and ( n32124 , n32118 , n32123 );
and ( n32125 , n32114 , n32123 );
or ( n32126 , n32119 , n32124 , n32125 );
and ( n32127 , n31307 , n30911 );
and ( n32128 , n31228 , n30909 );
nor ( n32129 , n32127 , n32128 );
xnor ( n32130 , n32129 , n30848 );
and ( n32131 , n32126 , n32130 );
and ( n32132 , n31476 , n30770 );
and ( n32133 , n31366 , n30768 );
nor ( n32134 , n32132 , n32133 );
xnor ( n32135 , n32134 , n30752 );
and ( n32136 , n32130 , n32135 );
and ( n32137 , n32126 , n32135 );
or ( n32138 , n32131 , n32136 , n32137 );
xor ( n32139 , n31996 , n32000 );
xor ( n32140 , n32139 , n32005 );
and ( n32141 , n32138 , n32140 );
xor ( n32142 , n31970 , n31974 );
xor ( n32143 , n32142 , n31977 );
and ( n32144 , n32140 , n32143 );
and ( n32145 , n32138 , n32143 );
or ( n32146 , n32141 , n32144 , n32145 );
and ( n32147 , n32097 , n32146 );
xor ( n32148 , n31980 , n31984 );
xor ( n32149 , n32148 , n31989 );
and ( n32150 , n32146 , n32149 );
and ( n32151 , n32097 , n32149 );
or ( n32152 , n32147 , n32150 , n32151 );
xor ( n32153 , n31992 , n32028 );
xor ( n32154 , n32153 , n32031 );
and ( n32155 , n32152 , n32154 );
xor ( n32156 , n32038 , n32040 );
xor ( n32157 , n32156 , n32043 );
and ( n32158 , n32154 , n32157 );
and ( n32159 , n32152 , n32157 );
or ( n32160 , n32155 , n32158 , n32159 );
and ( n32161 , n32058 , n32160 );
xor ( n32162 , n31953 , n32052 );
and ( n32163 , n32161 , n32162 );
xor ( n32164 , n32161 , n32162 );
xor ( n32165 , n32152 , n32154 );
xor ( n32166 , n32165 , n32157 );
and ( n32167 , n30858 , n31354 );
and ( n32168 , n30816 , n31351 );
nor ( n32169 , n32167 , n32168 );
xnor ( n32170 , n32169 , n31146 );
and ( n32171 , n30967 , n31220 );
and ( n32172 , n30903 , n31218 );
nor ( n32173 , n32171 , n32172 );
xnor ( n32174 , n32173 , n31154 );
and ( n32175 , n32170 , n32174 );
and ( n32176 , n31160 , n30975 );
and ( n32177 , n31053 , n30973 );
nor ( n32178 , n32176 , n32177 );
xnor ( n32179 , n32178 , n30957 );
and ( n32180 , n32174 , n32179 );
and ( n32181 , n32170 , n32179 );
or ( n32182 , n32175 , n32180 , n32181 );
and ( n32183 , n31823 , n30691 );
and ( n32184 , n31741 , n30689 );
nor ( n32185 , n32183 , n32184 );
xnor ( n32186 , n32185 , n30696 );
and ( n32187 , n32110 , n30605 );
and ( n32188 , n32071 , n30603 );
nor ( n32189 , n32187 , n32188 );
xnor ( n32190 , n32189 , n30610 );
and ( n32191 , n32186 , n32190 );
xor ( n32192 , n30551 , n30553 );
buf ( n32193 , n32192 );
buf ( n32194 , n32193 );
buf ( n32195 , n32194 );
and ( n32196 , n32195 , n30597 );
and ( n32197 , n32190 , n32196 );
and ( n32198 , n32186 , n32196 );
or ( n32199 , n32191 , n32197 , n32198 );
and ( n32200 , n31645 , n30770 );
and ( n32201 , n31560 , n30768 );
nor ( n32202 , n32200 , n32201 );
xnor ( n32203 , n32202 , n30752 );
and ( n32204 , n32199 , n32203 );
and ( n32205 , n31741 , n30691 );
and ( n32206 , n31684 , n30689 );
nor ( n32207 , n32205 , n32206 );
xnor ( n32208 , n32207 , n30696 );
and ( n32209 , n32203 , n32208 );
and ( n32210 , n32199 , n32208 );
or ( n32211 , n32204 , n32209 , n32210 );
and ( n32212 , n31366 , n30911 );
and ( n32213 , n31307 , n30909 );
nor ( n32214 , n32212 , n32213 );
xnor ( n32215 , n32214 , n30848 );
and ( n32216 , n32211 , n32215 );
xor ( n32217 , n32062 , n32066 );
xor ( n32218 , n32217 , n32072 );
and ( n32219 , n32215 , n32218 );
and ( n32220 , n32211 , n32218 );
or ( n32221 , n32216 , n32219 , n32220 );
xor ( n32222 , n32126 , n32130 );
xor ( n32223 , n32222 , n32135 );
and ( n32224 , n32221 , n32223 );
xor ( n32225 , n32075 , n32079 );
xor ( n32226 , n32225 , n32082 );
and ( n32227 , n32223 , n32226 );
and ( n32228 , n32221 , n32226 );
or ( n32229 , n32224 , n32227 , n32228 );
and ( n32230 , n32182 , n32229 );
xor ( n32231 , n32085 , n32089 );
xor ( n32232 , n32231 , n32094 );
and ( n32233 , n32229 , n32232 );
and ( n32234 , n32182 , n32232 );
or ( n32235 , n32230 , n32233 , n32234 );
xor ( n32236 , n32097 , n32146 );
xor ( n32237 , n32236 , n32149 );
and ( n32238 , n32235 , n32237 );
xor ( n32239 , n32008 , n32022 );
xor ( n32240 , n32239 , n32025 );
and ( n32241 , n32237 , n32240 );
and ( n32242 , n32235 , n32240 );
or ( n32243 , n32238 , n32241 , n32242 );
and ( n32244 , n32166 , n32243 );
xor ( n32245 , n32058 , n32160 );
and ( n32246 , n32244 , n32245 );
xor ( n32247 , n32244 , n32245 );
xor ( n32248 , n32235 , n32237 );
xor ( n32249 , n32248 , n32240 );
and ( n32250 , n30903 , n31354 );
and ( n32251 , n30858 , n31351 );
nor ( n32252 , n32250 , n32251 );
xnor ( n32253 , n32252 , n31146 );
and ( n32254 , n31053 , n31220 );
and ( n32255 , n30967 , n31218 );
nor ( n32256 , n32254 , n32255 );
xnor ( n32257 , n32256 , n31154 );
and ( n32258 , n32253 , n32257 );
and ( n32259 , n31228 , n30975 );
and ( n32260 , n31160 , n30973 );
nor ( n32261 , n32259 , n32260 );
xnor ( n32262 , n32261 , n30957 );
and ( n32263 , n32257 , n32262 );
and ( n32264 , n32253 , n32262 );
or ( n32265 , n32258 , n32263 , n32264 );
and ( n32266 , n32071 , n30645 );
and ( n32267 , n31966 , n30643 );
nor ( n32268 , n32266 , n32267 );
xnor ( n32269 , n32268 , n30619 );
and ( n32270 , n32195 , n30605 );
and ( n32271 , n32110 , n30603 );
nor ( n32272 , n32270 , n32271 );
xnor ( n32273 , n32272 , n30610 );
and ( n32274 , n32269 , n32273 );
not ( n32275 , n30553 );
buf ( n32276 , n32275 );
buf ( n32277 , n32276 );
buf ( n32278 , n32277 );
and ( n32279 , n32278 , n30597 );
and ( n32280 , n32273 , n32279 );
and ( n32281 , n32269 , n32279 );
or ( n32282 , n32274 , n32280 , n32281 );
and ( n32283 , n31684 , n30770 );
and ( n32284 , n31645 , n30768 );
nor ( n32285 , n32283 , n32284 );
xnor ( n32286 , n32285 , n30752 );
and ( n32287 , n32282 , n32286 );
and ( n32288 , n31966 , n30645 );
and ( n32289 , n31864 , n30643 );
nor ( n32290 , n32288 , n32289 );
xnor ( n32291 , n32290 , n30619 );
and ( n32292 , n32286 , n32291 );
and ( n32293 , n32282 , n32291 );
or ( n32294 , n32287 , n32292 , n32293 );
and ( n32295 , n31476 , n30911 );
and ( n32296 , n31366 , n30909 );
nor ( n32297 , n32295 , n32296 );
xnor ( n32298 , n32297 , n30848 );
and ( n32299 , n32294 , n32298 );
xor ( n32300 , n32101 , n32105 );
xor ( n32301 , n32300 , n32111 );
and ( n32302 , n32298 , n32301 );
and ( n32303 , n32294 , n32301 );
or ( n32304 , n32299 , n32302 , n32303 );
xor ( n32305 , n32114 , n32118 );
xor ( n32306 , n32305 , n32123 );
and ( n32307 , n32304 , n32306 );
xor ( n32308 , n32211 , n32215 );
xor ( n32309 , n32308 , n32218 );
and ( n32310 , n32306 , n32309 );
and ( n32311 , n32304 , n32309 );
or ( n32312 , n32307 , n32310 , n32311 );
and ( n32313 , n32265 , n32312 );
xor ( n32314 , n32170 , n32174 );
xor ( n32315 , n32314 , n32179 );
and ( n32316 , n32312 , n32315 );
and ( n32317 , n32265 , n32315 );
or ( n32318 , n32313 , n32316 , n32317 );
xor ( n32319 , n32182 , n32229 );
xor ( n32320 , n32319 , n32232 );
and ( n32321 , n32318 , n32320 );
xor ( n32322 , n32138 , n32140 );
xor ( n32323 , n32322 , n32143 );
and ( n32324 , n32320 , n32323 );
and ( n32325 , n32318 , n32323 );
or ( n32326 , n32321 , n32324 , n32325 );
and ( n32327 , n32249 , n32326 );
xor ( n32328 , n32166 , n32243 );
and ( n32329 , n32327 , n32328 );
xor ( n32330 , n32327 , n32328 );
xor ( n32331 , n32318 , n32320 );
xor ( n32332 , n32331 , n32323 );
and ( n32333 , n32110 , n30645 );
and ( n32334 , n32071 , n30643 );
nor ( n32335 , n32333 , n32334 );
xnor ( n32336 , n32335 , n30619 );
and ( n32337 , n32278 , n30605 );
and ( n32338 , n32195 , n30603 );
nor ( n32339 , n32337 , n32338 );
xnor ( n32340 , n32339 , n30610 );
and ( n32341 , n32336 , n32340 );
xnor ( n32342 , n30543 , n30545 );
buf ( n32343 , n32342 );
buf ( n32344 , n32343 );
buf ( n32345 , n32344 );
and ( n32346 , n32345 , n30597 );
and ( n32347 , n32340 , n32346 );
and ( n32348 , n32336 , n32346 );
or ( n32349 , n32341 , n32347 , n32348 );
and ( n32350 , n31741 , n30770 );
and ( n32351 , n31684 , n30768 );
nor ( n32352 , n32350 , n32351 );
xnor ( n32353 , n32352 , n30752 );
and ( n32354 , n32349 , n32353 );
and ( n32355 , n31864 , n30691 );
and ( n32356 , n31823 , n30689 );
nor ( n32357 , n32355 , n32356 );
xnor ( n32358 , n32357 , n30696 );
and ( n32359 , n32353 , n32358 );
and ( n32360 , n32349 , n32358 );
or ( n32361 , n32354 , n32359 , n32360 );
and ( n32362 , n31560 , n30911 );
and ( n32363 , n31476 , n30909 );
nor ( n32364 , n32362 , n32363 );
xnor ( n32365 , n32364 , n30848 );
and ( n32366 , n32361 , n32365 );
xor ( n32367 , n32186 , n32190 );
xor ( n32368 , n32367 , n32196 );
and ( n32369 , n32365 , n32368 );
and ( n32370 , n32361 , n32368 );
or ( n32371 , n32366 , n32369 , n32370 );
and ( n32372 , n31228 , n31220 );
and ( n32373 , n31160 , n31218 );
nor ( n32374 , n32372 , n32373 );
xnor ( n32375 , n32374 , n31154 );
and ( n32376 , n31366 , n30975 );
and ( n32377 , n31307 , n30973 );
nor ( n32378 , n32376 , n32377 );
xnor ( n32379 , n32378 , n30957 );
and ( n32380 , n32375 , n32379 );
xor ( n32381 , n32282 , n32286 );
xor ( n32382 , n32381 , n32291 );
and ( n32383 , n32379 , n32382 );
and ( n32384 , n32375 , n32382 );
or ( n32385 , n32380 , n32383 , n32384 );
and ( n32386 , n32371 , n32385 );
and ( n32387 , n30967 , n31354 );
and ( n32388 , n30903 , n31351 );
nor ( n32389 , n32387 , n32388 );
xnor ( n32390 , n32389 , n31146 );
and ( n32391 , n32385 , n32390 );
and ( n32392 , n32371 , n32390 );
or ( n32393 , n32386 , n32391 , n32392 );
and ( n32394 , n31160 , n31220 );
and ( n32395 , n31053 , n31218 );
nor ( n32396 , n32394 , n32395 );
xnor ( n32397 , n32396 , n31154 );
and ( n32398 , n31307 , n30975 );
and ( n32399 , n31228 , n30973 );
nor ( n32400 , n32398 , n32399 );
xnor ( n32401 , n32400 , n30957 );
and ( n32402 , n32397 , n32401 );
xor ( n32403 , n32199 , n32203 );
xor ( n32404 , n32403 , n32208 );
and ( n32405 , n32401 , n32404 );
and ( n32406 , n32397 , n32404 );
or ( n32407 , n32402 , n32405 , n32406 );
and ( n32408 , n32393 , n32407 );
xor ( n32409 , n32253 , n32257 );
xor ( n32410 , n32409 , n32262 );
and ( n32411 , n32407 , n32410 );
and ( n32412 , n32393 , n32410 );
or ( n32413 , n32408 , n32411 , n32412 );
xor ( n32414 , n32265 , n32312 );
xor ( n32415 , n32414 , n32315 );
and ( n32416 , n32413 , n32415 );
xor ( n32417 , n32221 , n32223 );
xor ( n32418 , n32417 , n32226 );
and ( n32419 , n32415 , n32418 );
and ( n32420 , n32413 , n32418 );
or ( n32421 , n32416 , n32419 , n32420 );
and ( n32422 , n32332 , n32421 );
xor ( n32423 , n32249 , n32326 );
and ( n32424 , n32422 , n32423 );
xor ( n32425 , n32422 , n32423 );
xor ( n32426 , n32413 , n32415 );
xor ( n32427 , n32426 , n32418 );
and ( n32428 , n32195 , n30645 );
and ( n32429 , n32110 , n30643 );
nor ( n32430 , n32428 , n32429 );
xnor ( n32431 , n32430 , n30619 );
and ( n32432 , n32345 , n30605 );
and ( n32433 , n32278 , n30603 );
nor ( n32434 , n32432 , n32433 );
xnor ( n32435 , n32434 , n30610 );
and ( n32436 , n32431 , n32435 );
xnor ( n32437 , n30541 , n30542 );
buf ( n32438 , n32437 );
buf ( n32439 , n32438 );
buf ( n32440 , n32439 );
and ( n32441 , n32440 , n30597 );
and ( n32442 , n32435 , n32441 );
and ( n32443 , n32431 , n32441 );
or ( n32444 , n32436 , n32442 , n32443 );
and ( n32445 , n31966 , n30691 );
and ( n32446 , n31864 , n30689 );
nor ( n32447 , n32445 , n32446 );
xnor ( n32448 , n32447 , n30696 );
and ( n32449 , n32444 , n32448 );
xor ( n32450 , n32336 , n32340 );
xor ( n32451 , n32450 , n32346 );
and ( n32452 , n32448 , n32451 );
and ( n32453 , n32444 , n32451 );
or ( n32454 , n32449 , n32452 , n32453 );
and ( n32455 , n31645 , n30911 );
and ( n32456 , n31560 , n30909 );
nor ( n32457 , n32455 , n32456 );
xnor ( n32458 , n32457 , n30848 );
and ( n32459 , n32454 , n32458 );
xor ( n32460 , n32269 , n32273 );
xor ( n32461 , n32460 , n32279 );
and ( n32462 , n32458 , n32461 );
and ( n32463 , n32454 , n32461 );
or ( n32464 , n32459 , n32462 , n32463 );
and ( n32465 , n31053 , n31354 );
and ( n32466 , n30967 , n31351 );
nor ( n32467 , n32465 , n32466 );
xnor ( n32468 , n32467 , n31146 );
and ( n32469 , n32464 , n32468 );
xor ( n32470 , n32361 , n32365 );
xor ( n32471 , n32470 , n32368 );
and ( n32472 , n32468 , n32471 );
and ( n32473 , n32464 , n32471 );
or ( n32474 , n32469 , n32472 , n32473 );
xor ( n32475 , n32294 , n32298 );
xor ( n32476 , n32475 , n32301 );
and ( n32477 , n32474 , n32476 );
xor ( n32478 , n32397 , n32401 );
xor ( n32479 , n32478 , n32404 );
and ( n32480 , n32476 , n32479 );
and ( n32481 , n32474 , n32479 );
or ( n32482 , n32477 , n32480 , n32481 );
xor ( n32483 , n32393 , n32407 );
xor ( n32484 , n32483 , n32410 );
and ( n32485 , n32482 , n32484 );
xor ( n32486 , n32304 , n32306 );
xor ( n32487 , n32486 , n32309 );
and ( n32488 , n32484 , n32487 );
and ( n32489 , n32482 , n32487 );
or ( n32490 , n32485 , n32488 , n32489 );
and ( n32491 , n32427 , n32490 );
xor ( n32492 , n32332 , n32421 );
and ( n32493 , n32491 , n32492 );
xor ( n32494 , n32491 , n32492 );
xor ( n32495 , n32427 , n32490 );
xor ( n32496 , n32482 , n32484 );
xor ( n32497 , n32496 , n32487 );
buf ( n32498 , n29289 );
buf ( n32499 , n32498 );
buf ( n32500 , n32499 );
buf ( n32501 , n32500 );
and ( n32502 , n32501 , n30603 );
not ( n32503 , n32502 );
and ( n32504 , n32503 , n30610 );
buf ( n32505 , n794 );
buf ( n32506 , n32505 );
and ( n32507 , n32504 , n32506 );
and ( n32508 , n32501 , n30597 );
and ( n32509 , n32507 , n32508 );
and ( n32510 , n32278 , n30645 );
and ( n32511 , n32195 , n30643 );
nor ( n32512 , n32510 , n32511 );
xnor ( n32513 , n32512 , n30619 );
and ( n32514 , n32509 , n32513 );
and ( n32515 , n32440 , n30605 );
and ( n32516 , n32345 , n30603 );
nor ( n32517 , n32515 , n32516 );
xnor ( n32518 , n32517 , n30610 );
and ( n32519 , n32513 , n32518 );
and ( n32520 , n32509 , n32518 );
or ( n32521 , n32514 , n32519 , n32520 );
and ( n32522 , n32071 , n30691 );
and ( n32523 , n31966 , n30689 );
nor ( n32524 , n32522 , n32523 );
xnor ( n32525 , n32524 , n30696 );
and ( n32526 , n32521 , n32525 );
xor ( n32527 , n32431 , n32435 );
xor ( n32528 , n32527 , n32441 );
and ( n32529 , n32525 , n32528 );
and ( n32530 , n32521 , n32528 );
or ( n32531 , n32526 , n32529 , n32530 );
and ( n32532 , n31684 , n30911 );
and ( n32533 , n31645 , n30909 );
nor ( n32534 , n32532 , n32533 );
xnor ( n32535 , n32534 , n30848 );
and ( n32536 , n32531 , n32535 );
and ( n32537 , n31823 , n30770 );
and ( n32538 , n31741 , n30768 );
nor ( n32539 , n32537 , n32538 );
xnor ( n32540 , n32539 , n30752 );
and ( n32541 , n32535 , n32540 );
and ( n32542 , n32531 , n32540 );
or ( n32543 , n32536 , n32541 , n32542 );
and ( n32544 , n31476 , n30975 );
and ( n32545 , n31366 , n30973 );
nor ( n32546 , n32544 , n32545 );
xnor ( n32547 , n32546 , n30957 );
and ( n32548 , n32543 , n32547 );
xor ( n32549 , n32349 , n32353 );
xor ( n32550 , n32549 , n32358 );
and ( n32551 , n32547 , n32550 );
and ( n32552 , n32543 , n32550 );
or ( n32553 , n32548 , n32551 , n32552 );
xor ( n32554 , n32507 , n32508 );
xor ( n32555 , n32504 , n32506 );
and ( n32556 , n32440 , n30645 );
and ( n32557 , n32345 , n30643 );
nor ( n32558 , n32556 , n32557 );
xnor ( n32559 , n32558 , n30619 );
and ( n32560 , n32555 , n32559 );
and ( n32561 , n32501 , n30605 );
not ( n32562 , n32561 );
xnor ( n32563 , n32562 , n30610 );
and ( n32564 , n32559 , n32563 );
and ( n32565 , n32555 , n32563 );
or ( n32566 , n32560 , n32564 , n32565 );
and ( n32567 , n32554 , n32566 );
and ( n32568 , n32440 , n30603 );
not ( n32569 , n32568 );
xnor ( n32570 , n32569 , n30610 );
and ( n32571 , n32566 , n32570 );
and ( n32572 , n32554 , n32570 );
or ( n32573 , n32567 , n32571 , n32572 );
and ( n32574 , n32110 , n30691 );
and ( n32575 , n32071 , n30689 );
nor ( n32576 , n32574 , n32575 );
xnor ( n32577 , n32576 , n30696 );
and ( n32578 , n32573 , n32577 );
xor ( n32579 , n32509 , n32513 );
xor ( n32580 , n32579 , n32518 );
and ( n32581 , n32577 , n32580 );
and ( n32582 , n32573 , n32580 );
or ( n32583 , n32578 , n32581 , n32582 );
and ( n32584 , n31741 , n30911 );
and ( n32585 , n31684 , n30909 );
nor ( n32586 , n32584 , n32585 );
xnor ( n32587 , n32586 , n30848 );
and ( n32588 , n32583 , n32587 );
and ( n32589 , n31864 , n30770 );
and ( n32590 , n31823 , n30768 );
nor ( n32591 , n32589 , n32590 );
xnor ( n32592 , n32591 , n30752 );
and ( n32593 , n32587 , n32592 );
and ( n32594 , n32583 , n32592 );
or ( n32595 , n32588 , n32593 , n32594 );
and ( n32596 , n31560 , n30975 );
and ( n32597 , n31476 , n30973 );
nor ( n32598 , n32596 , n32597 );
xnor ( n32599 , n32598 , n30957 );
and ( n32600 , n32595 , n32599 );
xor ( n32601 , n32444 , n32448 );
xor ( n32602 , n32601 , n32451 );
and ( n32603 , n32599 , n32602 );
and ( n32604 , n32595 , n32602 );
or ( n32605 , n32600 , n32603 , n32604 );
and ( n32606 , n31307 , n31220 );
and ( n32607 , n31228 , n31218 );
nor ( n32608 , n32606 , n32607 );
xnor ( n32609 , n32608 , n31154 );
and ( n32610 , n32605 , n32609 );
xor ( n32611 , n32454 , n32458 );
xor ( n32612 , n32611 , n32461 );
and ( n32613 , n32609 , n32612 );
and ( n32614 , n32605 , n32612 );
or ( n32615 , n32610 , n32613 , n32614 );
and ( n32616 , n32553 , n32615 );
xor ( n32617 , n32375 , n32379 );
xor ( n32618 , n32617 , n32382 );
and ( n32619 , n32615 , n32618 );
and ( n32620 , n32553 , n32618 );
or ( n32621 , n32616 , n32619 , n32620 );
xor ( n32622 , n32371 , n32385 );
xor ( n32623 , n32622 , n32390 );
and ( n32624 , n32621 , n32623 );
xor ( n32625 , n32474 , n32476 );
xor ( n32626 , n32625 , n32479 );
and ( n32627 , n32623 , n32626 );
and ( n32628 , n32621 , n32626 );
or ( n32629 , n32624 , n32627 , n32628 );
and ( n32630 , n32497 , n32629 );
and ( n32631 , n32495 , n32630 );
xor ( n32632 , n32495 , n32630 );
xor ( n32633 , n32621 , n32623 );
xor ( n32634 , n32633 , n32626 );
and ( n32635 , n32195 , n30691 );
and ( n32636 , n32110 , n30689 );
nor ( n32637 , n32635 , n32636 );
xnor ( n32638 , n32637 , n30696 );
and ( n32639 , n32345 , n30645 );
and ( n32640 , n32278 , n30643 );
nor ( n32641 , n32639 , n32640 );
xnor ( n32642 , n32641 , n30619 );
and ( n32643 , n32638 , n32642 );
xor ( n32644 , n32554 , n32566 );
xor ( n32645 , n32644 , n32570 );
and ( n32646 , n32642 , n32645 );
and ( n32647 , n32638 , n32645 );
or ( n32648 , n32643 , n32646 , n32647 );
and ( n32649 , n31823 , n30911 );
and ( n32650 , n31741 , n30909 );
nor ( n32651 , n32649 , n32650 );
xnor ( n32652 , n32651 , n30848 );
and ( n32653 , n32648 , n32652 );
and ( n32654 , n31966 , n30770 );
and ( n32655 , n31864 , n30768 );
nor ( n32656 , n32654 , n32655 );
xnor ( n32657 , n32656 , n30752 );
and ( n32658 , n32652 , n32657 );
and ( n32659 , n32648 , n32657 );
or ( n32660 , n32653 , n32658 , n32659 );
and ( n32661 , n31645 , n30975 );
and ( n32662 , n31560 , n30973 );
nor ( n32663 , n32661 , n32662 );
xnor ( n32664 , n32663 , n30957 );
and ( n32665 , n32660 , n32664 );
xor ( n32666 , n32521 , n32525 );
xor ( n32667 , n32666 , n32528 );
and ( n32668 , n32664 , n32667 );
and ( n32669 , n32660 , n32667 );
or ( n32670 , n32665 , n32668 , n32669 );
and ( n32671 , n31228 , n31354 );
and ( n32672 , n31160 , n31351 );
nor ( n32673 , n32671 , n32672 );
xnor ( n32674 , n32673 , n31146 );
and ( n32675 , n32670 , n32674 );
xor ( n32676 , n32531 , n32535 );
xor ( n32677 , n32676 , n32540 );
and ( n32678 , n32674 , n32677 );
and ( n32679 , n32670 , n32677 );
or ( n32680 , n32675 , n32678 , n32679 );
and ( n32681 , n31160 , n31354 );
and ( n32682 , n31053 , n31351 );
nor ( n32683 , n32681 , n32682 );
xnor ( n32684 , n32683 , n31146 );
and ( n32685 , n32680 , n32684 );
xor ( n32686 , n32543 , n32547 );
xor ( n32687 , n32686 , n32550 );
and ( n32688 , n32684 , n32687 );
and ( n32689 , n32680 , n32687 );
or ( n32690 , n32685 , n32688 , n32689 );
xor ( n32691 , n32464 , n32468 );
xor ( n32692 , n32691 , n32471 );
and ( n32693 , n32690 , n32692 );
xor ( n32694 , n32553 , n32615 );
xor ( n32695 , n32694 , n32618 );
and ( n32696 , n32692 , n32695 );
and ( n32697 , n32690 , n32695 );
or ( n32698 , n32693 , n32696 , n32697 );
and ( n32699 , n32634 , n32698 );
xor ( n32700 , n32497 , n32629 );
and ( n32701 , n32699 , n32700 );
xor ( n32702 , n32699 , n32700 );
xor ( n32703 , n32690 , n32692 );
xor ( n32704 , n32703 , n32695 );
and ( n32705 , n32501 , n30643 );
not ( n32706 , n32705 );
and ( n32707 , n32706 , n30619 );
buf ( n32708 , n796 );
buf ( n32709 , n32708 );
and ( n32710 , n32707 , n32709 );
and ( n32711 , n32710 , n32502 );
buf ( n32712 , n795 );
buf ( n32713 , n32712 );
and ( n32714 , n32502 , n32713 );
and ( n32715 , n32710 , n32713 );
or ( n32716 , n32711 , n32714 , n32715 );
and ( n32717 , n32278 , n30691 );
and ( n32718 , n32195 , n30689 );
nor ( n32719 , n32717 , n32718 );
xnor ( n32720 , n32719 , n30696 );
and ( n32721 , n32716 , n32720 );
xor ( n32722 , n32555 , n32559 );
xor ( n32723 , n32722 , n32563 );
and ( n32724 , n32720 , n32723 );
and ( n32725 , n32716 , n32723 );
or ( n32726 , n32721 , n32724 , n32725 );
and ( n32727 , n32071 , n30770 );
and ( n32728 , n31966 , n30768 );
nor ( n32729 , n32727 , n32728 );
xnor ( n32730 , n32729 , n30752 );
and ( n32731 , n32726 , n32730 );
xor ( n32732 , n32638 , n32642 );
xor ( n32733 , n32732 , n32645 );
and ( n32734 , n32730 , n32733 );
and ( n32735 , n32726 , n32733 );
or ( n32736 , n32731 , n32734 , n32735 );
and ( n32737 , n31684 , n30975 );
and ( n32738 , n31645 , n30973 );
nor ( n32739 , n32737 , n32738 );
xnor ( n32740 , n32739 , n30957 );
and ( n32741 , n32736 , n32740 );
xor ( n32742 , n32573 , n32577 );
xor ( n32743 , n32742 , n32580 );
and ( n32744 , n32740 , n32743 );
and ( n32745 , n32736 , n32743 );
or ( n32746 , n32741 , n32744 , n32745 );
and ( n32747 , n31476 , n31220 );
and ( n32748 , n31366 , n31218 );
nor ( n32749 , n32747 , n32748 );
xnor ( n32750 , n32749 , n31154 );
and ( n32751 , n32746 , n32750 );
xor ( n32752 , n32583 , n32587 );
xor ( n32753 , n32752 , n32592 );
and ( n32754 , n32750 , n32753 );
and ( n32755 , n32746 , n32753 );
or ( n32756 , n32751 , n32754 , n32755 );
and ( n32757 , n31366 , n31220 );
and ( n32758 , n31307 , n31218 );
nor ( n32759 , n32757 , n32758 );
xnor ( n32760 , n32759 , n31154 );
and ( n32761 , n32756 , n32760 );
xor ( n32762 , n32595 , n32599 );
xor ( n32763 , n32762 , n32602 );
and ( n32764 , n32760 , n32763 );
and ( n32765 , n32756 , n32763 );
or ( n32766 , n32761 , n32764 , n32765 );
xor ( n32767 , n32605 , n32609 );
xor ( n32768 , n32767 , n32612 );
and ( n32769 , n32766 , n32768 );
xor ( n32770 , n32680 , n32684 );
xor ( n32771 , n32770 , n32687 );
and ( n32772 , n32768 , n32771 );
and ( n32773 , n32766 , n32771 );
or ( n32774 , n32769 , n32772 , n32773 );
and ( n32775 , n32704 , n32774 );
xor ( n32776 , n32634 , n32698 );
and ( n32777 , n32775 , n32776 );
xor ( n32778 , n32775 , n32776 );
xor ( n32779 , n32766 , n32768 );
xor ( n32780 , n32779 , n32771 );
and ( n32781 , n32345 , n30691 );
and ( n32782 , n32278 , n30689 );
nor ( n32783 , n32781 , n32782 );
xnor ( n32784 , n32783 , n30696 );
and ( n32785 , n32440 , n30643 );
not ( n32786 , n32785 );
xnor ( n32787 , n32786 , n30619 );
and ( n32788 , n32784 , n32787 );
xor ( n32789 , n32710 , n32502 );
xor ( n32790 , n32789 , n32713 );
and ( n32791 , n32787 , n32790 );
and ( n32792 , n32784 , n32790 );
or ( n32793 , n32788 , n32791 , n32792 );
and ( n32794 , n32110 , n30770 );
and ( n32795 , n32071 , n30768 );
nor ( n32796 , n32794 , n32795 );
xnor ( n32797 , n32796 , n30752 );
and ( n32798 , n32793 , n32797 );
xor ( n32799 , n32716 , n32720 );
xor ( n32800 , n32799 , n32723 );
and ( n32801 , n32797 , n32800 );
and ( n32802 , n32793 , n32800 );
or ( n32803 , n32798 , n32801 , n32802 );
and ( n32804 , n31741 , n30975 );
and ( n32805 , n31684 , n30973 );
nor ( n32806 , n32804 , n32805 );
xnor ( n32807 , n32806 , n30957 );
and ( n32808 , n32803 , n32807 );
and ( n32809 , n31864 , n30911 );
and ( n32810 , n31823 , n30909 );
nor ( n32811 , n32809 , n32810 );
xnor ( n32812 , n32811 , n30848 );
and ( n32813 , n32807 , n32812 );
and ( n32814 , n32803 , n32812 );
or ( n32815 , n32808 , n32813 , n32814 );
and ( n32816 , n31560 , n31220 );
and ( n32817 , n31476 , n31218 );
nor ( n32818 , n32816 , n32817 );
xnor ( n32819 , n32818 , n31154 );
and ( n32820 , n32815 , n32819 );
xor ( n32821 , n32648 , n32652 );
xor ( n32822 , n32821 , n32657 );
and ( n32823 , n32819 , n32822 );
and ( n32824 , n32815 , n32822 );
or ( n32825 , n32820 , n32823 , n32824 );
and ( n32826 , n31307 , n31354 );
and ( n32827 , n31228 , n31351 );
nor ( n32828 , n32826 , n32827 );
xnor ( n32829 , n32828 , n31146 );
and ( n32830 , n32825 , n32829 );
xor ( n32831 , n32660 , n32664 );
xor ( n32832 , n32831 , n32667 );
and ( n32833 , n32829 , n32832 );
and ( n32834 , n32825 , n32832 );
or ( n32835 , n32830 , n32833 , n32834 );
xor ( n32836 , n32670 , n32674 );
xor ( n32837 , n32836 , n32677 );
and ( n32838 , n32835 , n32837 );
xor ( n32839 , n32756 , n32760 );
xor ( n32840 , n32839 , n32763 );
and ( n32841 , n32837 , n32840 );
and ( n32842 , n32835 , n32840 );
or ( n32843 , n32838 , n32841 , n32842 );
and ( n32844 , n32780 , n32843 );
xor ( n32845 , n32704 , n32774 );
and ( n32846 , n32844 , n32845 );
xor ( n32847 , n32844 , n32845 );
xor ( n32848 , n32707 , n32709 );
and ( n32849 , n32440 , n30691 );
and ( n32850 , n32345 , n30689 );
nor ( n32851 , n32849 , n32850 );
xnor ( n32852 , n32851 , n30696 );
and ( n32853 , n32848 , n32852 );
and ( n32854 , n32501 , n30645 );
not ( n32855 , n32854 );
xnor ( n32856 , n32855 , n30619 );
and ( n32857 , n32852 , n32856 );
and ( n32858 , n32848 , n32856 );
or ( n32859 , n32853 , n32857 , n32858 );
and ( n32860 , n32195 , n30770 );
and ( n32861 , n32110 , n30768 );
nor ( n32862 , n32860 , n32861 );
xnor ( n32863 , n32862 , n30752 );
and ( n32864 , n32859 , n32863 );
xor ( n32865 , n32784 , n32787 );
xor ( n32866 , n32865 , n32790 );
and ( n32867 , n32863 , n32866 );
and ( n32868 , n32859 , n32866 );
or ( n32869 , n32864 , n32867 , n32868 );
and ( n32870 , n31823 , n30975 );
and ( n32871 , n31741 , n30973 );
nor ( n32872 , n32870 , n32871 );
xnor ( n32873 , n32872 , n30957 );
and ( n32874 , n32869 , n32873 );
xor ( n32875 , n32793 , n32797 );
xor ( n32876 , n32875 , n32800 );
and ( n32877 , n32873 , n32876 );
and ( n32878 , n32869 , n32876 );
or ( n32879 , n32874 , n32877 , n32878 );
and ( n32880 , n31645 , n31220 );
and ( n32881 , n31560 , n31218 );
nor ( n32882 , n32880 , n32881 );
xnor ( n32883 , n32882 , n31154 );
and ( n32884 , n32879 , n32883 );
xor ( n32885 , n32726 , n32730 );
xor ( n32886 , n32885 , n32733 );
and ( n32887 , n32883 , n32886 );
and ( n32888 , n32879 , n32886 );
or ( n32889 , n32884 , n32887 , n32888 );
and ( n32890 , n31366 , n31354 );
and ( n32891 , n31307 , n31351 );
nor ( n32892 , n32890 , n32891 );
xnor ( n32893 , n32892 , n31146 );
and ( n32894 , n32889 , n32893 );
xor ( n32895 , n32736 , n32740 );
xor ( n32896 , n32895 , n32743 );
and ( n32897 , n32893 , n32896 );
and ( n32898 , n32889 , n32896 );
or ( n32899 , n32894 , n32897 , n32898 );
xor ( n32900 , n32746 , n32750 );
xor ( n32901 , n32900 , n32753 );
and ( n32902 , n32899 , n32901 );
xor ( n32903 , n32825 , n32829 );
xor ( n32904 , n32903 , n32832 );
and ( n32905 , n32901 , n32904 );
and ( n32906 , n32899 , n32904 );
or ( n32907 , n32902 , n32905 , n32906 );
xor ( n32908 , n32835 , n32837 );
xor ( n32909 , n32908 , n32840 );
and ( n32910 , n32907 , n32909 );
xor ( n32911 , n32780 , n32843 );
and ( n32912 , n32910 , n32911 );
xor ( n32913 , n32910 , n32911 );
xor ( n32914 , n32899 , n32901 );
xor ( n32915 , n32914 , n32904 );
and ( n32916 , n32501 , n30689 );
not ( n32917 , n32916 );
and ( n32918 , n32917 , n30696 );
buf ( n32919 , n798 );
buf ( n32920 , n32919 );
and ( n32921 , n32918 , n32920 );
and ( n32922 , n32921 , n32705 );
buf ( n32923 , n797 );
buf ( n32924 , n32923 );
and ( n32925 , n32705 , n32924 );
and ( n32926 , n32921 , n32924 );
or ( n32927 , n32922 , n32925 , n32926 );
and ( n32928 , n32278 , n30770 );
and ( n32929 , n32195 , n30768 );
nor ( n32930 , n32928 , n32929 );
xnor ( n32931 , n32930 , n30752 );
and ( n32932 , n32927 , n32931 );
xor ( n32933 , n32848 , n32852 );
xor ( n32934 , n32933 , n32856 );
and ( n32935 , n32931 , n32934 );
and ( n32936 , n32927 , n32934 );
or ( n32937 , n32932 , n32935 , n32936 );
and ( n32938 , n32071 , n30911 );
and ( n32939 , n31966 , n30909 );
nor ( n32940 , n32938 , n32939 );
xnor ( n32941 , n32940 , n30848 );
and ( n32942 , n32937 , n32941 );
xor ( n32943 , n32859 , n32863 );
xor ( n32944 , n32943 , n32866 );
and ( n32945 , n32941 , n32944 );
and ( n32946 , n32937 , n32944 );
or ( n32947 , n32942 , n32945 , n32946 );
and ( n32948 , n31684 , n31220 );
and ( n32949 , n31645 , n31218 );
nor ( n32950 , n32948 , n32949 );
xnor ( n32951 , n32950 , n31154 );
and ( n32952 , n32947 , n32951 );
and ( n32953 , n31966 , n30911 );
and ( n32954 , n31864 , n30909 );
nor ( n32955 , n32953 , n32954 );
xnor ( n32956 , n32955 , n30848 );
and ( n32957 , n32951 , n32956 );
and ( n32958 , n32947 , n32956 );
or ( n32959 , n32952 , n32957 , n32958 );
and ( n32960 , n31476 , n31354 );
and ( n32961 , n31366 , n31351 );
nor ( n32962 , n32960 , n32961 );
xnor ( n32963 , n32962 , n31146 );
and ( n32964 , n32959 , n32963 );
xor ( n32965 , n32803 , n32807 );
xor ( n32966 , n32965 , n32812 );
and ( n32967 , n32963 , n32966 );
and ( n32968 , n32959 , n32966 );
or ( n32969 , n32964 , n32967 , n32968 );
xor ( n32970 , n32815 , n32819 );
xor ( n32971 , n32970 , n32822 );
and ( n32972 , n32969 , n32971 );
xor ( n32973 , n32889 , n32893 );
xor ( n32974 , n32973 , n32896 );
and ( n32975 , n32971 , n32974 );
and ( n32976 , n32969 , n32974 );
or ( n32977 , n32972 , n32975 , n32976 );
and ( n32978 , n32915 , n32977 );
xor ( n32979 , n32907 , n32909 );
and ( n32980 , n32978 , n32979 );
xor ( n32981 , n32978 , n32979 );
xor ( n32982 , n32969 , n32971 );
xor ( n32983 , n32982 , n32974 );
and ( n32984 , n32345 , n30770 );
and ( n32985 , n32278 , n30768 );
nor ( n32986 , n32984 , n32985 );
xnor ( n32987 , n32986 , n30752 );
and ( n32988 , n32440 , n30689 );
not ( n32989 , n32988 );
xnor ( n32990 , n32989 , n30696 );
and ( n32991 , n32987 , n32990 );
xor ( n32992 , n32921 , n32705 );
xor ( n32993 , n32992 , n32924 );
and ( n32994 , n32990 , n32993 );
and ( n32995 , n32987 , n32993 );
or ( n32996 , n32991 , n32994 , n32995 );
and ( n32997 , n32110 , n30911 );
and ( n32998 , n32071 , n30909 );
nor ( n32999 , n32997 , n32998 );
xnor ( n33000 , n32999 , n30848 );
and ( n33001 , n32996 , n33000 );
xor ( n33002 , n32927 , n32931 );
xor ( n33003 , n33002 , n32934 );
and ( n33004 , n33000 , n33003 );
and ( n33005 , n32996 , n33003 );
or ( n33006 , n33001 , n33004 , n33005 );
and ( n33007 , n31741 , n31220 );
and ( n33008 , n31684 , n31218 );
nor ( n33009 , n33007 , n33008 );
xnor ( n33010 , n33009 , n31154 );
and ( n33011 , n33006 , n33010 );
and ( n33012 , n31864 , n30975 );
and ( n33013 , n31823 , n30973 );
nor ( n33014 , n33012 , n33013 );
xnor ( n33015 , n33014 , n30957 );
and ( n33016 , n33010 , n33015 );
and ( n33017 , n33006 , n33015 );
or ( n33018 , n33011 , n33016 , n33017 );
and ( n33019 , n31560 , n31354 );
and ( n33020 , n31476 , n31351 );
nor ( n33021 , n33019 , n33020 );
xnor ( n33022 , n33021 , n31146 );
and ( n33023 , n33018 , n33022 );
xor ( n33024 , n32869 , n32873 );
xor ( n33025 , n33024 , n32876 );
and ( n33026 , n33022 , n33025 );
and ( n33027 , n33018 , n33025 );
or ( n33028 , n33023 , n33026 , n33027 );
xor ( n33029 , n32959 , n32963 );
xor ( n33030 , n33029 , n32966 );
and ( n33031 , n33028 , n33030 );
xor ( n33032 , n32879 , n32883 );
xor ( n33033 , n33032 , n32886 );
and ( n33034 , n33030 , n33033 );
and ( n33035 , n33028 , n33033 );
or ( n33036 , n33031 , n33034 , n33035 );
and ( n33037 , n32983 , n33036 );
xor ( n33038 , n32915 , n32977 );
and ( n33039 , n33037 , n33038 );
xor ( n33040 , n33037 , n33038 );
xor ( n33041 , n32918 , n32920 );
and ( n33042 , n32440 , n30770 );
and ( n33043 , n32345 , n30768 );
nor ( n33044 , n33042 , n33043 );
xnor ( n33045 , n33044 , n30752 );
and ( n33046 , n33041 , n33045 );
and ( n33047 , n32501 , n30691 );
not ( n33048 , n33047 );
xnor ( n33049 , n33048 , n30696 );
and ( n33050 , n33045 , n33049 );
and ( n33051 , n33041 , n33049 );
or ( n33052 , n33046 , n33050 , n33051 );
and ( n33053 , n32195 , n30911 );
and ( n33054 , n32110 , n30909 );
nor ( n33055 , n33053 , n33054 );
xnor ( n33056 , n33055 , n30848 );
and ( n33057 , n33052 , n33056 );
xor ( n33058 , n32987 , n32990 );
xor ( n33059 , n33058 , n32993 );
and ( n33060 , n33056 , n33059 );
and ( n33061 , n33052 , n33059 );
or ( n33062 , n33057 , n33060 , n33061 );
and ( n33063 , n31823 , n31220 );
and ( n33064 , n31741 , n31218 );
nor ( n33065 , n33063 , n33064 );
xnor ( n33066 , n33065 , n31154 );
and ( n33067 , n33062 , n33066 );
xor ( n33068 , n32996 , n33000 );
xor ( n33069 , n33068 , n33003 );
and ( n33070 , n33066 , n33069 );
and ( n33071 , n33062 , n33069 );
or ( n33072 , n33067 , n33070 , n33071 );
and ( n33073 , n31645 , n31354 );
and ( n33074 , n31560 , n31351 );
nor ( n33075 , n33073 , n33074 );
xnor ( n33076 , n33075 , n31146 );
and ( n33077 , n33072 , n33076 );
xor ( n33078 , n32937 , n32941 );
xor ( n33079 , n33078 , n32944 );
and ( n33080 , n33076 , n33079 );
and ( n33081 , n33072 , n33079 );
or ( n33082 , n33077 , n33080 , n33081 );
xor ( n33083 , n32947 , n32951 );
xor ( n33084 , n33083 , n32956 );
and ( n33085 , n33082 , n33084 );
xor ( n33086 , n33018 , n33022 );
xor ( n33087 , n33086 , n33025 );
and ( n33088 , n33084 , n33087 );
and ( n33089 , n33082 , n33087 );
or ( n33090 , n33085 , n33088 , n33089 );
xor ( n33091 , n33028 , n33030 );
xor ( n33092 , n33091 , n33033 );
and ( n33093 , n33090 , n33092 );
xor ( n33094 , n32983 , n33036 );
and ( n33095 , n33093 , n33094 );
xor ( n33096 , n33093 , n33094 );
xor ( n33097 , n33090 , n33092 );
xor ( n33098 , n33082 , n33084 );
xor ( n33099 , n33098 , n33087 );
and ( n33100 , n32501 , n30768 );
not ( n33101 , n33100 );
and ( n33102 , n33101 , n30752 );
buf ( n33103 , n800 );
buf ( n33104 , n33103 );
and ( n33105 , n33102 , n33104 );
and ( n33106 , n33105 , n32916 );
buf ( n33107 , n799 );
buf ( n33108 , n33107 );
and ( n33109 , n32916 , n33108 );
and ( n33110 , n33105 , n33108 );
or ( n33111 , n33106 , n33109 , n33110 );
and ( n33112 , n32278 , n30911 );
and ( n33113 , n32195 , n30909 );
nor ( n33114 , n33112 , n33113 );
xnor ( n33115 , n33114 , n30848 );
and ( n33116 , n33111 , n33115 );
xor ( n33117 , n33041 , n33045 );
xor ( n33118 , n33117 , n33049 );
and ( n33119 , n33115 , n33118 );
and ( n33120 , n33111 , n33118 );
or ( n33121 , n33116 , n33119 , n33120 );
and ( n33122 , n32071 , n30975 );
and ( n33123 , n31966 , n30973 );
nor ( n33124 , n33122 , n33123 );
xnor ( n33125 , n33124 , n30957 );
and ( n33126 , n33121 , n33125 );
xor ( n33127 , n33052 , n33056 );
xor ( n33128 , n33127 , n33059 );
and ( n33129 , n33125 , n33128 );
and ( n33130 , n33121 , n33128 );
or ( n33131 , n33126 , n33129 , n33130 );
and ( n33132 , n31684 , n31354 );
and ( n33133 , n31645 , n31351 );
nor ( n33134 , n33132 , n33133 );
xnor ( n33135 , n33134 , n31146 );
and ( n33136 , n33131 , n33135 );
and ( n33137 , n31966 , n30975 );
and ( n33138 , n31864 , n30973 );
nor ( n33139 , n33137 , n33138 );
xnor ( n33140 , n33139 , n30957 );
and ( n33141 , n33135 , n33140 );
and ( n33142 , n33131 , n33140 );
or ( n33143 , n33136 , n33141 , n33142 );
xor ( n33144 , n33006 , n33010 );
xor ( n33145 , n33144 , n33015 );
and ( n33146 , n33143 , n33145 );
xor ( n33147 , n33072 , n33076 );
xor ( n33148 , n33147 , n33079 );
and ( n33149 , n33145 , n33148 );
and ( n33150 , n33143 , n33148 );
or ( n33151 , n33146 , n33149 , n33150 );
and ( n33152 , n33099 , n33151 );
xor ( n33153 , n33099 , n33151 );
xor ( n33154 , n33143 , n33145 );
xor ( n33155 , n33154 , n33148 );
and ( n33156 , n32345 , n30911 );
and ( n33157 , n32278 , n30909 );
nor ( n33158 , n33156 , n33157 );
xnor ( n33159 , n33158 , n30848 );
and ( n33160 , n32440 , n30768 );
not ( n33161 , n33160 );
xnor ( n33162 , n33161 , n30752 );
and ( n33163 , n33159 , n33162 );
xor ( n33164 , n33105 , n32916 );
xor ( n33165 , n33164 , n33108 );
and ( n33166 , n33162 , n33165 );
and ( n33167 , n33159 , n33165 );
or ( n33168 , n33163 , n33166 , n33167 );
and ( n33169 , n32110 , n30975 );
and ( n33170 , n32071 , n30973 );
nor ( n33171 , n33169 , n33170 );
xnor ( n33172 , n33171 , n30957 );
and ( n33173 , n33168 , n33172 );
xor ( n33174 , n33111 , n33115 );
xor ( n33175 , n33174 , n33118 );
and ( n33176 , n33172 , n33175 );
and ( n33177 , n33168 , n33175 );
or ( n33178 , n33173 , n33176 , n33177 );
and ( n33179 , n31741 , n31354 );
and ( n33180 , n31684 , n31351 );
nor ( n33181 , n33179 , n33180 );
xnor ( n33182 , n33181 , n31146 );
and ( n33183 , n33178 , n33182 );
and ( n33184 , n31864 , n31220 );
and ( n33185 , n31823 , n31218 );
nor ( n33186 , n33184 , n33185 );
xnor ( n33187 , n33186 , n31154 );
and ( n33188 , n33182 , n33187 );
and ( n33189 , n33178 , n33187 );
or ( n33190 , n33183 , n33188 , n33189 );
xor ( n33191 , n33131 , n33135 );
xor ( n33192 , n33191 , n33140 );
and ( n33193 , n33190 , n33192 );
xor ( n33194 , n33062 , n33066 );
xor ( n33195 , n33194 , n33069 );
and ( n33196 , n33192 , n33195 );
and ( n33197 , n33190 , n33195 );
or ( n33198 , n33193 , n33196 , n33197 );
and ( n33199 , n33155 , n33198 );
xor ( n33200 , n33155 , n33198 );
xor ( n33201 , n33102 , n33104 );
and ( n33202 , n32501 , n30909 );
not ( n33203 , n33202 );
and ( n33204 , n33203 , n30848 );
buf ( n33205 , n802 );
buf ( n33206 , n33205 );
and ( n33207 , n33204 , n33206 );
and ( n33208 , n33207 , n33100 );
buf ( n33209 , n801 );
buf ( n33210 , n33209 );
and ( n33211 , n33100 , n33210 );
and ( n33212 , n33207 , n33210 );
or ( n33213 , n33208 , n33211 , n33212 );
and ( n33214 , n33201 , n33213 );
and ( n33215 , n32501 , n30770 );
not ( n33216 , n33215 );
xnor ( n33217 , n33216 , n30752 );
and ( n33218 , n33213 , n33217 );
and ( n33219 , n33201 , n33217 );
or ( n33220 , n33214 , n33218 , n33219 );
and ( n33221 , n32195 , n30975 );
and ( n33222 , n32110 , n30973 );
nor ( n33223 , n33221 , n33222 );
xnor ( n33224 , n33223 , n30957 );
and ( n33225 , n33220 , n33224 );
xor ( n33226 , n33159 , n33162 );
xor ( n33227 , n33226 , n33165 );
and ( n33228 , n33224 , n33227 );
and ( n33229 , n33220 , n33227 );
or ( n33230 , n33225 , n33228 , n33229 );
and ( n33231 , n31966 , n31220 );
and ( n33232 , n31864 , n31218 );
nor ( n33233 , n33231 , n33232 );
xnor ( n33234 , n33233 , n31154 );
and ( n33235 , n33230 , n33234 );
xor ( n33236 , n33168 , n33172 );
xor ( n33237 , n33236 , n33175 );
and ( n33238 , n33234 , n33237 );
and ( n33239 , n33230 , n33237 );
or ( n33240 , n33235 , n33238 , n33239 );
xor ( n33241 , n33178 , n33182 );
xor ( n33242 , n33241 , n33187 );
and ( n33243 , n33240 , n33242 );
xor ( n33244 , n33121 , n33125 );
xor ( n33245 , n33244 , n33128 );
and ( n33246 , n33242 , n33245 );
and ( n33247 , n33240 , n33245 );
or ( n33248 , n33243 , n33246 , n33247 );
xor ( n33249 , n33190 , n33192 );
xor ( n33250 , n33249 , n33195 );
and ( n33251 , n33248 , n33250 );
xor ( n33252 , n33248 , n33250 );
xor ( n33253 , n33240 , n33242 );
xor ( n33254 , n33253 , n33245 );
and ( n33255 , n32278 , n30975 );
and ( n33256 , n32195 , n30973 );
nor ( n33257 , n33255 , n33256 );
xnor ( n33258 , n33257 , n30957 );
and ( n33259 , n32440 , n30911 );
and ( n33260 , n32345 , n30909 );
nor ( n33261 , n33259 , n33260 );
xnor ( n33262 , n33261 , n30848 );
and ( n33263 , n33258 , n33262 );
xor ( n33264 , n33201 , n33213 );
xor ( n33265 , n33264 , n33217 );
and ( n33266 , n33262 , n33265 );
and ( n33267 , n33258 , n33265 );
or ( n33268 , n33263 , n33266 , n33267 );
and ( n33269 , n32071 , n31220 );
and ( n33270 , n31966 , n31218 );
nor ( n33271 , n33269 , n33270 );
xnor ( n33272 , n33271 , n31154 );
and ( n33273 , n33268 , n33272 );
xor ( n33274 , n33220 , n33224 );
xor ( n33275 , n33274 , n33227 );
and ( n33276 , n33272 , n33275 );
and ( n33277 , n33268 , n33275 );
or ( n33278 , n33273 , n33276 , n33277 );
and ( n33279 , n31823 , n31354 );
and ( n33280 , n31741 , n31351 );
nor ( n33281 , n33279 , n33280 );
xnor ( n33282 , n33281 , n31146 );
and ( n33283 , n33278 , n33282 );
xor ( n33284 , n33230 , n33234 );
xor ( n33285 , n33284 , n33237 );
and ( n33286 , n33282 , n33285 );
and ( n33287 , n33278 , n33285 );
or ( n33288 , n33283 , n33286 , n33287 );
and ( n33289 , n33254 , n33288 );
xor ( n33290 , n33254 , n33288 );
xor ( n33291 , n33278 , n33282 );
xor ( n33292 , n33291 , n33285 );
and ( n33293 , n32345 , n30975 );
and ( n33294 , n32278 , n30973 );
nor ( n33295 , n33293 , n33294 );
xnor ( n33296 , n33295 , n30957 );
and ( n33297 , n32440 , n30909 );
not ( n33298 , n33297 );
xnor ( n33299 , n33298 , n30848 );
and ( n33300 , n33296 , n33299 );
xor ( n33301 , n33207 , n33100 );
xor ( n33302 , n33301 , n33210 );
and ( n33303 , n33299 , n33302 );
and ( n33304 , n33296 , n33302 );
or ( n33305 , n33300 , n33303 , n33304 );
and ( n33306 , n32110 , n31220 );
and ( n33307 , n32071 , n31218 );
nor ( n33308 , n33306 , n33307 );
xnor ( n33309 , n33308 , n31154 );
and ( n33310 , n33305 , n33309 );
xor ( n33311 , n33258 , n33262 );
xor ( n33312 , n33311 , n33265 );
and ( n33313 , n33309 , n33312 );
and ( n33314 , n33305 , n33312 );
or ( n33315 , n33310 , n33313 , n33314 );
and ( n33316 , n31864 , n31354 );
and ( n33317 , n31823 , n31351 );
nor ( n33318 , n33316 , n33317 );
xnor ( n33319 , n33318 , n31146 );
and ( n33320 , n33315 , n33319 );
xor ( n33321 , n33268 , n33272 );
xor ( n33322 , n33321 , n33275 );
and ( n33323 , n33319 , n33322 );
and ( n33324 , n33315 , n33322 );
or ( n33325 , n33320 , n33323 , n33324 );
and ( n33326 , n33292 , n33325 );
xor ( n33327 , n33292 , n33325 );
xor ( n33328 , n33315 , n33319 );
xor ( n33329 , n33328 , n33322 );
xor ( n33330 , n33204 , n33206 );
and ( n33331 , n32440 , n30975 );
and ( n33332 , n32345 , n30973 );
nor ( n33333 , n33331 , n33332 );
xnor ( n33334 , n33333 , n30957 );
and ( n33335 , n33330 , n33334 );
and ( n33336 , n32501 , n30911 );
not ( n33337 , n33336 );
xnor ( n33338 , n33337 , n30848 );
and ( n33339 , n33334 , n33338 );
and ( n33340 , n33330 , n33338 );
or ( n33341 , n33335 , n33339 , n33340 );
and ( n33342 , n32195 , n31220 );
and ( n33343 , n32110 , n31218 );
nor ( n33344 , n33342 , n33343 );
xnor ( n33345 , n33344 , n31154 );
and ( n33346 , n33341 , n33345 );
xor ( n33347 , n33296 , n33299 );
xor ( n33348 , n33347 , n33302 );
and ( n33349 , n33345 , n33348 );
and ( n33350 , n33341 , n33348 );
or ( n33351 , n33346 , n33349 , n33350 );
and ( n33352 , n31966 , n31354 );
and ( n33353 , n31864 , n31351 );
nor ( n33354 , n33352 , n33353 );
xnor ( n33355 , n33354 , n31146 );
and ( n33356 , n33351 , n33355 );
xor ( n33357 , n33305 , n33309 );
xor ( n33358 , n33357 , n33312 );
and ( n33359 , n33355 , n33358 );
and ( n33360 , n33351 , n33358 );
or ( n33361 , n33356 , n33359 , n33360 );
and ( n33362 , n33329 , n33361 );
xor ( n33363 , n33329 , n33361 );
and ( n33364 , n32501 , n30973 );
not ( n33365 , n33364 );
and ( n33366 , n33365 , n30957 );
buf ( n33367 , n804 );
buf ( n33368 , n33367 );
and ( n33369 , n33366 , n33368 );
and ( n33370 , n33369 , n33202 );
buf ( n33371 , n803 );
buf ( n33372 , n33371 );
and ( n33373 , n33202 , n33372 );
and ( n33374 , n33369 , n33372 );
or ( n33375 , n33370 , n33373 , n33374 );
and ( n33376 , n32278 , n31220 );
and ( n33377 , n32195 , n31218 );
nor ( n33378 , n33376 , n33377 );
xnor ( n33379 , n33378 , n31154 );
and ( n33380 , n33375 , n33379 );
xor ( n33381 , n33330 , n33334 );
xor ( n33382 , n33381 , n33338 );
and ( n33383 , n33379 , n33382 );
and ( n33384 , n33375 , n33382 );
or ( n33385 , n33380 , n33383 , n33384 );
and ( n33386 , n32071 , n31354 );
and ( n33387 , n31966 , n31351 );
nor ( n33388 , n33386 , n33387 );
xnor ( n33389 , n33388 , n31146 );
and ( n33390 , n33385 , n33389 );
xor ( n33391 , n33341 , n33345 );
xor ( n33392 , n33391 , n33348 );
and ( n33393 , n33389 , n33392 );
and ( n33394 , n33385 , n33392 );
or ( n33395 , n33390 , n33393 , n33394 );
xor ( n33396 , n33351 , n33355 );
xor ( n33397 , n33396 , n33358 );
and ( n33398 , n33395 , n33397 );
xor ( n33399 , n33395 , n33397 );
and ( n33400 , n32345 , n31220 );
and ( n33401 , n32278 , n31218 );
nor ( n33402 , n33400 , n33401 );
xnor ( n33403 , n33402 , n31154 );
and ( n33404 , n32440 , n30973 );
not ( n33405 , n33404 );
xnor ( n33406 , n33405 , n30957 );
and ( n33407 , n33403 , n33406 );
xor ( n33408 , n33369 , n33202 );
xor ( n33409 , n33408 , n33372 );
and ( n33410 , n33406 , n33409 );
and ( n33411 , n33403 , n33409 );
or ( n33412 , n33407 , n33410 , n33411 );
and ( n33413 , n32110 , n31354 );
and ( n33414 , n32071 , n31351 );
nor ( n33415 , n33413 , n33414 );
xnor ( n33416 , n33415 , n31146 );
and ( n33417 , n33412 , n33416 );
xor ( n33418 , n33375 , n33379 );
xor ( n33419 , n33418 , n33382 );
and ( n33420 , n33416 , n33419 );
and ( n33421 , n33412 , n33419 );
or ( n33422 , n33417 , n33420 , n33421 );
xor ( n33423 , n33385 , n33389 );
xor ( n33424 , n33423 , n33392 );
and ( n33425 , n33422 , n33424 );
xor ( n33426 , n33422 , n33424 );
xor ( n33427 , n33412 , n33416 );
xor ( n33428 , n33427 , n33419 );
xor ( n33429 , n33366 , n33368 );
and ( n33430 , n32501 , n31218 );
not ( n33431 , n33430 );
and ( n33432 , n33431 , n31154 );
buf ( n33433 , n806 );
buf ( n33434 , n33433 );
and ( n33435 , n33432 , n33434 );
and ( n33436 , n33435 , n33364 );
buf ( n33437 , n805 );
buf ( n33438 , n33437 );
and ( n33439 , n33364 , n33438 );
and ( n33440 , n33435 , n33438 );
or ( n33441 , n33436 , n33439 , n33440 );
and ( n33442 , n33429 , n33441 );
and ( n33443 , n32501 , n30975 );
not ( n33444 , n33443 );
xnor ( n33445 , n33444 , n30957 );
and ( n33446 , n33441 , n33445 );
and ( n33447 , n33429 , n33445 );
or ( n33448 , n33442 , n33446 , n33447 );
and ( n33449 , n32195 , n31354 );
and ( n33450 , n32110 , n31351 );
nor ( n33451 , n33449 , n33450 );
xnor ( n33452 , n33451 , n31146 );
and ( n33453 , n33448 , n33452 );
xor ( n33454 , n33403 , n33406 );
xor ( n33455 , n33454 , n33409 );
and ( n33456 , n33452 , n33455 );
and ( n33457 , n33448 , n33455 );
or ( n33458 , n33453 , n33456 , n33457 );
and ( n33459 , n33428 , n33458 );
xor ( n33460 , n33428 , n33458 );
xor ( n33461 , n33448 , n33452 );
xor ( n33462 , n33461 , n33455 );
and ( n33463 , n32278 , n31354 );
and ( n33464 , n32195 , n31351 );
nor ( n33465 , n33463 , n33464 );
xnor ( n33466 , n33465 , n31146 );
and ( n33467 , n32440 , n31220 );
and ( n33468 , n32345 , n31218 );
nor ( n33469 , n33467 , n33468 );
xnor ( n33470 , n33469 , n31154 );
and ( n33471 , n33466 , n33470 );
xor ( n33472 , n33429 , n33441 );
xor ( n33473 , n33472 , n33445 );
and ( n33474 , n33470 , n33473 );
and ( n33475 , n33466 , n33473 );
or ( n33476 , n33471 , n33474 , n33475 );
and ( n33477 , n33462 , n33476 );
xor ( n33478 , n33462 , n33476 );
and ( n33479 , n32345 , n31354 );
and ( n33480 , n32278 , n31351 );
nor ( n33481 , n33479 , n33480 );
xnor ( n33482 , n33481 , n31146 );
and ( n33483 , n32440 , n31218 );
not ( n33484 , n33483 );
xnor ( n33485 , n33484 , n31154 );
and ( n33486 , n33482 , n33485 );
xor ( n33487 , n33435 , n33364 );
xor ( n33488 , n33487 , n33438 );
and ( n33489 , n33485 , n33488 );
and ( n33490 , n33482 , n33488 );
or ( n33491 , n33486 , n33489 , n33490 );
xor ( n33492 , n33466 , n33470 );
xor ( n33493 , n33492 , n33473 );
and ( n33494 , n33491 , n33493 );
xor ( n33495 , n33491 , n33493 );
xor ( n33496 , n33432 , n33434 );
and ( n33497 , n32440 , n31354 );
and ( n33498 , n32345 , n31351 );
nor ( n33499 , n33497 , n33498 );
xnor ( n33500 , n33499 , n31146 );
and ( n33501 , n33496 , n33500 );
and ( n33502 , n32501 , n31220 );
not ( n33503 , n33502 );
xnor ( n33504 , n33503 , n31154 );
and ( n33505 , n33500 , n33504 );
and ( n33506 , n33496 , n33504 );
or ( n33507 , n33501 , n33505 , n33506 );
xor ( n33508 , n33482 , n33485 );
xor ( n33509 , n33508 , n33488 );
and ( n33510 , n33507 , n33509 );
xor ( n33511 , n33507 , n33509 );
xor ( n33512 , n33496 , n33500 );
xor ( n33513 , n33512 , n33504 );
buf ( n33514 , n32501 );
not ( n33515 , n33514 );
and ( n33516 , n33515 , n31146 );
buf ( n33517 , n808 );
buf ( n33518 , n33517 );
and ( n33519 , n33516 , n33518 );
and ( n33520 , n33519 , n33430 );
buf ( n33521 , n807 );
buf ( n33522 , n33521 );
and ( n33523 , n33430 , n33522 );
and ( n33524 , n33519 , n33522 );
or ( n33525 , n33520 , n33523 , n33524 );
and ( n33526 , n33513 , n33525 );
xor ( n33527 , n33513 , n33525 );
and ( n33528 , n32440 , n31351 );
not ( n33529 , n33528 );
xnor ( n33530 , n33529 , n31146 );
xor ( n33531 , n33519 , n33430 );
xor ( n33532 , n33531 , n33522 );
and ( n33533 , n33530 , n33532 );
xor ( n33534 , n33530 , n33532 );
and ( n33535 , n32501 , n31354 );
not ( n33536 , n33535 );
xnor ( n33537 , n33536 , n31146 );
xor ( n33538 , n33516 , n33518 );
and ( n33539 , n33537 , n33538 );
xor ( n33540 , n33537 , n33538 );
buf ( n33541 , n809 );
buf ( n33542 , n33541 );
and ( n33543 , n33514 , n33542 );
and ( n33544 , n33540 , n33543 );
or ( n33545 , n33539 , n33544 );
and ( n33546 , n33534 , n33545 );
or ( n33547 , n33533 , n33546 );
and ( n33548 , n33527 , n33547 );
or ( n33549 , n33526 , n33548 );
and ( n33550 , n33511 , n33549 );
or ( n33551 , n33510 , n33550 );
and ( n33552 , n33495 , n33551 );
or ( n33553 , n33494 , n33552 );
and ( n33554 , n33478 , n33553 );
or ( n33555 , n33477 , n33554 );
and ( n33556 , n33460 , n33555 );
or ( n33557 , n33459 , n33556 );
and ( n33558 , n33426 , n33557 );
or ( n33559 , n33425 , n33558 );
and ( n33560 , n33399 , n33559 );
or ( n33561 , n33398 , n33560 );
and ( n33562 , n33363 , n33561 );
or ( n33563 , n33362 , n33562 );
and ( n33564 , n33327 , n33563 );
or ( n33565 , n33326 , n33564 );
and ( n33566 , n33290 , n33565 );
or ( n33567 , n33289 , n33566 );
and ( n33568 , n33252 , n33567 );
or ( n33569 , n33251 , n33568 );
and ( n33570 , n33200 , n33569 );
or ( n33571 , n33199 , n33570 );
and ( n33572 , n33153 , n33571 );
or ( n33573 , n33152 , n33572 );
and ( n33574 , n33097 , n33573 );
and ( n33575 , n33096 , n33574 );
or ( n33576 , n33095 , n33575 );
and ( n33577 , n33040 , n33576 );
or ( n33578 , n33039 , n33577 );
and ( n33579 , n32981 , n33578 );
or ( n33580 , n32980 , n33579 );
and ( n33581 , n32913 , n33580 );
or ( n33582 , n32912 , n33581 );
and ( n33583 , n32847 , n33582 );
or ( n33584 , n32846 , n33583 );
and ( n33585 , n32778 , n33584 );
or ( n33586 , n32777 , n33585 );
and ( n33587 , n32702 , n33586 );
or ( n33588 , n32701 , n33587 );
and ( n33589 , n32632 , n33588 );
or ( n33590 , n32631 , n33589 );
and ( n33591 , n32494 , n33590 );
or ( n33592 , n32493 , n33591 );
and ( n33593 , n32425 , n33592 );
or ( n33594 , n32424 , n33593 );
and ( n33595 , n32330 , n33594 );
or ( n33596 , n32329 , n33595 );
and ( n33597 , n32247 , n33596 );
or ( n33598 , n32246 , n33597 );
and ( n33599 , n32164 , n33598 );
or ( n33600 , n32163 , n33599 );
and ( n33601 , n32056 , n33600 );
or ( n33602 , n32055 , n33601 );
and ( n33603 , n31951 , n33602 );
or ( n33604 , n31950 , n33603 );
and ( n33605 , n31927 , n33604 );
or ( n33606 , n31926 , n33605 );
and ( n33607 , n31807 , n33606 );
or ( n33608 , n31806 , n33607 );
and ( n33609 , n31726 , n33608 );
or ( n33610 , n31725 , n33609 );
and ( n33611 , n31630 , n33610 );
or ( n33612 , n31629 , n33611 );
and ( n33613 , n31547 , n33612 );
or ( n33614 , n31546 , n33613 );
and ( n33615 , n31463 , n33614 );
and ( n33616 , n31461 , n33615 );
and ( n33617 , n31459 , n33616 );
and ( n33618 , n31457 , n33617 );
and ( n33619 , n31455 , n33618 );
and ( n33620 , n31453 , n33619 );
and ( n33621 , n31451 , n33620 );
and ( n33622 , n31449 , n33621 );
and ( n33623 , n31447 , n33622 );
and ( n33624 , n31445 , n33623 );
xor ( n33625 , n31443 , n33624 );
buf ( n33626 , n33625 );
buf ( n33627 , n33626 );
buf ( n33628 , n33627 );
xor ( n33629 , n28117 , n28119 );
xor ( n33630 , n28119 , n28121 );
not ( n33631 , n33630 );
and ( n33632 , n33629 , n33631 );
and ( n33633 , n33628 , n33632 );
not ( n33634 , n33633 );
xnor ( n33635 , n33634 , n28124 );
and ( n33636 , n28536 , n33635 );
and ( n33637 , n28535 , n33635 );
or ( n33638 , n28537 , n33636 , n33637 );
and ( n33639 , n28534 , n33638 );
xor ( n33640 , n28316 , n28317 );
xor ( n33641 , n33640 , n28319 );
and ( n33642 , n33638 , n33641 );
and ( n33643 , n28534 , n33641 );
or ( n33644 , n33639 , n33642 , n33643 );
and ( n33645 , n28524 , n33644 );
xor ( n33646 , n28289 , n28291 );
xor ( n33647 , n33646 , n28293 );
and ( n33648 , n33644 , n33647 );
and ( n33649 , n28524 , n33647 );
or ( n33650 , n33645 , n33648 , n33649 );
and ( n33651 , n28509 , n33650 );
and ( n33652 , n28493 , n33650 );
or ( n33653 , n28510 , n33651 , n33652 );
and ( n33654 , n28485 , n33653 );
xor ( n33655 , n28255 , n28257 );
xor ( n33656 , n33655 , n28260 );
and ( n33657 , n33653 , n33656 );
and ( n33658 , n28485 , n33656 );
or ( n33659 , n33654 , n33657 , n33658 );
and ( n33660 , n28475 , n33659 );
xor ( n33661 , n28158 , n28160 );
xor ( n33662 , n33661 , n28163 );
and ( n33663 , n33659 , n33662 );
and ( n33664 , n28475 , n33662 );
or ( n33665 , n33660 , n33663 , n33664 );
xor ( n33666 , n28097 , n28098 );
xor ( n33667 , n33666 , n28166 );
and ( n33668 , n33665 , n33667 );
xor ( n33669 , n28235 , n28352 );
xor ( n33670 , n33669 , n28355 );
and ( n33671 , n33667 , n33670 );
and ( n33672 , n33665 , n33670 );
or ( n33673 , n33668 , n33671 , n33672 );
xor ( n33674 , n28169 , n28358 );
xor ( n33675 , n33674 , n28361 );
and ( n33676 , n33673 , n33675 );
xor ( n33677 , n28170 , n28171 );
xor ( n33678 , n33677 , n28232 );
xor ( n33679 , n28253 , n28263 );
xor ( n33680 , n33679 , n28349 );
and ( n33681 , n33678 , n33680 );
xor ( n33682 , n28277 , n28299 );
xor ( n33683 , n33682 , n28346 );
xor ( n33684 , n28279 , n28287 );
xor ( n33685 , n33684 , n28296 );
xor ( n33686 , n28325 , n28340 );
xor ( n33687 , n33686 , n28343 );
and ( n33688 , n33685 , n33687 );
xor ( n33689 , n28458 , n28460 );
xor ( n33690 , n33689 , n28463 );
and ( n33691 , n33687 , n33690 );
and ( n33692 , n33685 , n33690 );
or ( n33693 , n33688 , n33691 , n33692 );
and ( n33694 , n33683 , n33693 );
xnor ( n33695 , n28469 , n28471 );
xor ( n33696 , n28307 , n28314 );
xor ( n33697 , n33696 , n28322 );
xor ( n33698 , n28332 , n28334 );
xor ( n33699 , n33698 , n28337 );
and ( n33700 , n33697 , n33699 );
xor ( n33701 , n28486 , n28487 );
xor ( n33702 , n33701 , n28490 );
and ( n33703 , n33699 , n33702 );
and ( n33704 , n33697 , n33702 );
or ( n33705 , n33700 , n33703 , n33704 );
and ( n33706 , n33695 , n33705 );
xor ( n33707 , n28451 , n28452 );
xor ( n33708 , n33707 , n28455 );
and ( n33709 , n24052 , n25026 );
and ( n33710 , n23620 , n26229 );
and ( n33711 , n33709 , n33710 );
and ( n33712 , n23483 , n26376 );
and ( n33713 , n33710 , n33712 );
and ( n33714 , n33709 , n33712 );
or ( n33715 , n33711 , n33713 , n33714 );
and ( n33716 , n25742 , n22172 );
xor ( n33717 , n33715 , n33716 );
and ( n33718 , n25623 , n22337 );
xor ( n33719 , n33717 , n33718 );
xor ( n33720 , n28444 , n28445 );
xor ( n33721 , n33720 , n28448 );
and ( n33722 , n33719 , n33721 );
and ( n33723 , n26980 , n21178 );
and ( n33724 , n26678 , n21527 );
xor ( n33725 , n33723 , n33724 );
xor ( n33726 , n28205 , n28206 );
xor ( n33727 , n33726 , n28211 );
xor ( n33728 , n33725 , n33727 );
and ( n33729 , n33721 , n33728 );
and ( n33730 , n33719 , n33728 );
or ( n33731 , n33722 , n33729 , n33730 );
and ( n33732 , n33708 , n33731 );
xor ( n33733 , n28326 , n28327 );
xor ( n33734 , n33733 , n28329 );
and ( n33735 , n23742 , n26229 );
and ( n33736 , n23483 , n26876 );
and ( n33737 , n33735 , n33736 );
buf ( n33738 , n11378 );
buf ( n33739 , n33738 );
and ( n33740 , n22936 , n33739 );
not ( n33741 , n33740 );
and ( n33742 , n33736 , n33741 );
and ( n33743 , n33735 , n33741 );
or ( n33744 , n33737 , n33742 , n33743 );
and ( n33745 , n25959 , n22172 );
and ( n33746 , n33744 , n33745 );
and ( n33747 , n25742 , n22337 );
and ( n33748 , n33745 , n33747 );
and ( n33749 , n33744 , n33747 );
or ( n33750 , n33746 , n33748 , n33749 );
and ( n33751 , n33734 , n33750 );
and ( n33752 , n26980 , n21296 );
and ( n33753 , n26399 , n21827 );
and ( n33754 , n33752 , n33753 );
xor ( n33755 , n33709 , n33710 );
xor ( n33756 , n33755 , n33712 );
and ( n33757 , n33753 , n33756 );
and ( n33758 , n33752 , n33756 );
or ( n33759 , n33754 , n33757 , n33758 );
and ( n33760 , n33750 , n33759 );
and ( n33761 , n33734 , n33759 );
or ( n33762 , n33751 , n33760 , n33761 );
and ( n33763 , n33731 , n33762 );
and ( n33764 , n33708 , n33762 );
or ( n33765 , n33732 , n33763 , n33764 );
and ( n33766 , n33705 , n33765 );
and ( n33767 , n33695 , n33765 );
or ( n33768 , n33706 , n33766 , n33767 );
and ( n33769 , n33693 , n33768 );
and ( n33770 , n33683 , n33768 );
or ( n33771 , n33694 , n33769 , n33770 );
and ( n33772 , n33680 , n33771 );
and ( n33773 , n33678 , n33771 );
or ( n33774 , n33681 , n33772 , n33773 );
and ( n33775 , n23215 , n27246 );
xnor ( n33776 , n28519 , n28520 );
or ( n33777 , n33775 , n33776 );
and ( n33778 , n22824 , n33739 );
not ( n33779 , n33778 );
xor ( n33780 , n28525 , n28533 );
and ( n33781 , n33779 , n33780 );
and ( n33782 , n33777 , n33781 );
buf ( n33783 , n33778 );
and ( n33784 , n33781 , n33783 );
and ( n33785 , n33777 , n33783 );
or ( n33786 , n33782 , n33784 , n33785 );
xor ( n33787 , n28511 , n28512 );
xor ( n33788 , n33787 , n28514 );
and ( n33789 , n27591 , n21178 );
and ( n33790 , n26933 , n21527 );
and ( n33791 , n33789 , n33790 );
and ( n33792 , n26782 , n21666 );
and ( n33793 , n33790 , n33792 );
and ( n33794 , n33789 , n33792 );
or ( n33795 , n33791 , n33793 , n33794 );
and ( n33796 , n33788 , n33795 );
and ( n33797 , n27389 , n21296 );
and ( n33798 , n26980 , n21429 );
and ( n33799 , n33797 , n33798 );
and ( n33800 , n26678 , n21827 );
and ( n33801 , n33798 , n33800 );
and ( n33802 , n33797 , n33800 );
or ( n33803 , n33799 , n33801 , n33802 );
and ( n33804 , n33795 , n33803 );
and ( n33805 , n33788 , n33803 );
or ( n33806 , n33796 , n33804 , n33805 );
xor ( n33807 , n28124 , n28517 );
xor ( n33808 , n33807 , n28521 );
and ( n33809 , n33806 , n33808 );
xor ( n33810 , n28534 , n33638 );
xor ( n33811 , n33810 , n33641 );
and ( n33812 , n33808 , n33811 );
and ( n33813 , n33806 , n33811 );
or ( n33814 , n33809 , n33812 , n33813 );
and ( n33815 , n33786 , n33814 );
xor ( n33816 , n28495 , n28497 );
xor ( n33817 , n33816 , n28506 );
and ( n33818 , n33814 , n33817 );
and ( n33819 , n33786 , n33817 );
or ( n33820 , n33815 , n33818 , n33819 );
xor ( n33821 , n28477 , n28479 );
xor ( n33822 , n33821 , n28482 );
and ( n33823 , n33820 , n33822 );
xor ( n33824 , n28493 , n28509 );
xor ( n33825 , n33824 , n33650 );
and ( n33826 , n33822 , n33825 );
and ( n33827 , n33820 , n33825 );
or ( n33828 , n33823 , n33826 , n33827 );
xor ( n33829 , n28389 , n28391 );
xor ( n33830 , n33829 , n28394 );
and ( n33831 , n33828 , n33830 );
xor ( n33832 , n28443 , n28466 );
xor ( n33833 , n33832 , n28472 );
and ( n33834 , n33830 , n33833 );
and ( n33835 , n33828 , n33833 );
or ( n33836 , n33831 , n33834 , n33835 );
xor ( n33837 , n28384 , n28386 );
xor ( n33838 , n33837 , n28397 );
and ( n33839 , n33836 , n33838 );
xor ( n33840 , n28475 , n33659 );
xor ( n33841 , n33840 , n33662 );
and ( n33842 , n33838 , n33841 );
and ( n33843 , n33836 , n33841 );
or ( n33844 , n33839 , n33842 , n33843 );
and ( n33845 , n33774 , n33844 );
xor ( n33846 , n28379 , n28381 );
xor ( n33847 , n33846 , n28400 );
and ( n33848 , n33844 , n33847 );
and ( n33849 , n33774 , n33847 );
or ( n33850 , n33845 , n33848 , n33849 );
and ( n33851 , n33675 , n33850 );
and ( n33852 , n33673 , n33850 );
or ( n33853 , n33676 , n33851 , n33852 );
xor ( n33854 , n28372 , n28406 );
xor ( n33855 , n33854 , n28409 );
and ( n33856 , n33853 , n33855 );
xor ( n33857 , n28374 , n28376 );
xor ( n33858 , n33857 , n28403 );
xor ( n33859 , n33665 , n33667 );
xor ( n33860 , n33859 , n33670 );
xor ( n33861 , n28485 , n33653 );
xor ( n33862 , n33861 , n33656 );
and ( n33863 , n33715 , n33716 );
and ( n33864 , n33716 , n33718 );
and ( n33865 , n33715 , n33718 );
or ( n33866 , n33863 , n33864 , n33865 );
buf ( n33867 , n33740 );
and ( n33868 , n23742 , n25617 );
and ( n33869 , n33867 , n33868 );
and ( n33870 , n23336 , n26876 );
and ( n33871 , n33868 , n33870 );
and ( n33872 , n33867 , n33870 );
or ( n33873 , n33869 , n33871 , n33872 );
and ( n33874 , n26933 , n21296 );
and ( n33875 , n33873 , n33874 );
and ( n33876 , n26148 , n21827 );
and ( n33877 , n33874 , n33876 );
and ( n33878 , n33873 , n33876 );
or ( n33879 , n33875 , n33877 , n33878 );
and ( n33880 , n33866 , n33879 );
xor ( n33881 , n28173 , n28174 );
xor ( n33882 , n33881 , n28176 );
and ( n33883 , n33879 , n33882 );
and ( n33884 , n33866 , n33882 );
or ( n33885 , n33880 , n33883 , n33884 );
and ( n33886 , n24337 , n24540 );
and ( n33887 , n23903 , n25284 );
and ( n33888 , n33886 , n33887 );
xor ( n33889 , n33779 , n33780 );
not ( n33890 , n33889 );
and ( n33891 , n33887 , n33890 );
and ( n33892 , n33886 , n33890 );
or ( n33893 , n33888 , n33891 , n33892 );
and ( n33894 , n28129 , n20890 );
and ( n33895 , n33893 , n33894 );
and ( n33896 , n27962 , n20909 );
and ( n33897 , n33894 , n33896 );
and ( n33898 , n33893 , n33896 );
or ( n33899 , n33895 , n33897 , n33898 );
and ( n33900 , n33723 , n33724 );
and ( n33901 , n33724 , n33727 );
and ( n33902 , n33723 , n33727 );
or ( n33903 , n33900 , n33901 , n33902 );
and ( n33904 , n33899 , n33903 );
xor ( n33905 , n28214 , n28215 );
xor ( n33906 , n33905 , n28217 );
and ( n33907 , n33903 , n33906 );
and ( n33908 , n33899 , n33906 );
or ( n33909 , n33904 , n33907 , n33908 );
and ( n33910 , n33885 , n33909 );
xor ( n33911 , n28204 , n28220 );
xor ( n33912 , n33911 , n28223 );
and ( n33913 , n33909 , n33912 );
and ( n33914 , n33885 , n33912 );
or ( n33915 , n33910 , n33913 , n33914 );
and ( n33916 , n33862 , n33915 );
and ( n33917 , n24993 , n23322 );
and ( n33918 , n24731 , n23508 );
and ( n33919 , n33917 , n33918 );
and ( n33920 , n24546 , n24064 );
and ( n33921 , n33918 , n33920 );
and ( n33922 , n33917 , n33920 );
or ( n33923 , n33919 , n33921 , n33922 );
and ( n33924 , n24337 , n25026 );
and ( n33925 , n23336 , n27246 );
and ( n33926 , n33924 , n33925 );
and ( n33927 , n23089 , n28209 );
and ( n33928 , n33925 , n33927 );
and ( n33929 , n33924 , n33927 );
or ( n33930 , n33926 , n33928 , n33929 );
and ( n33931 , n25623 , n22562 );
and ( n33932 , n33930 , n33931 );
and ( n33933 , n25220 , n22987 );
and ( n33934 , n33931 , n33933 );
and ( n33935 , n33930 , n33933 );
or ( n33936 , n33932 , n33934 , n33935 );
and ( n33937 , n33923 , n33936 );
and ( n33938 , n27389 , n21085 );
and ( n33939 , n33936 , n33938 );
and ( n33940 , n33923 , n33938 );
or ( n33941 , n33937 , n33939 , n33940 );
and ( n33942 , n23903 , n25617 );
and ( n33943 , n23620 , n26376 );
and ( n33944 , n33942 , n33943 );
and ( n33945 , n23215 , n27558 );
and ( n33946 , n33943 , n33945 );
and ( n33947 , n33942 , n33945 );
or ( n33948 , n33944 , n33946 , n33947 );
and ( n33949 , n28129 , n20909 );
and ( n33950 , n33948 , n33949 );
and ( n33951 , n25451 , n22784 );
and ( n33952 , n33949 , n33951 );
and ( n33953 , n33948 , n33951 );
or ( n33954 , n33950 , n33952 , n33953 );
xnor ( n33955 , n33775 , n33776 );
and ( n33956 , n27962 , n20949 );
and ( n33957 , n33955 , n33956 );
and ( n33958 , n24624 , n23758 );
and ( n33959 , n33956 , n33958 );
and ( n33960 , n33955 , n33958 );
or ( n33961 , n33957 , n33959 , n33960 );
and ( n33962 , n33954 , n33961 );
xor ( n33963 , n28308 , n28309 );
xor ( n33964 , n33963 , n28311 );
and ( n33965 , n33961 , n33964 );
and ( n33966 , n33954 , n33964 );
or ( n33967 , n33962 , n33965 , n33966 );
or ( n33968 , n33941 , n33967 );
xor ( n33969 , n28524 , n33644 );
xor ( n33970 , n33969 , n33647 );
xor ( n33971 , n33866 , n33879 );
xor ( n33972 , n33971 , n33882 );
and ( n33973 , n33970 , n33972 );
and ( n33974 , n28129 , n20949 );
and ( n33975 , n25220 , n23322 );
and ( n33976 , n33974 , n33975 );
and ( n33977 , n24731 , n23758 );
and ( n33978 , n33975 , n33977 );
and ( n33979 , n33974 , n33977 );
or ( n33980 , n33976 , n33978 , n33979 );
and ( n33981 , n23742 , n26376 );
and ( n33982 , n23215 , n28209 );
and ( n33983 , n33981 , n33982 );
and ( n33984 , n23089 , n33739 );
and ( n33985 , n33982 , n33984 );
and ( n33986 , n33981 , n33984 );
or ( n33987 , n33983 , n33985 , n33986 );
and ( n33988 , n24546 , n25026 );
and ( n33989 , n23483 , n27246 );
and ( n33990 , n33988 , n33989 );
and ( n33991 , n23336 , n27558 );
and ( n33992 , n33989 , n33991 );
and ( n33993 , n33988 , n33991 );
or ( n33994 , n33990 , n33992 , n33993 );
and ( n33995 , n33987 , n33994 );
and ( n33996 , n25742 , n22562 );
and ( n33997 , n33994 , n33996 );
and ( n33998 , n33987 , n33996 );
or ( n33999 , n33995 , n33997 , n33998 );
and ( n34000 , n33980 , n33999 );
and ( n34001 , n26933 , n21429 );
and ( n34002 , n33999 , n34001 );
and ( n34003 , n33980 , n34001 );
or ( n34004 , n34000 , n34002 , n34003 );
and ( n34005 , n25451 , n22987 );
and ( n34006 , n24993 , n23508 );
and ( n34007 , n34005 , n34006 );
and ( n34008 , n24624 , n24064 );
and ( n34009 , n34006 , n34008 );
and ( n34010 , n34005 , n34008 );
or ( n34011 , n34007 , n34009 , n34010 );
and ( n34012 , n27863 , n21039 );
and ( n34013 , n34011 , n34012 );
xor ( n34014 , n33867 , n33868 );
xor ( n34015 , n34014 , n33870 );
and ( n34016 , n34012 , n34015 );
and ( n34017 , n34011 , n34015 );
or ( n34018 , n34013 , n34016 , n34017 );
and ( n34019 , n34004 , n34018 );
xor ( n34020 , n28499 , n28500 );
xor ( n34021 , n34020 , n28503 );
and ( n34022 , n34018 , n34021 );
and ( n34023 , n34004 , n34021 );
or ( n34024 , n34019 , n34022 , n34023 );
and ( n34025 , n33972 , n34024 );
and ( n34026 , n33970 , n34024 );
or ( n34027 , n33973 , n34025 , n34026 );
and ( n34028 , n33968 , n34027 );
and ( n34029 , n33628 , n28117 );
xor ( n34030 , n33873 , n33874 );
xor ( n34031 , n34030 , n33876 );
or ( n34032 , n34029 , n34031 );
xor ( n34033 , n33719 , n33721 );
xor ( n34034 , n34033 , n33728 );
xor ( n34035 , n31445 , n33623 );
buf ( n34036 , n34035 );
buf ( n34037 , n34036 );
buf ( n34038 , n34037 );
and ( n34039 , n34038 , n28117 );
xor ( n34040 , n33752 , n33753 );
xor ( n34041 , n34040 , n33756 );
or ( n34042 , n34039 , n34041 );
and ( n34043 , n34034 , n34042 );
buf ( n34044 , n33889 );
and ( n34045 , n34042 , n34044 );
and ( n34046 , n34034 , n34044 );
or ( n34047 , n34043 , n34045 , n34046 );
and ( n34048 , n34032 , n34047 );
and ( n34049 , n26148 , n22172 );
and ( n34050 , n24546 , n24540 );
and ( n34051 , n34049 , n34050 );
and ( n34052 , n24052 , n25284 );
and ( n34053 , n34050 , n34052 );
and ( n34054 , n34049 , n34052 );
or ( n34055 , n34051 , n34053 , n34054 );
xor ( n34056 , n28535 , n28536 );
xor ( n34057 , n34056 , n33635 );
and ( n34058 , n34055 , n34057 );
and ( n34059 , n24731 , n24064 );
and ( n34060 , n24624 , n24540 );
and ( n34061 , n34059 , n34060 );
and ( n34062 , n24337 , n25284 );
and ( n34063 , n34060 , n34062 );
and ( n34064 , n34059 , n34062 );
or ( n34065 , n34061 , n34063 , n34064 );
and ( n34066 , n26399 , n21990 );
and ( n34067 , n34065 , n34066 );
xor ( n34068 , n33735 , n33736 );
xor ( n34069 , n34068 , n33741 );
and ( n34070 , n34066 , n34069 );
and ( n34071 , n34065 , n34069 );
or ( n34072 , n34067 , n34070 , n34071 );
and ( n34073 , n34057 , n34072 );
and ( n34074 , n34055 , n34072 );
or ( n34075 , n34058 , n34073 , n34074 );
xor ( n34076 , n31447 , n33622 );
buf ( n34077 , n34076 );
buf ( n34078 , n34077 );
buf ( n34079 , n34078 );
and ( n34080 , n34079 , n28117 );
and ( n34081 , n28532 , n34080 );
xor ( n34082 , n33942 , n33943 );
xor ( n34083 , n34082 , n33945 );
and ( n34084 , n34080 , n34083 );
and ( n34085 , n28532 , n34083 );
or ( n34086 , n34081 , n34084 , n34085 );
xor ( n34087 , n34005 , n34006 );
xor ( n34088 , n34087 , n34008 );
and ( n34089 , n27863 , n21178 );
and ( n34090 , n26980 , n21527 );
and ( n34091 , n34089 , n34090 );
and ( n34092 , n26933 , n21666 );
and ( n34093 , n34090 , n34092 );
and ( n34094 , n34089 , n34092 );
or ( n34095 , n34091 , n34093 , n34094 );
and ( n34096 , n34088 , n34095 );
buf ( n34097 , n22824 );
buf ( n34098 , n767 );
buf ( n34099 , n34098 );
buf ( n34100 , n768 );
buf ( n34101 , n34100 );
and ( n34102 , n34099 , n34101 );
not ( n34103 , n34102 );
and ( n34104 , n28529 , n34103 );
not ( n34105 , n34104 );
and ( n34106 , n34097 , n34105 );
and ( n34107 , n34095 , n34106 );
and ( n34108 , n34088 , n34106 );
or ( n34109 , n34096 , n34107 , n34108 );
and ( n34110 , n34086 , n34109 );
and ( n34111 , n28129 , n21039 );
and ( n34112 , n27389 , n21429 );
and ( n34113 , n34111 , n34112 );
and ( n34114 , n26678 , n21990 );
and ( n34115 , n34112 , n34114 );
and ( n34116 , n34111 , n34114 );
or ( n34117 , n34113 , n34115 , n34116 );
and ( n34118 , n25220 , n23508 );
and ( n34119 , n23620 , n26876 );
and ( n34120 , n34118 , n34119 );
buf ( n34121 , n11708 );
buf ( n34122 , n34121 );
and ( n34123 , n22936 , n34122 );
and ( n34124 , n34119 , n34123 );
and ( n34125 , n34118 , n34123 );
or ( n34126 , n34120 , n34124 , n34125 );
and ( n34127 , n34117 , n34126 );
xor ( n34128 , n33797 , n33798 );
xor ( n34129 , n34128 , n33800 );
and ( n34130 , n34126 , n34129 );
and ( n34131 , n34117 , n34129 );
or ( n34132 , n34127 , n34130 , n34131 );
and ( n34133 , n34109 , n34132 );
and ( n34134 , n34086 , n34132 );
or ( n34135 , n34110 , n34133 , n34134 );
and ( n34136 , n34075 , n34135 );
xor ( n34137 , n33734 , n33750 );
xor ( n34138 , n34137 , n33759 );
and ( n34139 , n34135 , n34138 );
and ( n34140 , n34075 , n34138 );
or ( n34141 , n34136 , n34139 , n34140 );
and ( n34142 , n34047 , n34141 );
and ( n34143 , n34032 , n34141 );
or ( n34144 , n34048 , n34142 , n34143 );
and ( n34145 , n34027 , n34144 );
and ( n34146 , n33968 , n34144 );
or ( n34147 , n34028 , n34145 , n34146 );
and ( n34148 , n33915 , n34147 );
and ( n34149 , n33862 , n34147 );
or ( n34150 , n33916 , n34148 , n34149 );
xor ( n34151 , n33697 , n33699 );
xor ( n34152 , n34151 , n33702 );
xor ( n34153 , n33708 , n33731 );
xor ( n34154 , n34153 , n33762 );
and ( n34155 , n34152 , n34154 );
xor ( n34156 , n33786 , n33814 );
xor ( n34157 , n34156 , n33817 );
and ( n34158 , n34154 , n34157 );
and ( n34159 , n34152 , n34157 );
or ( n34160 , n34155 , n34158 , n34159 );
xor ( n34161 , n33685 , n33687 );
xor ( n34162 , n34161 , n33690 );
and ( n34163 , n34160 , n34162 );
xor ( n34164 , n33695 , n33705 );
xor ( n34165 , n34164 , n33765 );
and ( n34166 , n34162 , n34165 );
and ( n34167 , n34160 , n34165 );
or ( n34168 , n34163 , n34166 , n34167 );
xor ( n34169 , n33683 , n33693 );
xor ( n34170 , n34169 , n33768 );
and ( n34171 , n34168 , n34170 );
xor ( n34172 , n33828 , n33830 );
xor ( n34173 , n34172 , n33833 );
and ( n34174 , n34170 , n34173 );
and ( n34175 , n34168 , n34173 );
or ( n34176 , n34171 , n34174 , n34175 );
and ( n34177 , n34150 , n34176 );
xor ( n34178 , n33678 , n33680 );
xor ( n34179 , n34178 , n33771 );
and ( n34180 , n34176 , n34179 );
and ( n34181 , n34150 , n34179 );
or ( n34182 , n34177 , n34180 , n34181 );
and ( n34183 , n33860 , n34182 );
xor ( n34184 , n33774 , n33844 );
xor ( n34185 , n34184 , n33847 );
and ( n34186 , n34182 , n34185 );
and ( n34187 , n33860 , n34185 );
or ( n34188 , n34183 , n34186 , n34187 );
and ( n34189 , n33858 , n34188 );
xor ( n34190 , n33673 , n33675 );
xor ( n34191 , n34190 , n33850 );
and ( n34192 , n34188 , n34191 );
and ( n34193 , n33858 , n34191 );
or ( n34194 , n34189 , n34192 , n34193 );
and ( n34195 , n33855 , n34194 );
and ( n34196 , n33853 , n34194 );
or ( n34197 , n33856 , n34195 , n34196 );
or ( n34198 , n28442 , n34197 );
or ( n34199 , n28440 , n34198 );
and ( n34200 , n28438 , n34199 );
xor ( n34201 , n28438 , n34199 );
xnor ( n34202 , n28440 , n34198 );
xnor ( n34203 , n28442 , n34197 );
xor ( n34204 , n33853 , n33855 );
xor ( n34205 , n34204 , n34194 );
not ( n34206 , n34205 );
xor ( n34207 , n33858 , n34188 );
xor ( n34208 , n34207 , n34191 );
xor ( n34209 , n33836 , n33838 );
xor ( n34210 , n34209 , n33841 );
xor ( n34211 , n33820 , n33822 );
xor ( n34212 , n34211 , n33825 );
xor ( n34213 , n33885 , n33909 );
xor ( n34214 , n34213 , n33912 );
and ( n34215 , n34212 , n34214 );
xor ( n34216 , n33899 , n33903 );
xor ( n34217 , n34216 , n33906 );
xnor ( n34218 , n33941 , n33967 );
and ( n34219 , n34217 , n34218 );
xor ( n34220 , n33923 , n33936 );
xor ( n34221 , n34220 , n33938 );
xor ( n34222 , n33954 , n33961 );
xor ( n34223 , n34222 , n33964 );
or ( n34224 , n34221 , n34223 );
and ( n34225 , n34218 , n34224 );
and ( n34226 , n34217 , n34224 );
or ( n34227 , n34219 , n34225 , n34226 );
and ( n34228 , n34214 , n34227 );
and ( n34229 , n34212 , n34227 );
or ( n34230 , n34215 , n34228 , n34229 );
xor ( n34231 , n33777 , n33781 );
xor ( n34232 , n34231 , n33783 );
xor ( n34233 , n33806 , n33808 );
xor ( n34234 , n34233 , n33811 );
and ( n34235 , n34232 , n34234 );
xor ( n34236 , n33893 , n33894 );
xor ( n34237 , n34236 , n33896 );
and ( n34238 , n34234 , n34237 );
and ( n34239 , n34232 , n34237 );
or ( n34240 , n34235 , n34238 , n34239 );
xor ( n34241 , n34004 , n34018 );
xor ( n34242 , n34241 , n34021 );
xnor ( n34243 , n34029 , n34031 );
and ( n34244 , n34242 , n34243 );
and ( n34245 , n23483 , n27558 );
and ( n34246 , n23336 , n28209 );
and ( n34247 , n34245 , n34246 );
and ( n34248 , n23215 , n33739 );
and ( n34249 , n34246 , n34248 );
and ( n34250 , n34245 , n34248 );
or ( n34251 , n34247 , n34249 , n34250 );
and ( n34252 , n24624 , n25026 );
and ( n34253 , n23903 , n26376 );
and ( n34254 , n34252 , n34253 );
and ( n34255 , n23620 , n27246 );
and ( n34256 , n34253 , n34255 );
and ( n34257 , n34252 , n34255 );
or ( n34258 , n34254 , n34256 , n34257 );
and ( n34259 , n34251 , n34258 );
and ( n34260 , n25959 , n22562 );
and ( n34261 , n34258 , n34260 );
and ( n34262 , n34251 , n34260 );
or ( n34263 , n34259 , n34261 , n34262 );
and ( n34264 , n25623 , n22987 );
and ( n34265 , n25451 , n23322 );
and ( n34266 , n34264 , n34265 );
xor ( n34267 , n33981 , n33982 );
xor ( n34268 , n34267 , n33984 );
and ( n34269 , n34265 , n34268 );
and ( n34270 , n34264 , n34268 );
or ( n34271 , n34266 , n34269 , n34270 );
and ( n34272 , n34263 , n34271 );
and ( n34273 , n27863 , n21085 );
and ( n34274 , n34271 , n34273 );
and ( n34275 , n34263 , n34273 );
or ( n34276 , n34272 , n34274 , n34275 );
xor ( n34277 , n33948 , n33949 );
xor ( n34278 , n34277 , n33951 );
and ( n34279 , n34276 , n34278 );
xor ( n34280 , n33744 , n33745 );
xor ( n34281 , n34280 , n33747 );
and ( n34282 , n34278 , n34281 );
and ( n34283 , n34276 , n34281 );
or ( n34284 , n34279 , n34282 , n34283 );
and ( n34285 , n34243 , n34284 );
and ( n34286 , n34242 , n34284 );
or ( n34287 , n34244 , n34285 , n34286 );
and ( n34288 , n34240 , n34287 );
xor ( n34289 , n33930 , n33931 );
xor ( n34290 , n34289 , n33933 );
xor ( n34291 , n33955 , n33956 );
xor ( n34292 , n34291 , n33958 );
and ( n34293 , n34290 , n34292 );
and ( n34294 , n25959 , n22337 );
and ( n34295 , n25623 , n22784 );
and ( n34296 , n34294 , n34295 );
xor ( n34297 , n33924 , n33925 );
xor ( n34298 , n34297 , n33927 );
and ( n34299 , n34295 , n34298 );
and ( n34300 , n34294 , n34298 );
or ( n34301 , n34296 , n34299 , n34300 );
xor ( n34302 , n33917 , n33918 );
xor ( n34303 , n34302 , n33920 );
and ( n34304 , n34301 , n34303 );
xor ( n34305 , n33886 , n33887 );
xor ( n34306 , n34305 , n33890 );
and ( n34307 , n34303 , n34306 );
and ( n34308 , n34301 , n34306 );
or ( n34309 , n34304 , n34307 , n34308 );
and ( n34310 , n34293 , n34309 );
xor ( n34311 , n33788 , n33795 );
xor ( n34312 , n34311 , n33803 );
xor ( n34313 , n34011 , n34012 );
xor ( n34314 , n34313 , n34015 );
and ( n34315 , n34312 , n34314 );
xnor ( n34316 , n34039 , n34041 );
and ( n34317 , n34314 , n34316 );
and ( n34318 , n34312 , n34316 );
or ( n34319 , n34315 , n34317 , n34318 );
and ( n34320 , n34309 , n34319 );
and ( n34321 , n34293 , n34319 );
or ( n34322 , n34310 , n34320 , n34321 );
and ( n34323 , n34287 , n34322 );
and ( n34324 , n34240 , n34322 );
or ( n34325 , n34288 , n34323 , n34324 );
and ( n34326 , n34038 , n33632 );
and ( n34327 , n33628 , n33630 );
nor ( n34328 , n34326 , n34327 );
xnor ( n34329 , n34328 , n28124 );
xor ( n34330 , n33974 , n33975 );
xor ( n34331 , n34330 , n33977 );
and ( n34332 , n34329 , n34331 );
xor ( n34333 , n33987 , n33994 );
xor ( n34334 , n34333 , n33996 );
and ( n34335 , n34331 , n34334 );
and ( n34336 , n34329 , n34334 );
or ( n34337 , n34332 , n34335 , n34336 );
xor ( n34338 , n34049 , n34050 );
xor ( n34339 , n34338 , n34052 );
and ( n34340 , n23089 , n34122 );
buf ( n34341 , n34340 );
and ( n34342 , n24052 , n25617 );
and ( n34343 , n34341 , n34342 );
and ( n34344 , n23903 , n26229 );
and ( n34345 , n34342 , n34344 );
and ( n34346 , n34341 , n34344 );
or ( n34347 , n34343 , n34345 , n34346 );
and ( n34348 , n34339 , n34347 );
xor ( n34349 , n28121 , n28527 );
xor ( n34350 , n28527 , n28529 );
not ( n34351 , n34350 );
and ( n34352 , n34349 , n34351 );
and ( n34353 , n33628 , n34352 );
not ( n34354 , n34353 );
xnor ( n34355 , n34354 , n28532 );
xor ( n34356 , n34059 , n34060 );
xor ( n34357 , n34356 , n34062 );
and ( n34358 , n34355 , n34357 );
and ( n34359 , n26782 , n21827 );
and ( n34360 , n26399 , n22172 );
xor ( n34361 , n34359 , n34360 );
and ( n34362 , n26148 , n22337 );
xor ( n34363 , n34361 , n34362 );
and ( n34364 , n34357 , n34363 );
and ( n34365 , n34355 , n34363 );
or ( n34366 , n34358 , n34364 , n34365 );
and ( n34367 , n34347 , n34366 );
and ( n34368 , n34339 , n34366 );
or ( n34369 , n34348 , n34367 , n34368 );
and ( n34370 , n34337 , n34369 );
xor ( n34371 , n34089 , n34090 );
xor ( n34372 , n34371 , n34092 );
xor ( n34373 , n34097 , n34105 );
and ( n34374 , n34372 , n34373 );
and ( n34375 , n24993 , n24064 );
and ( n34376 , n24731 , n24540 );
and ( n34377 , n34375 , n34376 );
and ( n34378 , n24546 , n25284 );
and ( n34379 , n34376 , n34378 );
and ( n34380 , n34375 , n34378 );
or ( n34381 , n34377 , n34379 , n34380 );
and ( n34382 , n34373 , n34381 );
and ( n34383 , n34372 , n34381 );
or ( n34384 , n34374 , n34382 , n34383 );
and ( n34385 , n26933 , n21827 );
and ( n34386 , n26678 , n22172 );
and ( n34387 , n34385 , n34386 );
and ( n34388 , n26399 , n22337 );
and ( n34389 , n34386 , n34388 );
and ( n34390 , n34385 , n34388 );
or ( n34391 , n34387 , n34389 , n34390 );
and ( n34392 , n28129 , n21085 );
and ( n34393 , n27962 , n21178 );
and ( n34394 , n34392 , n34393 );
and ( n34395 , n27389 , n21527 );
and ( n34396 , n34393 , n34395 );
and ( n34397 , n34392 , n34395 );
or ( n34398 , n34394 , n34396 , n34397 );
and ( n34399 , n34391 , n34398 );
and ( n34400 , n27863 , n21296 );
and ( n34401 , n27591 , n21429 );
and ( n34402 , n34400 , n34401 );
and ( n34403 , n23742 , n26876 );
and ( n34404 , n34401 , n34403 );
and ( n34405 , n34400 , n34403 );
or ( n34406 , n34402 , n34404 , n34405 );
and ( n34407 , n34398 , n34406 );
and ( n34408 , n34391 , n34406 );
or ( n34409 , n34399 , n34407 , n34408 );
and ( n34410 , n34384 , n34409 );
and ( n34411 , n34038 , n34352 );
and ( n34412 , n33628 , n34350 );
nor ( n34413 , n34411 , n34412 );
xnor ( n34414 , n34413 , n28532 );
and ( n34415 , n34104 , n34414 );
xor ( n34416 , n31449 , n33621 );
buf ( n34417 , n34416 );
buf ( n34418 , n34417 );
buf ( n34419 , n34418 );
and ( n34420 , n34419 , n33632 );
and ( n34421 , n34079 , n33630 );
nor ( n34422 , n34420 , n34421 );
xnor ( n34423 , n34422 , n28124 );
and ( n34424 , n34414 , n34423 );
and ( n34425 , n34104 , n34423 );
or ( n34426 , n34415 , n34424 , n34425 );
xor ( n34427 , n34111 , n34112 );
xor ( n34428 , n34427 , n34114 );
and ( n34429 , n34426 , n34428 );
xor ( n34430 , n34118 , n34119 );
xor ( n34431 , n34430 , n34123 );
and ( n34432 , n34428 , n34431 );
and ( n34433 , n34426 , n34431 );
or ( n34434 , n34429 , n34432 , n34433 );
and ( n34435 , n34409 , n34434 );
and ( n34436 , n34384 , n34434 );
or ( n34437 , n34410 , n34435 , n34436 );
and ( n34438 , n34369 , n34437 );
and ( n34439 , n34337 , n34437 );
or ( n34440 , n34370 , n34438 , n34439 );
xor ( n34441 , n28532 , n34080 );
xor ( n34442 , n34441 , n34083 );
xor ( n34443 , n34088 , n34095 );
xor ( n34444 , n34443 , n34106 );
and ( n34445 , n34442 , n34444 );
xor ( n34446 , n34117 , n34126 );
xor ( n34447 , n34446 , n34129 );
and ( n34448 , n34444 , n34447 );
and ( n34449 , n34442 , n34447 );
or ( n34450 , n34445 , n34448 , n34449 );
xor ( n34451 , n34055 , n34057 );
xor ( n34452 , n34451 , n34072 );
and ( n34453 , n34450 , n34452 );
xor ( n34454 , n34086 , n34109 );
xor ( n34455 , n34454 , n34132 );
and ( n34456 , n34452 , n34455 );
and ( n34457 , n34450 , n34455 );
or ( n34458 , n34453 , n34456 , n34457 );
and ( n34459 , n34440 , n34458 );
xor ( n34460 , n34034 , n34042 );
xor ( n34461 , n34460 , n34044 );
and ( n34462 , n34458 , n34461 );
and ( n34463 , n34440 , n34461 );
or ( n34464 , n34459 , n34462 , n34463 );
xor ( n34465 , n33970 , n33972 );
xor ( n34466 , n34465 , n34024 );
and ( n34467 , n34464 , n34466 );
xor ( n34468 , n34032 , n34047 );
xor ( n34469 , n34468 , n34141 );
and ( n34470 , n34466 , n34469 );
and ( n34471 , n34464 , n34469 );
or ( n34472 , n34467 , n34470 , n34471 );
and ( n34473 , n34325 , n34472 );
xor ( n34474 , n33968 , n34027 );
xor ( n34475 , n34474 , n34144 );
and ( n34476 , n34472 , n34475 );
and ( n34477 , n34325 , n34475 );
or ( n34478 , n34473 , n34476 , n34477 );
and ( n34479 , n34230 , n34478 );
xor ( n34480 , n33862 , n33915 );
xor ( n34481 , n34480 , n34147 );
and ( n34482 , n34478 , n34481 );
and ( n34483 , n34230 , n34481 );
or ( n34484 , n34479 , n34482 , n34483 );
and ( n34485 , n34210 , n34484 );
xor ( n34486 , n34150 , n34176 );
xor ( n34487 , n34486 , n34179 );
and ( n34488 , n34484 , n34487 );
and ( n34489 , n34210 , n34487 );
or ( n34490 , n34485 , n34488 , n34489 );
xor ( n34491 , n33860 , n34182 );
xor ( n34492 , n34491 , n34185 );
and ( n34493 , n34490 , n34492 );
xor ( n34494 , n34168 , n34170 );
xor ( n34495 , n34494 , n34173 );
xor ( n34496 , n34160 , n34162 );
xor ( n34497 , n34496 , n34165 );
xor ( n34498 , n34152 , n34154 );
xor ( n34499 , n34498 , n34157 );
xor ( n34500 , n34075 , n34135 );
xor ( n34501 , n34500 , n34138 );
xnor ( n34502 , n34221 , n34223 );
and ( n34503 , n34501 , n34502 );
and ( n34504 , n34359 , n34360 );
and ( n34505 , n34360 , n34362 );
and ( n34506 , n34359 , n34362 );
or ( n34507 , n34504 , n34505 , n34506 );
and ( n34508 , n24337 , n25617 );
and ( n34509 , n24052 , n26229 );
and ( n34510 , n34508 , n34509 );
not ( n34511 , n34340 );
and ( n34512 , n34509 , n34511 );
and ( n34513 , n34508 , n34511 );
or ( n34514 , n34510 , n34512 , n34513 );
and ( n34515 , n25742 , n22784 );
and ( n34516 , n34514 , n34515 );
and ( n34517 , n24993 , n23758 );
and ( n34518 , n34515 , n34517 );
and ( n34519 , n34514 , n34517 );
or ( n34520 , n34516 , n34518 , n34519 );
and ( n34521 , n34507 , n34520 );
and ( n34522 , n27962 , n21039 );
and ( n34523 , n34520 , n34522 );
and ( n34524 , n34507 , n34522 );
or ( n34525 , n34521 , n34523 , n34524 );
xor ( n34526 , n33980 , n33999 );
xor ( n34527 , n34526 , n34001 );
and ( n34528 , n34525 , n34527 );
xor ( n34529 , n34301 , n34303 );
xor ( n34530 , n34529 , n34306 );
and ( n34531 , n34527 , n34530 );
and ( n34532 , n34525 , n34530 );
or ( n34533 , n34528 , n34531 , n34532 );
and ( n34534 , n34502 , n34533 );
and ( n34535 , n34501 , n34533 );
or ( n34536 , n34503 , n34534 , n34535 );
and ( n34537 , n34499 , n34536 );
xor ( n34538 , n34276 , n34278 );
xor ( n34539 , n34538 , n34281 );
xor ( n34540 , n34290 , n34292 );
and ( n34541 , n34539 , n34540 );
and ( n34542 , n24731 , n25026 );
and ( n34543 , n24052 , n26376 );
and ( n34544 , n34542 , n34543 );
and ( n34545 , n23620 , n27558 );
and ( n34546 , n34543 , n34545 );
and ( n34547 , n34542 , n34545 );
or ( n34548 , n34544 , n34546 , n34547 );
and ( n34549 , n26148 , n22562 );
and ( n34550 , n34548 , n34549 );
and ( n34551 , n25742 , n22987 );
and ( n34552 , n34549 , n34551 );
and ( n34553 , n34548 , n34551 );
or ( n34554 , n34550 , n34552 , n34553 );
and ( n34555 , n25623 , n23322 );
and ( n34556 , n25451 , n23508 );
and ( n34557 , n34555 , n34556 );
xor ( n34558 , n34245 , n34246 );
xor ( n34559 , n34558 , n34248 );
and ( n34560 , n34556 , n34559 );
and ( n34561 , n34555 , n34559 );
or ( n34562 , n34557 , n34560 , n34561 );
and ( n34563 , n34554 , n34562 );
and ( n34564 , n27962 , n21085 );
and ( n34565 , n34562 , n34564 );
and ( n34566 , n34554 , n34564 );
or ( n34567 , n34563 , n34565 , n34566 );
xor ( n34568 , n33789 , n33790 );
xor ( n34569 , n34568 , n33792 );
and ( n34570 , n34567 , n34569 );
xor ( n34571 , n34065 , n34066 );
xor ( n34572 , n34571 , n34069 );
and ( n34573 , n34569 , n34572 );
and ( n34574 , n34567 , n34572 );
or ( n34575 , n34570 , n34573 , n34574 );
and ( n34576 , n34540 , n34575 );
and ( n34577 , n34539 , n34575 );
or ( n34578 , n34541 , n34576 , n34577 );
and ( n34579 , n27591 , n21296 );
xor ( n34580 , n33988 , n33989 );
xor ( n34581 , n34580 , n33991 );
and ( n34582 , n34579 , n34581 );
xor ( n34583 , n34341 , n34342 );
xor ( n34584 , n34583 , n34344 );
and ( n34585 , n34581 , n34584 );
and ( n34586 , n34579 , n34584 );
or ( n34587 , n34582 , n34585 , n34586 );
xor ( n34588 , n34294 , n34295 );
xor ( n34589 , n34588 , n34298 );
or ( n34590 , n34587 , n34589 );
xor ( n34591 , n34507 , n34520 );
xor ( n34592 , n34591 , n34522 );
xor ( n34593 , n34263 , n34271 );
xor ( n34594 , n34593 , n34273 );
and ( n34595 , n34592 , n34594 );
xor ( n34596 , n34329 , n34331 );
xor ( n34597 , n34596 , n34334 );
and ( n34598 , n34594 , n34597 );
and ( n34599 , n34592 , n34597 );
or ( n34600 , n34595 , n34598 , n34599 );
and ( n34601 , n34590 , n34600 );
xor ( n34602 , n34251 , n34258 );
xor ( n34603 , n34602 , n34260 );
xor ( n34604 , n34264 , n34265 );
xor ( n34605 , n34604 , n34268 );
and ( n34606 , n34603 , n34605 );
xor ( n34607 , n34375 , n34376 );
xor ( n34608 , n34607 , n34378 );
xor ( n34609 , n34252 , n34253 );
xor ( n34610 , n34609 , n34255 );
and ( n34611 , n34608 , n34610 );
xor ( n34612 , n34385 , n34386 );
xor ( n34613 , n34612 , n34388 );
and ( n34614 , n34610 , n34613 );
and ( n34615 , n34608 , n34613 );
or ( n34616 , n34611 , n34614 , n34615 );
and ( n34617 , n34605 , n34616 );
and ( n34618 , n34603 , n34616 );
or ( n34619 , n34606 , n34617 , n34618 );
xor ( n34620 , n34392 , n34393 );
xor ( n34621 , n34620 , n34395 );
and ( n34622 , n23483 , n28209 );
and ( n34623 , n23336 , n33739 );
and ( n34624 , n34622 , n34623 );
and ( n34625 , n23215 , n34122 );
and ( n34626 , n34623 , n34625 );
and ( n34627 , n34622 , n34625 );
or ( n34628 , n34624 , n34626 , n34627 );
and ( n34629 , n34621 , n34628 );
and ( n34630 , n34079 , n34352 );
and ( n34631 , n34038 , n34350 );
nor ( n34632 , n34630 , n34631 );
xnor ( n34633 , n34632 , n28532 );
xor ( n34634 , n31451 , n33620 );
buf ( n34635 , n34634 );
buf ( n34636 , n34635 );
buf ( n34637 , n34636 );
and ( n34638 , n34637 , n33632 );
and ( n34639 , n34419 , n33630 );
nor ( n34640 , n34638 , n34639 );
xnor ( n34641 , n34640 , n28124 );
and ( n34642 , n34633 , n34641 );
xor ( n34643 , n31453 , n33619 );
buf ( n34644 , n34643 );
buf ( n34645 , n34644 );
buf ( n34646 , n34645 );
and ( n34647 , n34646 , n28117 );
and ( n34648 , n34641 , n34647 );
and ( n34649 , n34633 , n34647 );
or ( n34650 , n34642 , n34648 , n34649 );
and ( n34651 , n34628 , n34650 );
and ( n34652 , n34621 , n34650 );
or ( n34653 , n34629 , n34651 , n34652 );
buf ( n34654 , n22936 );
buf ( n34655 , n769 );
buf ( n34656 , n34655 );
buf ( n34657 , n770 );
buf ( n34658 , n34657 );
and ( n34659 , n34656 , n34658 );
not ( n34660 , n34659 );
and ( n34661 , n34101 , n34660 );
not ( n34662 , n34661 );
and ( n34663 , n34654 , n34662 );
and ( n34664 , n28129 , n21178 );
and ( n34665 , n24546 , n25617 );
and ( n34666 , n34664 , n34665 );
and ( n34667 , n24337 , n26229 );
and ( n34668 , n34665 , n34667 );
and ( n34669 , n34664 , n34667 );
or ( n34670 , n34666 , n34668 , n34669 );
and ( n34671 , n34663 , n34670 );
xor ( n34672 , n34400 , n34401 );
xor ( n34673 , n34672 , n34403 );
and ( n34674 , n34670 , n34673 );
and ( n34675 , n34663 , n34673 );
or ( n34676 , n34671 , n34674 , n34675 );
and ( n34677 , n34653 , n34676 );
xor ( n34678 , n34355 , n34357 );
xor ( n34679 , n34678 , n34363 );
and ( n34680 , n34676 , n34679 );
and ( n34681 , n34653 , n34679 );
or ( n34682 , n34677 , n34680 , n34681 );
and ( n34683 , n34619 , n34682 );
xor ( n34684 , n34372 , n34373 );
xor ( n34685 , n34684 , n34381 );
xor ( n34686 , n34391 , n34398 );
xor ( n34687 , n34686 , n34406 );
and ( n34688 , n34685 , n34687 );
xor ( n34689 , n34426 , n34428 );
xor ( n34690 , n34689 , n34431 );
and ( n34691 , n34687 , n34690 );
and ( n34692 , n34685 , n34690 );
or ( n34693 , n34688 , n34691 , n34692 );
and ( n34694 , n34682 , n34693 );
and ( n34695 , n34619 , n34693 );
or ( n34696 , n34683 , n34694 , n34695 );
and ( n34697 , n34600 , n34696 );
and ( n34698 , n34590 , n34696 );
or ( n34699 , n34601 , n34697 , n34698 );
and ( n34700 , n34578 , n34699 );
xor ( n34701 , n34339 , n34347 );
xor ( n34702 , n34701 , n34366 );
xor ( n34703 , n34384 , n34409 );
xor ( n34704 , n34703 , n34434 );
and ( n34705 , n34702 , n34704 );
xor ( n34706 , n34442 , n34444 );
xor ( n34707 , n34706 , n34447 );
and ( n34708 , n34704 , n34707 );
and ( n34709 , n34702 , n34707 );
or ( n34710 , n34705 , n34708 , n34709 );
xor ( n34711 , n34312 , n34314 );
xor ( n34712 , n34711 , n34316 );
and ( n34713 , n34710 , n34712 );
xor ( n34714 , n34337 , n34369 );
xor ( n34715 , n34714 , n34437 );
and ( n34716 , n34712 , n34715 );
and ( n34717 , n34710 , n34715 );
or ( n34718 , n34713 , n34716 , n34717 );
and ( n34719 , n34699 , n34718 );
and ( n34720 , n34578 , n34718 );
or ( n34721 , n34700 , n34719 , n34720 );
and ( n34722 , n34536 , n34721 );
and ( n34723 , n34499 , n34721 );
or ( n34724 , n34537 , n34722 , n34723 );
and ( n34725 , n34497 , n34724 );
xor ( n34726 , n34232 , n34234 );
xor ( n34727 , n34726 , n34237 );
xor ( n34728 , n34242 , n34243 );
xor ( n34729 , n34728 , n34284 );
and ( n34730 , n34727 , n34729 );
xor ( n34731 , n34293 , n34309 );
xor ( n34732 , n34731 , n34319 );
and ( n34733 , n34729 , n34732 );
and ( n34734 , n34727 , n34732 );
or ( n34735 , n34730 , n34733 , n34734 );
xor ( n34736 , n34217 , n34218 );
xor ( n34737 , n34736 , n34224 );
and ( n34738 , n34735 , n34737 );
xor ( n34739 , n34240 , n34287 );
xor ( n34740 , n34739 , n34322 );
and ( n34741 , n34737 , n34740 );
and ( n34742 , n34735 , n34740 );
or ( n34743 , n34738 , n34741 , n34742 );
and ( n34744 , n34724 , n34743 );
and ( n34745 , n34497 , n34743 );
or ( n34746 , n34725 , n34744 , n34745 );
and ( n34747 , n34495 , n34746 );
xor ( n34748 , n34230 , n34478 );
xor ( n34749 , n34748 , n34481 );
and ( n34750 , n34746 , n34749 );
and ( n34751 , n34495 , n34749 );
or ( n34752 , n34747 , n34750 , n34751 );
xor ( n34753 , n34210 , n34484 );
xor ( n34754 , n34753 , n34487 );
and ( n34755 , n34752 , n34754 );
xor ( n34756 , n34212 , n34214 );
xor ( n34757 , n34756 , n34227 );
xor ( n34758 , n34325 , n34472 );
xor ( n34759 , n34758 , n34475 );
and ( n34760 , n34757 , n34759 );
xor ( n34761 , n34464 , n34466 );
xor ( n34762 , n34761 , n34469 );
xor ( n34763 , n34440 , n34458 );
xor ( n34764 , n34763 , n34461 );
xor ( n34765 , n34450 , n34452 );
xor ( n34766 , n34765 , n34455 );
xor ( n34767 , n34525 , n34527 );
xor ( n34768 , n34767 , n34530 );
and ( n34769 , n34766 , n34768 );
xor ( n34770 , n34567 , n34569 );
xor ( n34771 , n34770 , n34572 );
xnor ( n34772 , n34587 , n34589 );
and ( n34773 , n34771 , n34772 );
and ( n34774 , n34079 , n33632 );
and ( n34775 , n34038 , n33630 );
nor ( n34776 , n34774 , n34775 );
xnor ( n34777 , n34776 , n28124 );
and ( n34778 , n34419 , n28117 );
and ( n34779 , n34777 , n34778 );
xor ( n34780 , n34579 , n34581 );
xor ( n34781 , n34780 , n34584 );
and ( n34782 , n34778 , n34781 );
and ( n34783 , n34777 , n34781 );
or ( n34784 , n34779 , n34782 , n34783 );
and ( n34785 , n34772 , n34784 );
and ( n34786 , n34771 , n34784 );
or ( n34787 , n34773 , n34785 , n34786 );
and ( n34788 , n34768 , n34787 );
and ( n34789 , n34766 , n34787 );
or ( n34790 , n34769 , n34788 , n34789 );
and ( n34791 , n34764 , n34790 );
and ( n34792 , n23620 , n28209 );
and ( n34793 , n23483 , n33739 );
and ( n34794 , n34792 , n34793 );
and ( n34795 , n23336 , n34122 );
and ( n34796 , n34793 , n34795 );
and ( n34797 , n34792 , n34795 );
or ( n34798 , n34794 , n34796 , n34797 );
and ( n34799 , n25623 , n23508 );
and ( n34800 , n34798 , n34799 );
and ( n34801 , n24624 , n25284 );
and ( n34802 , n34799 , n34801 );
and ( n34803 , n34798 , n34801 );
or ( n34804 , n34800 , n34802 , n34803 );
and ( n34805 , n26980 , n21666 );
and ( n34806 , n34804 , n34805 );
and ( n34807 , n26782 , n21990 );
and ( n34808 , n34805 , n34807 );
and ( n34809 , n34804 , n34807 );
or ( n34810 , n34806 , n34808 , n34809 );
xor ( n34811 , n34514 , n34515 );
xor ( n34812 , n34811 , n34517 );
or ( n34813 , n34810 , n34812 );
xor ( n34814 , n34554 , n34562 );
xor ( n34815 , n34814 , n34564 );
buf ( n34816 , n11835 );
buf ( n34817 , n34816 );
and ( n34818 , n23215 , n34817 );
buf ( n34819 , n34818 );
and ( n34820 , n23903 , n26876 );
and ( n34821 , n34819 , n34820 );
and ( n34822 , n23742 , n27246 );
and ( n34823 , n34820 , n34822 );
and ( n34824 , n34819 , n34822 );
or ( n34825 , n34821 , n34823 , n34824 );
and ( n34826 , n25959 , n22784 );
and ( n34827 , n34825 , n34826 );
and ( n34828 , n25220 , n23758 );
and ( n34829 , n34826 , n34828 );
and ( n34830 , n34825 , n34828 );
or ( n34831 , n34827 , n34829 , n34830 );
and ( n34832 , n34815 , n34831 );
and ( n34833 , n25451 , n23758 );
and ( n34834 , n25220 , n24064 );
and ( n34835 , n34833 , n34834 );
and ( n34836 , n24993 , n24540 );
and ( n34837 , n34834 , n34836 );
and ( n34838 , n34833 , n34836 );
or ( n34839 , n34835 , n34837 , n34838 );
and ( n34840 , n25959 , n22987 );
and ( n34841 , n25742 , n23322 );
and ( n34842 , n34840 , n34841 );
xor ( n34843 , n34622 , n34623 );
xor ( n34844 , n34843 , n34625 );
and ( n34845 , n34841 , n34844 );
and ( n34846 , n34840 , n34844 );
or ( n34847 , n34842 , n34845 , n34846 );
and ( n34848 , n34839 , n34847 );
xor ( n34849 , n34508 , n34509 );
xor ( n34850 , n34849 , n34511 );
and ( n34851 , n34847 , n34850 );
and ( n34852 , n34839 , n34850 );
or ( n34853 , n34848 , n34851 , n34852 );
and ( n34854 , n34831 , n34853 );
and ( n34855 , n34815 , n34853 );
or ( n34856 , n34832 , n34854 , n34855 );
and ( n34857 , n34813 , n34856 );
and ( n34858 , n26782 , n22172 );
and ( n34859 , n26678 , n22337 );
and ( n34860 , n34858 , n34859 );
and ( n34861 , n26148 , n22784 );
and ( n34862 , n34859 , n34861 );
and ( n34863 , n34858 , n34861 );
or ( n34864 , n34860 , n34862 , n34863 );
and ( n34865 , n24337 , n26376 );
and ( n34866 , n23903 , n27246 );
and ( n34867 , n34865 , n34866 );
and ( n34868 , n23742 , n27558 );
and ( n34869 , n34866 , n34868 );
and ( n34870 , n34865 , n34868 );
or ( n34871 , n34867 , n34869 , n34870 );
and ( n34872 , n24993 , n25026 );
and ( n34873 , n24546 , n26229 );
and ( n34874 , n34872 , n34873 );
not ( n34875 , n34818 );
and ( n34876 , n34873 , n34875 );
and ( n34877 , n34872 , n34875 );
or ( n34878 , n34874 , n34876 , n34877 );
and ( n34879 , n34871 , n34878 );
and ( n34880 , n26399 , n22562 );
and ( n34881 , n34878 , n34880 );
and ( n34882 , n34871 , n34880 );
or ( n34883 , n34879 , n34881 , n34882 );
and ( n34884 , n34864 , n34883 );
xor ( n34885 , n34548 , n34549 );
xor ( n34886 , n34885 , n34551 );
and ( n34887 , n34883 , n34886 );
and ( n34888 , n34864 , n34886 );
or ( n34889 , n34884 , n34887 , n34888 );
xor ( n34890 , n34104 , n34414 );
xor ( n34891 , n34890 , n34423 );
xor ( n34892 , n34555 , n34556 );
xor ( n34893 , n34892 , n34559 );
and ( n34894 , n34891 , n34893 );
and ( n34895 , n27962 , n21296 );
and ( n34896 , n26980 , n21827 );
and ( n34897 , n34895 , n34896 );
xor ( n34898 , n34542 , n34543 );
xor ( n34899 , n34898 , n34545 );
and ( n34900 , n34896 , n34899 );
and ( n34901 , n34895 , n34899 );
or ( n34902 , n34897 , n34900 , n34901 );
and ( n34903 , n34893 , n34902 );
and ( n34904 , n34891 , n34902 );
or ( n34905 , n34894 , n34903 , n34904 );
and ( n34906 , n34889 , n34905 );
and ( n34907 , n23089 , n34817 );
xor ( n34908 , n28529 , n34099 );
xor ( n34909 , n34099 , n34101 );
not ( n34910 , n34909 );
and ( n34911 , n34908 , n34910 );
and ( n34912 , n33628 , n34911 );
not ( n34913 , n34912 );
xnor ( n34914 , n34913 , n34104 );
and ( n34915 , n34907 , n34914 );
xor ( n34916 , n34858 , n34859 );
xor ( n34917 , n34916 , n34861 );
and ( n34918 , n34914 , n34917 );
and ( n34919 , n34907 , n34917 );
or ( n34920 , n34915 , n34918 , n34919 );
xor ( n34921 , n34833 , n34834 );
xor ( n34922 , n34921 , n34836 );
and ( n34923 , n27591 , n21527 );
and ( n34924 , n27389 , n21666 );
xor ( n34925 , n34923 , n34924 );
and ( n34926 , n26933 , n21990 );
xor ( n34927 , n34925 , n34926 );
and ( n34928 , n34922 , n34927 );
xor ( n34929 , n34633 , n34641 );
xor ( n34930 , n34929 , n34647 );
and ( n34931 , n34927 , n34930 );
and ( n34932 , n34922 , n34930 );
or ( n34933 , n34928 , n34931 , n34932 );
and ( n34934 , n34920 , n34933 );
xor ( n34935 , n34654 , n34662 );
and ( n34936 , n24731 , n25284 );
and ( n34937 , n34936 , n34661 );
and ( n34938 , n34646 , n33632 );
and ( n34939 , n34637 , n33630 );
nor ( n34940 , n34938 , n34939 );
xnor ( n34941 , n34940 , n28124 );
and ( n34942 , n34661 , n34941 );
and ( n34943 , n34936 , n34941 );
or ( n34944 , n34937 , n34942 , n34943 );
and ( n34945 , n34935 , n34944 );
xor ( n34946 , n34664 , n34665 );
xor ( n34947 , n34946 , n34667 );
and ( n34948 , n34944 , n34947 );
and ( n34949 , n34935 , n34947 );
or ( n34950 , n34945 , n34948 , n34949 );
and ( n34951 , n34933 , n34950 );
and ( n34952 , n34920 , n34950 );
or ( n34953 , n34934 , n34951 , n34952 );
and ( n34954 , n34905 , n34953 );
and ( n34955 , n34889 , n34953 );
or ( n34956 , n34906 , n34954 , n34955 );
and ( n34957 , n34856 , n34956 );
and ( n34958 , n34813 , n34956 );
or ( n34959 , n34857 , n34957 , n34958 );
xor ( n34960 , n34608 , n34610 );
xor ( n34961 , n34960 , n34613 );
xor ( n34962 , n34621 , n34628 );
xor ( n34963 , n34962 , n34650 );
and ( n34964 , n34961 , n34963 );
xor ( n34965 , n34663 , n34670 );
xor ( n34966 , n34965 , n34673 );
and ( n34967 , n34963 , n34966 );
and ( n34968 , n34961 , n34966 );
or ( n34969 , n34964 , n34967 , n34968 );
xor ( n34970 , n34603 , n34605 );
xor ( n34971 , n34970 , n34616 );
and ( n34972 , n34969 , n34971 );
xor ( n34973 , n34653 , n34676 );
xor ( n34974 , n34973 , n34679 );
and ( n34975 , n34971 , n34974 );
and ( n34976 , n34969 , n34974 );
or ( n34977 , n34972 , n34975 , n34976 );
xor ( n34978 , n34592 , n34594 );
xor ( n34979 , n34978 , n34597 );
and ( n34980 , n34977 , n34979 );
xor ( n34981 , n34619 , n34682 );
xor ( n34982 , n34981 , n34693 );
and ( n34983 , n34979 , n34982 );
and ( n34984 , n34977 , n34982 );
or ( n34985 , n34980 , n34983 , n34984 );
and ( n34986 , n34959 , n34985 );
xor ( n34987 , n34539 , n34540 );
xor ( n34988 , n34987 , n34575 );
and ( n34989 , n34985 , n34988 );
and ( n34990 , n34959 , n34988 );
or ( n34991 , n34986 , n34989 , n34990 );
and ( n34992 , n34790 , n34991 );
and ( n34993 , n34764 , n34991 );
or ( n34994 , n34791 , n34992 , n34993 );
and ( n34995 , n34762 , n34994 );
xor ( n34996 , n34501 , n34502 );
xor ( n34997 , n34996 , n34533 );
xor ( n34998 , n34578 , n34699 );
xor ( n34999 , n34998 , n34718 );
and ( n35000 , n34997 , n34999 );
xor ( n35001 , n34727 , n34729 );
xor ( n35002 , n35001 , n34732 );
and ( n35003 , n34999 , n35002 );
and ( n35004 , n34997 , n35002 );
or ( n35005 , n35000 , n35003 , n35004 );
and ( n35006 , n34994 , n35005 );
and ( n35007 , n34762 , n35005 );
or ( n35008 , n34995 , n35006 , n35007 );
and ( n35009 , n34759 , n35008 );
and ( n35010 , n34757 , n35008 );
or ( n35011 , n34760 , n35009 , n35010 );
xor ( n35012 , n34495 , n34746 );
xor ( n35013 , n35012 , n34749 );
and ( n35014 , n35011 , n35013 );
xor ( n35015 , n34497 , n34724 );
xor ( n35016 , n35015 , n34743 );
xor ( n35017 , n34499 , n34536 );
xor ( n35018 , n35017 , n34721 );
xor ( n35019 , n34735 , n34737 );
xor ( n35020 , n35019 , n34740 );
and ( n35021 , n35018 , n35020 );
xor ( n35022 , n34590 , n34600 );
xor ( n35023 , n35022 , n34696 );
xor ( n35024 , n34710 , n34712 );
xor ( n35025 , n35024 , n34715 );
and ( n35026 , n35023 , n35025 );
xor ( n35027 , n34702 , n34704 );
xor ( n35028 , n35027 , n34707 );
xor ( n35029 , n34685 , n34687 );
xor ( n35030 , n35029 , n34690 );
xor ( n35031 , n34777 , n34778 );
xor ( n35032 , n35031 , n34781 );
and ( n35033 , n35030 , n35032 );
xnor ( n35034 , n34810 , n34812 );
and ( n35035 , n35032 , n35034 );
and ( n35036 , n35030 , n35034 );
or ( n35037 , n35033 , n35035 , n35036 );
and ( n35038 , n35028 , n35037 );
xor ( n35039 , n34825 , n34826 );
xor ( n35040 , n35039 , n34828 );
xor ( n35041 , n34804 , n34805 );
xor ( n35042 , n35041 , n34807 );
and ( n35043 , n35040 , n35042 );
xor ( n35044 , n34839 , n34847 );
xor ( n35045 , n35044 , n34850 );
and ( n35046 , n35042 , n35045 );
and ( n35047 , n35040 , n35045 );
or ( n35048 , n35043 , n35046 , n35047 );
xor ( n35049 , n34864 , n34883 );
xor ( n35050 , n35049 , n34886 );
and ( n35051 , n28129 , n21296 );
and ( n35052 , n27389 , n21827 );
and ( n35053 , n35051 , n35052 );
and ( n35054 , n26933 , n22172 );
and ( n35055 , n35052 , n35054 );
and ( n35056 , n35051 , n35054 );
or ( n35057 , n35053 , n35055 , n35056 );
xor ( n35058 , n34871 , n34878 );
xor ( n35059 , n35058 , n34880 );
and ( n35060 , n35057 , n35059 );
xor ( n35061 , n34840 , n34841 );
xor ( n35062 , n35061 , n34844 );
and ( n35063 , n35059 , n35062 );
and ( n35064 , n35057 , n35062 );
or ( n35065 , n35060 , n35063 , n35064 );
and ( n35066 , n35050 , n35065 );
and ( n35067 , n25742 , n23508 );
and ( n35068 , n24624 , n25617 );
and ( n35069 , n35067 , n35068 );
and ( n35070 , n24052 , n26876 );
and ( n35071 , n35068 , n35070 );
and ( n35072 , n35067 , n35070 );
or ( n35073 , n35069 , n35071 , n35072 );
xor ( n35074 , n34819 , n34820 );
xor ( n35075 , n35074 , n34822 );
or ( n35076 , n35073 , n35075 );
and ( n35077 , n35065 , n35076 );
and ( n35078 , n35050 , n35076 );
or ( n35079 , n35066 , n35077 , n35078 );
and ( n35080 , n35048 , n35079 );
and ( n35081 , n27863 , n21429 );
xor ( n35082 , n34798 , n34799 );
xor ( n35083 , n35082 , n34801 );
or ( n35084 , n35081 , n35083 );
and ( n35085 , n27863 , n21527 );
and ( n35086 , n27591 , n21666 );
and ( n35087 , n35085 , n35086 );
and ( n35088 , n26980 , n21990 );
and ( n35089 , n35086 , n35088 );
and ( n35090 , n35085 , n35088 );
or ( n35091 , n35087 , n35089 , n35090 );
xor ( n35092 , n34895 , n34896 );
xor ( n35093 , n35092 , n34899 );
and ( n35094 , n35091 , n35093 );
and ( n35095 , n35084 , n35094 );
and ( n35096 , n24731 , n25617 );
and ( n35097 , n24624 , n26229 );
and ( n35098 , n35096 , n35097 );
and ( n35099 , n24337 , n26876 );
and ( n35100 , n35097 , n35099 );
and ( n35101 , n35096 , n35099 );
or ( n35102 , n35098 , n35100 , n35101 );
and ( n35103 , n26782 , n22337 );
and ( n35104 , n35102 , n35103 );
and ( n35105 , n26399 , n22784 );
and ( n35106 , n35103 , n35105 );
and ( n35107 , n35102 , n35105 );
or ( n35108 , n35104 , n35106 , n35107 );
and ( n35109 , n34419 , n34352 );
and ( n35110 , n34079 , n34350 );
nor ( n35111 , n35109 , n35110 );
xnor ( n35112 , n35111 , n28532 );
xor ( n35113 , n35051 , n35052 );
xor ( n35114 , n35113 , n35054 );
or ( n35115 , n35112 , n35114 );
and ( n35116 , n35108 , n35115 );
xor ( n35117 , n34865 , n34866 );
xor ( n35118 , n35117 , n34868 );
xor ( n35119 , n35085 , n35086 );
xor ( n35120 , n35119 , n35088 );
and ( n35121 , n35118 , n35120 );
and ( n35122 , n23742 , n28209 );
and ( n35123 , n23620 , n33739 );
and ( n35124 , n35122 , n35123 );
and ( n35125 , n23483 , n34122 );
and ( n35126 , n35123 , n35125 );
and ( n35127 , n35122 , n35125 );
or ( n35128 , n35124 , n35126 , n35127 );
and ( n35129 , n35120 , n35128 );
and ( n35130 , n35118 , n35128 );
or ( n35131 , n35121 , n35129 , n35130 );
and ( n35132 , n35115 , n35131 );
and ( n35133 , n35108 , n35131 );
or ( n35134 , n35116 , n35132 , n35133 );
and ( n35135 , n35094 , n35134 );
and ( n35136 , n35084 , n35134 );
or ( n35137 , n35095 , n35135 , n35136 );
and ( n35138 , n35079 , n35137 );
and ( n35139 , n35048 , n35137 );
or ( n35140 , n35080 , n35138 , n35139 );
and ( n35141 , n35037 , n35140 );
and ( n35142 , n35028 , n35140 );
or ( n35143 , n35038 , n35141 , n35142 );
and ( n35144 , n35025 , n35143 );
and ( n35145 , n35023 , n35143 );
or ( n35146 , n35026 , n35144 , n35145 );
and ( n35147 , n27591 , n21827 );
and ( n35148 , n26980 , n22172 );
and ( n35149 , n35147 , n35148 );
and ( n35150 , n26933 , n22337 );
and ( n35151 , n35148 , n35150 );
and ( n35152 , n35147 , n35150 );
or ( n35153 , n35149 , n35151 , n35152 );
buf ( n35154 , n23089 );
buf ( n35155 , n771 );
buf ( n35156 , n35155 );
buf ( n35157 , n772 );
buf ( n35158 , n35157 );
and ( n35159 , n35156 , n35158 );
not ( n35160 , n35159 );
and ( n35161 , n34658 , n35160 );
not ( n35162 , n35161 );
or ( n35163 , n35154 , n35162 );
and ( n35164 , n35153 , n35163 );
and ( n35165 , n25959 , n23508 );
and ( n35166 , n25623 , n24064 );
and ( n35167 , n35165 , n35166 );
buf ( n35168 , n12120 );
buf ( n35169 , n35168 );
and ( n35170 , n23215 , n35169 );
and ( n35171 , n35166 , n35170 );
and ( n35172 , n35165 , n35170 );
or ( n35173 , n35167 , n35171 , n35172 );
and ( n35174 , n35163 , n35173 );
and ( n35175 , n35153 , n35173 );
or ( n35176 , n35164 , n35174 , n35175 );
xor ( n35177 , n34907 , n34914 );
xor ( n35178 , n35177 , n34917 );
and ( n35179 , n35176 , n35178 );
xor ( n35180 , n34922 , n34927 );
xor ( n35181 , n35180 , n34930 );
and ( n35182 , n35178 , n35181 );
and ( n35183 , n35176 , n35181 );
or ( n35184 , n35179 , n35182 , n35183 );
xor ( n35185 , n34891 , n34893 );
xor ( n35186 , n35185 , n34902 );
and ( n35187 , n35184 , n35186 );
xor ( n35188 , n34920 , n34933 );
xor ( n35189 , n35188 , n34950 );
and ( n35190 , n35186 , n35189 );
and ( n35191 , n35184 , n35189 );
or ( n35192 , n35187 , n35190 , n35191 );
xor ( n35193 , n34815 , n34831 );
xor ( n35194 , n35193 , n34853 );
and ( n35195 , n35192 , n35194 );
xor ( n35196 , n34889 , n34905 );
xor ( n35197 , n35196 , n34953 );
and ( n35198 , n35194 , n35197 );
and ( n35199 , n35192 , n35197 );
or ( n35200 , n35195 , n35198 , n35199 );
xor ( n35201 , n34771 , n34772 );
xor ( n35202 , n35201 , n34784 );
and ( n35203 , n35200 , n35202 );
xor ( n35204 , n34813 , n34856 );
xor ( n35205 , n35204 , n34956 );
and ( n35206 , n35202 , n35205 );
and ( n35207 , n35200 , n35205 );
or ( n35208 , n35203 , n35206 , n35207 );
xor ( n35209 , n34766 , n34768 );
xor ( n35210 , n35209 , n34787 );
and ( n35211 , n35208 , n35210 );
xor ( n35212 , n34959 , n34985 );
xor ( n35213 , n35212 , n34988 );
and ( n35214 , n35210 , n35213 );
and ( n35215 , n35208 , n35213 );
or ( n35216 , n35211 , n35214 , n35215 );
and ( n35217 , n35146 , n35216 );
xor ( n35218 , n34764 , n34790 );
xor ( n35219 , n35218 , n34991 );
and ( n35220 , n35216 , n35219 );
and ( n35221 , n35146 , n35219 );
or ( n35222 , n35217 , n35220 , n35221 );
and ( n35223 , n35020 , n35222 );
and ( n35224 , n35018 , n35222 );
or ( n35225 , n35021 , n35223 , n35224 );
and ( n35226 , n35016 , n35225 );
xor ( n35227 , n34757 , n34759 );
xor ( n35228 , n35227 , n35008 );
and ( n35229 , n35225 , n35228 );
and ( n35230 , n35016 , n35228 );
or ( n35231 , n35226 , n35229 , n35230 );
and ( n35232 , n35013 , n35231 );
and ( n35233 , n35011 , n35231 );
or ( n35234 , n35014 , n35232 , n35233 );
and ( n35235 , n34754 , n35234 );
and ( n35236 , n34752 , n35234 );
or ( n35237 , n34755 , n35235 , n35236 );
and ( n35238 , n34492 , n35237 );
and ( n35239 , n34490 , n35237 );
or ( n35240 , n34493 , n35238 , n35239 );
and ( n35241 , n34208 , n35240 );
xor ( n35242 , n34208 , n35240 );
xor ( n35243 , n34490 , n34492 );
xor ( n35244 , n35243 , n35237 );
xor ( n35245 , n34752 , n34754 );
xor ( n35246 , n35245 , n35234 );
xor ( n35247 , n35011 , n35013 );
xor ( n35248 , n35247 , n35231 );
xor ( n35249 , n34762 , n34994 );
xor ( n35250 , n35249 , n35005 );
xor ( n35251 , n34997 , n34999 );
xor ( n35252 , n35251 , n35002 );
xor ( n35253 , n34977 , n34979 );
xor ( n35254 , n35253 , n34982 );
xor ( n35255 , n34969 , n34971 );
xor ( n35256 , n35255 , n34974 );
and ( n35257 , n34923 , n34924 );
and ( n35258 , n34924 , n34926 );
and ( n35259 , n34923 , n34926 );
or ( n35260 , n35257 , n35258 , n35259 );
and ( n35261 , n25220 , n25026 );
and ( n35262 , n24546 , n26376 );
and ( n35263 , n35261 , n35262 );
and ( n35264 , n23903 , n27558 );
and ( n35265 , n35262 , n35264 );
and ( n35266 , n35261 , n35264 );
or ( n35267 , n35263 , n35265 , n35266 );
and ( n35268 , n26678 , n22562 );
and ( n35269 , n35267 , n35268 );
and ( n35270 , n25623 , n23758 );
and ( n35271 , n35268 , n35270 );
and ( n35272 , n35267 , n35270 );
or ( n35273 , n35269 , n35271 , n35272 );
and ( n35274 , n23336 , n35169 );
buf ( n35275 , n35274 );
and ( n35276 , n24052 , n27246 );
and ( n35277 , n35275 , n35276 );
and ( n35278 , n23336 , n34817 );
and ( n35279 , n35276 , n35278 );
and ( n35280 , n35275 , n35278 );
or ( n35281 , n35277 , n35279 , n35280 );
and ( n35282 , n26148 , n22987 );
and ( n35283 , n35281 , n35282 );
and ( n35284 , n25959 , n23322 );
and ( n35285 , n35282 , n35284 );
and ( n35286 , n35281 , n35284 );
or ( n35287 , n35283 , n35285 , n35286 );
and ( n35288 , n35273 , n35287 );
and ( n35289 , n25451 , n24064 );
and ( n35290 , n25220 , n24540 );
and ( n35291 , n35289 , n35290 );
xor ( n35292 , n34792 , n34793 );
xor ( n35293 , n35292 , n34795 );
and ( n35294 , n35290 , n35293 );
and ( n35295 , n35289 , n35293 );
or ( n35296 , n35291 , n35294 , n35295 );
and ( n35297 , n35287 , n35296 );
and ( n35298 , n35273 , n35296 );
or ( n35299 , n35288 , n35297 , n35298 );
and ( n35300 , n35260 , n35299 );
and ( n35301 , n34637 , n28117 );
and ( n35302 , n35299 , n35301 );
and ( n35303 , n35260 , n35301 );
or ( n35304 , n35300 , n35302 , n35303 );
and ( n35305 , n35256 , n35304 );
xor ( n35306 , n34961 , n34963 );
xor ( n35307 , n35306 , n34966 );
xor ( n35308 , n34935 , n34944 );
xor ( n35309 , n35308 , n34947 );
xnor ( n35310 , n35073 , n35075 );
and ( n35311 , n35309 , n35310 );
xnor ( n35312 , n35081 , n35083 );
and ( n35313 , n35310 , n35312 );
and ( n35314 , n35309 , n35312 );
or ( n35315 , n35311 , n35313 , n35314 );
and ( n35316 , n35307 , n35315 );
xor ( n35317 , n35091 , n35093 );
and ( n35318 , n25451 , n25026 );
and ( n35319 , n24337 , n27246 );
and ( n35320 , n35318 , n35319 );
and ( n35321 , n24052 , n27558 );
and ( n35322 , n35319 , n35321 );
and ( n35323 , n35318 , n35321 );
or ( n35324 , n35320 , n35322 , n35323 );
and ( n35325 , n24624 , n26376 );
and ( n35326 , n23620 , n34122 );
and ( n35327 , n35325 , n35326 );
not ( n35328 , n35274 );
and ( n35329 , n35326 , n35328 );
and ( n35330 , n35325 , n35328 );
or ( n35331 , n35327 , n35329 , n35330 );
and ( n35332 , n35324 , n35331 );
and ( n35333 , n26399 , n22987 );
and ( n35334 , n35331 , n35333 );
and ( n35335 , n35324 , n35333 );
or ( n35336 , n35332 , n35334 , n35335 );
and ( n35337 , n26148 , n23322 );
and ( n35338 , n25742 , n23758 );
and ( n35339 , n35337 , n35338 );
xor ( n35340 , n35122 , n35123 );
xor ( n35341 , n35340 , n35125 );
and ( n35342 , n35338 , n35341 );
and ( n35343 , n35337 , n35341 );
or ( n35344 , n35339 , n35342 , n35343 );
and ( n35345 , n35336 , n35344 );
and ( n35346 , n27962 , n21429 );
and ( n35347 , n35344 , n35346 );
and ( n35348 , n35336 , n35346 );
or ( n35349 , n35345 , n35347 , n35348 );
and ( n35350 , n35317 , n35349 );
xor ( n35351 , n35067 , n35068 );
xor ( n35352 , n35351 , n35070 );
xor ( n35353 , n34872 , n34873 );
xor ( n35354 , n35353 , n34875 );
and ( n35355 , n35352 , n35354 );
xor ( n35356 , n35289 , n35290 );
xor ( n35357 , n35356 , n35293 );
and ( n35358 , n35354 , n35357 );
and ( n35359 , n35352 , n35357 );
or ( n35360 , n35355 , n35358 , n35359 );
and ( n35361 , n35349 , n35360 );
and ( n35362 , n35317 , n35360 );
or ( n35363 , n35350 , n35361 , n35362 );
and ( n35364 , n35315 , n35363 );
and ( n35365 , n35307 , n35363 );
or ( n35366 , n35316 , n35364 , n35365 );
and ( n35367 , n35304 , n35366 );
and ( n35368 , n35256 , n35366 );
or ( n35369 , n35305 , n35367 , n35368 );
and ( n35370 , n35254 , n35369 );
xor ( n35371 , n34101 , n34656 );
xor ( n35372 , n34656 , n34658 );
not ( n35373 , n35372 );
and ( n35374 , n35371 , n35373 );
and ( n35375 , n33628 , n35374 );
not ( n35376 , n35375 );
xnor ( n35377 , n35376 , n34661 );
and ( n35378 , n34637 , n34352 );
and ( n35379 , n34419 , n34350 );
nor ( n35380 , n35378 , n35379 );
xnor ( n35381 , n35380 , n28532 );
and ( n35382 , n35377 , n35381 );
xor ( n35383 , n31455 , n33618 );
buf ( n35384 , n35383 );
buf ( n35385 , n35384 );
buf ( n35386 , n35385 );
and ( n35387 , n35386 , n33632 );
and ( n35388 , n34646 , n33630 );
nor ( n35389 , n35387 , n35388 );
xnor ( n35390 , n35389 , n28124 );
and ( n35391 , n35381 , n35390 );
and ( n35392 , n35377 , n35390 );
or ( n35393 , n35382 , n35391 , n35392 );
xor ( n35394 , n34936 , n34661 );
xor ( n35395 , n35394 , n34941 );
and ( n35396 , n35393 , n35395 );
xnor ( n35397 , n35112 , n35114 );
and ( n35398 , n35395 , n35397 );
and ( n35399 , n35393 , n35397 );
or ( n35400 , n35396 , n35398 , n35399 );
and ( n35401 , n23903 , n28209 );
and ( n35402 , n23742 , n33739 );
and ( n35403 , n35401 , n35402 );
and ( n35404 , n23483 , n34817 );
and ( n35405 , n35402 , n35404 );
and ( n35406 , n35401 , n35404 );
or ( n35407 , n35403 , n35405 , n35406 );
and ( n35408 , n25451 , n24540 );
and ( n35409 , n35407 , n35408 );
and ( n35410 , n24993 , n25284 );
and ( n35411 , n35408 , n35410 );
and ( n35412 , n35407 , n35410 );
or ( n35413 , n35409 , n35411 , n35412 );
and ( n35414 , n25742 , n24064 );
and ( n35415 , n25623 , n24540 );
and ( n35416 , n35414 , n35415 );
and ( n35417 , n25220 , n25284 );
and ( n35418 , n35415 , n35417 );
and ( n35419 , n35414 , n35417 );
or ( n35420 , n35416 , n35418 , n35419 );
and ( n35421 , n27863 , n21666 );
and ( n35422 , n35420 , n35421 );
and ( n35423 , n27389 , n21990 );
and ( n35424 , n35421 , n35423 );
and ( n35425 , n35420 , n35423 );
or ( n35426 , n35422 , n35424 , n35425 );
and ( n35427 , n35413 , n35426 );
xnor ( n35428 , n35154 , n35162 );
and ( n35429 , n27863 , n21827 );
and ( n35430 , n27389 , n22172 );
and ( n35431 , n35429 , n35430 );
and ( n35432 , n26980 , n22337 );
and ( n35433 , n35430 , n35432 );
and ( n35434 , n35429 , n35432 );
or ( n35435 , n35431 , n35433 , n35434 );
and ( n35436 , n35428 , n35435 );
and ( n35437 , n26678 , n22987 );
and ( n35438 , n35437 , n35161 );
and ( n35439 , n34419 , n34911 );
and ( n35440 , n34079 , n34909 );
nor ( n35441 , n35439 , n35440 );
xnor ( n35442 , n35441 , n34104 );
and ( n35443 , n35161 , n35442 );
and ( n35444 , n35437 , n35442 );
or ( n35445 , n35438 , n35443 , n35444 );
and ( n35446 , n35435 , n35445 );
and ( n35447 , n35428 , n35445 );
or ( n35448 , n35436 , n35446 , n35447 );
and ( n35449 , n35426 , n35448 );
and ( n35450 , n35413 , n35448 );
or ( n35451 , n35427 , n35449 , n35450 );
and ( n35452 , n35400 , n35451 );
xor ( n35453 , n35108 , n35115 );
xor ( n35454 , n35453 , n35131 );
and ( n35455 , n35451 , n35454 );
and ( n35456 , n35400 , n35454 );
or ( n35457 , n35452 , n35455 , n35456 );
xor ( n35458 , n35040 , n35042 );
xor ( n35459 , n35458 , n35045 );
and ( n35460 , n35457 , n35459 );
xor ( n35461 , n35050 , n35065 );
xor ( n35462 , n35461 , n35076 );
and ( n35463 , n35459 , n35462 );
and ( n35464 , n35457 , n35462 );
or ( n35465 , n35460 , n35463 , n35464 );
xor ( n35466 , n35030 , n35032 );
xor ( n35467 , n35466 , n35034 );
and ( n35468 , n35465 , n35467 );
xor ( n35469 , n35048 , n35079 );
xor ( n35470 , n35469 , n35137 );
and ( n35471 , n35467 , n35470 );
and ( n35472 , n35465 , n35470 );
or ( n35473 , n35468 , n35471 , n35472 );
and ( n35474 , n35369 , n35473 );
and ( n35475 , n35254 , n35473 );
or ( n35476 , n35370 , n35474 , n35475 );
xor ( n35477 , n35023 , n35025 );
xor ( n35478 , n35477 , n35143 );
and ( n35479 , n35476 , n35478 );
xor ( n35480 , n35208 , n35210 );
xor ( n35481 , n35480 , n35213 );
and ( n35482 , n35478 , n35481 );
and ( n35483 , n35476 , n35481 );
or ( n35484 , n35479 , n35482 , n35483 );
and ( n35485 , n35252 , n35484 );
xor ( n35486 , n35146 , n35216 );
xor ( n35487 , n35486 , n35219 );
and ( n35488 , n35484 , n35487 );
and ( n35489 , n35252 , n35487 );
or ( n35490 , n35485 , n35488 , n35489 );
and ( n35491 , n35250 , n35490 );
xor ( n35492 , n35018 , n35020 );
xor ( n35493 , n35492 , n35222 );
and ( n35494 , n35490 , n35493 );
and ( n35495 , n35250 , n35493 );
or ( n35496 , n35491 , n35494 , n35495 );
xor ( n35497 , n35016 , n35225 );
xor ( n35498 , n35497 , n35228 );
and ( n35499 , n35496 , n35498 );
xor ( n35500 , n35496 , n35498 );
xor ( n35501 , n35250 , n35490 );
xor ( n35502 , n35501 , n35493 );
xor ( n35503 , n35252 , n35484 );
xor ( n35504 , n35503 , n35487 );
xor ( n35505 , n35028 , n35037 );
xor ( n35506 , n35505 , n35140 );
xor ( n35507 , n35200 , n35202 );
xor ( n35508 , n35507 , n35205 );
and ( n35509 , n35506 , n35508 );
xor ( n35510 , n35192 , n35194 );
xor ( n35511 , n35510 , n35197 );
xor ( n35512 , n35084 , n35094 );
xor ( n35513 , n35512 , n35134 );
xor ( n35514 , n35184 , n35186 );
xor ( n35515 , n35514 , n35189 );
and ( n35516 , n35513 , n35515 );
xor ( n35517 , n35260 , n35299 );
xor ( n35518 , n35517 , n35301 );
and ( n35519 , n35515 , n35518 );
and ( n35520 , n35513 , n35518 );
or ( n35521 , n35516 , n35519 , n35520 );
and ( n35522 , n35511 , n35521 );
and ( n35523 , n35386 , n28117 );
xor ( n35524 , n35267 , n35268 );
xor ( n35525 , n35524 , n35270 );
and ( n35526 , n35523 , n35525 );
xor ( n35527 , n35281 , n35282 );
xor ( n35528 , n35527 , n35284 );
and ( n35529 , n35525 , n35528 );
and ( n35530 , n35523 , n35528 );
or ( n35531 , n35526 , n35529 , n35530 );
xor ( n35532 , n35057 , n35059 );
xor ( n35533 , n35532 , n35062 );
and ( n35534 , n35531 , n35533 );
xor ( n35535 , n35176 , n35178 );
xor ( n35536 , n35535 , n35181 );
xor ( n35537 , n35273 , n35287 );
xor ( n35538 , n35537 , n35296 );
and ( n35539 , n35536 , n35538 );
and ( n35540 , n23742 , n34122 );
and ( n35541 , n23620 , n34817 );
and ( n35542 , n35540 , n35541 );
buf ( n35543 , n12619 );
buf ( n35544 , n35543 );
and ( n35545 , n23336 , n35544 );
and ( n35546 , n35541 , n35545 );
and ( n35547 , n35540 , n35545 );
or ( n35548 , n35542 , n35546 , n35547 );
and ( n35549 , n26148 , n23508 );
and ( n35550 , n35548 , n35549 );
and ( n35551 , n24993 , n25617 );
and ( n35552 , n35549 , n35551 );
and ( n35553 , n35548 , n35551 );
or ( n35554 , n35550 , n35552 , n35553 );
xor ( n35555 , n35261 , n35262 );
xor ( n35556 , n35555 , n35264 );
and ( n35557 , n35554 , n35556 );
xor ( n35558 , n35275 , n35276 );
xor ( n35559 , n35558 , n35278 );
and ( n35560 , n35556 , n35559 );
and ( n35561 , n35554 , n35559 );
or ( n35562 , n35557 , n35560 , n35561 );
and ( n35563 , n34038 , n34911 );
and ( n35564 , n33628 , n34909 );
nor ( n35565 , n35563 , n35564 );
xnor ( n35566 , n35565 , n34104 );
and ( n35567 , n35562 , n35566 );
xor ( n35568 , n35102 , n35103 );
xor ( n35569 , n35568 , n35105 );
and ( n35570 , n35566 , n35569 );
and ( n35571 , n35562 , n35569 );
or ( n35572 , n35567 , n35570 , n35571 );
and ( n35573 , n35538 , n35572 );
and ( n35574 , n35536 , n35572 );
or ( n35575 , n35539 , n35573 , n35574 );
and ( n35576 , n35534 , n35575 );
and ( n35577 , n28129 , n21429 );
and ( n35578 , n27962 , n21527 );
and ( n35579 , n35577 , n35578 );
xor ( n35580 , n35096 , n35097 );
xor ( n35581 , n35580 , n35099 );
and ( n35582 , n35578 , n35581 );
and ( n35583 , n35577 , n35581 );
or ( n35584 , n35579 , n35582 , n35583 );
xor ( n35585 , n35336 , n35344 );
xor ( n35586 , n35585 , n35346 );
or ( n35587 , n35584 , n35586 );
xor ( n35588 , n35118 , n35120 );
xor ( n35589 , n35588 , n35128 );
xor ( n35590 , n35153 , n35163 );
xor ( n35591 , n35590 , n35173 );
and ( n35592 , n35589 , n35591 );
xor ( n35593 , n35352 , n35354 );
xor ( n35594 , n35593 , n35357 );
and ( n35595 , n35591 , n35594 );
and ( n35596 , n35589 , n35594 );
or ( n35597 , n35592 , n35595 , n35596 );
and ( n35598 , n35587 , n35597 );
and ( n35599 , n23483 , n35169 );
buf ( n35600 , n23215 );
and ( n35601 , n35599 , n35600 );
buf ( n35602 , n773 );
buf ( n35603 , n35602 );
buf ( n35604 , n774 );
buf ( n35605 , n35604 );
and ( n35606 , n35603 , n35605 );
not ( n35607 , n35606 );
and ( n35608 , n35158 , n35607 );
not ( n35609 , n35608 );
and ( n35610 , n35600 , n35609 );
and ( n35611 , n35599 , n35609 );
or ( n35612 , n35601 , n35610 , n35611 );
and ( n35613 , n24731 , n26229 );
and ( n35614 , n35612 , n35613 );
and ( n35615 , n24546 , n26876 );
and ( n35616 , n35613 , n35615 );
and ( n35617 , n35612 , n35615 );
or ( n35618 , n35614 , n35616 , n35617 );
and ( n35619 , n26782 , n22562 );
and ( n35620 , n35618 , n35619 );
and ( n35621 , n26678 , n22784 );
and ( n35622 , n35619 , n35621 );
and ( n35623 , n35618 , n35621 );
or ( n35624 , n35620 , n35622 , n35623 );
xor ( n35625 , n35165 , n35166 );
xor ( n35626 , n35625 , n35170 );
xor ( n35627 , n35377 , n35381 );
xor ( n35628 , n35627 , n35390 );
and ( n35629 , n35626 , n35628 );
xor ( n35630 , n35407 , n35408 );
xor ( n35631 , n35630 , n35410 );
and ( n35632 , n35628 , n35631 );
and ( n35633 , n35626 , n35631 );
or ( n35634 , n35629 , n35632 , n35633 );
and ( n35635 , n35624 , n35634 );
xor ( n35636 , n35420 , n35421 );
xor ( n35637 , n35636 , n35423 );
xor ( n35638 , n35577 , n35578 );
xor ( n35639 , n35638 , n35581 );
and ( n35640 , n35637 , n35639 );
and ( n35641 , n25623 , n25026 );
and ( n35642 , n24993 , n26229 );
and ( n35643 , n35641 , n35642 );
and ( n35644 , n24624 , n26876 );
and ( n35645 , n35642 , n35644 );
and ( n35646 , n35641 , n35644 );
or ( n35647 , n35643 , n35645 , n35646 );
and ( n35648 , n26933 , n22562 );
and ( n35649 , n35647 , n35648 );
and ( n35650 , n26782 , n22784 );
and ( n35651 , n35648 , n35650 );
and ( n35652 , n35647 , n35650 );
or ( n35653 , n35649 , n35651 , n35652 );
and ( n35654 , n35639 , n35653 );
and ( n35655 , n35637 , n35653 );
or ( n35656 , n35640 , n35654 , n35655 );
and ( n35657 , n35634 , n35656 );
and ( n35658 , n35624 , n35656 );
or ( n35659 , n35635 , n35657 , n35658 );
and ( n35660 , n35597 , n35659 );
and ( n35661 , n35587 , n35659 );
or ( n35662 , n35598 , n35660 , n35661 );
and ( n35663 , n35575 , n35662 );
and ( n35664 , n35534 , n35662 );
or ( n35665 , n35576 , n35663 , n35664 );
and ( n35666 , n35521 , n35665 );
and ( n35667 , n35511 , n35665 );
or ( n35668 , n35522 , n35666 , n35667 );
and ( n35669 , n35508 , n35668 );
and ( n35670 , n35506 , n35668 );
or ( n35671 , n35509 , n35669 , n35670 );
xor ( n35672 , n35476 , n35478 );
xor ( n35673 , n35672 , n35481 );
and ( n35674 , n35671 , n35673 );
and ( n35675 , n26399 , n23322 );
and ( n35676 , n25959 , n23758 );
and ( n35677 , n35675 , n35676 );
xor ( n35678 , n35401 , n35402 );
xor ( n35679 , n35678 , n35404 );
and ( n35680 , n35676 , n35679 );
and ( n35681 , n35675 , n35679 );
or ( n35682 , n35677 , n35680 , n35681 );
and ( n35683 , n34646 , n34352 );
and ( n35684 , n34637 , n34350 );
nor ( n35685 , n35683 , n35684 );
xnor ( n35686 , n35685 , n28532 );
xor ( n35687 , n31459 , n33616 );
buf ( n35688 , n35687 );
buf ( n35689 , n35688 );
buf ( n35690 , n35689 );
and ( n35691 , n35690 , n28117 );
and ( n35692 , n35686 , n35691 );
xor ( n35693 , n35429 , n35430 );
xor ( n35694 , n35693 , n35432 );
and ( n35695 , n35691 , n35694 );
and ( n35696 , n35686 , n35694 );
or ( n35697 , n35692 , n35695 , n35696 );
and ( n35698 , n35682 , n35697 );
and ( n35699 , n24337 , n27558 );
and ( n35700 , n24052 , n28209 );
and ( n35701 , n35699 , n35700 );
and ( n35702 , n23903 , n33739 );
and ( n35703 , n35700 , n35702 );
and ( n35704 , n35699 , n35702 );
or ( n35705 , n35701 , n35703 , n35704 );
and ( n35706 , n34079 , n35374 );
and ( n35707 , n34038 , n35372 );
nor ( n35708 , n35706 , n35707 );
xnor ( n35709 , n35708 , n34661 );
and ( n35710 , n34637 , n34911 );
and ( n35711 , n34419 , n34909 );
nor ( n35712 , n35710 , n35711 );
xnor ( n35713 , n35712 , n34104 );
and ( n35714 , n35709 , n35713 );
xor ( n35715 , n31461 , n33615 );
buf ( n35716 , n35715 );
buf ( n35717 , n35716 );
buf ( n35718 , n35717 );
and ( n35719 , n35718 , n28117 );
and ( n35720 , n35713 , n35719 );
and ( n35721 , n35709 , n35719 );
or ( n35722 , n35714 , n35720 , n35721 );
and ( n35723 , n35705 , n35722 );
and ( n35724 , n27962 , n21827 );
and ( n35725 , n27591 , n22172 );
and ( n35726 , n35724 , n35725 );
and ( n35727 , n26678 , n23322 );
and ( n35728 , n35725 , n35727 );
and ( n35729 , n35724 , n35727 );
or ( n35730 , n35726 , n35728 , n35729 );
and ( n35731 , n35722 , n35730 );
and ( n35732 , n35705 , n35730 );
or ( n35733 , n35723 , n35731 , n35732 );
and ( n35734 , n35697 , n35733 );
and ( n35735 , n35682 , n35733 );
or ( n35736 , n35698 , n35734 , n35735 );
xor ( n35737 , n35393 , n35395 );
xor ( n35738 , n35737 , n35397 );
and ( n35739 , n35736 , n35738 );
xor ( n35740 , n35413 , n35426 );
xor ( n35741 , n35740 , n35448 );
and ( n35742 , n35738 , n35741 );
and ( n35743 , n35736 , n35741 );
or ( n35744 , n35739 , n35742 , n35743 );
xor ( n35745 , n35309 , n35310 );
xor ( n35746 , n35745 , n35312 );
and ( n35747 , n35744 , n35746 );
xor ( n35748 , n35317 , n35349 );
xor ( n35749 , n35748 , n35360 );
and ( n35750 , n35746 , n35749 );
and ( n35751 , n35744 , n35749 );
or ( n35752 , n35747 , n35750 , n35751 );
xor ( n35753 , n35307 , n35315 );
xor ( n35754 , n35753 , n35363 );
and ( n35755 , n35752 , n35754 );
xor ( n35756 , n35457 , n35459 );
xor ( n35757 , n35756 , n35462 );
and ( n35758 , n35754 , n35757 );
and ( n35759 , n35752 , n35757 );
or ( n35760 , n35755 , n35758 , n35759 );
xor ( n35761 , n35256 , n35304 );
xor ( n35762 , n35761 , n35366 );
and ( n35763 , n35760 , n35762 );
xor ( n35764 , n35465 , n35467 );
xor ( n35765 , n35764 , n35470 );
and ( n35766 , n35762 , n35765 );
and ( n35767 , n35760 , n35765 );
or ( n35768 , n35763 , n35766 , n35767 );
xor ( n35769 , n35254 , n35369 );
xor ( n35770 , n35769 , n35473 );
and ( n35771 , n35768 , n35770 );
xor ( n35772 , n35400 , n35451 );
xor ( n35773 , n35772 , n35454 );
xor ( n35774 , n35531 , n35533 );
and ( n35775 , n35773 , n35774 );
and ( n35776 , n34079 , n34911 );
and ( n35777 , n34038 , n34909 );
nor ( n35778 , n35776 , n35777 );
xnor ( n35779 , n35778 , n34104 );
xor ( n35780 , n35324 , n35331 );
xor ( n35781 , n35780 , n35333 );
and ( n35782 , n35779 , n35781 );
xor ( n35783 , n35337 , n35338 );
xor ( n35784 , n35783 , n35341 );
and ( n35785 , n35781 , n35784 );
and ( n35786 , n35779 , n35784 );
or ( n35787 , n35782 , n35785 , n35786 );
xor ( n35788 , n35523 , n35525 );
xor ( n35789 , n35788 , n35528 );
or ( n35790 , n35787 , n35789 );
and ( n35791 , n35774 , n35790 );
and ( n35792 , n35773 , n35790 );
or ( n35793 , n35775 , n35791 , n35792 );
xor ( n35794 , n35562 , n35566 );
xor ( n35795 , n35794 , n35569 );
xnor ( n35796 , n35584 , n35586 );
and ( n35797 , n35795 , n35796 );
xor ( n35798 , n35147 , n35148 );
xor ( n35799 , n35798 , n35150 );
xor ( n35800 , n35618 , n35619 );
xor ( n35801 , n35800 , n35621 );
and ( n35802 , n35799 , n35801 );
xor ( n35803 , n35554 , n35556 );
xor ( n35804 , n35803 , n35559 );
and ( n35805 , n35801 , n35804 );
and ( n35806 , n35799 , n35804 );
or ( n35807 , n35802 , n35805 , n35806 );
and ( n35808 , n35796 , n35807 );
and ( n35809 , n35795 , n35807 );
or ( n35810 , n35797 , n35808 , n35809 );
and ( n35811 , n34038 , n35374 );
and ( n35812 , n33628 , n35372 );
nor ( n35813 , n35811 , n35812 );
xnor ( n35814 , n35813 , n34661 );
xor ( n35815 , n31457 , n33617 );
buf ( n35816 , n35815 );
buf ( n35817 , n35816 );
buf ( n35818 , n35817 );
and ( n35819 , n35818 , n33632 );
and ( n35820 , n35386 , n33630 );
nor ( n35821 , n35819 , n35820 );
xnor ( n35822 , n35821 , n28124 );
and ( n35823 , n35814 , n35822 );
xor ( n35824 , n35647 , n35648 );
xor ( n35825 , n35824 , n35650 );
and ( n35826 , n35822 , n35825 );
and ( n35827 , n35814 , n35825 );
or ( n35828 , n35823 , n35826 , n35827 );
xor ( n35829 , n35779 , n35781 );
xor ( n35830 , n35829 , n35784 );
or ( n35831 , n35828 , n35830 );
and ( n35832 , n25742 , n24540 );
and ( n35833 , n25220 , n25617 );
and ( n35834 , n35832 , n35833 );
xor ( n35835 , n35599 , n35600 );
xor ( n35836 , n35835 , n35609 );
and ( n35837 , n35833 , n35836 );
and ( n35838 , n35832 , n35836 );
or ( n35839 , n35834 , n35837 , n35838 );
xor ( n35840 , n35318 , n35319 );
xor ( n35841 , n35840 , n35321 );
and ( n35842 , n35839 , n35841 );
xor ( n35843 , n35325 , n35326 );
xor ( n35844 , n35843 , n35328 );
and ( n35845 , n35841 , n35844 );
and ( n35846 , n35839 , n35844 );
or ( n35847 , n35842 , n35845 , n35846 );
and ( n35848 , n35818 , n28117 );
and ( n35849 , n35847 , n35848 );
and ( n35850 , n35831 , n35849 );
xor ( n35851 , n35428 , n35435 );
xor ( n35852 , n35851 , n35445 );
and ( n35853 , n24052 , n33739 );
and ( n35854 , n23903 , n34122 );
and ( n35855 , n35853 , n35854 );
and ( n35856 , n23483 , n35544 );
and ( n35857 , n35854 , n35856 );
and ( n35858 , n35853 , n35856 );
or ( n35859 , n35855 , n35857 , n35858 );
and ( n35860 , n26399 , n23508 );
and ( n35861 , n35859 , n35860 );
and ( n35862 , n25959 , n24064 );
and ( n35863 , n35860 , n35862 );
and ( n35864 , n35859 , n35862 );
or ( n35865 , n35861 , n35863 , n35864 );
and ( n35866 , n27962 , n21666 );
and ( n35867 , n35865 , n35866 );
and ( n35868 , n27591 , n21990 );
and ( n35869 , n35866 , n35868 );
and ( n35870 , n35865 , n35868 );
or ( n35871 , n35867 , n35869 , n35870 );
and ( n35872 , n35852 , n35871 );
and ( n35873 , n28129 , n21527 );
xor ( n35874 , n35414 , n35415 );
xor ( n35875 , n35874 , n35417 );
and ( n35876 , n35873 , n35875 );
xor ( n35877 , n35612 , n35613 );
xor ( n35878 , n35877 , n35615 );
and ( n35879 , n35875 , n35878 );
and ( n35880 , n35873 , n35878 );
or ( n35881 , n35876 , n35879 , n35880 );
and ( n35882 , n35871 , n35881 );
and ( n35883 , n35852 , n35881 );
or ( n35884 , n35872 , n35882 , n35883 );
and ( n35885 , n35849 , n35884 );
and ( n35886 , n35831 , n35884 );
or ( n35887 , n35850 , n35885 , n35886 );
and ( n35888 , n35810 , n35887 );
and ( n35889 , n25742 , n25026 );
and ( n35890 , n24731 , n26876 );
and ( n35891 , n35889 , n35890 );
and ( n35892 , n24546 , n27558 );
and ( n35893 , n35890 , n35892 );
and ( n35894 , n35889 , n35892 );
or ( n35895 , n35891 , n35893 , n35894 );
and ( n35896 , n27389 , n22337 );
and ( n35897 , n35895 , n35896 );
and ( n35898 , n26933 , n22784 );
and ( n35899 , n35896 , n35898 );
and ( n35900 , n35895 , n35898 );
or ( n35901 , n35897 , n35899 , n35900 );
xor ( n35902 , n35548 , n35549 );
xor ( n35903 , n35902 , n35551 );
or ( n35904 , n35901 , n35903 );
and ( n35905 , n24731 , n26376 );
and ( n35906 , n24546 , n27246 );
and ( n35907 , n35905 , n35906 );
xor ( n35908 , n34658 , n35156 );
xor ( n35909 , n35156 , n35158 );
not ( n35910 , n35909 );
and ( n35911 , n35908 , n35910 );
and ( n35912 , n33628 , n35911 );
not ( n35913 , n35912 );
xnor ( n35914 , n35913 , n35161 );
and ( n35915 , n35906 , n35914 );
and ( n35916 , n35905 , n35914 );
or ( n35917 , n35907 , n35915 , n35916 );
xor ( n35918 , n35437 , n35161 );
xor ( n35919 , n35918 , n35442 );
and ( n35920 , n35917 , n35919 );
xor ( n35921 , n35675 , n35676 );
xor ( n35922 , n35921 , n35679 );
and ( n35923 , n35919 , n35922 );
and ( n35924 , n35917 , n35922 );
or ( n35925 , n35920 , n35923 , n35924 );
and ( n35926 , n35904 , n35925 );
and ( n35927 , n26980 , n22562 );
and ( n35928 , n26782 , n22987 );
and ( n35929 , n35927 , n35928 );
xor ( n35930 , n35699 , n35700 );
xor ( n35931 , n35930 , n35702 );
and ( n35932 , n35928 , n35931 );
and ( n35933 , n35927 , n35931 );
or ( n35934 , n35929 , n35932 , n35933 );
and ( n35935 , n26148 , n23758 );
and ( n35936 , n25451 , n25284 );
and ( n35937 , n35935 , n35936 );
xor ( n35938 , n35540 , n35541 );
xor ( n35939 , n35938 , n35545 );
and ( n35940 , n35936 , n35939 );
and ( n35941 , n35935 , n35939 );
or ( n35942 , n35937 , n35940 , n35941 );
and ( n35943 , n35934 , n35942 );
and ( n35944 , n35386 , n34352 );
and ( n35945 , n34646 , n34350 );
nor ( n35946 , n35944 , n35945 );
xnor ( n35947 , n35946 , n28532 );
and ( n35948 , n35690 , n33632 );
and ( n35949 , n35818 , n33630 );
nor ( n35950 , n35948 , n35949 );
xnor ( n35951 , n35950 , n28124 );
and ( n35952 , n35947 , n35951 );
xor ( n35953 , n35709 , n35713 );
xor ( n35954 , n35953 , n35719 );
and ( n35955 , n35951 , n35954 );
and ( n35956 , n35947 , n35954 );
or ( n35957 , n35952 , n35955 , n35956 );
and ( n35958 , n35942 , n35957 );
and ( n35959 , n35934 , n35957 );
or ( n35960 , n35943 , n35958 , n35959 );
and ( n35961 , n35925 , n35960 );
and ( n35962 , n35904 , n35960 );
or ( n35963 , n35926 , n35961 , n35962 );
and ( n35964 , n24624 , n27246 );
and ( n35965 , n24337 , n28209 );
and ( n35966 , n35964 , n35965 );
and ( n35967 , n23742 , n34817 );
and ( n35968 , n35965 , n35967 );
and ( n35969 , n35964 , n35967 );
or ( n35970 , n35966 , n35968 , n35969 );
and ( n35971 , n28129 , n21827 );
and ( n35972 , n27863 , n22172 );
and ( n35973 , n35971 , n35972 );
and ( n35974 , n27591 , n22337 );
and ( n35975 , n35972 , n35974 );
and ( n35976 , n35971 , n35974 );
or ( n35977 , n35973 , n35975 , n35976 );
and ( n35978 , n35970 , n35977 );
and ( n35979 , n26782 , n23322 );
and ( n35980 , n26399 , n23758 );
and ( n35981 , n35979 , n35980 );
and ( n35982 , n24993 , n26376 );
and ( n35983 , n35980 , n35982 );
and ( n35984 , n35979 , n35982 );
or ( n35985 , n35981 , n35983 , n35984 );
and ( n35986 , n35977 , n35985 );
and ( n35987 , n35970 , n35985 );
or ( n35988 , n35978 , n35986 , n35987 );
and ( n35989 , n23620 , n35169 );
and ( n35990 , n35989 , n35608 );
and ( n35991 , n34038 , n35911 );
and ( n35992 , n33628 , n35909 );
nor ( n35993 , n35991 , n35992 );
xnor ( n35994 , n35993 , n35161 );
and ( n35995 , n35608 , n35994 );
and ( n35996 , n35989 , n35994 );
or ( n35997 , n35990 , n35995 , n35996 );
and ( n35998 , n34419 , n35374 );
and ( n35999 , n34079 , n35372 );
nor ( n36000 , n35998 , n35999 );
xnor ( n36001 , n36000 , n34661 );
and ( n36002 , n34646 , n34911 );
and ( n36003 , n34637 , n34909 );
nor ( n36004 , n36002 , n36003 );
xnor ( n36005 , n36004 , n34104 );
and ( n36006 , n36001 , n36005 );
and ( n36007 , n35818 , n34352 );
and ( n36008 , n35386 , n34350 );
nor ( n36009 , n36007 , n36008 );
xnor ( n36010 , n36009 , n28532 );
and ( n36011 , n36005 , n36010 );
and ( n36012 , n36001 , n36010 );
or ( n36013 , n36006 , n36011 , n36012 );
and ( n36014 , n35997 , n36013 );
xor ( n36015 , n35724 , n35725 );
xor ( n36016 , n36015 , n35727 );
and ( n36017 , n36013 , n36016 );
and ( n36018 , n35997 , n36016 );
or ( n36019 , n36014 , n36017 , n36018 );
and ( n36020 , n35988 , n36019 );
xor ( n36021 , n35686 , n35691 );
xor ( n36022 , n36021 , n35694 );
and ( n36023 , n36019 , n36022 );
and ( n36024 , n35988 , n36022 );
or ( n36025 , n36020 , n36023 , n36024 );
xor ( n36026 , n35626 , n35628 );
xor ( n36027 , n36026 , n35631 );
and ( n36028 , n36025 , n36027 );
xor ( n36029 , n35637 , n35639 );
xor ( n36030 , n36029 , n35653 );
and ( n36031 , n36027 , n36030 );
and ( n36032 , n36025 , n36030 );
or ( n36033 , n36028 , n36031 , n36032 );
and ( n36034 , n35963 , n36033 );
xor ( n36035 , n35589 , n35591 );
xor ( n36036 , n36035 , n35594 );
and ( n36037 , n36033 , n36036 );
and ( n36038 , n35963 , n36036 );
or ( n36039 , n36034 , n36037 , n36038 );
and ( n36040 , n35887 , n36039 );
and ( n36041 , n35810 , n36039 );
or ( n36042 , n35888 , n36040 , n36041 );
and ( n36043 , n35793 , n36042 );
xor ( n36044 , n35536 , n35538 );
xor ( n36045 , n36044 , n35572 );
xor ( n36046 , n35587 , n35597 );
xor ( n36047 , n36046 , n35659 );
and ( n36048 , n36045 , n36047 );
xor ( n36049 , n35744 , n35746 );
xor ( n36050 , n36049 , n35749 );
and ( n36051 , n36047 , n36050 );
and ( n36052 , n36045 , n36050 );
or ( n36053 , n36048 , n36051 , n36052 );
and ( n36054 , n36042 , n36053 );
and ( n36055 , n35793 , n36053 );
or ( n36056 , n36043 , n36054 , n36055 );
xor ( n36057 , n35513 , n35515 );
xor ( n36058 , n36057 , n35518 );
xor ( n36059 , n35534 , n35575 );
xor ( n36060 , n36059 , n35662 );
and ( n36061 , n36058 , n36060 );
xor ( n36062 , n35752 , n35754 );
xor ( n36063 , n36062 , n35757 );
and ( n36064 , n36060 , n36063 );
and ( n36065 , n36058 , n36063 );
or ( n36066 , n36061 , n36064 , n36065 );
and ( n36067 , n36056 , n36066 );
xor ( n36068 , n35511 , n35521 );
xor ( n36069 , n36068 , n35665 );
and ( n36070 , n36066 , n36069 );
and ( n36071 , n36056 , n36069 );
or ( n36072 , n36067 , n36070 , n36071 );
and ( n36073 , n35770 , n36072 );
and ( n36074 , n35768 , n36072 );
or ( n36075 , n35771 , n36073 , n36074 );
and ( n36076 , n35673 , n36075 );
and ( n36077 , n35671 , n36075 );
or ( n36078 , n35674 , n36076 , n36077 );
and ( n36079 , n35504 , n36078 );
xor ( n36080 , n35506 , n35508 );
xor ( n36081 , n36080 , n35668 );
xor ( n36082 , n35760 , n35762 );
xor ( n36083 , n36082 , n35765 );
xor ( n36084 , n35624 , n35634 );
xor ( n36085 , n36084 , n35656 );
xor ( n36086 , n35736 , n35738 );
xor ( n36087 , n36086 , n35741 );
and ( n36088 , n36085 , n36087 );
xnor ( n36089 , n35787 , n35789 );
and ( n36090 , n36087 , n36089 );
and ( n36091 , n36085 , n36089 );
or ( n36092 , n36088 , n36090 , n36091 );
xor ( n36093 , n35682 , n35697 );
xor ( n36094 , n36093 , n35733 );
xor ( n36095 , n35799 , n35801 );
xor ( n36096 , n36095 , n35804 );
and ( n36097 , n36094 , n36096 );
xnor ( n36098 , n35828 , n35830 );
and ( n36099 , n36096 , n36098 );
and ( n36100 , n36094 , n36098 );
or ( n36101 , n36097 , n36099 , n36100 );
xor ( n36102 , n35847 , n35848 );
xor ( n36103 , n35705 , n35722 );
xor ( n36104 , n36103 , n35730 );
xor ( n36105 , n35865 , n35866 );
xor ( n36106 , n36105 , n35868 );
and ( n36107 , n36104 , n36106 );
xor ( n36108 , n35839 , n35841 );
xor ( n36109 , n36108 , n35844 );
and ( n36110 , n36106 , n36109 );
and ( n36111 , n36104 , n36109 );
or ( n36112 , n36107 , n36110 , n36111 );
and ( n36113 , n36102 , n36112 );
xor ( n36114 , n35873 , n35875 );
xor ( n36115 , n36114 , n35878 );
xor ( n36116 , n35814 , n35822 );
xor ( n36117 , n36116 , n35825 );
and ( n36118 , n36115 , n36117 );
xnor ( n36119 , n35901 , n35903 );
and ( n36120 , n36117 , n36119 );
and ( n36121 , n36115 , n36119 );
or ( n36122 , n36118 , n36120 , n36121 );
and ( n36123 , n36112 , n36122 );
and ( n36124 , n36102 , n36122 );
or ( n36125 , n36113 , n36123 , n36124 );
and ( n36126 , n36101 , n36125 );
and ( n36127 , n25959 , n24540 );
and ( n36128 , n25623 , n25284 );
and ( n36129 , n36127 , n36128 );
xor ( n36130 , n35853 , n35854 );
xor ( n36131 , n36130 , n35856 );
and ( n36132 , n36128 , n36131 );
and ( n36133 , n36127 , n36131 );
or ( n36134 , n36129 , n36132 , n36133 );
and ( n36135 , n28129 , n21666 );
and ( n36136 , n36134 , n36135 );
xor ( n36137 , n35641 , n35642 );
xor ( n36138 , n36137 , n35644 );
and ( n36139 , n36135 , n36138 );
and ( n36140 , n36134 , n36138 );
or ( n36141 , n36136 , n36139 , n36140 );
and ( n36142 , n25623 , n25617 );
and ( n36143 , n25451 , n26229 );
and ( n36144 , n36142 , n36143 );
and ( n36145 , n24993 , n26876 );
and ( n36146 , n36143 , n36145 );
and ( n36147 , n36142 , n36145 );
or ( n36148 , n36144 , n36146 , n36147 );
and ( n36149 , n26980 , n22784 );
and ( n36150 , n36148 , n36149 );
xor ( n36151 , n35964 , n35965 );
xor ( n36152 , n36151 , n35967 );
and ( n36153 , n36149 , n36152 );
and ( n36154 , n36148 , n36152 );
or ( n36155 , n36150 , n36153 , n36154 );
xor ( n36156 , n35935 , n35936 );
xor ( n36157 , n36156 , n35939 );
and ( n36158 , n36155 , n36157 );
xor ( n36159 , n35832 , n35833 );
xor ( n36160 , n36159 , n35836 );
and ( n36161 , n36157 , n36160 );
and ( n36162 , n36155 , n36160 );
or ( n36163 , n36158 , n36161 , n36162 );
and ( n36164 , n36141 , n36163 );
xor ( n36165 , n35905 , n35906 );
xor ( n36166 , n36165 , n35914 );
xor ( n36167 , n35859 , n35860 );
xor ( n36168 , n36167 , n35862 );
and ( n36169 , n36166 , n36168 );
xor ( n36170 , n35895 , n35896 );
xor ( n36171 , n36170 , n35898 );
and ( n36172 , n36168 , n36171 );
and ( n36173 , n36166 , n36171 );
or ( n36174 , n36169 , n36172 , n36173 );
and ( n36175 , n36163 , n36174 );
and ( n36176 , n36141 , n36174 );
or ( n36177 , n36164 , n36175 , n36176 );
xor ( n36178 , n35927 , n35928 );
xor ( n36179 , n36178 , n35931 );
and ( n36180 , n25220 , n26376 );
and ( n36181 , n24731 , n27246 );
and ( n36182 , n36180 , n36181 );
and ( n36183 , n24624 , n27558 );
and ( n36184 , n36181 , n36183 );
and ( n36185 , n36180 , n36183 );
or ( n36186 , n36182 , n36184 , n36185 );
and ( n36187 , n27389 , n22562 );
and ( n36188 , n36186 , n36187 );
and ( n36189 , n26933 , n22987 );
and ( n36190 , n36187 , n36189 );
and ( n36191 , n36186 , n36189 );
or ( n36192 , n36188 , n36190 , n36191 );
and ( n36193 , n36179 , n36192 );
and ( n36194 , n35718 , n33632 );
and ( n36195 , n35690 , n33630 );
nor ( n36196 , n36194 , n36195 );
xnor ( n36197 , n36196 , n28124 );
xor ( n36198 , n31463 , n33614 );
buf ( n36199 , n36198 );
buf ( n36200 , n36199 );
buf ( n36201 , n36200 );
and ( n36202 , n36201 , n28117 );
and ( n36203 , n36197 , n36202 );
xor ( n36204 , n35889 , n35890 );
xor ( n36205 , n36204 , n35892 );
and ( n36206 , n36202 , n36205 );
and ( n36207 , n36197 , n36205 );
or ( n36208 , n36203 , n36206 , n36207 );
and ( n36209 , n36192 , n36208 );
and ( n36210 , n36179 , n36208 );
or ( n36211 , n36193 , n36209 , n36210 );
xor ( n36212 , n35971 , n35972 );
xor ( n36213 , n36212 , n35974 );
buf ( n36214 , n23336 );
buf ( n36215 , n775 );
buf ( n36216 , n36215 );
buf ( n36217 , n776 );
buf ( n36218 , n36217 );
and ( n36219 , n36216 , n36218 );
not ( n36220 , n36219 );
and ( n36221 , n35605 , n36220 );
not ( n36222 , n36221 );
and ( n36223 , n36214 , n36222 );
and ( n36224 , n36213 , n36223 );
and ( n36225 , n25959 , n25026 );
and ( n36226 , n24337 , n33739 );
and ( n36227 , n36225 , n36226 );
buf ( n36228 , n12668 );
buf ( n36229 , n36228 );
and ( n36230 , n23483 , n36229 );
and ( n36231 , n36226 , n36230 );
and ( n36232 , n36225 , n36230 );
or ( n36233 , n36227 , n36231 , n36232 );
and ( n36234 , n36223 , n36233 );
and ( n36235 , n36213 , n36233 );
or ( n36236 , n36224 , n36234 , n36235 );
xor ( n36237 , n35979 , n35980 );
xor ( n36238 , n36237 , n35982 );
xor ( n36239 , n35989 , n35608 );
xor ( n36240 , n36239 , n35994 );
and ( n36241 , n36238 , n36240 );
xor ( n36242 , n36001 , n36005 );
xor ( n36243 , n36242 , n36010 );
and ( n36244 , n36240 , n36243 );
and ( n36245 , n36238 , n36243 );
or ( n36246 , n36241 , n36244 , n36245 );
and ( n36247 , n36236 , n36246 );
xor ( n36248 , n35947 , n35951 );
xor ( n36249 , n36248 , n35954 );
and ( n36250 , n36246 , n36249 );
and ( n36251 , n36236 , n36249 );
or ( n36252 , n36247 , n36250 , n36251 );
and ( n36253 , n36211 , n36252 );
xor ( n36254 , n35917 , n35919 );
xor ( n36255 , n36254 , n35922 );
and ( n36256 , n36252 , n36255 );
and ( n36257 , n36211 , n36255 );
or ( n36258 , n36253 , n36256 , n36257 );
and ( n36259 , n36177 , n36258 );
xor ( n36260 , n35852 , n35871 );
xor ( n36261 , n36260 , n35881 );
and ( n36262 , n36258 , n36261 );
and ( n36263 , n36177 , n36261 );
or ( n36264 , n36259 , n36262 , n36263 );
and ( n36265 , n36125 , n36264 );
and ( n36266 , n36101 , n36264 );
or ( n36267 , n36126 , n36265 , n36266 );
and ( n36268 , n36092 , n36267 );
xor ( n36269 , n35795 , n35796 );
xor ( n36270 , n36269 , n35807 );
xor ( n36271 , n35831 , n35849 );
xor ( n36272 , n36271 , n35884 );
and ( n36273 , n36270 , n36272 );
xor ( n36274 , n35963 , n36033 );
xor ( n36275 , n36274 , n36036 );
and ( n36276 , n36272 , n36275 );
and ( n36277 , n36270 , n36275 );
or ( n36278 , n36273 , n36276 , n36277 );
and ( n36279 , n36267 , n36278 );
and ( n36280 , n36092 , n36278 );
or ( n36281 , n36268 , n36279 , n36280 );
xor ( n36282 , n35773 , n35774 );
xor ( n36283 , n36282 , n35790 );
xor ( n36284 , n35810 , n35887 );
xor ( n36285 , n36284 , n36039 );
and ( n36286 , n36283 , n36285 );
xor ( n36287 , n36045 , n36047 );
xor ( n36288 , n36287 , n36050 );
and ( n36289 , n36285 , n36288 );
and ( n36290 , n36283 , n36288 );
or ( n36291 , n36286 , n36289 , n36290 );
and ( n36292 , n36281 , n36291 );
xor ( n36293 , n35793 , n36042 );
xor ( n36294 , n36293 , n36053 );
and ( n36295 , n36291 , n36294 );
and ( n36296 , n36281 , n36294 );
or ( n36297 , n36292 , n36295 , n36296 );
and ( n36298 , n36083 , n36297 );
xor ( n36299 , n36056 , n36066 );
xor ( n36300 , n36299 , n36069 );
and ( n36301 , n36297 , n36300 );
and ( n36302 , n36083 , n36300 );
or ( n36303 , n36298 , n36301 , n36302 );
and ( n36304 , n36081 , n36303 );
xor ( n36305 , n35768 , n35770 );
xor ( n36306 , n36305 , n36072 );
and ( n36307 , n36303 , n36306 );
and ( n36308 , n36081 , n36306 );
or ( n36309 , n36304 , n36307 , n36308 );
xor ( n36310 , n35671 , n35673 );
xor ( n36311 , n36310 , n36075 );
and ( n36312 , n36309 , n36311 );
xor ( n36313 , n36081 , n36303 );
xor ( n36314 , n36313 , n36306 );
xor ( n36315 , n36058 , n36060 );
xor ( n36316 , n36315 , n36063 );
xor ( n36317 , n35904 , n35925 );
xor ( n36318 , n36317 , n35960 );
xor ( n36319 , n36025 , n36027 );
xor ( n36320 , n36319 , n36030 );
and ( n36321 , n36318 , n36320 );
xor ( n36322 , n35934 , n35942 );
xor ( n36323 , n36322 , n35957 );
xor ( n36324 , n35988 , n36019 );
xor ( n36325 , n36324 , n36022 );
and ( n36326 , n36323 , n36325 );
xor ( n36327 , n35970 , n35977 );
xor ( n36328 , n36327 , n35985 );
xor ( n36329 , n35997 , n36013 );
xor ( n36330 , n36329 , n36016 );
and ( n36331 , n36328 , n36330 );
xor ( n36332 , n36155 , n36157 );
xor ( n36333 , n36332 , n36160 );
and ( n36334 , n36330 , n36333 );
and ( n36335 , n36328 , n36333 );
or ( n36336 , n36331 , n36334 , n36335 );
and ( n36337 , n36325 , n36336 );
and ( n36338 , n36323 , n36336 );
or ( n36339 , n36326 , n36337 , n36338 );
and ( n36340 , n36320 , n36339 );
and ( n36341 , n36318 , n36339 );
or ( n36342 , n36321 , n36340 , n36341 );
xor ( n36343 , n36186 , n36187 );
xor ( n36344 , n36343 , n36189 );
xor ( n36345 , n36148 , n36149 );
xor ( n36346 , n36345 , n36152 );
and ( n36347 , n36344 , n36346 );
and ( n36348 , n24052 , n34817 );
and ( n36349 , n23903 , n35169 );
and ( n36350 , n36348 , n36349 );
and ( n36351 , n23742 , n35544 );
and ( n36352 , n36349 , n36351 );
and ( n36353 , n36348 , n36351 );
or ( n36354 , n36350 , n36352 , n36353 );
and ( n36355 , n26399 , n24064 );
and ( n36356 , n36354 , n36355 );
and ( n36357 , n26148 , n24540 );
and ( n36358 , n36355 , n36357 );
and ( n36359 , n36354 , n36357 );
or ( n36360 , n36356 , n36358 , n36359 );
and ( n36361 , n36346 , n36360 );
and ( n36362 , n36344 , n36360 );
or ( n36363 , n36347 , n36361 , n36362 );
xor ( n36364 , n35158 , n35603 );
xor ( n36365 , n35603 , n35605 );
not ( n36366 , n36365 );
and ( n36367 , n36364 , n36366 );
and ( n36368 , n33628 , n36367 );
not ( n36369 , n36368 );
xnor ( n36370 , n36369 , n35608 );
and ( n36371 , n35690 , n34352 );
and ( n36372 , n35818 , n34350 );
nor ( n36373 , n36371 , n36372 );
xnor ( n36374 , n36373 , n28532 );
and ( n36375 , n36370 , n36374 );
xor ( n36376 , n36180 , n36181 );
xor ( n36377 , n36376 , n36183 );
and ( n36378 , n36374 , n36377 );
and ( n36379 , n36370 , n36377 );
or ( n36380 , n36375 , n36378 , n36379 );
and ( n36381 , n27962 , n22172 );
and ( n36382 , n27863 , n22337 );
xor ( n36383 , n36381 , n36382 );
and ( n36384 , n27389 , n22784 );
xor ( n36385 , n36383 , n36384 );
xor ( n36386 , n36214 , n36222 );
and ( n36387 , n36385 , n36386 );
and ( n36388 , n26678 , n24064 );
and ( n36389 , n26399 , n24540 );
and ( n36390 , n36388 , n36389 );
and ( n36391 , n25742 , n25617 );
and ( n36392 , n36389 , n36391 );
and ( n36393 , n36388 , n36391 );
or ( n36394 , n36390 , n36392 , n36393 );
and ( n36395 , n36386 , n36394 );
and ( n36396 , n36385 , n36394 );
or ( n36397 , n36387 , n36395 , n36396 );
and ( n36398 , n36380 , n36397 );
and ( n36399 , n34038 , n36367 );
and ( n36400 , n33628 , n36365 );
nor ( n36401 , n36399 , n36400 );
xnor ( n36402 , n36401 , n35608 );
and ( n36403 , n34646 , n35374 );
and ( n36404 , n34637 , n35372 );
nor ( n36405 , n36403 , n36404 );
xnor ( n36406 , n36405 , n34661 );
and ( n36407 , n36402 , n36406 );
xor ( n36408 , n31547 , n33612 );
buf ( n36409 , n36408 );
buf ( n36410 , n36409 );
buf ( n36411 , n36410 );
and ( n36412 , n36411 , n33632 );
and ( n36413 , n36201 , n33630 );
nor ( n36414 , n36412 , n36413 );
xnor ( n36415 , n36414 , n28124 );
and ( n36416 , n36406 , n36415 );
and ( n36417 , n36402 , n36415 );
or ( n36418 , n36407 , n36416 , n36417 );
and ( n36419 , n34419 , n35911 );
and ( n36420 , n34079 , n35909 );
nor ( n36421 , n36419 , n36420 );
xnor ( n36422 , n36421 , n35161 );
and ( n36423 , n36221 , n36422 );
xor ( n36424 , n31630 , n33610 );
buf ( n36425 , n36424 );
buf ( n36426 , n36425 );
buf ( n36427 , n36426 );
and ( n36428 , n36427 , n28117 );
and ( n36429 , n36422 , n36428 );
and ( n36430 , n36221 , n36428 );
or ( n36431 , n36423 , n36429 , n36430 );
and ( n36432 , n36418 , n36431 );
xor ( n36433 , n36225 , n36226 );
xor ( n36434 , n36433 , n36230 );
and ( n36435 , n36431 , n36434 );
and ( n36436 , n36418 , n36434 );
or ( n36437 , n36432 , n36435 , n36436 );
and ( n36438 , n36397 , n36437 );
and ( n36439 , n36380 , n36437 );
or ( n36440 , n36398 , n36438 , n36439 );
and ( n36441 , n36363 , n36440 );
xor ( n36442 , n36197 , n36202 );
xor ( n36443 , n36442 , n36205 );
xor ( n36444 , n36213 , n36223 );
xor ( n36445 , n36444 , n36233 );
and ( n36446 , n36443 , n36445 );
xor ( n36447 , n36238 , n36240 );
xor ( n36448 , n36447 , n36243 );
and ( n36449 , n36445 , n36448 );
and ( n36450 , n36443 , n36448 );
or ( n36451 , n36446 , n36449 , n36450 );
and ( n36452 , n36440 , n36451 );
and ( n36453 , n36363 , n36451 );
or ( n36454 , n36441 , n36452 , n36453 );
xor ( n36455 , n36166 , n36168 );
xor ( n36456 , n36455 , n36171 );
xor ( n36457 , n36179 , n36192 );
xor ( n36458 , n36457 , n36208 );
and ( n36459 , n36456 , n36458 );
xor ( n36460 , n36236 , n36246 );
xor ( n36461 , n36460 , n36249 );
and ( n36462 , n36458 , n36461 );
and ( n36463 , n36456 , n36461 );
or ( n36464 , n36459 , n36462 , n36463 );
and ( n36465 , n36454 , n36464 );
xor ( n36466 , n36104 , n36106 );
xor ( n36467 , n36466 , n36109 );
and ( n36468 , n36464 , n36467 );
and ( n36469 , n36454 , n36467 );
or ( n36470 , n36465 , n36468 , n36469 );
xor ( n36471 , n36115 , n36117 );
xor ( n36472 , n36471 , n36119 );
xor ( n36473 , n36141 , n36163 );
xor ( n36474 , n36473 , n36174 );
and ( n36475 , n36472 , n36474 );
xor ( n36476 , n36211 , n36252 );
xor ( n36477 , n36476 , n36255 );
and ( n36478 , n36474 , n36477 );
and ( n36479 , n36472 , n36477 );
or ( n36480 , n36475 , n36478 , n36479 );
and ( n36481 , n36470 , n36480 );
xor ( n36482 , n36094 , n36096 );
xor ( n36483 , n36482 , n36098 );
and ( n36484 , n36480 , n36483 );
and ( n36485 , n36470 , n36483 );
or ( n36486 , n36481 , n36484 , n36485 );
and ( n36487 , n36342 , n36486 );
xor ( n36488 , n36085 , n36087 );
xor ( n36489 , n36488 , n36089 );
and ( n36490 , n36486 , n36489 );
and ( n36491 , n36342 , n36489 );
or ( n36492 , n36487 , n36490 , n36491 );
xor ( n36493 , n36092 , n36267 );
xor ( n36494 , n36493 , n36278 );
and ( n36495 , n36492 , n36494 );
xor ( n36496 , n36283 , n36285 );
xor ( n36497 , n36496 , n36288 );
and ( n36498 , n36494 , n36497 );
and ( n36499 , n36492 , n36497 );
or ( n36500 , n36495 , n36498 , n36499 );
and ( n36501 , n36316 , n36500 );
xor ( n36502 , n36281 , n36291 );
xor ( n36503 , n36502 , n36294 );
and ( n36504 , n36500 , n36503 );
and ( n36505 , n36316 , n36503 );
or ( n36506 , n36501 , n36504 , n36505 );
xor ( n36507 , n36083 , n36297 );
xor ( n36508 , n36507 , n36300 );
and ( n36509 , n36506 , n36508 );
xor ( n36510 , n36316 , n36500 );
xor ( n36511 , n36510 , n36503 );
xor ( n36512 , n36101 , n36125 );
xor ( n36513 , n36512 , n36264 );
xor ( n36514 , n36270 , n36272 );
xor ( n36515 , n36514 , n36275 );
and ( n36516 , n36513 , n36515 );
xor ( n36517 , n36102 , n36112 );
xor ( n36518 , n36517 , n36122 );
xor ( n36519 , n36177 , n36258 );
xor ( n36520 , n36519 , n36261 );
and ( n36521 , n36518 , n36520 );
and ( n36522 , n26148 , n24064 );
and ( n36523 , n25451 , n25617 );
and ( n36524 , n36522 , n36523 );
and ( n36525 , n25220 , n26229 );
and ( n36526 , n36523 , n36525 );
and ( n36527 , n36522 , n36525 );
or ( n36528 , n36524 , n36526 , n36527 );
and ( n36529 , n24052 , n34122 );
and ( n36530 , n23903 , n34817 );
and ( n36531 , n36529 , n36530 );
and ( n36532 , n23620 , n35544 );
and ( n36533 , n36530 , n36532 );
and ( n36534 , n36529 , n36532 );
or ( n36535 , n36531 , n36533 , n36534 );
and ( n36536 , n23620 , n36229 );
buf ( n36537 , n36536 );
and ( n36538 , n24546 , n28209 );
and ( n36539 , n36537 , n36538 );
and ( n36540 , n23742 , n35169 );
and ( n36541 , n36538 , n36540 );
and ( n36542 , n36537 , n36540 );
or ( n36543 , n36539 , n36541 , n36542 );
and ( n36544 , n36535 , n36543 );
and ( n36545 , n26678 , n23508 );
and ( n36546 , n36543 , n36545 );
and ( n36547 , n36535 , n36545 );
or ( n36548 , n36544 , n36546 , n36547 );
and ( n36549 , n36528 , n36548 );
and ( n36550 , n27863 , n21990 );
and ( n36551 , n36548 , n36550 );
and ( n36552 , n36528 , n36550 );
or ( n36553 , n36549 , n36551 , n36552 );
buf ( n36554 , n23483 );
not ( n36555 , n36218 );
or ( n36556 , n36554 , n36555 );
and ( n36557 , n24337 , n34122 );
and ( n36558 , n36556 , n36557 );
not ( n36559 , n36536 );
and ( n36560 , n36557 , n36559 );
and ( n36561 , n36556 , n36559 );
or ( n36562 , n36558 , n36560 , n36561 );
and ( n36563 , n26782 , n23508 );
and ( n36564 , n36562 , n36563 );
and ( n36565 , n25742 , n25284 );
and ( n36566 , n36563 , n36565 );
and ( n36567 , n36562 , n36565 );
or ( n36568 , n36564 , n36566 , n36567 );
and ( n36569 , n27962 , n21990 );
and ( n36570 , n36568 , n36569 );
xor ( n36571 , n36522 , n36523 );
xor ( n36572 , n36571 , n36525 );
and ( n36573 , n36569 , n36572 );
and ( n36574 , n36568 , n36572 );
or ( n36575 , n36570 , n36573 , n36574 );
xor ( n36576 , n36402 , n36406 );
xor ( n36577 , n36576 , n36415 );
and ( n36578 , n34079 , n36367 );
and ( n36579 , n34038 , n36365 );
nor ( n36580 , n36578 , n36579 );
xnor ( n36581 , n36580 , n35608 );
and ( n36582 , n36201 , n34352 );
and ( n36583 , n35718 , n34350 );
nor ( n36584 , n36582 , n36583 );
xnor ( n36585 , n36584 , n28532 );
and ( n36586 , n36581 , n36585 );
and ( n36587 , n36427 , n33632 );
and ( n36588 , n36411 , n33630 );
nor ( n36589 , n36587 , n36588 );
xnor ( n36590 , n36589 , n28124 );
and ( n36591 , n36585 , n36590 );
and ( n36592 , n36581 , n36590 );
or ( n36593 , n36586 , n36591 , n36592 );
and ( n36594 , n36577 , n36593 );
and ( n36595 , n26980 , n23508 );
and ( n36596 , n26782 , n24064 );
and ( n36597 , n36595 , n36596 );
and ( n36598 , n26678 , n24540 );
and ( n36599 , n36596 , n36598 );
and ( n36600 , n36595 , n36598 );
or ( n36601 , n36597 , n36599 , n36600 );
and ( n36602 , n36593 , n36601 );
and ( n36603 , n36577 , n36601 );
or ( n36604 , n36594 , n36602 , n36603 );
xor ( n36605 , n36370 , n36374 );
xor ( n36606 , n36605 , n36377 );
and ( n36607 , n36604 , n36606 );
xor ( n36608 , n36385 , n36386 );
xor ( n36609 , n36608 , n36394 );
and ( n36610 , n36606 , n36609 );
and ( n36611 , n36604 , n36609 );
or ( n36612 , n36607 , n36610 , n36611 );
xor ( n36613 , n36344 , n36346 );
xor ( n36614 , n36613 , n36360 );
and ( n36615 , n36612 , n36614 );
xor ( n36616 , n36380 , n36397 );
xor ( n36617 , n36616 , n36437 );
and ( n36618 , n36614 , n36617 );
and ( n36619 , n36612 , n36617 );
or ( n36620 , n36615 , n36618 , n36619 );
and ( n36621 , n36575 , n36620 );
xor ( n36622 , n36328 , n36330 );
xor ( n36623 , n36622 , n36333 );
and ( n36624 , n36620 , n36623 );
and ( n36625 , n36575 , n36623 );
or ( n36626 , n36621 , n36624 , n36625 );
and ( n36627 , n36553 , n36626 );
xor ( n36628 , n36323 , n36325 );
xor ( n36629 , n36628 , n36336 );
and ( n36630 , n36626 , n36629 );
and ( n36631 , n36553 , n36629 );
or ( n36632 , n36627 , n36630 , n36631 );
and ( n36633 , n36520 , n36632 );
and ( n36634 , n36518 , n36632 );
or ( n36635 , n36521 , n36633 , n36634 );
and ( n36636 , n36515 , n36635 );
and ( n36637 , n36513 , n36635 );
or ( n36638 , n36516 , n36636 , n36637 );
xor ( n36639 , n36492 , n36494 );
xor ( n36640 , n36639 , n36497 );
and ( n36641 , n36638 , n36640 );
xor ( n36642 , n36342 , n36486 );
xor ( n36643 , n36642 , n36489 );
xor ( n36644 , n36318 , n36320 );
xor ( n36645 , n36644 , n36339 );
xor ( n36646 , n36470 , n36480 );
xor ( n36647 , n36646 , n36483 );
and ( n36648 , n36645 , n36647 );
xor ( n36649 , n36454 , n36464 );
xor ( n36650 , n36649 , n36467 );
xor ( n36651 , n36472 , n36474 );
xor ( n36652 , n36651 , n36477 );
and ( n36653 , n36650 , n36652 );
xor ( n36654 , n36528 , n36548 );
xor ( n36655 , n36654 , n36550 );
xor ( n36656 , n36134 , n36135 );
xor ( n36657 , n36656 , n36138 );
or ( n36658 , n36655 , n36657 );
and ( n36659 , n36652 , n36658 );
and ( n36660 , n36650 , n36658 );
or ( n36661 , n36653 , n36659 , n36660 );
and ( n36662 , n36647 , n36661 );
and ( n36663 , n36645 , n36661 );
or ( n36664 , n36648 , n36662 , n36663 );
and ( n36665 , n36643 , n36664 );
xor ( n36666 , n36513 , n36515 );
xor ( n36667 , n36666 , n36635 );
and ( n36668 , n36664 , n36667 );
and ( n36669 , n36643 , n36667 );
or ( n36670 , n36665 , n36668 , n36669 );
and ( n36671 , n36640 , n36670 );
and ( n36672 , n36638 , n36670 );
or ( n36673 , n36641 , n36671 , n36672 );
and ( n36674 , n36511 , n36673 );
xor ( n36675 , n36638 , n36640 );
xor ( n36676 , n36675 , n36670 );
xor ( n36677 , n36363 , n36440 );
xor ( n36678 , n36677 , n36451 );
xor ( n36679 , n36456 , n36458 );
xor ( n36680 , n36679 , n36461 );
and ( n36681 , n36678 , n36680 );
and ( n36682 , n36381 , n36382 );
and ( n36683 , n36382 , n36384 );
and ( n36684 , n36381 , n36384 );
or ( n36685 , n36682 , n36683 , n36684 );
and ( n36686 , n24052 , n35169 );
and ( n36687 , n23742 , n36229 );
and ( n36688 , n36686 , n36687 );
buf ( n36689 , n12963 );
buf ( n36690 , n36689 );
and ( n36691 , n23620 , n36690 );
and ( n36692 , n36687 , n36691 );
and ( n36693 , n36686 , n36691 );
or ( n36694 , n36688 , n36692 , n36693 );
and ( n36695 , n25623 , n26229 );
and ( n36696 , n36694 , n36695 );
and ( n36697 , n25220 , n26876 );
and ( n36698 , n36695 , n36697 );
and ( n36699 , n36694 , n36697 );
or ( n36700 , n36696 , n36698 , n36699 );
and ( n36701 , n27591 , n22562 );
and ( n36702 , n36700 , n36701 );
xor ( n36703 , n36529 , n36530 );
xor ( n36704 , n36703 , n36532 );
and ( n36705 , n36701 , n36704 );
and ( n36706 , n36700 , n36704 );
or ( n36707 , n36702 , n36705 , n36706 );
and ( n36708 , n36685 , n36707 );
xor ( n36709 , n36535 , n36543 );
xor ( n36710 , n36709 , n36545 );
and ( n36711 , n36707 , n36710 );
and ( n36712 , n36685 , n36710 );
or ( n36713 , n36708 , n36711 , n36712 );
and ( n36714 , n36680 , n36713 );
and ( n36715 , n36678 , n36713 );
or ( n36716 , n36681 , n36714 , n36715 );
and ( n36717 , n26148 , n25026 );
and ( n36718 , n25451 , n26376 );
and ( n36719 , n36717 , n36718 );
and ( n36720 , n24993 , n27246 );
and ( n36721 , n36718 , n36720 );
and ( n36722 , n36717 , n36720 );
or ( n36723 , n36719 , n36721 , n36722 );
and ( n36724 , n26980 , n22987 );
and ( n36725 , n36723 , n36724 );
and ( n36726 , n26933 , n23322 );
and ( n36727 , n36724 , n36726 );
and ( n36728 , n36723 , n36726 );
or ( n36729 , n36725 , n36727 , n36728 );
and ( n36730 , n24731 , n27558 );
and ( n36731 , n24624 , n28209 );
and ( n36732 , n36730 , n36731 );
and ( n36733 , n24546 , n33739 );
and ( n36734 , n36731 , n36733 );
and ( n36735 , n36730 , n36733 );
or ( n36736 , n36732 , n36734 , n36735 );
and ( n36737 , n26678 , n23758 );
and ( n36738 , n36736 , n36737 );
xor ( n36739 , n36537 , n36538 );
xor ( n36740 , n36739 , n36540 );
and ( n36741 , n36737 , n36740 );
and ( n36742 , n36736 , n36740 );
or ( n36743 , n36738 , n36741 , n36742 );
and ( n36744 , n36729 , n36743 );
xor ( n36745 , n36127 , n36128 );
xor ( n36746 , n36745 , n36131 );
and ( n36747 , n36743 , n36746 );
and ( n36748 , n36729 , n36746 );
or ( n36749 , n36744 , n36747 , n36748 );
and ( n36750 , n34079 , n35911 );
and ( n36751 , n34038 , n35909 );
nor ( n36752 , n36750 , n36751 );
xnor ( n36753 , n36752 , n35161 );
and ( n36754 , n34637 , n35374 );
and ( n36755 , n34419 , n35372 );
nor ( n36756 , n36754 , n36755 );
xnor ( n36757 , n36756 , n34661 );
and ( n36758 , n36753 , n36757 );
and ( n36759 , n36411 , n28117 );
and ( n36760 , n36757 , n36759 );
and ( n36761 , n36753 , n36759 );
or ( n36762 , n36758 , n36760 , n36761 );
and ( n36763 , n35386 , n34911 );
and ( n36764 , n34646 , n34909 );
nor ( n36765 , n36763 , n36764 );
xnor ( n36766 , n36765 , n34104 );
and ( n36767 , n36201 , n33632 );
and ( n36768 , n35718 , n33630 );
nor ( n36769 , n36767 , n36768 );
xnor ( n36770 , n36769 , n28124 );
and ( n36771 , n36766 , n36770 );
xor ( n36772 , n36700 , n36701 );
xor ( n36773 , n36772 , n36704 );
and ( n36774 , n36770 , n36773 );
and ( n36775 , n36766 , n36773 );
or ( n36776 , n36771 , n36774 , n36775 );
or ( n36777 , n36762 , n36776 );
and ( n36778 , n36749 , n36777 );
xor ( n36779 , n36443 , n36445 );
xor ( n36780 , n36779 , n36448 );
xor ( n36781 , n36568 , n36569 );
xor ( n36782 , n36781 , n36572 );
and ( n36783 , n36780 , n36782 );
and ( n36784 , n23903 , n36229 );
and ( n36785 , n23742 , n36690 );
and ( n36786 , n36784 , n36785 );
and ( n36787 , n24731 , n28209 );
and ( n36788 , n36786 , n36787 );
and ( n36789 , n24337 , n34817 );
and ( n36790 , n36787 , n36789 );
and ( n36791 , n36786 , n36789 );
or ( n36792 , n36788 , n36790 , n36791 );
xnor ( n36793 , n36554 , n36555 );
and ( n36794 , n24624 , n33739 );
and ( n36795 , n36793 , n36794 );
and ( n36796 , n23903 , n35544 );
and ( n36797 , n36794 , n36796 );
and ( n36798 , n36793 , n36796 );
or ( n36799 , n36795 , n36797 , n36798 );
and ( n36800 , n36792 , n36799 );
and ( n36801 , n26933 , n23508 );
and ( n36802 , n36799 , n36801 );
and ( n36803 , n36792 , n36801 );
or ( n36804 , n36800 , n36802 , n36803 );
and ( n36805 , n28129 , n21990 );
and ( n36806 , n36804 , n36805 );
xor ( n36807 , n36142 , n36143 );
xor ( n36808 , n36807 , n36145 );
and ( n36809 , n36805 , n36808 );
and ( n36810 , n36804 , n36808 );
or ( n36811 , n36806 , n36809 , n36810 );
and ( n36812 , n36782 , n36811 );
and ( n36813 , n36780 , n36811 );
or ( n36814 , n36783 , n36812 , n36813 );
and ( n36815 , n36777 , n36814 );
and ( n36816 , n36749 , n36814 );
or ( n36817 , n36778 , n36815 , n36816 );
and ( n36818 , n36716 , n36817 );
xor ( n36819 , n36553 , n36626 );
xor ( n36820 , n36819 , n36629 );
and ( n36821 , n36817 , n36820 );
and ( n36822 , n36716 , n36820 );
or ( n36823 , n36818 , n36821 , n36822 );
xor ( n36824 , n36518 , n36520 );
xor ( n36825 , n36824 , n36632 );
and ( n36826 , n36823 , n36825 );
and ( n36827 , n27962 , n22562 );
and ( n36828 , n27591 , n22987 );
and ( n36829 , n36827 , n36828 );
and ( n36830 , n27389 , n23322 );
and ( n36831 , n36828 , n36830 );
and ( n36832 , n36827 , n36830 );
or ( n36833 , n36829 , n36831 , n36832 );
and ( n36834 , n26678 , n25026 );
and ( n36835 , n24731 , n33739 );
and ( n36836 , n36834 , n36835 );
and ( n36837 , n24624 , n34122 );
and ( n36838 , n36835 , n36837 );
and ( n36839 , n36834 , n36837 );
or ( n36840 , n36836 , n36838 , n36839 );
and ( n36841 , n25742 , n26376 );
and ( n36842 , n25451 , n27246 );
and ( n36843 , n36841 , n36842 );
and ( n36844 , n25220 , n27558 );
and ( n36845 , n36842 , n36844 );
and ( n36846 , n36841 , n36844 );
or ( n36847 , n36843 , n36845 , n36846 );
and ( n36848 , n36840 , n36847 );
and ( n36849 , n26933 , n23758 );
and ( n36850 , n36847 , n36849 );
and ( n36851 , n36840 , n36849 );
or ( n36852 , n36848 , n36850 , n36851 );
and ( n36853 , n36833 , n36852 );
xor ( n36854 , n36388 , n36389 );
xor ( n36855 , n36854 , n36391 );
and ( n36856 , n36852 , n36855 );
and ( n36857 , n36833 , n36855 );
or ( n36858 , n36853 , n36856 , n36857 );
and ( n36859 , n28129 , n22337 );
and ( n36860 , n27863 , n22784 );
and ( n36861 , n36859 , n36860 );
and ( n36862 , n26399 , n25026 );
and ( n36863 , n24993 , n27558 );
xor ( n36864 , n36862 , n36863 );
and ( n36865 , n24546 , n34122 );
xor ( n36866 , n36864 , n36865 );
and ( n36867 , n36860 , n36866 );
and ( n36868 , n36859 , n36866 );
or ( n36869 , n36861 , n36867 , n36868 );
and ( n36870 , n36862 , n36863 );
and ( n36871 , n36863 , n36865 );
and ( n36872 , n36862 , n36865 );
or ( n36873 , n36870 , n36871 , n36872 );
and ( n36874 , n27389 , n22987 );
xor ( n36875 , n36873 , n36874 );
and ( n36876 , n26980 , n23322 );
xor ( n36877 , n36875 , n36876 );
and ( n36878 , n36869 , n36877 );
and ( n36879 , n26782 , n23758 );
and ( n36880 , n25959 , n25284 );
xor ( n36881 , n36879 , n36880 );
xor ( n36882 , n36348 , n36349 );
xor ( n36883 , n36882 , n36351 );
xor ( n36884 , n36881 , n36883 );
and ( n36885 , n36877 , n36884 );
and ( n36886 , n36869 , n36884 );
or ( n36887 , n36878 , n36885 , n36886 );
and ( n36888 , n36858 , n36887 );
and ( n36889 , n36873 , n36874 );
and ( n36890 , n36874 , n36876 );
and ( n36891 , n36873 , n36876 );
or ( n36892 , n36889 , n36890 , n36891 );
and ( n36893 , n36879 , n36880 );
and ( n36894 , n36880 , n36883 );
and ( n36895 , n36879 , n36883 );
or ( n36896 , n36893 , n36894 , n36895 );
xor ( n36897 , n36892 , n36896 );
xor ( n36898 , n36354 , n36355 );
xor ( n36899 , n36898 , n36357 );
xor ( n36900 , n36897 , n36899 );
and ( n36901 , n36887 , n36900 );
and ( n36902 , n36858 , n36900 );
or ( n36903 , n36888 , n36901 , n36902 );
xor ( n36904 , n36418 , n36431 );
xor ( n36905 , n36904 , n36434 );
and ( n36906 , n26148 , n25284 );
xor ( n36907 , n35605 , n36216 );
xor ( n36908 , n36216 , n36218 );
not ( n36909 , n36908 );
and ( n36910 , n36907 , n36909 );
and ( n36911 , n33628 , n36910 );
not ( n36912 , n36911 );
xnor ( n36913 , n36912 , n36221 );
and ( n36914 , n36906 , n36913 );
and ( n36915 , n35386 , n35374 );
and ( n36916 , n34646 , n35372 );
nor ( n36917 , n36915 , n36916 );
xnor ( n36918 , n36917 , n34661 );
and ( n36919 , n36913 , n36918 );
and ( n36920 , n36906 , n36918 );
or ( n36921 , n36914 , n36919 , n36920 );
xor ( n36922 , n36221 , n36422 );
xor ( n36923 , n36922 , n36428 );
and ( n36924 , n36921 , n36923 );
xor ( n36925 , n36694 , n36695 );
xor ( n36926 , n36925 , n36697 );
and ( n36927 , n36923 , n36926 );
and ( n36928 , n36921 , n36926 );
or ( n36929 , n36924 , n36927 , n36928 );
and ( n36930 , n36905 , n36929 );
and ( n36931 , n28129 , n22172 );
and ( n36932 , n27962 , n22337 );
xor ( n36933 , n36931 , n36932 );
xor ( n36934 , n36717 , n36718 );
xor ( n36935 , n36934 , n36720 );
xor ( n36936 , n36933 , n36935 );
and ( n36937 , n35690 , n34911 );
and ( n36938 , n35818 , n34909 );
nor ( n36939 , n36937 , n36938 );
xnor ( n36940 , n36939 , n34104 );
xor ( n36941 , n36827 , n36828 );
xor ( n36942 , n36941 , n36830 );
and ( n36943 , n36940 , n36942 );
and ( n36944 , n26933 , n24064 );
and ( n36945 , n26782 , n24540 );
and ( n36946 , n36944 , n36945 );
and ( n36947 , n26148 , n25617 );
and ( n36948 , n36945 , n36947 );
and ( n36949 , n36944 , n36947 );
or ( n36950 , n36946 , n36948 , n36949 );
and ( n36951 , n36942 , n36950 );
and ( n36952 , n36940 , n36950 );
or ( n36953 , n36943 , n36951 , n36952 );
and ( n36954 , n36936 , n36953 );
and ( n36955 , n27389 , n23508 );
and ( n36956 , n24993 , n28209 );
and ( n36957 , n36955 , n36956 );
and ( n36958 , n24337 , n35169 );
and ( n36959 , n36956 , n36958 );
and ( n36960 , n36955 , n36958 );
or ( n36961 , n36957 , n36959 , n36960 );
and ( n36962 , n34038 , n36910 );
and ( n36963 , n33628 , n36908 );
nor ( n36964 , n36962 , n36963 );
xnor ( n36965 , n36964 , n36221 );
and ( n36966 , n36218 , n36965 );
and ( n36967 , n35818 , n35374 );
and ( n36968 , n35386 , n35372 );
nor ( n36969 , n36967 , n36968 );
xnor ( n36970 , n36969 , n34661 );
and ( n36971 , n36965 , n36970 );
and ( n36972 , n36218 , n36970 );
or ( n36973 , n36966 , n36971 , n36972 );
and ( n36974 , n36961 , n36973 );
xor ( n36975 , n36595 , n36596 );
xor ( n36976 , n36975 , n36598 );
and ( n36977 , n36973 , n36976 );
and ( n36978 , n36961 , n36976 );
or ( n36979 , n36974 , n36977 , n36978 );
and ( n36980 , n36953 , n36979 );
and ( n36981 , n36936 , n36979 );
or ( n36982 , n36954 , n36980 , n36981 );
and ( n36983 , n36929 , n36982 );
and ( n36984 , n36905 , n36982 );
or ( n36985 , n36930 , n36983 , n36984 );
and ( n36986 , n36903 , n36985 );
xor ( n36987 , n36612 , n36614 );
xor ( n36988 , n36987 , n36617 );
and ( n36989 , n36985 , n36988 );
and ( n36990 , n36903 , n36988 );
or ( n36991 , n36986 , n36989 , n36990 );
xor ( n36992 , n36575 , n36620 );
xor ( n36993 , n36992 , n36623 );
and ( n36994 , n36991 , n36993 );
xnor ( n36995 , n36655 , n36657 );
and ( n36996 , n36993 , n36995 );
and ( n36997 , n36991 , n36995 );
or ( n36998 , n36994 , n36996 , n36997 );
and ( n36999 , n36892 , n36896 );
and ( n37000 , n36896 , n36899 );
and ( n37001 , n36892 , n36899 );
or ( n37002 , n36999 , n37000 , n37001 );
and ( n37003 , n36931 , n36932 );
and ( n37004 , n36932 , n36935 );
and ( n37005 , n36931 , n36935 );
or ( n37006 , n37003 , n37004 , n37005 );
xor ( n37007 , n36723 , n36724 );
xor ( n37008 , n37007 , n36726 );
and ( n37009 , n37006 , n37008 );
xor ( n37010 , n36736 , n36737 );
xor ( n37011 , n37010 , n36740 );
and ( n37012 , n37008 , n37011 );
and ( n37013 , n37006 , n37011 );
or ( n37014 , n37009 , n37012 , n37013 );
and ( n37015 , n37002 , n37014 );
xor ( n37016 , n36729 , n36743 );
xor ( n37017 , n37016 , n36746 );
and ( n37018 , n37014 , n37017 );
and ( n37019 , n37002 , n37017 );
or ( n37020 , n37015 , n37018 , n37019 );
and ( n37021 , n25959 , n25617 );
and ( n37022 , n25742 , n26229 );
and ( n37023 , n37021 , n37022 );
and ( n37024 , n25451 , n26876 );
and ( n37025 , n37022 , n37024 );
and ( n37026 , n37021 , n37024 );
or ( n37027 , n37023 , n37025 , n37026 );
and ( n37028 , n25623 , n26376 );
and ( n37029 , n25220 , n27246 );
and ( n37030 , n37028 , n37029 );
xor ( n37031 , n36686 , n36687 );
xor ( n37032 , n37031 , n36691 );
and ( n37033 , n37029 , n37032 );
and ( n37034 , n37028 , n37032 );
or ( n37035 , n37030 , n37033 , n37034 );
and ( n37036 , n37027 , n37035 );
and ( n37037 , n27591 , n22784 );
and ( n37038 , n37035 , n37037 );
and ( n37039 , n37027 , n37037 );
or ( n37040 , n37036 , n37038 , n37039 );
and ( n37041 , n27863 , n22562 );
xor ( n37042 , n36730 , n36731 );
xor ( n37043 , n37042 , n36733 );
and ( n37044 , n37041 , n37043 );
xor ( n37045 , n36556 , n36557 );
xor ( n37046 , n37045 , n36559 );
and ( n37047 , n37043 , n37046 );
and ( n37048 , n37041 , n37046 );
or ( n37049 , n37044 , n37047 , n37048 );
and ( n37050 , n37040 , n37049 );
xor ( n37051 , n36562 , n36563 );
xor ( n37052 , n37051 , n36565 );
and ( n37053 , n37049 , n37052 );
and ( n37054 , n37040 , n37052 );
or ( n37055 , n37050 , n37053 , n37054 );
xor ( n37056 , n36685 , n36707 );
xor ( n37057 , n37056 , n36710 );
or ( n37058 , n37055 , n37057 );
and ( n37059 , n37020 , n37058 );
xnor ( n37060 , n36762 , n36776 );
and ( n37061 , n28129 , n22562 );
and ( n37062 , n27863 , n22987 );
and ( n37063 , n37061 , n37062 );
and ( n37064 , n27591 , n23322 );
and ( n37065 , n37062 , n37064 );
and ( n37066 , n37061 , n37064 );
or ( n37067 , n37063 , n37065 , n37066 );
and ( n37068 , n26782 , n25026 );
and ( n37069 , n25451 , n27558 );
and ( n37070 , n37068 , n37069 );
and ( n37071 , n24624 , n34817 );
and ( n37072 , n37069 , n37071 );
and ( n37073 , n37068 , n37071 );
or ( n37074 , n37070 , n37072 , n37073 );
and ( n37075 , n26980 , n23758 );
and ( n37076 , n37074 , n37075 );
and ( n37077 , n26399 , n25284 );
and ( n37078 , n37075 , n37077 );
and ( n37079 , n37074 , n37077 );
or ( n37080 , n37076 , n37078 , n37079 );
and ( n37081 , n37067 , n37080 );
xor ( n37082 , n37021 , n37022 );
xor ( n37083 , n37082 , n37024 );
and ( n37084 , n37080 , n37083 );
and ( n37085 , n37067 , n37083 );
or ( n37086 , n37081 , n37084 , n37085 );
and ( n37087 , n35818 , n34911 );
and ( n37088 , n35386 , n34909 );
nor ( n37089 , n37087 , n37088 );
xnor ( n37090 , n37089 , n34104 );
and ( n37091 , n37086 , n37090 );
and ( n37092 , n35718 , n34352 );
and ( n37093 , n35690 , n34350 );
nor ( n37094 , n37092 , n37093 );
xnor ( n37095 , n37094 , n28532 );
and ( n37096 , n37090 , n37095 );
and ( n37097 , n37086 , n37095 );
or ( n37098 , n37091 , n37096 , n37097 );
xor ( n37099 , n36753 , n36757 );
xor ( n37100 , n37099 , n36759 );
and ( n37101 , n37098 , n37100 );
xor ( n37102 , n36766 , n36770 );
xor ( n37103 , n37102 , n36773 );
and ( n37104 , n37100 , n37103 );
and ( n37105 , n37098 , n37103 );
or ( n37106 , n37101 , n37104 , n37105 );
and ( n37107 , n37060 , n37106 );
xor ( n37108 , n36604 , n36606 );
xor ( n37109 , n37108 , n36609 );
xor ( n37110 , n36804 , n36805 );
xor ( n37111 , n37110 , n36808 );
and ( n37112 , n37109 , n37111 );
xor ( n37113 , n36858 , n36887 );
xor ( n37114 , n37113 , n36900 );
and ( n37115 , n37111 , n37114 );
and ( n37116 , n37109 , n37114 );
or ( n37117 , n37112 , n37115 , n37116 );
and ( n37118 , n37106 , n37117 );
and ( n37119 , n37060 , n37117 );
or ( n37120 , n37107 , n37118 , n37119 );
and ( n37121 , n37058 , n37120 );
and ( n37122 , n37020 , n37120 );
or ( n37123 , n37059 , n37121 , n37122 );
and ( n37124 , n36998 , n37123 );
xor ( n37125 , n36577 , n36593 );
xor ( n37126 , n37125 , n36601 );
xor ( n37127 , n37027 , n37035 );
xor ( n37128 , n37127 , n37037 );
and ( n37129 , n37126 , n37128 );
xor ( n37130 , n36906 , n36913 );
xor ( n37131 , n37130 , n36918 );
xor ( n37132 , n37028 , n37029 );
xor ( n37133 , n37132 , n37032 );
and ( n37134 , n37131 , n37133 );
xor ( n37135 , n36784 , n36785 );
and ( n37136 , n24546 , n34817 );
and ( n37137 , n37135 , n37136 );
and ( n37138 , n24052 , n35544 );
and ( n37139 , n37136 , n37138 );
and ( n37140 , n37135 , n37138 );
or ( n37141 , n37137 , n37139 , n37140 );
and ( n37142 , n37133 , n37141 );
and ( n37143 , n37131 , n37141 );
or ( n37144 , n37134 , n37142 , n37143 );
and ( n37145 , n37128 , n37144 );
and ( n37146 , n37126 , n37144 );
or ( n37147 , n37129 , n37145 , n37146 );
xor ( n37148 , n31726 , n33608 );
buf ( n37149 , n37148 );
buf ( n37150 , n37149 );
buf ( n37151 , n37150 );
and ( n37152 , n37151 , n33632 );
and ( n37153 , n36427 , n33630 );
nor ( n37154 , n37152 , n37153 );
xnor ( n37155 , n37154 , n28124 );
xor ( n37156 , n31807 , n33606 );
buf ( n37157 , n37156 );
buf ( n37158 , n37157 );
buf ( n37159 , n37158 );
and ( n37160 , n37159 , n28117 );
and ( n37161 , n37155 , n37160 );
xor ( n37162 , n36834 , n36835 );
xor ( n37163 , n37162 , n36837 );
and ( n37164 , n37160 , n37163 );
and ( n37165 , n37155 , n37163 );
or ( n37166 , n37161 , n37164 , n37165 );
xor ( n37167 , n37061 , n37062 );
xor ( n37168 , n37167 , n37064 );
xor ( n37169 , n36944 , n36945 );
xor ( n37170 , n37169 , n36947 );
and ( n37171 , n37168 , n37170 );
and ( n37172 , n25220 , n28209 );
and ( n37173 , n24993 , n33739 );
and ( n37174 , n37172 , n37173 );
and ( n37175 , n24337 , n35544 );
and ( n37176 , n37173 , n37175 );
and ( n37177 , n37172 , n37175 );
or ( n37178 , n37174 , n37176 , n37177 );
and ( n37179 , n37170 , n37178 );
and ( n37180 , n37168 , n37178 );
or ( n37181 , n37171 , n37179 , n37180 );
and ( n37182 , n37166 , n37181 );
and ( n37183 , n28129 , n22784 );
and ( n37184 , n24731 , n34122 );
and ( n37185 , n37183 , n37184 );
buf ( n37186 , n13411 );
buf ( n37187 , n37186 );
and ( n37188 , n23742 , n37187 );
and ( n37189 , n37184 , n37188 );
and ( n37190 , n37183 , n37188 );
or ( n37191 , n37185 , n37189 , n37190 );
buf ( n37192 , n23620 );
buf ( n37193 , n777 );
buf ( n37194 , n37193 );
xor ( n37195 , n36218 , n37194 );
not ( n37196 , n37194 );
and ( n37197 , n37195 , n37196 );
and ( n37198 , n33628 , n37197 );
not ( n37199 , n37198 );
xnor ( n37200 , n37199 , n36218 );
and ( n37201 , n37192 , n37200 );
and ( n37202 , n34079 , n36910 );
and ( n37203 , n34038 , n36908 );
nor ( n37204 , n37202 , n37203 );
xnor ( n37205 , n37204 , n36221 );
and ( n37206 , n37200 , n37205 );
and ( n37207 , n37192 , n37205 );
or ( n37208 , n37201 , n37206 , n37207 );
and ( n37209 , n37191 , n37208 );
and ( n37210 , n34637 , n36367 );
and ( n37211 , n34419 , n36365 );
nor ( n37212 , n37210 , n37211 );
xnor ( n37213 , n37212 , n35608 );
and ( n37214 , n35386 , n35911 );
and ( n37215 , n34646 , n35909 );
nor ( n37216 , n37214 , n37215 );
xnor ( n37217 , n37216 , n35161 );
and ( n37218 , n37213 , n37217 );
and ( n37219 , n36427 , n34352 );
and ( n37220 , n36411 , n34350 );
nor ( n37221 , n37219 , n37220 );
xnor ( n37222 , n37221 , n28532 );
and ( n37223 , n37217 , n37222 );
and ( n37224 , n37213 , n37222 );
or ( n37225 , n37218 , n37223 , n37224 );
and ( n37226 , n37208 , n37225 );
and ( n37227 , n37191 , n37225 );
or ( n37228 , n37209 , n37226 , n37227 );
and ( n37229 , n37181 , n37228 );
and ( n37230 , n37166 , n37228 );
or ( n37231 , n37182 , n37229 , n37230 );
xor ( n37232 , n36921 , n36923 );
xor ( n37233 , n37232 , n36926 );
and ( n37234 , n37231 , n37233 );
xor ( n37235 , n36936 , n36953 );
xor ( n37236 , n37235 , n36979 );
and ( n37237 , n37233 , n37236 );
and ( n37238 , n37231 , n37236 );
or ( n37239 , n37234 , n37237 , n37238 );
and ( n37240 , n37147 , n37239 );
xor ( n37241 , n36905 , n36929 );
xor ( n37242 , n37241 , n36982 );
and ( n37243 , n37239 , n37242 );
and ( n37244 , n37147 , n37242 );
or ( n37245 , n37240 , n37243 , n37244 );
xor ( n37246 , n36780 , n36782 );
xor ( n37247 , n37246 , n36811 );
and ( n37248 , n37245 , n37247 );
xor ( n37249 , n36903 , n36985 );
xor ( n37250 , n37249 , n36988 );
and ( n37251 , n37247 , n37250 );
and ( n37252 , n37245 , n37250 );
or ( n37253 , n37248 , n37251 , n37252 );
xor ( n37254 , n36678 , n36680 );
xor ( n37255 , n37254 , n36713 );
and ( n37256 , n37253 , n37255 );
xor ( n37257 , n36749 , n36777 );
xor ( n37258 , n37257 , n36814 );
and ( n37259 , n37255 , n37258 );
and ( n37260 , n37253 , n37258 );
or ( n37261 , n37256 , n37259 , n37260 );
and ( n37262 , n37123 , n37261 );
and ( n37263 , n36998 , n37261 );
or ( n37264 , n37124 , n37262 , n37263 );
and ( n37265 , n36825 , n37264 );
and ( n37266 , n36823 , n37264 );
or ( n37267 , n36826 , n37265 , n37266 );
xor ( n37268 , n36643 , n36664 );
xor ( n37269 , n37268 , n36667 );
and ( n37270 , n37267 , n37269 );
xor ( n37271 , n36645 , n36647 );
xor ( n37272 , n37271 , n36661 );
xor ( n37273 , n36650 , n36652 );
xor ( n37274 , n37273 , n36658 );
xor ( n37275 , n36716 , n36817 );
xor ( n37276 , n37275 , n36820 );
and ( n37277 , n37274 , n37276 );
and ( n37278 , n24546 , n35169 );
and ( n37279 , n24052 , n36229 );
and ( n37280 , n37278 , n37279 );
and ( n37281 , n23903 , n36690 );
and ( n37282 , n37279 , n37281 );
and ( n37283 , n37278 , n37281 );
or ( n37284 , n37280 , n37282 , n37283 );
and ( n37285 , n25959 , n26229 );
and ( n37286 , n37284 , n37285 );
and ( n37287 , n25623 , n26876 );
and ( n37288 , n37285 , n37287 );
and ( n37289 , n37284 , n37287 );
or ( n37290 , n37286 , n37288 , n37289 );
xor ( n37291 , n36786 , n36787 );
xor ( n37292 , n37291 , n36789 );
and ( n37293 , n37290 , n37292 );
xor ( n37294 , n36793 , n36794 );
xor ( n37295 , n37294 , n36796 );
and ( n37296 , n37292 , n37295 );
and ( n37297 , n37290 , n37295 );
or ( n37298 , n37293 , n37296 , n37297 );
xor ( n37299 , n36792 , n36799 );
xor ( n37300 , n37299 , n36801 );
and ( n37301 , n37298 , n37300 );
xor ( n37302 , n37041 , n37043 );
xor ( n37303 , n37302 , n37046 );
and ( n37304 , n37300 , n37303 );
and ( n37305 , n37298 , n37303 );
or ( n37306 , n37301 , n37304 , n37305 );
xor ( n37307 , n37040 , n37049 );
xor ( n37308 , n37307 , n37052 );
and ( n37309 , n37306 , n37308 );
xor ( n37310 , n37006 , n37008 );
xor ( n37311 , n37310 , n37011 );
and ( n37312 , n37308 , n37311 );
and ( n37313 , n37306 , n37311 );
or ( n37314 , n37309 , n37312 , n37313 );
xor ( n37315 , n37002 , n37014 );
xor ( n37316 , n37315 , n37017 );
and ( n37317 , n37314 , n37316 );
xnor ( n37318 , n37055 , n37057 );
xor ( n37319 , n37098 , n37100 );
xor ( n37320 , n37319 , n37103 );
xor ( n37321 , n37086 , n37090 );
xor ( n37322 , n37321 , n37095 );
xor ( n37323 , n37298 , n37300 );
xor ( n37324 , n37323 , n37303 );
and ( n37325 , n37322 , n37324 );
and ( n37326 , n37151 , n28117 );
xor ( n37327 , n36840 , n36847 );
xor ( n37328 , n37327 , n36849 );
and ( n37329 , n37326 , n37328 );
xor ( n37330 , n37290 , n37292 );
xor ( n37331 , n37330 , n37295 );
and ( n37332 , n37328 , n37331 );
and ( n37333 , n37326 , n37331 );
or ( n37334 , n37329 , n37332 , n37333 );
and ( n37335 , n37324 , n37334 );
and ( n37336 , n37322 , n37334 );
or ( n37337 , n37325 , n37335 , n37336 );
and ( n37338 , n37320 , n37337 );
xor ( n37339 , n36940 , n36942 );
xor ( n37340 , n37339 , n36950 );
xor ( n37341 , n36961 , n36973 );
xor ( n37342 , n37341 , n36976 );
and ( n37343 , n37340 , n37342 );
xor ( n37344 , n37067 , n37080 );
xor ( n37345 , n37344 , n37083 );
and ( n37346 , n37342 , n37345 );
and ( n37347 , n37340 , n37345 );
or ( n37348 , n37343 , n37346 , n37347 );
xor ( n37349 , n36955 , n36956 );
xor ( n37350 , n37349 , n36958 );
xor ( n37351 , n36218 , n36965 );
xor ( n37352 , n37351 , n36970 );
and ( n37353 , n37350 , n37352 );
xor ( n37354 , n37074 , n37075 );
xor ( n37355 , n37354 , n37077 );
and ( n37356 , n37352 , n37355 );
and ( n37357 , n37350 , n37355 );
or ( n37358 , n37353 , n37356 , n37357 );
xor ( n37359 , n37135 , n37136 );
xor ( n37360 , n37359 , n37138 );
and ( n37361 , n26782 , n25284 );
and ( n37362 , n26678 , n25617 );
and ( n37363 , n37361 , n37362 );
and ( n37364 , n26399 , n26229 );
and ( n37365 , n37362 , n37364 );
and ( n37366 , n37361 , n37364 );
or ( n37367 , n37363 , n37365 , n37366 );
and ( n37368 , n26399 , n25617 );
and ( n37369 , n25959 , n26376 );
xor ( n37370 , n37368 , n37369 );
and ( n37371 , n25623 , n27246 );
xor ( n37372 , n37370 , n37371 );
and ( n37373 , n37367 , n37372 );
xor ( n37374 , n37068 , n37069 );
xor ( n37375 , n37374 , n37071 );
and ( n37376 , n37372 , n37375 );
and ( n37377 , n37367 , n37375 );
or ( n37378 , n37373 , n37376 , n37377 );
and ( n37379 , n37360 , n37378 );
and ( n37380 , n37159 , n33632 );
and ( n37381 , n37151 , n33630 );
nor ( n37382 , n37380 , n37381 );
xnor ( n37383 , n37382 , n28124 );
xor ( n37384 , n31927 , n33604 );
buf ( n37385 , n37384 );
buf ( n37386 , n37385 );
buf ( n37387 , n37386 );
and ( n37388 , n37387 , n28117 );
and ( n37389 , n37383 , n37388 );
and ( n37390 , n26148 , n26376 );
and ( n37391 , n25959 , n26876 );
and ( n37392 , n37390 , n37391 );
and ( n37393 , n25742 , n27246 );
and ( n37394 , n37391 , n37393 );
and ( n37395 , n37390 , n37393 );
or ( n37396 , n37392 , n37394 , n37395 );
and ( n37397 , n37388 , n37396 );
and ( n37398 , n37383 , n37396 );
or ( n37399 , n37389 , n37397 , n37398 );
and ( n37400 , n37378 , n37399 );
and ( n37401 , n37360 , n37399 );
or ( n37402 , n37379 , n37400 , n37401 );
and ( n37403 , n37358 , n37402 );
and ( n37404 , n34038 , n37197 );
and ( n37405 , n33628 , n37194 );
nor ( n37406 , n37404 , n37405 );
xnor ( n37407 , n37406 , n36218 );
and ( n37408 , n34646 , n36367 );
and ( n37409 , n34637 , n36365 );
nor ( n37410 , n37408 , n37409 );
xnor ( n37411 , n37410 , n35608 );
and ( n37412 , n37407 , n37411 );
and ( n37413 , n35818 , n35911 );
and ( n37414 , n35386 , n35909 );
nor ( n37415 , n37413 , n37414 );
xnor ( n37416 , n37415 , n35161 );
and ( n37417 , n37411 , n37416 );
and ( n37418 , n37407 , n37416 );
or ( n37419 , n37412 , n37417 , n37418 );
and ( n37420 , n24052 , n36690 );
and ( n37421 , n23903 , n37187 );
and ( n37422 , n37420 , n37421 );
and ( n37423 , n37419 , n37422 );
and ( n37424 , n34419 , n36910 );
and ( n37425 , n34079 , n36908 );
nor ( n37426 , n37424 , n37425 );
xnor ( n37427 , n37426 , n36221 );
and ( n37428 , n37151 , n34352 );
and ( n37429 , n36427 , n34350 );
nor ( n37430 , n37428 , n37429 );
xnor ( n37431 , n37430 , n28532 );
and ( n37432 , n37427 , n37431 );
and ( n37433 , n37387 , n33632 );
and ( n37434 , n37159 , n33630 );
nor ( n37435 , n37433 , n37434 );
xnor ( n37436 , n37435 , n28124 );
and ( n37437 , n37431 , n37436 );
and ( n37438 , n37427 , n37436 );
or ( n37439 , n37432 , n37437 , n37438 );
and ( n37440 , n37422 , n37439 );
and ( n37441 , n37419 , n37439 );
or ( n37442 , n37423 , n37440 , n37441 );
xor ( n37443 , n37183 , n37184 );
xor ( n37444 , n37443 , n37188 );
xor ( n37445 , n37192 , n37200 );
xor ( n37446 , n37445 , n37205 );
and ( n37447 , n37444 , n37446 );
xor ( n37448 , n37213 , n37217 );
xor ( n37449 , n37448 , n37222 );
and ( n37450 , n37446 , n37449 );
and ( n37451 , n37444 , n37449 );
or ( n37452 , n37447 , n37450 , n37451 );
and ( n37453 , n37442 , n37452 );
xor ( n37454 , n37155 , n37160 );
xor ( n37455 , n37454 , n37163 );
and ( n37456 , n37452 , n37455 );
and ( n37457 , n37442 , n37455 );
or ( n37458 , n37453 , n37456 , n37457 );
and ( n37459 , n37402 , n37458 );
and ( n37460 , n37358 , n37458 );
or ( n37461 , n37403 , n37459 , n37460 );
and ( n37462 , n37348 , n37461 );
xor ( n37463 , n37126 , n37128 );
xor ( n37464 , n37463 , n37144 );
and ( n37465 , n37461 , n37464 );
and ( n37466 , n37348 , n37464 );
or ( n37467 , n37462 , n37465 , n37466 );
and ( n37468 , n37337 , n37467 );
and ( n37469 , n37320 , n37467 );
or ( n37470 , n37338 , n37468 , n37469 );
and ( n37471 , n37318 , n37470 );
xor ( n37472 , n37060 , n37106 );
xor ( n37473 , n37472 , n37117 );
and ( n37474 , n37470 , n37473 );
and ( n37475 , n37318 , n37473 );
or ( n37476 , n37471 , n37474 , n37475 );
and ( n37477 , n37317 , n37476 );
xor ( n37478 , n36991 , n36993 );
xor ( n37479 , n37478 , n36995 );
and ( n37480 , n37476 , n37479 );
and ( n37481 , n37317 , n37479 );
or ( n37482 , n37477 , n37480 , n37481 );
and ( n37483 , n37276 , n37482 );
and ( n37484 , n37274 , n37482 );
or ( n37485 , n37277 , n37483 , n37484 );
and ( n37486 , n37272 , n37485 );
xor ( n37487 , n36823 , n36825 );
xor ( n37488 , n37487 , n37264 );
and ( n37489 , n37485 , n37488 );
and ( n37490 , n37272 , n37488 );
or ( n37491 , n37486 , n37489 , n37490 );
and ( n37492 , n37269 , n37491 );
and ( n37493 , n37267 , n37491 );
or ( n37494 , n37270 , n37492 , n37493 );
and ( n37495 , n36676 , n37494 );
xor ( n37496 , n37267 , n37269 );
xor ( n37497 , n37496 , n37491 );
xor ( n37498 , n36998 , n37123 );
xor ( n37499 , n37498 , n37261 );
xor ( n37500 , n37020 , n37058 );
xor ( n37501 , n37500 , n37120 );
xor ( n37502 , n37253 , n37255 );
xor ( n37503 , n37502 , n37258 );
and ( n37504 , n37501 , n37503 );
xor ( n37505 , n37245 , n37247 );
xor ( n37506 , n37505 , n37250 );
xor ( n37507 , n37314 , n37316 );
and ( n37508 , n37506 , n37507 );
xor ( n37509 , n37420 , n37421 );
and ( n37510 , n24993 , n34122 );
and ( n37511 , n37509 , n37510 );
and ( n37512 , n24731 , n34817 );
and ( n37513 , n37510 , n37512 );
and ( n37514 , n37509 , n37512 );
or ( n37515 , n37511 , n37513 , n37514 );
and ( n37516 , n26980 , n24064 );
and ( n37517 , n37515 , n37516 );
and ( n37518 , n26933 , n24540 );
and ( n37519 , n37516 , n37518 );
and ( n37520 , n37515 , n37518 );
or ( n37521 , n37517 , n37519 , n37520 );
and ( n37522 , n25451 , n28209 );
and ( n37523 , n25220 , n33739 );
and ( n37524 , n37522 , n37523 );
and ( n37525 , n24546 , n35544 );
and ( n37526 , n37523 , n37525 );
and ( n37527 , n37522 , n37525 );
or ( n37528 , n37524 , n37526 , n37527 );
and ( n37529 , n26678 , n25284 );
and ( n37530 , n37528 , n37529 );
xor ( n37531 , n37278 , n37279 );
xor ( n37532 , n37531 , n37281 );
and ( n37533 , n37529 , n37532 );
and ( n37534 , n37528 , n37532 );
or ( n37535 , n37530 , n37533 , n37534 );
and ( n37536 , n37521 , n37535 );
xor ( n37537 , n36841 , n36842 );
xor ( n37538 , n37537 , n36844 );
and ( n37539 , n37535 , n37538 );
and ( n37540 , n37521 , n37538 );
or ( n37541 , n37536 , n37539 , n37540 );
and ( n37542 , n34637 , n35911 );
and ( n37543 , n34419 , n35909 );
nor ( n37544 , n37542 , n37543 );
xnor ( n37545 , n37544 , n35161 );
and ( n37546 , n37541 , n37545 );
xor ( n37547 , n36859 , n36860 );
xor ( n37548 , n37547 , n36866 );
and ( n37549 , n37545 , n37548 );
and ( n37550 , n37541 , n37548 );
or ( n37551 , n37546 , n37549 , n37550 );
xor ( n37552 , n36833 , n36852 );
xor ( n37553 , n37552 , n36855 );
and ( n37554 , n37551 , n37553 );
xor ( n37555 , n36869 , n36877 );
xor ( n37556 , n37555 , n36884 );
and ( n37557 , n37553 , n37556 );
and ( n37558 , n37551 , n37556 );
or ( n37559 , n37554 , n37557 , n37558 );
xor ( n37560 , n37306 , n37308 );
xor ( n37561 , n37560 , n37311 );
or ( n37562 , n37559 , n37561 );
and ( n37563 , n37507 , n37562 );
and ( n37564 , n37506 , n37562 );
or ( n37565 , n37508 , n37563 , n37564 );
and ( n37566 , n37503 , n37565 );
and ( n37567 , n37501 , n37565 );
or ( n37568 , n37504 , n37566 , n37567 );
and ( n37569 , n37499 , n37568 );
xor ( n37570 , n37274 , n37276 );
xor ( n37571 , n37570 , n37482 );
and ( n37572 , n37568 , n37571 );
and ( n37573 , n37499 , n37571 );
or ( n37574 , n37569 , n37572 , n37573 );
xor ( n37575 , n37272 , n37485 );
xor ( n37576 , n37575 , n37488 );
and ( n37577 , n37574 , n37576 );
xor ( n37578 , n37317 , n37476 );
xor ( n37579 , n37578 , n37479 );
xor ( n37580 , n37109 , n37111 );
xor ( n37581 , n37580 , n37114 );
xor ( n37582 , n37147 , n37239 );
xor ( n37583 , n37582 , n37242 );
and ( n37584 , n37581 , n37583 );
xor ( n37585 , n37231 , n37233 );
xor ( n37586 , n37585 , n37236 );
xor ( n37587 , n37131 , n37133 );
xor ( n37588 , n37587 , n37141 );
xor ( n37589 , n37166 , n37181 );
xor ( n37590 , n37589 , n37228 );
and ( n37591 , n37588 , n37590 );
xor ( n37592 , n37326 , n37328 );
xor ( n37593 , n37592 , n37331 );
and ( n37594 , n37590 , n37593 );
and ( n37595 , n37588 , n37593 );
or ( n37596 , n37591 , n37594 , n37595 );
and ( n37597 , n37586 , n37596 );
and ( n37598 , n37368 , n37369 );
and ( n37599 , n37369 , n37371 );
and ( n37600 , n37368 , n37371 );
or ( n37601 , n37598 , n37599 , n37600 );
and ( n37602 , n24052 , n37187 );
buf ( n37603 , n23742 );
and ( n37604 , n37602 , n37603 );
and ( n37605 , n24624 , n35169 );
and ( n37606 , n37604 , n37605 );
and ( n37607 , n24337 , n36229 );
and ( n37608 , n37605 , n37607 );
and ( n37609 , n37604 , n37607 );
or ( n37610 , n37606 , n37608 , n37609 );
and ( n37611 , n26148 , n26229 );
and ( n37612 , n37610 , n37611 );
and ( n37613 , n25742 , n26876 );
and ( n37614 , n37611 , n37613 );
and ( n37615 , n37610 , n37613 );
or ( n37616 , n37612 , n37614 , n37615 );
and ( n37617 , n37601 , n37616 );
and ( n37618 , n27962 , n22784 );
and ( n37619 , n37616 , n37618 );
and ( n37620 , n37601 , n37618 );
or ( n37621 , n37617 , n37619 , n37620 );
and ( n37622 , n24546 , n36229 );
and ( n37623 , n24337 , n36690 );
and ( n37624 , n37622 , n37623 );
buf ( n37625 , n13689 );
buf ( n37626 , n37625 );
and ( n37627 , n23903 , n37626 );
and ( n37628 , n37623 , n37627 );
and ( n37629 , n37622 , n37627 );
or ( n37630 , n37624 , n37628 , n37629 );
and ( n37631 , n26933 , n25026 );
and ( n37632 , n37630 , n37631 );
and ( n37633 , n25623 , n27558 );
and ( n37634 , n37631 , n37633 );
and ( n37635 , n37630 , n37633 );
or ( n37636 , n37632 , n37634 , n37635 );
and ( n37637 , n27591 , n23508 );
and ( n37638 , n37636 , n37637 );
and ( n37639 , n27389 , n23758 );
and ( n37640 , n37637 , n37639 );
and ( n37641 , n37636 , n37639 );
or ( n37642 , n37638 , n37640 , n37641 );
and ( n37643 , n27962 , n22987 );
and ( n37644 , n27863 , n23322 );
and ( n37645 , n37643 , n37644 );
xor ( n37646 , n37172 , n37173 );
xor ( n37647 , n37646 , n37175 );
and ( n37648 , n37644 , n37647 );
and ( n37649 , n37643 , n37647 );
or ( n37650 , n37645 , n37648 , n37649 );
and ( n37651 , n37642 , n37650 );
xor ( n37652 , n37284 , n37285 );
xor ( n37653 , n37652 , n37287 );
and ( n37654 , n37650 , n37653 );
and ( n37655 , n37642 , n37653 );
or ( n37656 , n37651 , n37654 , n37655 );
and ( n37657 , n37621 , n37656 );
xor ( n37658 , n37168 , n37170 );
xor ( n37659 , n37658 , n37178 );
xor ( n37660 , n37191 , n37208 );
xor ( n37661 , n37660 , n37225 );
and ( n37662 , n37659 , n37661 );
xor ( n37663 , n37643 , n37644 );
xor ( n37664 , n37663 , n37647 );
xor ( n37665 , n37407 , n37411 );
xor ( n37666 , n37665 , n37416 );
and ( n37667 , n26782 , n25617 );
and ( n37668 , n26678 , n26229 );
and ( n37669 , n37667 , n37668 );
and ( n37670 , n34079 , n37197 );
and ( n37671 , n34038 , n37194 );
nor ( n37672 , n37670 , n37671 );
xnor ( n37673 , n37672 , n36218 );
and ( n37674 , n37668 , n37673 );
and ( n37675 , n37667 , n37673 );
or ( n37676 , n37669 , n37674 , n37675 );
and ( n37677 , n37666 , n37676 );
and ( n37678 , n35386 , n36367 );
and ( n37679 , n34646 , n36365 );
nor ( n37680 , n37678 , n37679 );
xnor ( n37681 , n37680 , n35608 );
and ( n37682 , n35690 , n35911 );
and ( n37683 , n35818 , n35909 );
nor ( n37684 , n37682 , n37683 );
xnor ( n37685 , n37684 , n35161 );
and ( n37686 , n37681 , n37685 );
and ( n37687 , n36201 , n35374 );
and ( n37688 , n35718 , n35372 );
nor ( n37689 , n37687 , n37688 );
xnor ( n37690 , n37689 , n34661 );
and ( n37691 , n37685 , n37690 );
and ( n37692 , n37681 , n37690 );
or ( n37693 , n37686 , n37691 , n37692 );
and ( n37694 , n37676 , n37693 );
and ( n37695 , n37666 , n37693 );
or ( n37696 , n37677 , n37694 , n37695 );
and ( n37697 , n37664 , n37696 );
xor ( n37698 , n37383 , n37388 );
xor ( n37699 , n37698 , n37396 );
and ( n37700 , n37696 , n37699 );
and ( n37701 , n37664 , n37699 );
or ( n37702 , n37697 , n37700 , n37701 );
and ( n37703 , n37661 , n37702 );
and ( n37704 , n37659 , n37702 );
or ( n37705 , n37662 , n37703 , n37704 );
and ( n37706 , n37656 , n37705 );
and ( n37707 , n37621 , n37705 );
or ( n37708 , n37657 , n37706 , n37707 );
and ( n37709 , n37596 , n37708 );
and ( n37710 , n37586 , n37708 );
or ( n37711 , n37597 , n37709 , n37710 );
and ( n37712 , n37583 , n37711 );
and ( n37713 , n37581 , n37711 );
or ( n37714 , n37584 , n37712 , n37713 );
xor ( n37715 , n37318 , n37470 );
xor ( n37716 , n37715 , n37473 );
and ( n37717 , n37714 , n37716 );
xor ( n37718 , n37350 , n37352 );
xor ( n37719 , n37718 , n37355 );
xor ( n37720 , n37360 , n37378 );
xor ( n37721 , n37720 , n37399 );
and ( n37722 , n37719 , n37721 );
xor ( n37723 , n37442 , n37452 );
xor ( n37724 , n37723 , n37455 );
and ( n37725 , n37721 , n37724 );
and ( n37726 , n37719 , n37724 );
or ( n37727 , n37722 , n37725 , n37726 );
xor ( n37728 , n37340 , n37342 );
xor ( n37729 , n37728 , n37345 );
and ( n37730 , n37727 , n37729 );
xor ( n37731 , n37358 , n37402 );
xor ( n37732 , n37731 , n37458 );
and ( n37733 , n37729 , n37732 );
and ( n37734 , n37727 , n37732 );
or ( n37735 , n37730 , n37733 , n37734 );
xor ( n37736 , n37322 , n37324 );
xor ( n37737 , n37736 , n37334 );
and ( n37738 , n37735 , n37737 );
xor ( n37739 , n37348 , n37461 );
xor ( n37740 , n37739 , n37464 );
and ( n37741 , n37737 , n37740 );
and ( n37742 , n37735 , n37740 );
or ( n37743 , n37738 , n37741 , n37742 );
xor ( n37744 , n37320 , n37337 );
xor ( n37745 , n37744 , n37467 );
and ( n37746 , n37743 , n37745 );
xnor ( n37747 , n37559 , n37561 );
and ( n37748 , n37745 , n37747 );
and ( n37749 , n37743 , n37747 );
or ( n37750 , n37746 , n37748 , n37749 );
and ( n37751 , n37716 , n37750 );
and ( n37752 , n37714 , n37750 );
or ( n37753 , n37717 , n37751 , n37752 );
and ( n37754 , n37579 , n37753 );
xor ( n37755 , n37501 , n37503 );
xor ( n37756 , n37755 , n37565 );
and ( n37757 , n37753 , n37756 );
and ( n37758 , n37579 , n37756 );
or ( n37759 , n37754 , n37757 , n37758 );
xor ( n37760 , n37499 , n37568 );
xor ( n37761 , n37760 , n37571 );
and ( n37762 , n37759 , n37761 );
xor ( n37763 , n37551 , n37553 );
xor ( n37764 , n37763 , n37556 );
and ( n37765 , n34419 , n36367 );
and ( n37766 , n34079 , n36365 );
nor ( n37767 , n37765 , n37766 );
xnor ( n37768 , n37767 , n35608 );
and ( n37769 , n36411 , n34352 );
and ( n37770 , n36201 , n34350 );
nor ( n37771 , n37769 , n37770 );
xnor ( n37772 , n37771 , n28532 );
and ( n37773 , n37768 , n37772 );
xor ( n37774 , n37601 , n37616 );
xor ( n37775 , n37774 , n37618 );
and ( n37776 , n37772 , n37775 );
and ( n37777 , n37768 , n37775 );
or ( n37778 , n37773 , n37776 , n37777 );
xor ( n37779 , n36581 , n36585 );
xor ( n37780 , n37779 , n36590 );
and ( n37781 , n37778 , n37780 );
xor ( n37782 , n37541 , n37545 );
xor ( n37783 , n37782 , n37548 );
and ( n37784 , n37780 , n37783 );
and ( n37785 , n37778 , n37783 );
or ( n37786 , n37781 , n37784 , n37785 );
and ( n37787 , n37764 , n37786 );
and ( n37788 , n24337 , n37187 );
and ( n37789 , n24052 , n37626 );
and ( n37790 , n37788 , n37789 );
and ( n37791 , n25451 , n33739 );
and ( n37792 , n37790 , n37791 );
and ( n37793 , n25220 , n34122 );
and ( n37794 , n37791 , n37793 );
and ( n37795 , n37790 , n37793 );
or ( n37796 , n37792 , n37794 , n37795 );
xor ( n37797 , n37602 , n37603 );
and ( n37798 , n24993 , n34817 );
and ( n37799 , n37797 , n37798 );
and ( n37800 , n24731 , n35169 );
and ( n37801 , n37798 , n37800 );
and ( n37802 , n37797 , n37800 );
or ( n37803 , n37799 , n37801 , n37802 );
and ( n37804 , n37796 , n37803 );
and ( n37805 , n26980 , n24540 );
and ( n37806 , n37803 , n37805 );
and ( n37807 , n37796 , n37805 );
or ( n37808 , n37804 , n37806 , n37807 );
and ( n37809 , n27863 , n23508 );
and ( n37810 , n27389 , n24064 );
and ( n37811 , n37809 , n37810 );
xor ( n37812 , n37604 , n37605 );
xor ( n37813 , n37812 , n37607 );
and ( n37814 , n37810 , n37813 );
and ( n37815 , n37809 , n37813 );
or ( n37816 , n37811 , n37814 , n37815 );
and ( n37817 , n37808 , n37816 );
xor ( n37818 , n37610 , n37611 );
xor ( n37819 , n37818 , n37613 );
and ( n37820 , n37816 , n37819 );
and ( n37821 , n37808 , n37819 );
or ( n37822 , n37817 , n37820 , n37821 );
and ( n37823 , n26980 , n25026 );
and ( n37824 , n25623 , n28209 );
and ( n37825 , n37823 , n37824 );
and ( n37826 , n24624 , n35544 );
and ( n37827 , n37824 , n37826 );
and ( n37828 , n37823 , n37826 );
or ( n37829 , n37825 , n37827 , n37828 );
and ( n37830 , n26399 , n26376 );
and ( n37831 , n25959 , n27246 );
and ( n37832 , n37830 , n37831 );
and ( n37833 , n25742 , n27558 );
and ( n37834 , n37831 , n37833 );
and ( n37835 , n37830 , n37833 );
or ( n37836 , n37832 , n37834 , n37835 );
and ( n37837 , n37829 , n37836 );
and ( n37838 , n27591 , n23758 );
and ( n37839 , n37836 , n37838 );
and ( n37840 , n37829 , n37838 );
or ( n37841 , n37837 , n37839 , n37840 );
and ( n37842 , n28129 , n22987 );
and ( n37843 , n27962 , n23322 );
and ( n37844 , n37842 , n37843 );
xor ( n37845 , n37522 , n37523 );
xor ( n37846 , n37845 , n37525 );
and ( n37847 , n37843 , n37846 );
and ( n37848 , n37842 , n37846 );
or ( n37849 , n37844 , n37847 , n37848 );
and ( n37850 , n37841 , n37849 );
xor ( n37851 , n37528 , n37529 );
xor ( n37852 , n37851 , n37532 );
and ( n37853 , n37849 , n37852 );
and ( n37854 , n37841 , n37852 );
or ( n37855 , n37850 , n37853 , n37854 );
and ( n37856 , n37822 , n37855 );
and ( n37857 , n34646 , n35911 );
and ( n37858 , n34637 , n35909 );
nor ( n37859 , n37857 , n37858 );
xnor ( n37860 , n37859 , n35161 );
and ( n37861 , n37855 , n37860 );
and ( n37862 , n37822 , n37860 );
or ( n37863 , n37856 , n37861 , n37862 );
and ( n37864 , n35718 , n34911 );
and ( n37865 , n35690 , n34909 );
nor ( n37866 , n37864 , n37865 );
xnor ( n37867 , n37866 , n34104 );
xor ( n37868 , n37521 , n37535 );
xor ( n37869 , n37868 , n37538 );
or ( n37870 , n37867 , n37869 );
and ( n37871 , n37863 , n37870 );
xor ( n37872 , n37642 , n37650 );
xor ( n37873 , n37872 , n37653 );
and ( n37874 , n25623 , n33739 );
and ( n37875 , n25451 , n34122 );
and ( n37876 , n37874 , n37875 );
and ( n37877 , n24993 , n35169 );
and ( n37878 , n37875 , n37877 );
and ( n37879 , n37874 , n37877 );
or ( n37880 , n37876 , n37878 , n37879 );
and ( n37881 , n25742 , n28209 );
and ( n37882 , n25220 , n34817 );
and ( n37883 , n37881 , n37882 );
and ( n37884 , n24731 , n35544 );
and ( n37885 , n37882 , n37884 );
and ( n37886 , n37881 , n37884 );
or ( n37887 , n37883 , n37885 , n37886 );
and ( n37888 , n37880 , n37887 );
and ( n37889 , n27389 , n24540 );
and ( n37890 , n37887 , n37889 );
and ( n37891 , n37880 , n37889 );
or ( n37892 , n37888 , n37890 , n37891 );
and ( n37893 , n26933 , n25284 );
and ( n37894 , n26148 , n26876 );
and ( n37895 , n37893 , n37894 );
xor ( n37896 , n37622 , n37623 );
xor ( n37897 , n37896 , n37627 );
and ( n37898 , n37894 , n37897 );
and ( n37899 , n37893 , n37897 );
or ( n37900 , n37895 , n37898 , n37899 );
and ( n37901 , n37892 , n37900 );
xor ( n37902 , n37390 , n37391 );
xor ( n37903 , n37902 , n37393 );
and ( n37904 , n37900 , n37903 );
and ( n37905 , n37892 , n37903 );
or ( n37906 , n37901 , n37904 , n37905 );
and ( n37907 , n36201 , n34911 );
and ( n37908 , n35718 , n34909 );
nor ( n37909 , n37907 , n37908 );
xnor ( n37910 , n37909 , n34104 );
and ( n37911 , n37906 , n37910 );
xor ( n37912 , n37367 , n37372 );
xor ( n37913 , n37912 , n37375 );
and ( n37914 , n37910 , n37913 );
and ( n37915 , n37906 , n37913 );
or ( n37916 , n37911 , n37914 , n37915 );
and ( n37917 , n37873 , n37916 );
xor ( n37918 , n37419 , n37422 );
xor ( n37919 , n37918 , n37439 );
xor ( n37920 , n37444 , n37446 );
xor ( n37921 , n37920 , n37449 );
and ( n37922 , n37919 , n37921 );
xor ( n37923 , n37515 , n37516 );
xor ( n37924 , n37923 , n37518 );
and ( n37925 , n37921 , n37924 );
and ( n37926 , n37919 , n37924 );
or ( n37927 , n37922 , n37925 , n37926 );
and ( n37928 , n37916 , n37927 );
and ( n37929 , n37873 , n37927 );
or ( n37930 , n37917 , n37928 , n37929 );
and ( n37931 , n37870 , n37930 );
and ( n37932 , n37863 , n37930 );
or ( n37933 , n37871 , n37931 , n37932 );
and ( n37934 , n37786 , n37933 );
and ( n37935 , n37764 , n37933 );
or ( n37936 , n37787 , n37934 , n37935 );
xor ( n37937 , n37636 , n37637 );
xor ( n37938 , n37937 , n37639 );
xor ( n37939 , n37427 , n37431 );
xor ( n37940 , n37939 , n37436 );
xor ( n37941 , n37630 , n37631 );
xor ( n37942 , n37941 , n37633 );
and ( n37943 , n37940 , n37942 );
xor ( n37944 , n37509 , n37510 );
xor ( n37945 , n37944 , n37512 );
and ( n37946 , n37942 , n37945 );
and ( n37947 , n37940 , n37945 );
or ( n37948 , n37943 , n37946 , n37947 );
and ( n37949 , n37938 , n37948 );
and ( n37950 , n37159 , n34352 );
and ( n37951 , n37151 , n34350 );
nor ( n37952 , n37950 , n37951 );
xnor ( n37953 , n37952 , n28532 );
and ( n37954 , n27591 , n24540 );
and ( n37955 , n26980 , n25284 );
and ( n37956 , n37954 , n37955 );
and ( n37957 , n26782 , n26229 );
and ( n37958 , n37955 , n37957 );
and ( n37959 , n37954 , n37957 );
or ( n37960 , n37956 , n37958 , n37959 );
and ( n37961 , n37953 , n37960 );
and ( n37962 , n24624 , n36229 );
and ( n37963 , n24546 , n36690 );
and ( n37964 , n37962 , n37963 );
and ( n37965 , n34419 , n37197 );
and ( n37966 , n34079 , n37194 );
nor ( n37967 , n37965 , n37966 );
xnor ( n37968 , n37967 , n36218 );
and ( n37969 , n37963 , n37968 );
and ( n37970 , n37962 , n37968 );
or ( n37971 , n37964 , n37969 , n37970 );
and ( n37972 , n37960 , n37971 );
and ( n37973 , n37953 , n37971 );
or ( n37974 , n37961 , n37972 , n37973 );
and ( n37975 , n34646 , n36910 );
and ( n37976 , n34637 , n36908 );
nor ( n37977 , n37975 , n37976 );
xnor ( n37978 , n37977 , n36221 );
and ( n37979 , n35718 , n35911 );
and ( n37980 , n35690 , n35909 );
nor ( n37981 , n37979 , n37980 );
xnor ( n37982 , n37981 , n35161 );
and ( n37983 , n37978 , n37982 );
and ( n37984 , n36411 , n35374 );
and ( n37985 , n36201 , n35372 );
nor ( n37986 , n37984 , n37985 );
xnor ( n37987 , n37986 , n34661 );
and ( n37988 , n37982 , n37987 );
and ( n37989 , n37978 , n37987 );
or ( n37990 , n37983 , n37988 , n37989 );
and ( n37991 , n37151 , n34911 );
and ( n37992 , n36427 , n34909 );
nor ( n37993 , n37991 , n37992 );
xnor ( n37994 , n37993 , n34104 );
and ( n37995 , n37387 , n34352 );
and ( n37996 , n37159 , n34350 );
nor ( n37997 , n37995 , n37996 );
xnor ( n37998 , n37997 , n28532 );
and ( n37999 , n37994 , n37998 );
xor ( n38000 , n32164 , n33598 );
buf ( n38001 , n38000 );
buf ( n38002 , n38001 );
buf ( n38003 , n38002 );
and ( n38004 , n38003 , n28117 );
and ( n38005 , n37998 , n38004 );
and ( n38006 , n37994 , n38004 );
or ( n38007 , n37999 , n38005 , n38006 );
and ( n38008 , n37990 , n38007 );
xor ( n38009 , n37667 , n37668 );
xor ( n38010 , n38009 , n37673 );
and ( n38011 , n38007 , n38010 );
and ( n38012 , n37990 , n38010 );
or ( n38013 , n38008 , n38011 , n38012 );
and ( n38014 , n37974 , n38013 );
xor ( n38015 , n37666 , n37676 );
xor ( n38016 , n38015 , n37693 );
and ( n38017 , n38013 , n38016 );
and ( n38018 , n37974 , n38016 );
or ( n38019 , n38014 , n38017 , n38018 );
and ( n38020 , n37948 , n38019 );
and ( n38021 , n37938 , n38019 );
or ( n38022 , n37949 , n38020 , n38021 );
xor ( n38023 , n37659 , n37661 );
xor ( n38024 , n38023 , n37702 );
and ( n38025 , n38022 , n38024 );
xor ( n38026 , n37719 , n37721 );
xor ( n38027 , n38026 , n37724 );
and ( n38028 , n38024 , n38027 );
and ( n38029 , n38022 , n38027 );
or ( n38030 , n38025 , n38028 , n38029 );
xor ( n38031 , n37588 , n37590 );
xor ( n38032 , n38031 , n37593 );
and ( n38033 , n38030 , n38032 );
xor ( n38034 , n37621 , n37656 );
xor ( n38035 , n38034 , n37705 );
and ( n38036 , n38032 , n38035 );
and ( n38037 , n38030 , n38035 );
or ( n38038 , n38033 , n38036 , n38037 );
xor ( n38039 , n37586 , n37596 );
xor ( n38040 , n38039 , n37708 );
and ( n38041 , n38038 , n38040 );
xor ( n38042 , n37735 , n37737 );
xor ( n38043 , n38042 , n37740 );
and ( n38044 , n38040 , n38043 );
and ( n38045 , n38038 , n38043 );
or ( n38046 , n38041 , n38044 , n38045 );
and ( n38047 , n37936 , n38046 );
xor ( n38048 , n37581 , n37583 );
xor ( n38049 , n38048 , n37711 );
and ( n38050 , n38046 , n38049 );
and ( n38051 , n37936 , n38049 );
or ( n38052 , n38047 , n38050 , n38051 );
xor ( n38053 , n37506 , n37507 );
xor ( n38054 , n38053 , n37562 );
and ( n38055 , n38052 , n38054 );
xor ( n38056 , n37727 , n37729 );
xor ( n38057 , n38056 , n37732 );
xor ( n38058 , n37778 , n37780 );
xor ( n38059 , n38058 , n37783 );
and ( n38060 , n38057 , n38059 );
and ( n38061 , n26678 , n26376 );
and ( n38062 , n26148 , n27246 );
and ( n38063 , n38061 , n38062 );
and ( n38064 , n25959 , n27558 );
and ( n38065 , n38062 , n38064 );
and ( n38066 , n38061 , n38064 );
or ( n38067 , n38063 , n38065 , n38066 );
xor ( n38068 , n37788 , n37789 );
and ( n38069 , n24624 , n36690 );
and ( n38070 , n24546 , n37187 );
and ( n38071 , n38069 , n38070 );
and ( n38072 , n24337 , n37626 );
and ( n38073 , n38070 , n38072 );
and ( n38074 , n38069 , n38072 );
or ( n38075 , n38071 , n38073 , n38074 );
and ( n38076 , n38068 , n38075 );
and ( n38077 , n27389 , n25026 );
and ( n38078 , n38075 , n38077 );
and ( n38079 , n38068 , n38077 );
or ( n38080 , n38076 , n38078 , n38079 );
and ( n38081 , n38067 , n38080 );
and ( n38082 , n27863 , n23758 );
and ( n38083 , n38080 , n38082 );
and ( n38084 , n38067 , n38082 );
or ( n38085 , n38081 , n38083 , n38084 );
xor ( n38086 , n37796 , n37803 );
xor ( n38087 , n38086 , n37805 );
and ( n38088 , n38085 , n38087 );
xor ( n38089 , n37809 , n37810 );
xor ( n38090 , n38089 , n37813 );
and ( n38091 , n38087 , n38090 );
and ( n38092 , n38085 , n38090 );
or ( n38093 , n38088 , n38091 , n38092 );
and ( n38094 , n35690 , n35374 );
and ( n38095 , n35818 , n35372 );
nor ( n38096 , n38094 , n38095 );
xnor ( n38097 , n38096 , n34661 );
and ( n38098 , n38093 , n38097 );
xor ( n38099 , n37808 , n37816 );
xor ( n38100 , n38099 , n37819 );
and ( n38101 , n38097 , n38100 );
and ( n38102 , n38093 , n38100 );
or ( n38103 , n38098 , n38101 , n38102 );
xor ( n38104 , n37822 , n37855 );
xor ( n38105 , n38104 , n37860 );
and ( n38106 , n38103 , n38105 );
xor ( n38107 , n37768 , n37772 );
xor ( n38108 , n38107 , n37775 );
and ( n38109 , n38105 , n38108 );
and ( n38110 , n38103 , n38108 );
or ( n38111 , n38106 , n38109 , n38110 );
and ( n38112 , n38059 , n38111 );
and ( n38113 , n38057 , n38111 );
or ( n38114 , n38060 , n38112 , n38113 );
xnor ( n38115 , n37867 , n37869 );
and ( n38116 , n28129 , n23322 );
xor ( n38117 , n37823 , n37824 );
xor ( n38118 , n38117 , n37826 );
and ( n38119 , n38116 , n38118 );
xor ( n38120 , n37790 , n37791 );
xor ( n38121 , n38120 , n37793 );
and ( n38122 , n38118 , n38121 );
and ( n38123 , n38116 , n38121 );
or ( n38124 , n38119 , n38122 , n38123 );
and ( n38125 , n27962 , n23508 );
and ( n38126 , n27591 , n24064 );
and ( n38127 , n38125 , n38126 );
xor ( n38128 , n37797 , n37798 );
xor ( n38129 , n38128 , n37800 );
and ( n38130 , n38126 , n38129 );
and ( n38131 , n38125 , n38129 );
or ( n38132 , n38127 , n38130 , n38131 );
and ( n38133 , n38124 , n38132 );
xor ( n38134 , n37361 , n37362 );
xor ( n38135 , n38134 , n37364 );
and ( n38136 , n38132 , n38135 );
and ( n38137 , n38124 , n38135 );
or ( n38138 , n38133 , n38136 , n38137 );
xor ( n38139 , n31951 , n33602 );
buf ( n38140 , n38139 );
buf ( n38141 , n38140 );
buf ( n38142 , n38141 );
and ( n38143 , n38142 , n28117 );
xor ( n38144 , n37829 , n37836 );
xor ( n38145 , n38144 , n37838 );
and ( n38146 , n38143 , n38145 );
xor ( n38147 , n37842 , n37843 );
xor ( n38148 , n38147 , n37846 );
and ( n38149 , n38145 , n38148 );
and ( n38150 , n38143 , n38148 );
or ( n38151 , n38146 , n38149 , n38150 );
and ( n38152 , n38138 , n38151 );
xor ( n38153 , n37841 , n37849 );
xor ( n38154 , n38153 , n37852 );
and ( n38155 , n38151 , n38154 );
and ( n38156 , n38138 , n38154 );
or ( n38157 , n38152 , n38155 , n38156 );
and ( n38158 , n38115 , n38157 );
xor ( n38159 , n37664 , n37696 );
xor ( n38160 , n38159 , n37699 );
xor ( n38161 , n37906 , n37910 );
xor ( n38162 , n38161 , n37913 );
and ( n38163 , n38160 , n38162 );
xor ( n38164 , n38143 , n38145 );
xor ( n38165 , n38164 , n38148 );
xor ( n38166 , n37681 , n37685 );
xor ( n38167 , n38166 , n37690 );
xor ( n38168 , n37893 , n37894 );
xor ( n38169 , n38168 , n37897 );
and ( n38170 , n38167 , n38169 );
xor ( n38171 , n38061 , n38062 );
xor ( n38172 , n38171 , n38064 );
and ( n38173 , n25959 , n28209 );
and ( n38174 , n25742 , n33739 );
and ( n38175 , n38173 , n38174 );
and ( n38176 , n24993 , n35544 );
and ( n38177 , n38174 , n38176 );
and ( n38178 , n38173 , n38176 );
or ( n38179 , n38175 , n38177 , n38178 );
and ( n38180 , n38172 , n38179 );
and ( n38181 , n26933 , n26229 );
and ( n38182 , n26399 , n27246 );
and ( n38183 , n38181 , n38182 );
and ( n38184 , n26148 , n27558 );
and ( n38185 , n38182 , n38184 );
and ( n38186 , n38181 , n38184 );
or ( n38187 , n38183 , n38185 , n38186 );
and ( n38188 , n38179 , n38187 );
and ( n38189 , n38172 , n38187 );
or ( n38190 , n38180 , n38188 , n38189 );
and ( n38191 , n38169 , n38190 );
and ( n38192 , n38167 , n38190 );
or ( n38193 , n38170 , n38191 , n38192 );
and ( n38194 , n38165 , n38193 );
and ( n38195 , n28129 , n23758 );
and ( n38196 , n26980 , n25617 );
and ( n38197 , n38195 , n38196 );
and ( n38198 , n25623 , n34122 );
and ( n38199 , n38196 , n38198 );
and ( n38200 , n38195 , n38198 );
or ( n38201 , n38197 , n38199 , n38200 );
and ( n38202 , n25451 , n34817 );
buf ( n38203 , n13781 );
buf ( n38204 , n38203 );
and ( n38205 , n24052 , n38204 );
and ( n38206 , n38202 , n38205 );
buf ( n38207 , n23903 );
and ( n38208 , n38205 , n38207 );
and ( n38209 , n38202 , n38207 );
or ( n38210 , n38206 , n38208 , n38209 );
and ( n38211 , n38201 , n38210 );
and ( n38212 , n34637 , n37197 );
and ( n38213 , n34419 , n37194 );
nor ( n38214 , n38212 , n38213 );
xnor ( n38215 , n38214 , n36218 );
and ( n38216 , n35386 , n36910 );
and ( n38217 , n34646 , n36908 );
nor ( n38218 , n38216 , n38217 );
xnor ( n38219 , n38218 , n36221 );
and ( n38220 , n38215 , n38219 );
and ( n38221 , n35690 , n36367 );
and ( n38222 , n35818 , n36365 );
nor ( n38223 , n38221 , n38222 );
xnor ( n38224 , n38223 , n35608 );
and ( n38225 , n38219 , n38224 );
and ( n38226 , n38215 , n38224 );
or ( n38227 , n38220 , n38225 , n38226 );
and ( n38228 , n38210 , n38227 );
and ( n38229 , n38201 , n38227 );
or ( n38230 , n38211 , n38228 , n38229 );
and ( n38231 , n36201 , n35911 );
and ( n38232 , n35718 , n35909 );
nor ( n38233 , n38231 , n38232 );
xnor ( n38234 , n38233 , n35161 );
and ( n38235 , n36427 , n35374 );
and ( n38236 , n36411 , n35372 );
nor ( n38237 , n38235 , n38236 );
xnor ( n38238 , n38237 , n34661 );
and ( n38239 , n38234 , n38238 );
and ( n38240 , n37159 , n34911 );
and ( n38241 , n37151 , n34909 );
nor ( n38242 , n38240 , n38241 );
xnor ( n38243 , n38242 , n34104 );
and ( n38244 , n38238 , n38243 );
and ( n38245 , n38234 , n38243 );
or ( n38246 , n38239 , n38244 , n38245 );
xor ( n38247 , n37954 , n37955 );
xor ( n38248 , n38247 , n37957 );
and ( n38249 , n38246 , n38248 );
xor ( n38250 , n37962 , n37963 );
xor ( n38251 , n38250 , n37968 );
and ( n38252 , n38248 , n38251 );
and ( n38253 , n38246 , n38251 );
or ( n38254 , n38249 , n38252 , n38253 );
and ( n38255 , n38230 , n38254 );
xor ( n38256 , n37953 , n37960 );
xor ( n38257 , n38256 , n37971 );
and ( n38258 , n38254 , n38257 );
and ( n38259 , n38230 , n38257 );
or ( n38260 , n38255 , n38258 , n38259 );
and ( n38261 , n38193 , n38260 );
and ( n38262 , n38165 , n38260 );
or ( n38263 , n38194 , n38261 , n38262 );
and ( n38264 , n38162 , n38263 );
and ( n38265 , n38160 , n38263 );
or ( n38266 , n38163 , n38264 , n38265 );
and ( n38267 , n38157 , n38266 );
and ( n38268 , n38115 , n38266 );
or ( n38269 , n38158 , n38267 , n38268 );
xor ( n38270 , n37863 , n37870 );
xor ( n38271 , n38270 , n37930 );
and ( n38272 , n38269 , n38271 );
xor ( n38273 , n38030 , n38032 );
xor ( n38274 , n38273 , n38035 );
and ( n38275 , n38271 , n38274 );
and ( n38276 , n38269 , n38274 );
or ( n38277 , n38272 , n38275 , n38276 );
and ( n38278 , n38114 , n38277 );
xor ( n38279 , n37764 , n37786 );
xor ( n38280 , n38279 , n37933 );
and ( n38281 , n38277 , n38280 );
and ( n38282 , n38114 , n38280 );
or ( n38283 , n38278 , n38281 , n38282 );
xor ( n38284 , n37743 , n37745 );
xor ( n38285 , n38284 , n37747 );
and ( n38286 , n38283 , n38285 );
xor ( n38287 , n37936 , n38046 );
xor ( n38288 , n38287 , n38049 );
and ( n38289 , n38285 , n38288 );
and ( n38290 , n38283 , n38288 );
or ( n38291 , n38286 , n38289 , n38290 );
and ( n38292 , n38054 , n38291 );
and ( n38293 , n38052 , n38291 );
or ( n38294 , n38055 , n38292 , n38293 );
xor ( n38295 , n37579 , n37753 );
xor ( n38296 , n38295 , n37756 );
and ( n38297 , n38294 , n38296 );
xor ( n38298 , n37714 , n37716 );
xor ( n38299 , n38298 , n37750 );
xor ( n38300 , n38052 , n38054 );
xor ( n38301 , n38300 , n38291 );
and ( n38302 , n38299 , n38301 );
xor ( n38303 , n38038 , n38040 );
xor ( n38304 , n38303 , n38043 );
xor ( n38305 , n37873 , n37916 );
xor ( n38306 , n38305 , n37927 );
xor ( n38307 , n38022 , n38024 );
xor ( n38308 , n38307 , n38027 );
and ( n38309 , n38306 , n38308 );
xor ( n38310 , n38103 , n38105 );
xor ( n38311 , n38310 , n38108 );
and ( n38312 , n38308 , n38311 );
and ( n38313 , n38306 , n38311 );
or ( n38314 , n38309 , n38312 , n38313 );
xor ( n38315 , n37919 , n37921 );
xor ( n38316 , n38315 , n37924 );
xor ( n38317 , n37938 , n37948 );
xor ( n38318 , n38317 , n38019 );
and ( n38319 , n38316 , n38318 );
xor ( n38320 , n38093 , n38097 );
xor ( n38321 , n38320 , n38100 );
and ( n38322 , n38318 , n38321 );
and ( n38323 , n38316 , n38321 );
or ( n38324 , n38319 , n38322 , n38323 );
xor ( n38325 , n38138 , n38151 );
xor ( n38326 , n38325 , n38154 );
and ( n38327 , n24993 , n36229 );
and ( n38328 , n24731 , n36690 );
and ( n38329 , n38327 , n38328 );
and ( n38330 , n24546 , n37626 );
and ( n38331 , n38328 , n38330 );
and ( n38332 , n38327 , n38330 );
or ( n38333 , n38329 , n38331 , n38332 );
and ( n38334 , n27591 , n25026 );
and ( n38335 , n38333 , n38334 );
and ( n38336 , n26782 , n26376 );
and ( n38337 , n38334 , n38336 );
and ( n38338 , n38333 , n38336 );
or ( n38339 , n38335 , n38337 , n38338 );
and ( n38340 , n28129 , n23508 );
and ( n38341 , n38339 , n38340 );
and ( n38342 , n27863 , n24064 );
and ( n38343 , n38340 , n38342 );
and ( n38344 , n38339 , n38342 );
or ( n38345 , n38341 , n38343 , n38344 );
and ( n38346 , n27962 , n23758 );
xor ( n38347 , n37874 , n37875 );
xor ( n38348 , n38347 , n37877 );
and ( n38349 , n38346 , n38348 );
xor ( n38350 , n37881 , n37882 );
xor ( n38351 , n38350 , n37884 );
and ( n38352 , n38348 , n38351 );
and ( n38353 , n38346 , n38351 );
or ( n38354 , n38349 , n38352 , n38353 );
and ( n38355 , n38345 , n38354 );
xor ( n38356 , n32056 , n33600 );
buf ( n38357 , n38356 );
buf ( n38358 , n38357 );
buf ( n38359 , n38358 );
and ( n38360 , n38359 , n28117 );
and ( n38361 , n38354 , n38360 );
and ( n38362 , n38345 , n38360 );
or ( n38363 , n38355 , n38361 , n38362 );
and ( n38364 , n36411 , n34911 );
and ( n38365 , n36201 , n34909 );
nor ( n38366 , n38364 , n38365 );
xnor ( n38367 , n38366 , n34104 );
and ( n38368 , n38363 , n38367 );
xor ( n38369 , n37892 , n37900 );
xor ( n38370 , n38369 , n37903 );
and ( n38371 , n38367 , n38370 );
and ( n38372 , n38363 , n38370 );
or ( n38373 , n38368 , n38371 , n38372 );
and ( n38374 , n38326 , n38373 );
and ( n38375 , n35718 , n35374 );
and ( n38376 , n35690 , n35372 );
nor ( n38377 , n38375 , n38376 );
xnor ( n38378 , n38377 , n34661 );
xor ( n38379 , n38124 , n38132 );
xor ( n38380 , n38379 , n38135 );
and ( n38381 , n38378 , n38380 );
xor ( n38382 , n38085 , n38087 );
xor ( n38383 , n38382 , n38090 );
and ( n38384 , n38380 , n38383 );
and ( n38385 , n38378 , n38383 );
or ( n38386 , n38381 , n38384 , n38385 );
and ( n38387 , n38373 , n38386 );
and ( n38388 , n38326 , n38386 );
or ( n38389 , n38374 , n38387 , n38388 );
and ( n38390 , n38324 , n38389 );
xor ( n38391 , n37940 , n37942 );
xor ( n38392 , n38391 , n37945 );
xor ( n38393 , n37974 , n38013 );
xor ( n38394 , n38393 , n38016 );
and ( n38395 , n38392 , n38394 );
and ( n38396 , n38142 , n33632 );
and ( n38397 , n37387 , n33630 );
nor ( n38398 , n38396 , n38397 );
xnor ( n38399 , n38398 , n28124 );
xor ( n38400 , n37880 , n37887 );
xor ( n38401 , n38400 , n37889 );
and ( n38402 , n38399 , n38401 );
xor ( n38403 , n38125 , n38126 );
xor ( n38404 , n38403 , n38129 );
and ( n38405 , n38401 , n38404 );
and ( n38406 , n38399 , n38404 );
or ( n38407 , n38402 , n38405 , n38406 );
and ( n38408 , n38394 , n38407 );
and ( n38409 , n38392 , n38407 );
or ( n38410 , n38395 , n38408 , n38409 );
and ( n38411 , n24624 , n37187 );
and ( n38412 , n24337 , n38204 );
and ( n38413 , n38411 , n38412 );
and ( n38414 , n25220 , n35169 );
and ( n38415 , n38413 , n38414 );
and ( n38416 , n24731 , n36229 );
and ( n38417 , n38414 , n38416 );
and ( n38418 , n38413 , n38416 );
or ( n38419 , n38415 , n38417 , n38418 );
and ( n38420 , n26933 , n25617 );
and ( n38421 , n38419 , n38420 );
and ( n38422 , n26399 , n26876 );
and ( n38423 , n38420 , n38422 );
and ( n38424 , n38419 , n38422 );
or ( n38425 , n38421 , n38423 , n38424 );
xor ( n38426 , n37830 , n37831 );
xor ( n38427 , n38426 , n37833 );
and ( n38428 , n38425 , n38427 );
xor ( n38429 , n37990 , n38007 );
xor ( n38430 , n38429 , n38010 );
xor ( n38431 , n38067 , n38080 );
xor ( n38432 , n38431 , n38082 );
and ( n38433 , n38430 , n38432 );
xor ( n38434 , n38116 , n38118 );
xor ( n38435 , n38434 , n38121 );
and ( n38436 , n38432 , n38435 );
and ( n38437 , n38430 , n38435 );
or ( n38438 , n38433 , n38436 , n38437 );
and ( n38439 , n38428 , n38438 );
and ( n38440 , n35818 , n36367 );
and ( n38441 , n35386 , n36365 );
nor ( n38442 , n38440 , n38441 );
xnor ( n38443 , n38442 , n35608 );
and ( n38444 , n38359 , n33632 );
and ( n38445 , n38142 , n33630 );
nor ( n38446 , n38444 , n38445 );
xnor ( n38447 , n38446 , n28124 );
and ( n38448 , n38443 , n38447 );
xor ( n38449 , n38346 , n38348 );
xor ( n38450 , n38449 , n38351 );
and ( n38451 , n38447 , n38450 );
and ( n38452 , n38443 , n38450 );
or ( n38453 , n38448 , n38451 , n38452 );
xor ( n38454 , n37978 , n37982 );
xor ( n38455 , n38454 , n37987 );
xor ( n38456 , n37994 , n37998 );
xor ( n38457 , n38456 , n38004 );
and ( n38458 , n38455 , n38457 );
xor ( n38459 , n32247 , n33596 );
buf ( n38460 , n38459 );
buf ( n38461 , n38460 );
buf ( n38462 , n38461 );
and ( n38463 , n38462 , n28117 );
xor ( n38464 , n38069 , n38070 );
xor ( n38465 , n38464 , n38072 );
and ( n38466 , n38463 , n38465 );
xor ( n38467 , n38173 , n38174 );
xor ( n38468 , n38467 , n38176 );
and ( n38469 , n38465 , n38468 );
and ( n38470 , n38463 , n38468 );
or ( n38471 , n38466 , n38469 , n38470 );
and ( n38472 , n38457 , n38471 );
and ( n38473 , n38455 , n38471 );
or ( n38474 , n38458 , n38472 , n38473 );
and ( n38475 , n38453 , n38474 );
and ( n38476 , n26980 , n26229 );
and ( n38477 , n26933 , n26376 );
and ( n38478 , n38476 , n38477 );
and ( n38479 , n26678 , n27246 );
and ( n38480 , n38477 , n38479 );
and ( n38481 , n38476 , n38479 );
or ( n38482 , n38478 , n38480 , n38481 );
and ( n38483 , n36411 , n35911 );
and ( n38484 , n36201 , n35909 );
nor ( n38485 , n38483 , n38484 );
xnor ( n38486 , n38485 , n35161 );
and ( n38487 , n37151 , n35374 );
and ( n38488 , n36427 , n35372 );
nor ( n38489 , n38487 , n38488 );
xnor ( n38490 , n38489 , n34661 );
and ( n38491 , n38486 , n38490 );
and ( n38492 , n38482 , n38491 );
and ( n38493 , n28129 , n24064 );
and ( n38494 , n27962 , n24540 );
and ( n38495 , n38493 , n38494 );
and ( n38496 , n27863 , n25026 );
and ( n38497 , n38494 , n38496 );
and ( n38498 , n38493 , n38496 );
or ( n38499 , n38495 , n38497 , n38498 );
and ( n38500 , n38491 , n38499 );
and ( n38501 , n38482 , n38499 );
or ( n38502 , n38492 , n38500 , n38501 );
and ( n38503 , n26399 , n27558 );
and ( n38504 , n25451 , n35169 );
and ( n38505 , n38503 , n38504 );
and ( n38506 , n34646 , n37197 );
and ( n38507 , n34637 , n37194 );
nor ( n38508 , n38506 , n38507 );
xnor ( n38509 , n38508 , n36218 );
and ( n38510 , n38504 , n38509 );
and ( n38511 , n38503 , n38509 );
or ( n38512 , n38505 , n38510 , n38511 );
and ( n38513 , n35818 , n36910 );
and ( n38514 , n35386 , n36908 );
nor ( n38515 , n38513 , n38514 );
xnor ( n38516 , n38515 , n36221 );
and ( n38517 , n37387 , n34911 );
and ( n38518 , n37159 , n34909 );
nor ( n38519 , n38517 , n38518 );
xnor ( n38520 , n38519 , n34104 );
and ( n38521 , n38516 , n38520 );
and ( n38522 , n38359 , n34352 );
and ( n38523 , n38142 , n34350 );
nor ( n38524 , n38522 , n38523 );
xnor ( n38525 , n38524 , n28532 );
and ( n38526 , n38520 , n38525 );
and ( n38527 , n38516 , n38525 );
or ( n38528 , n38521 , n38526 , n38527 );
and ( n38529 , n38512 , n38528 );
xor ( n38530 , n38195 , n38196 );
xor ( n38531 , n38530 , n38198 );
and ( n38532 , n38528 , n38531 );
and ( n38533 , n38512 , n38531 );
or ( n38534 , n38529 , n38532 , n38533 );
and ( n38535 , n38502 , n38534 );
xor ( n38536 , n38202 , n38205 );
xor ( n38537 , n38536 , n38207 );
xor ( n38538 , n38215 , n38219 );
xor ( n38539 , n38538 , n38224 );
and ( n38540 , n38537 , n38539 );
xor ( n38541 , n38234 , n38238 );
xor ( n38542 , n38541 , n38243 );
and ( n38543 , n38539 , n38542 );
and ( n38544 , n38537 , n38542 );
or ( n38545 , n38540 , n38543 , n38544 );
and ( n38546 , n38534 , n38545 );
and ( n38547 , n38502 , n38545 );
or ( n38548 , n38535 , n38546 , n38547 );
and ( n38549 , n38474 , n38548 );
and ( n38550 , n38453 , n38548 );
or ( n38551 , n38475 , n38549 , n38550 );
and ( n38552 , n38438 , n38551 );
and ( n38553 , n38428 , n38551 );
or ( n38554 , n38439 , n38552 , n38553 );
and ( n38555 , n38410 , n38554 );
xor ( n38556 , n38160 , n38162 );
xor ( n38557 , n38556 , n38263 );
and ( n38558 , n38554 , n38557 );
and ( n38559 , n38410 , n38557 );
or ( n38560 , n38555 , n38558 , n38559 );
and ( n38561 , n38389 , n38560 );
and ( n38562 , n38324 , n38560 );
or ( n38563 , n38390 , n38561 , n38562 );
and ( n38564 , n38314 , n38563 );
xor ( n38565 , n38057 , n38059 );
xor ( n38566 , n38565 , n38111 );
and ( n38567 , n38563 , n38566 );
and ( n38568 , n38314 , n38566 );
or ( n38569 , n38564 , n38567 , n38568 );
and ( n38570 , n38304 , n38569 );
xor ( n38571 , n38114 , n38277 );
xor ( n38572 , n38571 , n38280 );
and ( n38573 , n38569 , n38572 );
and ( n38574 , n38304 , n38572 );
or ( n38575 , n38570 , n38573 , n38574 );
xor ( n38576 , n38283 , n38285 );
xor ( n38577 , n38576 , n38288 );
and ( n38578 , n38575 , n38577 );
xor ( n38579 , n38269 , n38271 );
xor ( n38580 , n38579 , n38274 );
xor ( n38581 , n38115 , n38157 );
xor ( n38582 , n38581 , n38266 );
xor ( n38583 , n38172 , n38179 );
xor ( n38584 , n38583 , n38187 );
xor ( n38585 , n38201 , n38210 );
xor ( n38586 , n38585 , n38227 );
and ( n38587 , n38584 , n38586 );
xor ( n38588 , n38246 , n38248 );
xor ( n38589 , n38588 , n38251 );
and ( n38590 , n38586 , n38589 );
and ( n38591 , n38584 , n38589 );
or ( n38592 , n38587 , n38590 , n38591 );
xor ( n38593 , n38167 , n38169 );
xor ( n38594 , n38593 , n38190 );
and ( n38595 , n38592 , n38594 );
xor ( n38596 , n38230 , n38254 );
xor ( n38597 , n38596 , n38257 );
and ( n38598 , n38594 , n38597 );
and ( n38599 , n38592 , n38597 );
or ( n38600 , n38595 , n38598 , n38599 );
xor ( n38601 , n38165 , n38193 );
xor ( n38602 , n38601 , n38260 );
and ( n38603 , n38600 , n38602 );
xor ( n38604 , n38363 , n38367 );
xor ( n38605 , n38604 , n38370 );
and ( n38606 , n38602 , n38605 );
and ( n38607 , n38600 , n38605 );
or ( n38608 , n38603 , n38606 , n38607 );
xor ( n38609 , n38378 , n38380 );
xor ( n38610 , n38609 , n38383 );
and ( n38611 , n25959 , n33739 );
and ( n38612 , n25742 , n34122 );
and ( n38613 , n38611 , n38612 );
and ( n38614 , n25623 , n34817 );
and ( n38615 , n38612 , n38614 );
and ( n38616 , n38611 , n38614 );
or ( n38617 , n38613 , n38615 , n38616 );
and ( n38618 , n27389 , n25284 );
and ( n38619 , n38617 , n38618 );
and ( n38620 , n26678 , n26876 );
and ( n38621 , n38618 , n38620 );
and ( n38622 , n38617 , n38620 );
or ( n38623 , n38619 , n38621 , n38622 );
and ( n38624 , n27962 , n24064 );
and ( n38625 , n27863 , n24540 );
and ( n38626 , n38624 , n38625 );
xor ( n38627 , n38413 , n38414 );
xor ( n38628 , n38627 , n38416 );
and ( n38629 , n38625 , n38628 );
and ( n38630 , n38624 , n38628 );
or ( n38631 , n38626 , n38629 , n38630 );
and ( n38632 , n38623 , n38631 );
xor ( n38633 , n38068 , n38075 );
xor ( n38634 , n38633 , n38077 );
and ( n38635 , n38631 , n38634 );
and ( n38636 , n38623 , n38634 );
or ( n38637 , n38632 , n38635 , n38636 );
and ( n38638 , n34637 , n36910 );
and ( n38639 , n34419 , n36908 );
nor ( n38640 , n38638 , n38639 );
xnor ( n38641 , n38640 , n36221 );
and ( n38642 , n38637 , n38641 );
and ( n38643 , n36427 , n34911 );
and ( n38644 , n36411 , n34909 );
nor ( n38645 , n38643 , n38644 );
xnor ( n38646 , n38645 , n34104 );
and ( n38647 , n38641 , n38646 );
and ( n38648 , n38637 , n38646 );
or ( n38649 , n38642 , n38647 , n38648 );
and ( n38650 , n38610 , n38649 );
xor ( n38651 , n38345 , n38354 );
xor ( n38652 , n38651 , n38360 );
xor ( n38653 , n38399 , n38401 );
xor ( n38654 , n38653 , n38404 );
or ( n38655 , n38652 , n38654 );
and ( n38656 , n38649 , n38655 );
and ( n38657 , n38610 , n38655 );
or ( n38658 , n38650 , n38656 , n38657 );
and ( n38659 , n38608 , n38658 );
xor ( n38660 , n38425 , n38427 );
xor ( n38661 , n38339 , n38340 );
xor ( n38662 , n38661 , n38342 );
xor ( n38663 , n38419 , n38420 );
xor ( n38664 , n38663 , n38422 );
and ( n38665 , n38662 , n38664 );
xor ( n38666 , n38443 , n38447 );
xor ( n38667 , n38666 , n38450 );
and ( n38668 , n38664 , n38667 );
and ( n38669 , n38662 , n38667 );
or ( n38670 , n38665 , n38668 , n38669 );
and ( n38671 , n38660 , n38670 );
and ( n38672 , n27389 , n25617 );
and ( n38673 , n26782 , n26876 );
and ( n38674 , n38672 , n38673 );
xor ( n38675 , n38327 , n38328 );
xor ( n38676 , n38675 , n38330 );
and ( n38677 , n38673 , n38676 );
and ( n38678 , n38672 , n38676 );
or ( n38679 , n38674 , n38677 , n38678 );
xor ( n38680 , n38181 , n38182 );
xor ( n38681 , n38680 , n38184 );
and ( n38682 , n38679 , n38681 );
xor ( n38683 , n38333 , n38334 );
xor ( n38684 , n38683 , n38336 );
and ( n38685 , n38681 , n38684 );
and ( n38686 , n38679 , n38684 );
or ( n38687 , n38682 , n38685 , n38686 );
xor ( n38688 , n38617 , n38618 );
xor ( n38689 , n38688 , n38620 );
and ( n38690 , n24731 , n37187 );
and ( n38691 , n24624 , n37626 );
and ( n38692 , n38690 , n38691 );
and ( n38693 , n24546 , n38204 );
and ( n38694 , n38691 , n38693 );
and ( n38695 , n38690 , n38693 );
or ( n38696 , n38692 , n38694 , n38695 );
and ( n38697 , n26148 , n28209 );
and ( n38698 , n38696 , n38697 );
and ( n38699 , n25220 , n35544 );
and ( n38700 , n38697 , n38699 );
and ( n38701 , n38696 , n38699 );
or ( n38702 , n38698 , n38700 , n38701 );
and ( n38703 , n38689 , n38702 );
xor ( n38704 , n38611 , n38612 );
xor ( n38705 , n38704 , n38614 );
xor ( n38706 , n38476 , n38477 );
xor ( n38707 , n38706 , n38479 );
and ( n38708 , n38705 , n38707 );
xor ( n38709 , n38411 , n38412 );
and ( n38710 , n38707 , n38709 );
and ( n38711 , n38705 , n38709 );
or ( n38712 , n38708 , n38710 , n38711 );
and ( n38713 , n38702 , n38712 );
and ( n38714 , n38689 , n38712 );
or ( n38715 , n38703 , n38713 , n38714 );
and ( n38716 , n38687 , n38715 );
xor ( n38717 , n38486 , n38490 );
and ( n38718 , n27591 , n25617 );
and ( n38719 , n27389 , n26229 );
and ( n38720 , n38718 , n38719 );
and ( n38721 , n26933 , n26876 );
and ( n38722 , n38719 , n38721 );
and ( n38723 , n38718 , n38721 );
or ( n38724 , n38720 , n38722 , n38723 );
and ( n38725 , n38717 , n38724 );
and ( n38726 , n26782 , n27246 );
and ( n38727 , n25220 , n36229 );
and ( n38728 , n38726 , n38727 );
and ( n38729 , n24993 , n36690 );
and ( n38730 , n38727 , n38729 );
and ( n38731 , n38726 , n38729 );
or ( n38732 , n38728 , n38730 , n38731 );
and ( n38733 , n38724 , n38732 );
and ( n38734 , n38717 , n38732 );
or ( n38735 , n38725 , n38733 , n38734 );
buf ( n38736 , n14265 );
buf ( n38737 , n38736 );
and ( n38738 , n24337 , n38737 );
buf ( n38739 , n24052 );
and ( n38740 , n38738 , n38739 );
and ( n38741 , n35386 , n37197 );
and ( n38742 , n34646 , n37194 );
nor ( n38743 , n38741 , n38742 );
xnor ( n38744 , n38743 , n36218 );
and ( n38745 , n38739 , n38744 );
and ( n38746 , n38738 , n38744 );
or ( n38747 , n38740 , n38745 , n38746 );
and ( n38748 , n35690 , n36910 );
and ( n38749 , n35818 , n36908 );
nor ( n38750 , n38748 , n38749 );
xnor ( n38751 , n38750 , n36221 );
and ( n38752 , n36201 , n36367 );
and ( n38753 , n35718 , n36365 );
nor ( n38754 , n38752 , n38753 );
xnor ( n38755 , n38754 , n35608 );
and ( n38756 , n38751 , n38755 );
and ( n38757 , n36427 , n35911 );
and ( n38758 , n36411 , n35909 );
nor ( n38759 , n38757 , n38758 );
xnor ( n38760 , n38759 , n35161 );
and ( n38761 , n38755 , n38760 );
and ( n38762 , n38751 , n38760 );
or ( n38763 , n38756 , n38761 , n38762 );
and ( n38764 , n38747 , n38763 );
and ( n38765 , n37159 , n35374 );
and ( n38766 , n37151 , n35372 );
nor ( n38767 , n38765 , n38766 );
xnor ( n38768 , n38767 , n34661 );
and ( n38769 , n38142 , n34911 );
and ( n38770 , n37387 , n34909 );
nor ( n38771 , n38769 , n38770 );
xnor ( n38772 , n38771 , n34104 );
and ( n38773 , n38768 , n38772 );
xor ( n38774 , n32330 , n33594 );
buf ( n38775 , n38774 );
buf ( n38776 , n38775 );
buf ( n38777 , n38776 );
and ( n38778 , n38777 , n33632 );
and ( n38779 , n38462 , n33630 );
nor ( n38780 , n38778 , n38779 );
xnor ( n38781 , n38780 , n28124 );
and ( n38782 , n38772 , n38781 );
and ( n38783 , n38768 , n38781 );
or ( n38784 , n38773 , n38782 , n38783 );
and ( n38785 , n38763 , n38784 );
and ( n38786 , n38747 , n38784 );
or ( n38787 , n38764 , n38785 , n38786 );
and ( n38788 , n38735 , n38787 );
xor ( n38789 , n38493 , n38494 );
xor ( n38790 , n38789 , n38496 );
xor ( n38791 , n38503 , n38504 );
xor ( n38792 , n38791 , n38509 );
and ( n38793 , n38790 , n38792 );
xor ( n38794 , n38516 , n38520 );
xor ( n38795 , n38794 , n38525 );
and ( n38796 , n38792 , n38795 );
and ( n38797 , n38790 , n38795 );
or ( n38798 , n38793 , n38796 , n38797 );
and ( n38799 , n38787 , n38798 );
and ( n38800 , n38735 , n38798 );
or ( n38801 , n38788 , n38799 , n38800 );
and ( n38802 , n38715 , n38801 );
and ( n38803 , n38687 , n38801 );
or ( n38804 , n38716 , n38802 , n38803 );
and ( n38805 , n38670 , n38804 );
and ( n38806 , n38660 , n38804 );
or ( n38807 , n38671 , n38805 , n38806 );
xor ( n38808 , n38463 , n38465 );
xor ( n38809 , n38808 , n38468 );
xor ( n38810 , n38482 , n38491 );
xor ( n38811 , n38810 , n38499 );
and ( n38812 , n38809 , n38811 );
xor ( n38813 , n38512 , n38528 );
xor ( n38814 , n38813 , n38531 );
and ( n38815 , n38811 , n38814 );
and ( n38816 , n38809 , n38814 );
or ( n38817 , n38812 , n38815 , n38816 );
xor ( n38818 , n38455 , n38457 );
xor ( n38819 , n38818 , n38471 );
and ( n38820 , n38817 , n38819 );
xor ( n38821 , n38502 , n38534 );
xor ( n38822 , n38821 , n38545 );
and ( n38823 , n38819 , n38822 );
and ( n38824 , n38817 , n38822 );
or ( n38825 , n38820 , n38823 , n38824 );
xor ( n38826 , n38430 , n38432 );
xor ( n38827 , n38826 , n38435 );
and ( n38828 , n38825 , n38827 );
xor ( n38829 , n38453 , n38474 );
xor ( n38830 , n38829 , n38548 );
and ( n38831 , n38827 , n38830 );
and ( n38832 , n38825 , n38830 );
or ( n38833 , n38828 , n38831 , n38832 );
and ( n38834 , n38807 , n38833 );
xor ( n38835 , n38392 , n38394 );
xor ( n38836 , n38835 , n38407 );
and ( n38837 , n38833 , n38836 );
and ( n38838 , n38807 , n38836 );
or ( n38839 , n38834 , n38837 , n38838 );
and ( n38840 , n38658 , n38839 );
and ( n38841 , n38608 , n38839 );
or ( n38842 , n38659 , n38840 , n38841 );
and ( n38843 , n38582 , n38842 );
xor ( n38844 , n38316 , n38318 );
xor ( n38845 , n38844 , n38321 );
xor ( n38846 , n38326 , n38373 );
xor ( n38847 , n38846 , n38386 );
and ( n38848 , n38845 , n38847 );
xor ( n38849 , n38410 , n38554 );
xor ( n38850 , n38849 , n38557 );
and ( n38851 , n38847 , n38850 );
and ( n38852 , n38845 , n38850 );
or ( n38853 , n38848 , n38851 , n38852 );
and ( n38854 , n38842 , n38853 );
and ( n38855 , n38582 , n38853 );
or ( n38856 , n38843 , n38854 , n38855 );
and ( n38857 , n38580 , n38856 );
xor ( n38858 , n38314 , n38563 );
xor ( n38859 , n38858 , n38566 );
and ( n38860 , n38856 , n38859 );
and ( n38861 , n38580 , n38859 );
or ( n38862 , n38857 , n38860 , n38861 );
xor ( n38863 , n38304 , n38569 );
xor ( n38864 , n38863 , n38572 );
and ( n38865 , n38862 , n38864 );
xor ( n38866 , n38306 , n38308 );
xor ( n38867 , n38866 , n38311 );
xor ( n38868 , n38324 , n38389 );
xor ( n38869 , n38868 , n38560 );
and ( n38870 , n38867 , n38869 );
xor ( n38871 , n38428 , n38438 );
xor ( n38872 , n38871 , n38551 );
xor ( n38873 , n38592 , n38594 );
xor ( n38874 , n38873 , n38597 );
xor ( n38875 , n38637 , n38641 );
xor ( n38876 , n38875 , n38646 );
and ( n38877 , n38874 , n38876 );
xnor ( n38878 , n38652 , n38654 );
and ( n38879 , n38876 , n38878 );
and ( n38880 , n38874 , n38878 );
or ( n38881 , n38877 , n38879 , n38880 );
and ( n38882 , n38872 , n38881 );
xor ( n38883 , n38584 , n38586 );
xor ( n38884 , n38883 , n38589 );
xor ( n38885 , n38623 , n38631 );
xor ( n38886 , n38885 , n38634 );
and ( n38887 , n38884 , n38886 );
and ( n38888 , n25220 , n36690 );
and ( n38889 , n24993 , n37187 );
and ( n38890 , n38888 , n38889 );
and ( n38891 , n24731 , n37626 );
and ( n38892 , n38889 , n38891 );
and ( n38893 , n38888 , n38891 );
or ( n38894 , n38890 , n38892 , n38893 );
and ( n38895 , n26980 , n26376 );
and ( n38896 , n38894 , n38895 );
and ( n38897 , n26399 , n28209 );
and ( n38898 , n38895 , n38897 );
and ( n38899 , n38894 , n38897 );
or ( n38900 , n38896 , n38898 , n38899 );
and ( n38901 , n27962 , n25026 );
and ( n38902 , n26678 , n27558 );
and ( n38903 , n38901 , n38902 );
xor ( n38904 , n38690 , n38691 );
xor ( n38905 , n38904 , n38693 );
and ( n38906 , n38902 , n38905 );
and ( n38907 , n38901 , n38905 );
or ( n38908 , n38903 , n38906 , n38907 );
and ( n38909 , n38900 , n38908 );
xor ( n38910 , n38696 , n38697 );
xor ( n38911 , n38910 , n38699 );
and ( n38912 , n38908 , n38911 );
and ( n38913 , n38900 , n38911 );
or ( n38914 , n38909 , n38912 , n38913 );
and ( n38915 , n38142 , n34352 );
and ( n38916 , n37387 , n34350 );
nor ( n38917 , n38915 , n38916 );
xnor ( n38918 , n38917 , n28532 );
and ( n38919 , n38914 , n38918 );
and ( n38920 , n38003 , n33632 );
and ( n38921 , n38359 , n33630 );
nor ( n38922 , n38920 , n38921 );
xnor ( n38923 , n38922 , n28124 );
and ( n38924 , n38918 , n38923 );
and ( n38925 , n38914 , n38923 );
or ( n38926 , n38919 , n38924 , n38925 );
and ( n38927 , n38886 , n38926 );
and ( n38928 , n38884 , n38926 );
or ( n38929 , n38887 , n38927 , n38928 );
xor ( n38930 , n38537 , n38539 );
xor ( n38931 , n38930 , n38542 );
xor ( n38932 , n38624 , n38625 );
xor ( n38933 , n38932 , n38628 );
and ( n38934 , n38931 , n38933 );
xor ( n38935 , n38679 , n38681 );
xor ( n38936 , n38935 , n38684 );
and ( n38937 , n38933 , n38936 );
and ( n38938 , n38931 , n38936 );
or ( n38939 , n38934 , n38937 , n38938 );
and ( n38940 , n26148 , n33739 );
and ( n38941 , n25959 , n34122 );
and ( n38942 , n38940 , n38941 );
and ( n38943 , n25742 , n34817 );
and ( n38944 , n38941 , n38943 );
and ( n38945 , n38940 , n38943 );
or ( n38946 , n38942 , n38944 , n38945 );
and ( n38947 , n24624 , n38204 );
and ( n38948 , n24546 , n38737 );
and ( n38949 , n38947 , n38948 );
and ( n38950 , n25623 , n35169 );
and ( n38951 , n38949 , n38950 );
and ( n38952 , n25451 , n35544 );
and ( n38953 , n38950 , n38952 );
and ( n38954 , n38949 , n38952 );
or ( n38955 , n38951 , n38953 , n38954 );
and ( n38956 , n38946 , n38955 );
and ( n38957 , n27591 , n25284 );
and ( n38958 , n38955 , n38957 );
and ( n38959 , n38946 , n38957 );
or ( n38960 , n38956 , n38958 , n38959 );
and ( n38961 , n38777 , n28117 );
xor ( n38962 , n38672 , n38673 );
xor ( n38963 , n38962 , n38676 );
or ( n38964 , n38961 , n38963 );
and ( n38965 , n38960 , n38964 );
and ( n38966 , n28129 , n25026 );
and ( n38967 , n26933 , n27246 );
and ( n38968 , n38966 , n38967 );
and ( n38969 , n26782 , n27558 );
and ( n38970 , n38967 , n38969 );
and ( n38971 , n38966 , n38969 );
or ( n38972 , n38968 , n38970 , n38971 );
xor ( n38973 , n38940 , n38941 );
xor ( n38974 , n38973 , n38943 );
or ( n38975 , n38972 , n38974 );
xor ( n38976 , n32425 , n33592 );
buf ( n38977 , n38976 );
buf ( n38978 , n38977 );
buf ( n38979 , n38978 );
and ( n38980 , n38979 , n28117 );
and ( n38981 , n27962 , n25284 );
and ( n38982 , n27863 , n25617 );
and ( n38983 , n38981 , n38982 );
and ( n38984 , n27591 , n26229 );
and ( n38985 , n38982 , n38984 );
and ( n38986 , n38981 , n38984 );
or ( n38987 , n38983 , n38985 , n38986 );
and ( n38988 , n38980 , n38987 );
and ( n38989 , n26980 , n26876 );
and ( n38990 , n25742 , n35169 );
and ( n38991 , n38989 , n38990 );
and ( n38992 , n25451 , n36229 );
and ( n38993 , n38990 , n38992 );
and ( n38994 , n38989 , n38992 );
or ( n38995 , n38991 , n38993 , n38994 );
and ( n38996 , n38987 , n38995 );
and ( n38997 , n38980 , n38995 );
or ( n38998 , n38988 , n38996 , n38997 );
and ( n38999 , n38975 , n38998 );
and ( n39000 , n35818 , n37197 );
and ( n39001 , n35386 , n37194 );
nor ( n39002 , n39000 , n39001 );
xnor ( n39003 , n39002 , n36218 );
and ( n39004 , n35718 , n36910 );
and ( n39005 , n35690 , n36908 );
nor ( n39006 , n39004 , n39005 );
xnor ( n39007 , n39006 , n36221 );
and ( n39008 , n39003 , n39007 );
and ( n39009 , n36411 , n36367 );
and ( n39010 , n36201 , n36365 );
nor ( n39011 , n39009 , n39010 );
xnor ( n39012 , n39011 , n35608 );
and ( n39013 , n39007 , n39012 );
and ( n39014 , n39003 , n39012 );
or ( n39015 , n39008 , n39013 , n39014 );
xor ( n39016 , n38718 , n38719 );
xor ( n39017 , n39016 , n38721 );
and ( n39018 , n39015 , n39017 );
xor ( n39019 , n38726 , n38727 );
xor ( n39020 , n39019 , n38729 );
and ( n39021 , n39017 , n39020 );
and ( n39022 , n39015 , n39020 );
or ( n39023 , n39018 , n39021 , n39022 );
and ( n39024 , n38998 , n39023 );
and ( n39025 , n38975 , n39023 );
or ( n39026 , n38999 , n39024 , n39025 );
and ( n39027 , n38964 , n39026 );
and ( n39028 , n38960 , n39026 );
or ( n39029 , n38965 , n39027 , n39028 );
and ( n39030 , n38939 , n39029 );
xor ( n39031 , n38738 , n38739 );
xor ( n39032 , n39031 , n38744 );
xor ( n39033 , n38751 , n38755 );
xor ( n39034 , n39033 , n38760 );
and ( n39035 , n39032 , n39034 );
xor ( n39036 , n38768 , n38772 );
xor ( n39037 , n39036 , n38781 );
and ( n39038 , n39034 , n39037 );
and ( n39039 , n39032 , n39037 );
or ( n39040 , n39035 , n39038 , n39039 );
xor ( n39041 , n38705 , n38707 );
xor ( n39042 , n39041 , n38709 );
and ( n39043 , n39040 , n39042 );
xor ( n39044 , n38717 , n38724 );
xor ( n39045 , n39044 , n38732 );
and ( n39046 , n39042 , n39045 );
and ( n39047 , n39040 , n39045 );
or ( n39048 , n39043 , n39046 , n39047 );
xor ( n39049 , n38689 , n38702 );
xor ( n39050 , n39049 , n38712 );
and ( n39051 , n39048 , n39050 );
xor ( n39052 , n38735 , n38787 );
xor ( n39053 , n39052 , n38798 );
and ( n39054 , n39050 , n39053 );
and ( n39055 , n39048 , n39053 );
or ( n39056 , n39051 , n39054 , n39055 );
and ( n39057 , n39029 , n39056 );
and ( n39058 , n38939 , n39056 );
or ( n39059 , n39030 , n39057 , n39058 );
and ( n39060 , n38929 , n39059 );
xor ( n39061 , n38662 , n38664 );
xor ( n39062 , n39061 , n38667 );
xor ( n39063 , n38687 , n38715 );
xor ( n39064 , n39063 , n38801 );
and ( n39065 , n39062 , n39064 );
xor ( n39066 , n38817 , n38819 );
xor ( n39067 , n39066 , n38822 );
and ( n39068 , n39064 , n39067 );
and ( n39069 , n39062 , n39067 );
or ( n39070 , n39065 , n39068 , n39069 );
and ( n39071 , n39059 , n39070 );
and ( n39072 , n38929 , n39070 );
or ( n39073 , n39060 , n39071 , n39072 );
and ( n39074 , n38881 , n39073 );
and ( n39075 , n38872 , n39073 );
or ( n39076 , n38882 , n39074 , n39075 );
xor ( n39077 , n38600 , n38602 );
xor ( n39078 , n39077 , n38605 );
xor ( n39079 , n38610 , n38649 );
xor ( n39080 , n39079 , n38655 );
and ( n39081 , n39078 , n39080 );
xor ( n39082 , n38807 , n38833 );
xor ( n39083 , n39082 , n38836 );
and ( n39084 , n39080 , n39083 );
and ( n39085 , n39078 , n39083 );
or ( n39086 , n39081 , n39084 , n39085 );
and ( n39087 , n39076 , n39086 );
xor ( n39088 , n38608 , n38658 );
xor ( n39089 , n39088 , n38839 );
and ( n39090 , n39086 , n39089 );
and ( n39091 , n39076 , n39089 );
or ( n39092 , n39087 , n39090 , n39091 );
and ( n39093 , n38869 , n39092 );
and ( n39094 , n38867 , n39092 );
or ( n39095 , n38870 , n39093 , n39094 );
xor ( n39096 , n38580 , n38856 );
xor ( n39097 , n39096 , n38859 );
and ( n39098 , n39095 , n39097 );
xor ( n39099 , n38582 , n38842 );
xor ( n39100 , n39099 , n38853 );
xor ( n39101 , n38845 , n38847 );
xor ( n39102 , n39101 , n38850 );
xor ( n39103 , n38660 , n38670 );
xor ( n39104 , n39103 , n38804 );
xor ( n39105 , n38825 , n38827 );
xor ( n39106 , n39105 , n38830 );
and ( n39107 , n39104 , n39106 );
xor ( n39108 , n38809 , n38811 );
xor ( n39109 , n39108 , n38814 );
xor ( n39110 , n38914 , n38918 );
xor ( n39111 , n39110 , n38923 );
and ( n39112 , n39109 , n39111 );
and ( n39113 , n25220 , n37187 );
and ( n39114 , n24731 , n38204 );
and ( n39115 , n39113 , n39114 );
and ( n39116 , n24624 , n38737 );
and ( n39117 , n39114 , n39116 );
and ( n39118 , n39113 , n39116 );
or ( n39119 , n39115 , n39117 , n39118 );
and ( n39120 , n25623 , n36229 );
and ( n39121 , n25451 , n36690 );
and ( n39122 , n39120 , n39121 );
and ( n39123 , n24993 , n37626 );
and ( n39124 , n39121 , n39123 );
and ( n39125 , n39120 , n39123 );
or ( n39126 , n39122 , n39124 , n39125 );
and ( n39127 , n39119 , n39126 );
and ( n39128 , n27389 , n26376 );
and ( n39129 , n39126 , n39128 );
and ( n39130 , n39119 , n39128 );
or ( n39131 , n39127 , n39129 , n39130 );
and ( n39132 , n28129 , n24540 );
and ( n39133 , n39131 , n39132 );
xor ( n39134 , n38949 , n38950 );
xor ( n39135 , n39134 , n38952 );
and ( n39136 , n39132 , n39135 );
and ( n39137 , n39131 , n39135 );
or ( n39138 , n39133 , n39136 , n39137 );
and ( n39139 , n38462 , n33632 );
and ( n39140 , n38003 , n33630 );
nor ( n39141 , n39139 , n39140 );
xnor ( n39142 , n39141 , n28124 );
and ( n39143 , n39138 , n39142 );
xor ( n39144 , n38946 , n38955 );
xor ( n39145 , n39144 , n38957 );
and ( n39146 , n39142 , n39145 );
and ( n39147 , n39138 , n39145 );
or ( n39148 , n39143 , n39146 , n39147 );
and ( n39149 , n39111 , n39148 );
and ( n39150 , n39109 , n39148 );
or ( n39151 , n39112 , n39149 , n39150 );
xor ( n39152 , n38747 , n38763 );
xor ( n39153 , n39152 , n38784 );
xor ( n39154 , n38790 , n38792 );
xor ( n39155 , n39154 , n38795 );
and ( n39156 , n39153 , n39155 );
xor ( n39157 , n38900 , n38908 );
xor ( n39158 , n39157 , n38911 );
and ( n39159 , n39155 , n39158 );
and ( n39160 , n39153 , n39158 );
or ( n39161 , n39156 , n39159 , n39160 );
xnor ( n39162 , n38961 , n38963 );
and ( n39163 , n26678 , n28209 );
and ( n39164 , n26399 , n33739 );
and ( n39165 , n39163 , n39164 );
and ( n39166 , n25623 , n35544 );
and ( n39167 , n39164 , n39166 );
and ( n39168 , n39163 , n39166 );
or ( n39169 , n39165 , n39167 , n39168 );
xor ( n39170 , n38947 , n38948 );
and ( n39171 , n26148 , n34122 );
and ( n39172 , n39170 , n39171 );
and ( n39173 , n25959 , n34817 );
and ( n39174 , n39171 , n39173 );
and ( n39175 , n39170 , n39173 );
or ( n39176 , n39172 , n39174 , n39175 );
and ( n39177 , n39169 , n39176 );
and ( n39178 , n27863 , n25284 );
and ( n39179 , n39176 , n39178 );
and ( n39180 , n39169 , n39178 );
or ( n39181 , n39177 , n39179 , n39180 );
and ( n39182 , n39162 , n39181 );
xor ( n39183 , n38894 , n38895 );
xor ( n39184 , n39183 , n38897 );
xor ( n39185 , n38901 , n38902 );
xor ( n39186 , n39185 , n38905 );
and ( n39187 , n39184 , n39186 );
and ( n39188 , n39181 , n39187 );
and ( n39189 , n39162 , n39187 );
or ( n39190 , n39182 , n39188 , n39189 );
and ( n39191 , n39161 , n39190 );
xnor ( n39192 , n38972 , n38974 );
and ( n39193 , n38979 , n33632 );
and ( n39194 , n38777 , n33630 );
nor ( n39195 , n39193 , n39194 );
xnor ( n39196 , n39195 , n28124 );
xor ( n39197 , n32494 , n33590 );
buf ( n39198 , n39197 );
buf ( n39199 , n39198 );
buf ( n39200 , n39199 );
and ( n39201 , n39200 , n28117 );
and ( n39202 , n39196 , n39201 );
xor ( n39203 , n38966 , n38967 );
xor ( n39204 , n39203 , n38969 );
and ( n39205 , n39201 , n39204 );
and ( n39206 , n39196 , n39204 );
or ( n39207 , n39202 , n39205 , n39206 );
and ( n39208 , n39192 , n39207 );
and ( n39209 , n37151 , n35911 );
and ( n39210 , n36427 , n35909 );
nor ( n39211 , n39209 , n39210 );
xnor ( n39212 , n39211 , n35161 );
and ( n39213 , n37387 , n35374 );
and ( n39214 , n37159 , n35372 );
nor ( n39215 , n39213 , n39214 );
xnor ( n39216 , n39215 , n34661 );
and ( n39217 , n39212 , n39216 );
xor ( n39218 , n38888 , n38889 );
xor ( n39219 , n39218 , n38891 );
and ( n39220 , n39216 , n39219 );
and ( n39221 , n39212 , n39219 );
or ( n39222 , n39217 , n39220 , n39221 );
and ( n39223 , n39207 , n39222 );
and ( n39224 , n39192 , n39222 );
or ( n39225 , n39208 , n39223 , n39224 );
and ( n39226 , n37159 , n35911 );
and ( n39227 , n37151 , n35909 );
nor ( n39228 , n39226 , n39227 );
xnor ( n39229 , n39228 , n35161 );
and ( n39230 , n38142 , n35374 );
and ( n39231 , n37387 , n35372 );
nor ( n39232 , n39230 , n39231 );
xnor ( n39233 , n39232 , n34661 );
or ( n39234 , n39229 , n39233 );
and ( n39235 , n28129 , n25284 );
and ( n39236 , n27962 , n25617 );
and ( n39237 , n39235 , n39236 );
and ( n39238 , n27863 , n26229 );
and ( n39239 , n39236 , n39238 );
and ( n39240 , n39235 , n39238 );
or ( n39241 , n39237 , n39239 , n39240 );
and ( n39242 , n39234 , n39241 );
and ( n39243 , n26782 , n28209 );
and ( n39244 , n26678 , n33739 );
and ( n39245 , n39243 , n39244 );
and ( n39246 , n26399 , n34122 );
and ( n39247 , n39244 , n39246 );
and ( n39248 , n39243 , n39246 );
or ( n39249 , n39245 , n39247 , n39248 );
and ( n39250 , n39241 , n39249 );
and ( n39251 , n39234 , n39249 );
or ( n39252 , n39242 , n39250 , n39251 );
and ( n39253 , n26148 , n34817 );
and ( n39254 , n25959 , n35169 );
and ( n39255 , n39253 , n39254 );
and ( n39256 , n25742 , n35544 );
and ( n39257 , n39254 , n39256 );
and ( n39258 , n39253 , n39256 );
or ( n39259 , n39255 , n39257 , n39258 );
buf ( n39260 , n14507 );
buf ( n39261 , n39260 );
and ( n39262 , n24546 , n39261 );
buf ( n39263 , n24337 );
and ( n39264 , n39262 , n39263 );
and ( n39265 , n35690 , n37197 );
and ( n39266 , n35818 , n37194 );
nor ( n39267 , n39265 , n39266 );
xnor ( n39268 , n39267 , n36218 );
and ( n39269 , n39263 , n39268 );
and ( n39270 , n39262 , n39268 );
or ( n39271 , n39264 , n39269 , n39270 );
and ( n39272 , n39259 , n39271 );
xor ( n39273 , n38981 , n38982 );
xor ( n39274 , n39273 , n38984 );
and ( n39275 , n39271 , n39274 );
and ( n39276 , n39259 , n39274 );
or ( n39277 , n39272 , n39275 , n39276 );
and ( n39278 , n39252 , n39277 );
xor ( n39279 , n38980 , n38987 );
xor ( n39280 , n39279 , n38995 );
and ( n39281 , n39277 , n39280 );
and ( n39282 , n39252 , n39280 );
or ( n39283 , n39278 , n39281 , n39282 );
and ( n39284 , n39225 , n39283 );
xor ( n39285 , n38975 , n38998 );
xor ( n39286 , n39285 , n39023 );
and ( n39287 , n39283 , n39286 );
and ( n39288 , n39225 , n39286 );
or ( n39289 , n39284 , n39287 , n39288 );
and ( n39290 , n39190 , n39289 );
and ( n39291 , n39161 , n39289 );
or ( n39292 , n39191 , n39290 , n39291 );
and ( n39293 , n39151 , n39292 );
xor ( n39294 , n38931 , n38933 );
xor ( n39295 , n39294 , n38936 );
xor ( n39296 , n38960 , n38964 );
xor ( n39297 , n39296 , n39026 );
and ( n39298 , n39295 , n39297 );
xor ( n39299 , n39048 , n39050 );
xor ( n39300 , n39299 , n39053 );
and ( n39301 , n39297 , n39300 );
and ( n39302 , n39295 , n39300 );
or ( n39303 , n39298 , n39301 , n39302 );
and ( n39304 , n39292 , n39303 );
and ( n39305 , n39151 , n39303 );
or ( n39306 , n39293 , n39304 , n39305 );
and ( n39307 , n39106 , n39306 );
and ( n39308 , n39104 , n39306 );
or ( n39309 , n39107 , n39307 , n39308 );
xor ( n39310 , n38884 , n38886 );
xor ( n39311 , n39310 , n38926 );
xor ( n39312 , n38939 , n39029 );
xor ( n39313 , n39312 , n39056 );
and ( n39314 , n39311 , n39313 );
xor ( n39315 , n39062 , n39064 );
xor ( n39316 , n39315 , n39067 );
and ( n39317 , n39313 , n39316 );
and ( n39318 , n39311 , n39316 );
or ( n39319 , n39314 , n39317 , n39318 );
xor ( n39320 , n38874 , n38876 );
xor ( n39321 , n39320 , n38878 );
and ( n39322 , n39319 , n39321 );
xor ( n39323 , n38929 , n39059 );
xor ( n39324 , n39323 , n39070 );
and ( n39325 , n39321 , n39324 );
and ( n39326 , n39319 , n39324 );
or ( n39327 , n39322 , n39325 , n39326 );
and ( n39328 , n39309 , n39327 );
xor ( n39329 , n38872 , n38881 );
xor ( n39330 , n39329 , n39073 );
and ( n39331 , n39327 , n39330 );
and ( n39332 , n39309 , n39330 );
or ( n39333 , n39328 , n39331 , n39332 );
and ( n39334 , n39102 , n39333 );
xor ( n39335 , n39076 , n39086 );
xor ( n39336 , n39335 , n39089 );
and ( n39337 , n39333 , n39336 );
and ( n39338 , n39102 , n39336 );
or ( n39339 , n39334 , n39337 , n39338 );
and ( n39340 , n39100 , n39339 );
xor ( n39341 , n38867 , n38869 );
xor ( n39342 , n39341 , n39092 );
and ( n39343 , n39339 , n39342 );
and ( n39344 , n39100 , n39342 );
or ( n39345 , n39340 , n39343 , n39344 );
and ( n39346 , n39097 , n39345 );
and ( n39347 , n39095 , n39345 );
or ( n39348 , n39098 , n39346 , n39347 );
and ( n39349 , n38864 , n39348 );
and ( n39350 , n38862 , n39348 );
or ( n39351 , n38865 , n39349 , n39350 );
and ( n39352 , n38577 , n39351 );
and ( n39353 , n38575 , n39351 );
or ( n39354 , n38578 , n39352 , n39353 );
and ( n39355 , n38301 , n39354 );
and ( n39356 , n38299 , n39354 );
or ( n39357 , n38302 , n39355 , n39356 );
and ( n39358 , n38296 , n39357 );
and ( n39359 , n38294 , n39357 );
or ( n39360 , n38297 , n39358 , n39359 );
and ( n39361 , n37761 , n39360 );
and ( n39362 , n37759 , n39360 );
or ( n39363 , n37762 , n39361 , n39362 );
and ( n39364 , n37576 , n39363 );
and ( n39365 , n37574 , n39363 );
or ( n39366 , n37577 , n39364 , n39365 );
or ( n39367 , n37497 , n39366 );
and ( n39368 , n37494 , n39367 );
and ( n39369 , n36676 , n39367 );
or ( n39370 , n37495 , n39368 , n39369 );
and ( n39371 , n36673 , n39370 );
and ( n39372 , n36511 , n39370 );
or ( n39373 , n36674 , n39371 , n39372 );
and ( n39374 , n36508 , n39373 );
and ( n39375 , n36506 , n39373 );
or ( n39376 , n36509 , n39374 , n39375 );
or ( n39377 , n36314 , n39376 );
and ( n39378 , n36311 , n39377 );
and ( n39379 , n36309 , n39377 );
or ( n39380 , n36312 , n39378 , n39379 );
and ( n39381 , n36078 , n39380 );
and ( n39382 , n35504 , n39380 );
or ( n39383 , n36079 , n39381 , n39382 );
and ( n39384 , n35502 , n39383 );
xor ( n39385 , n35502 , n39383 );
xor ( n39386 , n35504 , n36078 );
xor ( n39387 , n39386 , n39380 );
xor ( n39388 , n36309 , n36311 );
xor ( n39389 , n39388 , n39377 );
not ( n39390 , n39389 );
xnor ( n39391 , n36314 , n39376 );
xor ( n39392 , n36506 , n36508 );
xor ( n39393 , n39392 , n39373 );
not ( n39394 , n39393 );
xor ( n39395 , n36511 , n36673 );
xor ( n39396 , n39395 , n39370 );
not ( n39397 , n39396 );
xor ( n39398 , n36676 , n37494 );
xor ( n39399 , n39398 , n39367 );
not ( n39400 , n39399 );
xnor ( n39401 , n37497 , n39366 );
xor ( n39402 , n37574 , n37576 );
xor ( n39403 , n39402 , n39363 );
not ( n39404 , n39403 );
xor ( n39405 , n37759 , n37761 );
xor ( n39406 , n39405 , n39360 );
xor ( n39407 , n38294 , n38296 );
xor ( n39408 , n39407 , n39357 );
xor ( n39409 , n38299 , n38301 );
xor ( n39410 , n39409 , n39354 );
xor ( n39411 , n38575 , n38577 );
xor ( n39412 , n39411 , n39351 );
xor ( n39413 , n38862 , n38864 );
xor ( n39414 , n39413 , n39348 );
not ( n39415 , n39414 );
xor ( n39416 , n39095 , n39097 );
xor ( n39417 , n39416 , n39345 );
not ( n39418 , n39417 );
xor ( n39419 , n39100 , n39339 );
xor ( n39420 , n39419 , n39342 );
xor ( n39421 , n39078 , n39080 );
xor ( n39422 , n39421 , n39083 );
and ( n39423 , n35718 , n36367 );
and ( n39424 , n35690 , n36365 );
nor ( n39425 , n39423 , n39424 );
xnor ( n39426 , n39425 , n35608 );
xor ( n39427 , n39138 , n39142 );
xor ( n39428 , n39427 , n39145 );
and ( n39429 , n39426 , n39428 );
xor ( n39430 , n39040 , n39042 );
xor ( n39431 , n39430 , n39045 );
xor ( n39432 , n39015 , n39017 );
xor ( n39433 , n39432 , n39020 );
xor ( n39434 , n39032 , n39034 );
xor ( n39435 , n39434 , n39037 );
and ( n39436 , n39433 , n39435 );
xor ( n39437 , n39131 , n39132 );
xor ( n39438 , n39437 , n39135 );
and ( n39439 , n39435 , n39438 );
and ( n39440 , n39433 , n39438 );
or ( n39441 , n39436 , n39439 , n39440 );
and ( n39442 , n39431 , n39441 );
xor ( n39443 , n39184 , n39186 );
and ( n39444 , n27389 , n26876 );
and ( n39445 , n26933 , n27558 );
and ( n39446 , n39444 , n39445 );
xor ( n39447 , n39113 , n39114 );
xor ( n39448 , n39447 , n39116 );
and ( n39449 , n39445 , n39448 );
and ( n39450 , n39444 , n39448 );
or ( n39451 , n39446 , n39449 , n39450 );
xor ( n39452 , n39119 , n39126 );
xor ( n39453 , n39452 , n39128 );
or ( n39454 , n39451 , n39453 );
and ( n39455 , n39443 , n39454 );
xor ( n39456 , n38989 , n38990 );
xor ( n39457 , n39456 , n38992 );
xor ( n39458 , n39003 , n39007 );
xor ( n39459 , n39458 , n39012 );
and ( n39460 , n39457 , n39459 );
xor ( n39461 , n39196 , n39201 );
xor ( n39462 , n39461 , n39204 );
and ( n39463 , n39459 , n39462 );
and ( n39464 , n39457 , n39462 );
or ( n39465 , n39460 , n39463 , n39464 );
and ( n39466 , n39454 , n39465 );
and ( n39467 , n39443 , n39465 );
or ( n39468 , n39455 , n39466 , n39467 );
and ( n39469 , n39441 , n39468 );
and ( n39470 , n39431 , n39468 );
or ( n39471 , n39442 , n39469 , n39470 );
and ( n39472 , n39429 , n39471 );
and ( n39473 , n26148 , n35169 );
and ( n39474 , n25959 , n35544 );
and ( n39475 , n39473 , n39474 );
and ( n39476 , n25742 , n36229 );
and ( n39477 , n39474 , n39476 );
and ( n39478 , n39473 , n39476 );
or ( n39479 , n39475 , n39477 , n39478 );
and ( n39480 , n26782 , n33739 );
and ( n39481 , n26678 , n34122 );
and ( n39482 , n39480 , n39481 );
and ( n39483 , n26399 , n34817 );
and ( n39484 , n39481 , n39483 );
and ( n39485 , n39480 , n39483 );
or ( n39486 , n39482 , n39484 , n39485 );
and ( n39487 , n39479 , n39486 );
xor ( n39488 , n39120 , n39121 );
xor ( n39489 , n39488 , n39123 );
and ( n39490 , n39486 , n39489 );
and ( n39491 , n39479 , n39489 );
or ( n39492 , n39487 , n39490 , n39491 );
and ( n39493 , n36427 , n36367 );
and ( n39494 , n36411 , n36365 );
nor ( n39495 , n39493 , n39494 );
xnor ( n39496 , n39495 , n35608 );
xor ( n39497 , n32632 , n33588 );
buf ( n39498 , n39497 );
buf ( n39499 , n39498 );
buf ( n39500 , n39499 );
and ( n39501 , n39500 , n28117 );
and ( n39502 , n39496 , n39501 );
xnor ( n39503 , n39229 , n39233 );
and ( n39504 , n39501 , n39503 );
and ( n39505 , n39496 , n39503 );
or ( n39506 , n39502 , n39504 , n39505 );
and ( n39507 , n39492 , n39506 );
and ( n39508 , n24731 , n38737 );
and ( n39509 , n24624 , n39261 );
and ( n39510 , n39508 , n39509 );
and ( n39511 , n27863 , n26376 );
and ( n39512 , n27591 , n26876 );
and ( n39513 , n39511 , n39512 );
and ( n39514 , n27389 , n27246 );
and ( n39515 , n39512 , n39514 );
and ( n39516 , n39511 , n39514 );
or ( n39517 , n39513 , n39515 , n39516 );
and ( n39518 , n39510 , n39517 );
and ( n39519 , n26980 , n27558 );
and ( n39520 , n25451 , n37187 );
and ( n39521 , n39519 , n39520 );
and ( n39522 , n24993 , n38204 );
and ( n39523 , n39520 , n39522 );
and ( n39524 , n39519 , n39522 );
or ( n39525 , n39521 , n39523 , n39524 );
and ( n39526 , n39517 , n39525 );
and ( n39527 , n39510 , n39525 );
or ( n39528 , n39518 , n39526 , n39527 );
and ( n39529 , n39506 , n39528 );
and ( n39530 , n39492 , n39528 );
or ( n39531 , n39507 , n39529 , n39530 );
and ( n39532 , n35718 , n37197 );
and ( n39533 , n35690 , n37194 );
nor ( n39534 , n39532 , n39533 );
xnor ( n39535 , n39534 , n36218 );
and ( n39536 , n36411 , n36910 );
and ( n39537 , n36201 , n36908 );
nor ( n39538 , n39536 , n39537 );
xnor ( n39539 , n39538 , n36221 );
and ( n39540 , n39535 , n39539 );
and ( n39541 , n37151 , n36367 );
and ( n39542 , n36427 , n36365 );
nor ( n39543 , n39541 , n39542 );
xnor ( n39544 , n39543 , n35608 );
and ( n39545 , n39539 , n39544 );
and ( n39546 , n39535 , n39544 );
or ( n39547 , n39540 , n39545 , n39546 );
and ( n39548 , n37387 , n35911 );
and ( n39549 , n37159 , n35909 );
nor ( n39550 , n39548 , n39549 );
xnor ( n39551 , n39550 , n35161 );
and ( n39552 , n38359 , n35374 );
and ( n39553 , n38142 , n35372 );
nor ( n39554 , n39552 , n39553 );
xnor ( n39555 , n39554 , n34661 );
and ( n39556 , n39551 , n39555 );
and ( n39557 , n39500 , n33632 );
and ( n39558 , n39200 , n33630 );
nor ( n39559 , n39557 , n39558 );
xnor ( n39560 , n39559 , n28124 );
and ( n39561 , n39555 , n39560 );
and ( n39562 , n39551 , n39560 );
or ( n39563 , n39556 , n39561 , n39562 );
and ( n39564 , n39547 , n39563 );
xor ( n39565 , n39235 , n39236 );
xor ( n39566 , n39565 , n39238 );
and ( n39567 , n39563 , n39566 );
and ( n39568 , n39547 , n39566 );
or ( n39569 , n39564 , n39567 , n39568 );
xor ( n39570 , n39243 , n39244 );
xor ( n39571 , n39570 , n39246 );
xor ( n39572 , n39253 , n39254 );
xor ( n39573 , n39572 , n39256 );
and ( n39574 , n39571 , n39573 );
xor ( n39575 , n39262 , n39263 );
xor ( n39576 , n39575 , n39268 );
and ( n39577 , n39573 , n39576 );
and ( n39578 , n39571 , n39576 );
or ( n39579 , n39574 , n39577 , n39578 );
and ( n39580 , n39569 , n39579 );
xor ( n39581 , n39212 , n39216 );
xor ( n39582 , n39581 , n39219 );
and ( n39583 , n39579 , n39582 );
and ( n39584 , n39569 , n39582 );
or ( n39585 , n39580 , n39583 , n39584 );
and ( n39586 , n39531 , n39585 );
xor ( n39587 , n39192 , n39207 );
xor ( n39588 , n39587 , n39222 );
and ( n39589 , n39585 , n39588 );
and ( n39590 , n39531 , n39588 );
or ( n39591 , n39586 , n39589 , n39590 );
xor ( n39592 , n39153 , n39155 );
xor ( n39593 , n39592 , n39158 );
and ( n39594 , n39591 , n39593 );
xor ( n39595 , n39162 , n39181 );
xor ( n39596 , n39595 , n39187 );
and ( n39597 , n39593 , n39596 );
and ( n39598 , n39591 , n39596 );
or ( n39599 , n39594 , n39597 , n39598 );
and ( n39600 , n39471 , n39599 );
and ( n39601 , n39429 , n39599 );
or ( n39602 , n39472 , n39600 , n39601 );
xor ( n39603 , n39109 , n39111 );
xor ( n39604 , n39603 , n39148 );
xor ( n39605 , n39161 , n39190 );
xor ( n39606 , n39605 , n39289 );
and ( n39607 , n39604 , n39606 );
xor ( n39608 , n39295 , n39297 );
xor ( n39609 , n39608 , n39300 );
and ( n39610 , n39606 , n39609 );
and ( n39611 , n39604 , n39609 );
or ( n39612 , n39607 , n39610 , n39611 );
and ( n39613 , n39602 , n39612 );
xor ( n39614 , n39151 , n39292 );
xor ( n39615 , n39614 , n39303 );
and ( n39616 , n39612 , n39615 );
and ( n39617 , n39602 , n39615 );
or ( n39618 , n39613 , n39616 , n39617 );
xor ( n39619 , n39104 , n39106 );
xor ( n39620 , n39619 , n39306 );
and ( n39621 , n39618 , n39620 );
xor ( n39622 , n39319 , n39321 );
xor ( n39623 , n39622 , n39324 );
and ( n39624 , n39620 , n39623 );
and ( n39625 , n39618 , n39623 );
or ( n39626 , n39621 , n39624 , n39625 );
and ( n39627 , n39422 , n39626 );
xor ( n39628 , n39309 , n39327 );
xor ( n39629 , n39628 , n39330 );
and ( n39630 , n39626 , n39629 );
and ( n39631 , n39422 , n39629 );
or ( n39632 , n39627 , n39630 , n39631 );
xor ( n39633 , n39102 , n39333 );
xor ( n39634 , n39633 , n39336 );
and ( n39635 , n39632 , n39634 );
xor ( n39636 , n39422 , n39626 );
xor ( n39637 , n39636 , n39629 );
xor ( n39638 , n39311 , n39313 );
xor ( n39639 , n39638 , n39316 );
xor ( n39640 , n39225 , n39283 );
xor ( n39641 , n39640 , n39286 );
xor ( n39642 , n39426 , n39428 );
and ( n39643 , n39641 , n39642 );
xor ( n39644 , n39508 , n39509 );
and ( n39645 , n25623 , n36690 );
and ( n39646 , n39644 , n39645 );
and ( n39647 , n25220 , n37626 );
and ( n39648 , n39645 , n39647 );
and ( n39649 , n39644 , n39647 );
or ( n39650 , n39646 , n39648 , n39649 );
and ( n39651 , n27591 , n26376 );
and ( n39652 , n39650 , n39651 );
and ( n39653 , n26980 , n27246 );
and ( n39654 , n39651 , n39653 );
and ( n39655 , n39650 , n39653 );
or ( n39656 , n39652 , n39654 , n39655 );
xor ( n39657 , n39163 , n39164 );
xor ( n39658 , n39657 , n39166 );
and ( n39659 , n39656 , n39658 );
xor ( n39660 , n39170 , n39171 );
xor ( n39661 , n39660 , n39173 );
and ( n39662 , n39658 , n39661 );
and ( n39663 , n39656 , n39661 );
or ( n39664 , n39659 , n39662 , n39663 );
and ( n39665 , n38003 , n34352 );
and ( n39666 , n38359 , n34350 );
nor ( n39667 , n39665 , n39666 );
xnor ( n39668 , n39667 , n28532 );
and ( n39669 , n39664 , n39668 );
xor ( n39670 , n39169 , n39176 );
xor ( n39671 , n39670 , n39178 );
and ( n39672 , n39668 , n39671 );
and ( n39673 , n39664 , n39671 );
or ( n39674 , n39669 , n39672 , n39673 );
and ( n39675 , n39642 , n39674 );
and ( n39676 , n39641 , n39674 );
or ( n39677 , n39643 , n39675 , n39676 );
xor ( n39678 , n39252 , n39277 );
xor ( n39679 , n39678 , n39280 );
xor ( n39680 , n39234 , n39241 );
xor ( n39681 , n39680 , n39249 );
xor ( n39682 , n39259 , n39271 );
xor ( n39683 , n39682 , n39274 );
and ( n39684 , n39681 , n39683 );
xnor ( n39685 , n39451 , n39453 );
and ( n39686 , n39683 , n39685 );
and ( n39687 , n39681 , n39685 );
or ( n39688 , n39684 , n39686 , n39687 );
and ( n39689 , n39679 , n39688 );
and ( n39690 , n38003 , n34911 );
and ( n39691 , n38359 , n34909 );
nor ( n39692 , n39690 , n39691 );
xnor ( n39693 , n39692 , n34104 );
xor ( n39694 , n39479 , n39486 );
xor ( n39695 , n39694 , n39489 );
or ( n39696 , n39693 , n39695 );
xor ( n39697 , n39444 , n39445 );
xor ( n39698 , n39697 , n39448 );
xor ( n39699 , n39480 , n39481 );
xor ( n39700 , n39699 , n39483 );
and ( n39701 , n27863 , n26876 );
and ( n39702 , n27389 , n27558 );
and ( n39703 , n39701 , n39702 );
and ( n39704 , n26980 , n28209 );
and ( n39705 , n39702 , n39704 );
and ( n39706 , n39701 , n39704 );
or ( n39707 , n39703 , n39705 , n39706 );
and ( n39708 , n39700 , n39707 );
and ( n39709 , n25742 , n36690 );
and ( n39710 , n25623 , n37187 );
and ( n39711 , n39709 , n39710 );
buf ( n39712 , n14700 );
buf ( n39713 , n39712 );
and ( n39714 , n24624 , n39713 );
and ( n39715 , n39710 , n39714 );
and ( n39716 , n39709 , n39714 );
or ( n39717 , n39711 , n39715 , n39716 );
and ( n39718 , n39707 , n39717 );
and ( n39719 , n39700 , n39717 );
or ( n39720 , n39708 , n39718 , n39719 );
and ( n39721 , n39698 , n39720 );
buf ( n39722 , n24546 );
and ( n39723 , n36201 , n37197 );
and ( n39724 , n35718 , n37194 );
nor ( n39725 , n39723 , n39724 );
xnor ( n39726 , n39725 , n36218 );
and ( n39727 , n39722 , n39726 );
and ( n39728 , n36427 , n36910 );
and ( n39729 , n36411 , n36908 );
nor ( n39730 , n39728 , n39729 );
xnor ( n39731 , n39730 , n36221 );
and ( n39732 , n39726 , n39731 );
and ( n39733 , n39722 , n39731 );
or ( n39734 , n39727 , n39732 , n39733 );
and ( n39735 , n37159 , n36367 );
and ( n39736 , n37151 , n36365 );
nor ( n39737 , n39735 , n39736 );
xnor ( n39738 , n39737 , n35608 );
and ( n39739 , n38142 , n35911 );
and ( n39740 , n37387 , n35909 );
nor ( n39741 , n39739 , n39740 );
xnor ( n39742 , n39741 , n35161 );
and ( n39743 , n39738 , n39742 );
and ( n39744 , n38003 , n35374 );
and ( n39745 , n38359 , n35372 );
nor ( n39746 , n39744 , n39745 );
xnor ( n39747 , n39746 , n34661 );
and ( n39748 , n39742 , n39747 );
and ( n39749 , n39738 , n39747 );
or ( n39750 , n39743 , n39748 , n39749 );
and ( n39751 , n39734 , n39750 );
and ( n39752 , n38777 , n34911 );
and ( n39753 , n38462 , n34909 );
nor ( n39754 , n39752 , n39753 );
xnor ( n39755 , n39754 , n34104 );
xor ( n39756 , n32702 , n33586 );
buf ( n39757 , n39756 );
buf ( n39758 , n39757 );
buf ( n39759 , n39758 );
and ( n39760 , n39759 , n33632 );
and ( n39761 , n39500 , n33630 );
nor ( n39762 , n39760 , n39761 );
xnor ( n39763 , n39762 , n28124 );
and ( n39764 , n39755 , n39763 );
xor ( n39765 , n32778 , n33584 );
buf ( n39766 , n39765 );
buf ( n39767 , n39766 );
buf ( n39768 , n39767 );
and ( n39769 , n39768 , n28117 );
and ( n39770 , n39763 , n39769 );
and ( n39771 , n39755 , n39769 );
or ( n39772 , n39764 , n39770 , n39771 );
and ( n39773 , n39750 , n39772 );
and ( n39774 , n39734 , n39772 );
or ( n39775 , n39751 , n39773 , n39774 );
and ( n39776 , n39720 , n39775 );
and ( n39777 , n39698 , n39775 );
or ( n39778 , n39721 , n39776 , n39777 );
and ( n39779 , n39696 , n39778 );
xor ( n39780 , n39511 , n39512 );
xor ( n39781 , n39780 , n39514 );
xor ( n39782 , n39519 , n39520 );
xor ( n39783 , n39782 , n39522 );
and ( n39784 , n39781 , n39783 );
xor ( n39785 , n39535 , n39539 );
xor ( n39786 , n39785 , n39544 );
and ( n39787 , n39783 , n39786 );
and ( n39788 , n39781 , n39786 );
or ( n39789 , n39784 , n39787 , n39788 );
xor ( n39790 , n39496 , n39501 );
xor ( n39791 , n39790 , n39503 );
and ( n39792 , n39789 , n39791 );
xor ( n39793 , n39510 , n39517 );
xor ( n39794 , n39793 , n39525 );
and ( n39795 , n39791 , n39794 );
and ( n39796 , n39789 , n39794 );
or ( n39797 , n39792 , n39795 , n39796 );
and ( n39798 , n39778 , n39797 );
and ( n39799 , n39696 , n39797 );
or ( n39800 , n39779 , n39798 , n39799 );
and ( n39801 , n39688 , n39800 );
and ( n39802 , n39679 , n39800 );
or ( n39803 , n39689 , n39801 , n39802 );
xor ( n39804 , n39457 , n39459 );
xor ( n39805 , n39804 , n39462 );
xor ( n39806 , n39492 , n39506 );
xor ( n39807 , n39806 , n39528 );
and ( n39808 , n39805 , n39807 );
xor ( n39809 , n39569 , n39579 );
xor ( n39810 , n39809 , n39582 );
and ( n39811 , n39807 , n39810 );
and ( n39812 , n39805 , n39810 );
or ( n39813 , n39808 , n39811 , n39812 );
xor ( n39814 , n39433 , n39435 );
xor ( n39815 , n39814 , n39438 );
and ( n39816 , n39813 , n39815 );
xor ( n39817 , n39443 , n39454 );
xor ( n39818 , n39817 , n39465 );
and ( n39819 , n39815 , n39818 );
and ( n39820 , n39813 , n39818 );
or ( n39821 , n39816 , n39819 , n39820 );
and ( n39822 , n39803 , n39821 );
xor ( n39823 , n39431 , n39441 );
xor ( n39824 , n39823 , n39468 );
and ( n39825 , n39821 , n39824 );
and ( n39826 , n39803 , n39824 );
or ( n39827 , n39822 , n39825 , n39826 );
and ( n39828 , n39677 , n39827 );
xor ( n39829 , n39429 , n39471 );
xor ( n39830 , n39829 , n39599 );
and ( n39831 , n39827 , n39830 );
and ( n39832 , n39677 , n39830 );
or ( n39833 , n39828 , n39831 , n39832 );
and ( n39834 , n39639 , n39833 );
xor ( n39835 , n39602 , n39612 );
xor ( n39836 , n39835 , n39615 );
and ( n39837 , n39833 , n39836 );
and ( n39838 , n39639 , n39836 );
or ( n39839 , n39834 , n39837 , n39838 );
xor ( n39840 , n39618 , n39620 );
xor ( n39841 , n39840 , n39623 );
and ( n39842 , n39839 , n39841 );
xor ( n39843 , n39604 , n39606 );
xor ( n39844 , n39843 , n39609 );
xor ( n39845 , n39591 , n39593 );
xor ( n39846 , n39845 , n39596 );
xor ( n39847 , n39531 , n39585 );
xor ( n39848 , n39847 , n39588 );
xor ( n39849 , n39664 , n39668 );
xor ( n39850 , n39849 , n39671 );
and ( n39851 , n39848 , n39850 );
and ( n39852 , n38359 , n34911 );
and ( n39853 , n38142 , n34909 );
nor ( n39854 , n39852 , n39853 );
xnor ( n39855 , n39854 , n34104 );
and ( n39856 , n38462 , n34352 );
and ( n39857 , n38003 , n34350 );
nor ( n39858 , n39856 , n39857 );
xnor ( n39859 , n39858 , n28532 );
and ( n39860 , n39855 , n39859 );
xor ( n39861 , n39656 , n39658 );
xor ( n39862 , n39861 , n39661 );
and ( n39863 , n39859 , n39862 );
and ( n39864 , n39855 , n39862 );
or ( n39865 , n39860 , n39863 , n39864 );
and ( n39866 , n39850 , n39865 );
and ( n39867 , n39848 , n39865 );
or ( n39868 , n39851 , n39866 , n39867 );
and ( n39869 , n39846 , n39868 );
and ( n39870 , n38777 , n34352 );
and ( n39871 , n38462 , n34350 );
nor ( n39872 , n39870 , n39871 );
xnor ( n39873 , n39872 , n28532 );
and ( n39874 , n39200 , n33632 );
and ( n39875 , n38979 , n33630 );
nor ( n39876 , n39874 , n39875 );
xnor ( n39877 , n39876 , n28124 );
and ( n39878 , n39873 , n39877 );
xor ( n39879 , n39650 , n39651 );
xor ( n39880 , n39879 , n39653 );
and ( n39881 , n39877 , n39880 );
and ( n39882 , n39873 , n39880 );
or ( n39883 , n39878 , n39881 , n39882 );
xor ( n39884 , n39547 , n39563 );
xor ( n39885 , n39884 , n39566 );
xor ( n39886 , n39571 , n39573 );
xor ( n39887 , n39886 , n39576 );
and ( n39888 , n39885 , n39887 );
xnor ( n39889 , n39693 , n39695 );
and ( n39890 , n39887 , n39889 );
and ( n39891 , n39885 , n39889 );
or ( n39892 , n39888 , n39890 , n39891 );
and ( n39893 , n39883 , n39892 );
and ( n39894 , n25220 , n38204 );
and ( n39895 , n24993 , n38737 );
and ( n39896 , n39894 , n39895 );
and ( n39897 , n24731 , n39261 );
and ( n39898 , n39895 , n39897 );
and ( n39899 , n39894 , n39897 );
or ( n39900 , n39896 , n39898 , n39899 );
and ( n39901 , n24993 , n39261 );
and ( n39902 , n24731 , n39713 );
and ( n39903 , n39901 , n39902 );
and ( n39904 , n25959 , n36229 );
and ( n39905 , n39903 , n39904 );
and ( n39906 , n25451 , n37626 );
and ( n39907 , n39904 , n39906 );
and ( n39908 , n39903 , n39906 );
or ( n39909 , n39905 , n39907 , n39908 );
and ( n39910 , n39900 , n39909 );
and ( n39911 , n26933 , n28209 );
and ( n39912 , n39909 , n39911 );
and ( n39913 , n39900 , n39911 );
or ( n39914 , n39910 , n39912 , n39913 );
and ( n39915 , n26678 , n34817 );
and ( n39916 , n26399 , n35169 );
and ( n39917 , n39915 , n39916 );
and ( n39918 , n26148 , n35544 );
and ( n39919 , n39916 , n39918 );
and ( n39920 , n39915 , n39918 );
or ( n39921 , n39917 , n39919 , n39920 );
and ( n39922 , n26933 , n33739 );
and ( n39923 , n26782 , n34122 );
and ( n39924 , n39922 , n39923 );
xor ( n39925 , n39894 , n39895 );
xor ( n39926 , n39925 , n39897 );
and ( n39927 , n39923 , n39926 );
and ( n39928 , n39922 , n39926 );
or ( n39929 , n39924 , n39927 , n39928 );
and ( n39930 , n39921 , n39929 );
xor ( n39931 , n39473 , n39474 );
xor ( n39932 , n39931 , n39476 );
and ( n39933 , n39929 , n39932 );
and ( n39934 , n39921 , n39932 );
or ( n39935 , n39930 , n39933 , n39934 );
and ( n39936 , n39914 , n39935 );
and ( n39937 , n28129 , n25617 );
and ( n39938 , n27962 , n26229 );
and ( n39939 , n39937 , n39938 );
xor ( n39940 , n39644 , n39645 );
xor ( n39941 , n39940 , n39647 );
and ( n39942 , n39938 , n39941 );
and ( n39943 , n39937 , n39941 );
or ( n39944 , n39939 , n39942 , n39943 );
and ( n39945 , n39935 , n39944 );
and ( n39946 , n39914 , n39944 );
or ( n39947 , n39936 , n39945 , n39946 );
and ( n39948 , n39892 , n39947 );
and ( n39949 , n39883 , n39947 );
or ( n39950 , n39893 , n39948 , n39949 );
xor ( n39951 , n39551 , n39555 );
xor ( n39952 , n39951 , n39560 );
and ( n39953 , n26148 , n36229 );
and ( n39954 , n25742 , n37187 );
and ( n39955 , n39953 , n39954 );
and ( n39956 , n25623 , n37626 );
and ( n39957 , n39954 , n39956 );
and ( n39958 , n39953 , n39956 );
or ( n39959 , n39955 , n39957 , n39958 );
and ( n39960 , n27962 , n26376 );
and ( n39961 , n39959 , n39960 );
and ( n39962 , n27591 , n27246 );
and ( n39963 , n39960 , n39962 );
and ( n39964 , n39959 , n39962 );
or ( n39965 , n39961 , n39963 , n39964 );
and ( n39966 , n39952 , n39965 );
xor ( n39967 , n39915 , n39916 );
xor ( n39968 , n39967 , n39918 );
and ( n39969 , n27962 , n26876 );
and ( n39970 , n27863 , n27246 );
and ( n39971 , n39969 , n39970 );
and ( n39972 , n27389 , n28209 );
and ( n39973 , n39970 , n39972 );
and ( n39974 , n39969 , n39972 );
or ( n39975 , n39971 , n39973 , n39974 );
and ( n39976 , n39968 , n39975 );
and ( n39977 , n26980 , n33739 );
and ( n39978 , n26933 , n34122 );
and ( n39979 , n39977 , n39978 );
and ( n39980 , n25451 , n38204 );
and ( n39981 , n39978 , n39980 );
and ( n39982 , n39977 , n39980 );
or ( n39983 , n39979 , n39981 , n39982 );
and ( n39984 , n39975 , n39983 );
and ( n39985 , n39968 , n39983 );
or ( n39986 , n39976 , n39984 , n39985 );
and ( n39987 , n39965 , n39986 );
and ( n39988 , n39952 , n39986 );
or ( n39989 , n39966 , n39987 , n39988 );
and ( n39990 , n25220 , n38737 );
and ( n39991 , n36411 , n37197 );
and ( n39992 , n36201 , n37194 );
nor ( n39993 , n39991 , n39992 );
xnor ( n39994 , n39993 , n36218 );
and ( n39995 , n39990 , n39994 );
and ( n39996 , n37151 , n36910 );
and ( n39997 , n36427 , n36908 );
nor ( n39998 , n39996 , n39997 );
xnor ( n39999 , n39998 , n36221 );
and ( n40000 , n39994 , n39999 );
and ( n40001 , n39990 , n39999 );
or ( n40002 , n39995 , n40000 , n40001 );
and ( n40003 , n37387 , n36367 );
and ( n40004 , n37159 , n36365 );
nor ( n40005 , n40003 , n40004 );
xnor ( n40006 , n40005 , n35608 );
and ( n40007 , n38359 , n35911 );
and ( n40008 , n38142 , n35909 );
nor ( n40009 , n40007 , n40008 );
xnor ( n40010 , n40009 , n35161 );
and ( n40011 , n40006 , n40010 );
and ( n40012 , n39500 , n34352 );
and ( n40013 , n39200 , n34350 );
nor ( n40014 , n40012 , n40013 );
xnor ( n40015 , n40014 , n28532 );
and ( n40016 , n40010 , n40015 );
and ( n40017 , n40006 , n40015 );
or ( n40018 , n40011 , n40016 , n40017 );
and ( n40019 , n40002 , n40018 );
xor ( n40020 , n39701 , n39702 );
xor ( n40021 , n40020 , n39704 );
and ( n40022 , n40018 , n40021 );
and ( n40023 , n40002 , n40021 );
or ( n40024 , n40019 , n40022 , n40023 );
xor ( n40025 , n39709 , n39710 );
xor ( n40026 , n40025 , n39714 );
xor ( n40027 , n39722 , n39726 );
xor ( n40028 , n40027 , n39731 );
and ( n40029 , n40026 , n40028 );
xor ( n40030 , n39738 , n39742 );
xor ( n40031 , n40030 , n39747 );
and ( n40032 , n40028 , n40031 );
and ( n40033 , n40026 , n40031 );
or ( n40034 , n40029 , n40032 , n40033 );
and ( n40035 , n40024 , n40034 );
xor ( n40036 , n39700 , n39707 );
xor ( n40037 , n40036 , n39717 );
and ( n40038 , n40034 , n40037 );
and ( n40039 , n40024 , n40037 );
or ( n40040 , n40035 , n40038 , n40039 );
and ( n40041 , n39989 , n40040 );
xor ( n40042 , n39698 , n39720 );
xor ( n40043 , n40042 , n39775 );
and ( n40044 , n40040 , n40043 );
and ( n40045 , n39989 , n40043 );
or ( n40046 , n40041 , n40044 , n40045 );
xor ( n40047 , n39681 , n39683 );
xor ( n40048 , n40047 , n39685 );
and ( n40049 , n40046 , n40048 );
xor ( n40050 , n39696 , n39778 );
xor ( n40051 , n40050 , n39797 );
and ( n40052 , n40048 , n40051 );
and ( n40053 , n40046 , n40051 );
or ( n40054 , n40049 , n40052 , n40053 );
and ( n40055 , n39950 , n40054 );
xor ( n40056 , n39679 , n39688 );
xor ( n40057 , n40056 , n39800 );
and ( n40058 , n40054 , n40057 );
and ( n40059 , n39950 , n40057 );
or ( n40060 , n40055 , n40058 , n40059 );
and ( n40061 , n39868 , n40060 );
and ( n40062 , n39846 , n40060 );
or ( n40063 , n39869 , n40061 , n40062 );
and ( n40064 , n39844 , n40063 );
xor ( n40065 , n39677 , n39827 );
xor ( n40066 , n40065 , n39830 );
and ( n40067 , n40063 , n40066 );
and ( n40068 , n39844 , n40066 );
or ( n40069 , n40064 , n40067 , n40068 );
xor ( n40070 , n39639 , n39833 );
xor ( n40071 , n40070 , n39836 );
and ( n40072 , n40069 , n40071 );
xor ( n40073 , n39641 , n39642 );
xor ( n40074 , n40073 , n39674 );
xor ( n40075 , n39803 , n39821 );
xor ( n40076 , n40075 , n39824 );
and ( n40077 , n40074 , n40076 );
xor ( n40078 , n39813 , n39815 );
xor ( n40079 , n40078 , n39818 );
xor ( n40080 , n39805 , n39807 );
xor ( n40081 , n40080 , n39810 );
xor ( n40082 , n39855 , n39859 );
xor ( n40083 , n40082 , n39862 );
and ( n40084 , n40081 , n40083 );
and ( n40085 , n25451 , n38737 );
and ( n40086 , n25220 , n39261 );
and ( n40087 , n40085 , n40086 );
and ( n40088 , n24993 , n39713 );
and ( n40089 , n40086 , n40088 );
and ( n40090 , n40085 , n40088 );
or ( n40091 , n40087 , n40089 , n40090 );
and ( n40092 , n26782 , n34817 );
and ( n40093 , n40091 , n40092 );
and ( n40094 , n26399 , n35544 );
and ( n40095 , n40092 , n40094 );
and ( n40096 , n40091 , n40094 );
or ( n40097 , n40093 , n40095 , n40096 );
and ( n40098 , n28129 , n26229 );
and ( n40099 , n40097 , n40098 );
xor ( n40100 , n39903 , n39904 );
xor ( n40101 , n40100 , n39906 );
and ( n40102 , n40098 , n40101 );
and ( n40103 , n40097 , n40101 );
or ( n40104 , n40099 , n40102 , n40103 );
and ( n40105 , n38979 , n34352 );
and ( n40106 , n38777 , n34350 );
nor ( n40107 , n40105 , n40106 );
xnor ( n40108 , n40107 , n28532 );
and ( n40109 , n40104 , n40108 );
xor ( n40110 , n39937 , n39938 );
xor ( n40111 , n40110 , n39941 );
and ( n40112 , n40108 , n40111 );
and ( n40113 , n40104 , n40111 );
or ( n40114 , n40109 , n40112 , n40113 );
and ( n40115 , n36201 , n36910 );
and ( n40116 , n35718 , n36908 );
nor ( n40117 , n40115 , n40116 );
xnor ( n40118 , n40117 , n36221 );
and ( n40119 , n40114 , n40118 );
xor ( n40120 , n39873 , n39877 );
xor ( n40121 , n40120 , n39880 );
and ( n40122 , n40118 , n40121 );
and ( n40123 , n40114 , n40121 );
or ( n40124 , n40119 , n40122 , n40123 );
and ( n40125 , n40083 , n40124 );
and ( n40126 , n40081 , n40124 );
or ( n40127 , n40084 , n40125 , n40126 );
and ( n40128 , n40079 , n40127 );
xor ( n40129 , n39789 , n39791 );
xor ( n40130 , n40129 , n39794 );
and ( n40131 , n39759 , n28117 );
xor ( n40132 , n39900 , n39909 );
xor ( n40133 , n40132 , n39911 );
or ( n40134 , n40131 , n40133 );
and ( n40135 , n40130 , n40134 );
and ( n40136 , n38462 , n34911 );
and ( n40137 , n38003 , n34909 );
nor ( n40138 , n40136 , n40137 );
xnor ( n40139 , n40138 , n34104 );
xor ( n40140 , n39921 , n39929 );
xor ( n40141 , n40140 , n39932 );
or ( n40142 , n40139 , n40141 );
and ( n40143 , n40134 , n40142 );
and ( n40144 , n40130 , n40142 );
or ( n40145 , n40135 , n40143 , n40144 );
xor ( n40146 , n39734 , n39750 );
xor ( n40147 , n40146 , n39772 );
xor ( n40148 , n39781 , n39783 );
xor ( n40149 , n40148 , n39786 );
and ( n40150 , n40147 , n40149 );
xor ( n40151 , n39755 , n39763 );
xor ( n40152 , n40151 , n39769 );
xor ( n40153 , n39922 , n39923 );
xor ( n40154 , n40153 , n39926 );
and ( n40155 , n40152 , n40154 );
xor ( n40156 , n39901 , n39902 );
and ( n40157 , n26678 , n35169 );
and ( n40158 , n40156 , n40157 );
and ( n40159 , n25959 , n36690 );
and ( n40160 , n40157 , n40159 );
and ( n40161 , n40156 , n40159 );
or ( n40162 , n40158 , n40160 , n40161 );
and ( n40163 , n40154 , n40162 );
and ( n40164 , n40152 , n40162 );
or ( n40165 , n40155 , n40163 , n40164 );
and ( n40166 , n40149 , n40165 );
and ( n40167 , n40147 , n40165 );
or ( n40168 , n40150 , n40166 , n40167 );
xor ( n40169 , n32847 , n33582 );
buf ( n40170 , n40169 );
buf ( n40171 , n40170 );
buf ( n40172 , n40171 );
and ( n40173 , n40172 , n28117 );
and ( n40174 , n27962 , n27246 );
xor ( n40175 , n32913 , n33580 );
buf ( n40176 , n40175 );
buf ( n40177 , n40176 );
buf ( n40178 , n40177 );
and ( n40179 , n40178 , n28117 );
or ( n40180 , n40174 , n40179 );
and ( n40181 , n40173 , n40180 );
and ( n40182 , n28129 , n26876 );
and ( n40183 , n26782 , n35169 );
and ( n40184 , n40182 , n40183 );
and ( n40185 , n25959 , n37187 );
and ( n40186 , n40183 , n40185 );
and ( n40187 , n40182 , n40185 );
or ( n40188 , n40184 , n40186 , n40187 );
and ( n40189 , n40180 , n40188 );
and ( n40190 , n40173 , n40188 );
or ( n40191 , n40181 , n40189 , n40190 );
and ( n40192 , n25742 , n37626 );
and ( n40193 , n25623 , n38204 );
and ( n40194 , n40192 , n40193 );
buf ( n40195 , n14989 );
buf ( n40196 , n40195 );
and ( n40197 , n24731 , n40196 );
and ( n40198 , n40193 , n40197 );
and ( n40199 , n40192 , n40197 );
or ( n40200 , n40194 , n40198 , n40199 );
buf ( n40201 , n24624 );
and ( n40202 , n36427 , n37197 );
and ( n40203 , n36411 , n37194 );
nor ( n40204 , n40202 , n40203 );
xnor ( n40205 , n40204 , n36218 );
and ( n40206 , n40201 , n40205 );
and ( n40207 , n38777 , n35374 );
and ( n40208 , n38462 , n35372 );
nor ( n40209 , n40207 , n40208 );
xnor ( n40210 , n40209 , n34661 );
and ( n40211 , n40205 , n40210 );
and ( n40212 , n40201 , n40210 );
or ( n40213 , n40206 , n40211 , n40212 );
and ( n40214 , n40200 , n40213 );
xor ( n40215 , n39969 , n39970 );
xor ( n40216 , n40215 , n39972 );
and ( n40217 , n40213 , n40216 );
and ( n40218 , n40200 , n40216 );
or ( n40219 , n40214 , n40217 , n40218 );
and ( n40220 , n40191 , n40219 );
xor ( n40221 , n39977 , n39978 );
xor ( n40222 , n40221 , n39980 );
xor ( n40223 , n39990 , n39994 );
xor ( n40224 , n40223 , n39999 );
and ( n40225 , n40222 , n40224 );
xor ( n40226 , n40006 , n40010 );
xor ( n40227 , n40226 , n40015 );
and ( n40228 , n40224 , n40227 );
and ( n40229 , n40222 , n40227 );
or ( n40230 , n40225 , n40228 , n40229 );
and ( n40231 , n40219 , n40230 );
and ( n40232 , n40191 , n40230 );
or ( n40233 , n40220 , n40231 , n40232 );
xor ( n40234 , n39968 , n39975 );
xor ( n40235 , n40234 , n39983 );
xor ( n40236 , n40002 , n40018 );
xor ( n40237 , n40236 , n40021 );
and ( n40238 , n40235 , n40237 );
xor ( n40239 , n40026 , n40028 );
xor ( n40240 , n40239 , n40031 );
and ( n40241 , n40237 , n40240 );
and ( n40242 , n40235 , n40240 );
or ( n40243 , n40238 , n40241 , n40242 );
and ( n40244 , n40233 , n40243 );
xor ( n40245 , n39952 , n39965 );
xor ( n40246 , n40245 , n39986 );
and ( n40247 , n40243 , n40246 );
and ( n40248 , n40233 , n40246 );
or ( n40249 , n40244 , n40247 , n40248 );
and ( n40250 , n40168 , n40249 );
xor ( n40251 , n39885 , n39887 );
xor ( n40252 , n40251 , n39889 );
and ( n40253 , n40249 , n40252 );
and ( n40254 , n40168 , n40252 );
or ( n40255 , n40250 , n40253 , n40254 );
and ( n40256 , n40145 , n40255 );
xor ( n40257 , n39883 , n39892 );
xor ( n40258 , n40257 , n39947 );
and ( n40259 , n40255 , n40258 );
and ( n40260 , n40145 , n40258 );
or ( n40261 , n40256 , n40259 , n40260 );
and ( n40262 , n40127 , n40261 );
and ( n40263 , n40079 , n40261 );
or ( n40264 , n40128 , n40262 , n40263 );
and ( n40265 , n40076 , n40264 );
and ( n40266 , n40074 , n40264 );
or ( n40267 , n40077 , n40265 , n40266 );
xor ( n40268 , n39844 , n40063 );
xor ( n40269 , n40268 , n40066 );
and ( n40270 , n40267 , n40269 );
xor ( n40271 , n39846 , n39868 );
xor ( n40272 , n40271 , n40060 );
xor ( n40273 , n39848 , n39850 );
xor ( n40274 , n40273 , n39865 );
xor ( n40275 , n39950 , n40054 );
xor ( n40276 , n40275 , n40057 );
and ( n40277 , n40274 , n40276 );
xor ( n40278 , n40046 , n40048 );
xor ( n40279 , n40278 , n40051 );
xor ( n40280 , n39914 , n39935 );
xor ( n40281 , n40280 , n39944 );
xor ( n40282 , n39989 , n40040 );
xor ( n40283 , n40282 , n40043 );
and ( n40284 , n40281 , n40283 );
xor ( n40285 , n40114 , n40118 );
xor ( n40286 , n40285 , n40121 );
and ( n40287 , n40283 , n40286 );
and ( n40288 , n40281 , n40286 );
or ( n40289 , n40284 , n40287 , n40288 );
and ( n40290 , n40279 , n40289 );
xor ( n40291 , n40024 , n40034 );
xor ( n40292 , n40291 , n40037 );
xor ( n40293 , n40104 , n40108 );
xor ( n40294 , n40293 , n40111 );
and ( n40295 , n40292 , n40294 );
xnor ( n40296 , n40131 , n40133 );
and ( n40297 , n40294 , n40296 );
and ( n40298 , n40292 , n40296 );
or ( n40299 , n40295 , n40297 , n40298 );
xnor ( n40300 , n40139 , n40141 );
and ( n40301 , n39200 , n34352 );
and ( n40302 , n38979 , n34350 );
nor ( n40303 , n40301 , n40302 );
xnor ( n40304 , n40303 , n28532 );
xor ( n40305 , n39959 , n39960 );
xor ( n40306 , n40305 , n39962 );
and ( n40307 , n40304 , n40306 );
xor ( n40308 , n40097 , n40098 );
xor ( n40309 , n40308 , n40101 );
and ( n40310 , n40306 , n40309 );
and ( n40311 , n40304 , n40309 );
or ( n40312 , n40307 , n40310 , n40311 );
and ( n40313 , n40300 , n40312 );
and ( n40314 , n25220 , n39713 );
and ( n40315 , n24993 , n40196 );
and ( n40316 , n40314 , n40315 );
and ( n40317 , n26399 , n36229 );
and ( n40318 , n40316 , n40317 );
and ( n40319 , n26148 , n36690 );
and ( n40320 , n40317 , n40319 );
and ( n40321 , n40316 , n40319 );
or ( n40322 , n40318 , n40320 , n40321 );
and ( n40323 , n28129 , n26376 );
and ( n40324 , n40322 , n40323 );
and ( n40325 , n27591 , n27558 );
and ( n40326 , n40323 , n40325 );
and ( n40327 , n40322 , n40325 );
or ( n40328 , n40324 , n40326 , n40327 );
and ( n40329 , n27389 , n33739 );
and ( n40330 , n26980 , n34122 );
and ( n40331 , n40329 , n40330 );
and ( n40332 , n26933 , n34817 );
and ( n40333 , n40330 , n40332 );
and ( n40334 , n40329 , n40332 );
or ( n40335 , n40331 , n40333 , n40334 );
and ( n40336 , n27591 , n28209 );
and ( n40337 , n26678 , n35544 );
and ( n40338 , n40336 , n40337 );
xor ( n40339 , n40085 , n40086 );
xor ( n40340 , n40339 , n40088 );
and ( n40341 , n40337 , n40340 );
and ( n40342 , n40336 , n40340 );
or ( n40343 , n40338 , n40341 , n40342 );
and ( n40344 , n40335 , n40343 );
xor ( n40345 , n39953 , n39954 );
xor ( n40346 , n40345 , n39956 );
and ( n40347 , n40343 , n40346 );
and ( n40348 , n40335 , n40346 );
or ( n40349 , n40344 , n40347 , n40348 );
and ( n40350 , n40328 , n40349 );
xor ( n40351 , n40091 , n40092 );
xor ( n40352 , n40351 , n40094 );
xor ( n40353 , n40156 , n40157 );
xor ( n40354 , n40353 , n40159 );
and ( n40355 , n40352 , n40354 );
and ( n40356 , n39200 , n34911 );
and ( n40357 , n38979 , n34909 );
nor ( n40358 , n40356 , n40357 );
xnor ( n40359 , n40358 , n34104 );
xnor ( n40360 , n40174 , n40179 );
and ( n40361 , n40359 , n40360 );
and ( n40362 , n27863 , n28209 );
and ( n40363 , n27591 , n33739 );
and ( n40364 , n40362 , n40363 );
and ( n40365 , n27389 , n34122 );
and ( n40366 , n40363 , n40365 );
and ( n40367 , n40362 , n40365 );
or ( n40368 , n40364 , n40366 , n40367 );
and ( n40369 , n40360 , n40368 );
and ( n40370 , n40359 , n40368 );
or ( n40371 , n40361 , n40369 , n40370 );
and ( n40372 , n40354 , n40371 );
and ( n40373 , n40352 , n40371 );
or ( n40374 , n40355 , n40372 , n40373 );
and ( n40375 , n40349 , n40374 );
and ( n40376 , n40328 , n40374 );
or ( n40377 , n40350 , n40375 , n40376 );
and ( n40378 , n40312 , n40377 );
and ( n40379 , n40300 , n40377 );
or ( n40380 , n40313 , n40378 , n40379 );
and ( n40381 , n40299 , n40380 );
and ( n40382 , n26980 , n34817 );
and ( n40383 , n26933 , n35169 );
and ( n40384 , n40382 , n40383 );
and ( n40385 , n26782 , n35544 );
and ( n40386 , n40383 , n40385 );
and ( n40387 , n40382 , n40385 );
or ( n40388 , n40384 , n40386 , n40387 );
and ( n40389 , n25623 , n38737 );
and ( n40390 , n25451 , n39261 );
and ( n40391 , n40389 , n40390 );
and ( n40392 , n37151 , n37197 );
and ( n40393 , n36427 , n37194 );
nor ( n40394 , n40392 , n40393 );
xnor ( n40395 , n40394 , n36218 );
and ( n40396 , n40390 , n40395 );
and ( n40397 , n40389 , n40395 );
or ( n40398 , n40391 , n40396 , n40397 );
and ( n40399 , n40388 , n40398 );
and ( n40400 , n37387 , n36910 );
and ( n40401 , n37159 , n36908 );
nor ( n40402 , n40400 , n40401 );
xnor ( n40403 , n40402 , n36221 );
and ( n40404 , n38359 , n36367 );
and ( n40405 , n38142 , n36365 );
nor ( n40406 , n40404 , n40405 );
xnor ( n40407 , n40406 , n35608 );
and ( n40408 , n40403 , n40407 );
and ( n40409 , n38462 , n35911 );
and ( n40410 , n38003 , n35909 );
nor ( n40411 , n40409 , n40410 );
xnor ( n40412 , n40411 , n35161 );
and ( n40413 , n40407 , n40412 );
and ( n40414 , n40403 , n40412 );
or ( n40415 , n40408 , n40413 , n40414 );
and ( n40416 , n40398 , n40415 );
and ( n40417 , n40388 , n40415 );
or ( n40418 , n40399 , n40416 , n40417 );
and ( n40419 , n38979 , n35374 );
and ( n40420 , n38777 , n35372 );
nor ( n40421 , n40419 , n40420 );
xnor ( n40422 , n40421 , n34661 );
and ( n40423 , n39500 , n34911 );
and ( n40424 , n39200 , n34909 );
nor ( n40425 , n40423 , n40424 );
xnor ( n40426 , n40425 , n34104 );
and ( n40427 , n40422 , n40426 );
and ( n40428 , n40178 , n33632 );
and ( n40429 , n40172 , n33630 );
nor ( n40430 , n40428 , n40429 );
xnor ( n40431 , n40430 , n28124 );
and ( n40432 , n40426 , n40431 );
and ( n40433 , n40422 , n40431 );
or ( n40434 , n40427 , n40432 , n40433 );
xor ( n40435 , n40182 , n40183 );
xor ( n40436 , n40435 , n40185 );
and ( n40437 , n40434 , n40436 );
xor ( n40438 , n40192 , n40193 );
xor ( n40439 , n40438 , n40197 );
and ( n40440 , n40436 , n40439 );
and ( n40441 , n40434 , n40439 );
or ( n40442 , n40437 , n40440 , n40441 );
and ( n40443 , n40418 , n40442 );
xor ( n40444 , n40173 , n40180 );
xor ( n40445 , n40444 , n40188 );
and ( n40446 , n40442 , n40445 );
and ( n40447 , n40418 , n40445 );
or ( n40448 , n40443 , n40446 , n40447 );
xor ( n40449 , n40152 , n40154 );
xor ( n40450 , n40449 , n40162 );
and ( n40451 , n40448 , n40450 );
xor ( n40452 , n40191 , n40219 );
xor ( n40453 , n40452 , n40230 );
and ( n40454 , n40450 , n40453 );
and ( n40455 , n40448 , n40453 );
or ( n40456 , n40451 , n40454 , n40455 );
xor ( n40457 , n40147 , n40149 );
xor ( n40458 , n40457 , n40165 );
and ( n40459 , n40456 , n40458 );
xor ( n40460 , n40233 , n40243 );
xor ( n40461 , n40460 , n40246 );
and ( n40462 , n40458 , n40461 );
and ( n40463 , n40456 , n40461 );
or ( n40464 , n40459 , n40462 , n40463 );
and ( n40465 , n40380 , n40464 );
and ( n40466 , n40299 , n40464 );
or ( n40467 , n40381 , n40465 , n40466 );
and ( n40468 , n40289 , n40467 );
and ( n40469 , n40279 , n40467 );
or ( n40470 , n40290 , n40468 , n40469 );
and ( n40471 , n40276 , n40470 );
and ( n40472 , n40274 , n40470 );
or ( n40473 , n40277 , n40471 , n40472 );
and ( n40474 , n40272 , n40473 );
xor ( n40475 , n40074 , n40076 );
xor ( n40476 , n40475 , n40264 );
and ( n40477 , n40473 , n40476 );
and ( n40478 , n40272 , n40476 );
or ( n40479 , n40474 , n40477 , n40478 );
and ( n40480 , n40269 , n40479 );
and ( n40481 , n40267 , n40479 );
or ( n40482 , n40270 , n40480 , n40481 );
and ( n40483 , n40071 , n40482 );
and ( n40484 , n40069 , n40482 );
or ( n40485 , n40072 , n40483 , n40484 );
and ( n40486 , n39841 , n40485 );
and ( n40487 , n39839 , n40485 );
or ( n40488 , n39842 , n40486 , n40487 );
or ( n40489 , n39637 , n40488 );
and ( n40490 , n39634 , n40489 );
and ( n40491 , n39632 , n40489 );
or ( n40492 , n39635 , n40490 , n40491 );
and ( n40493 , n39420 , n40492 );
xor ( n40494 , n39420 , n40492 );
xor ( n40495 , n39632 , n39634 );
xor ( n40496 , n40495 , n40489 );
not ( n40497 , n40496 );
xnor ( n40498 , n39637 , n40488 );
xor ( n40499 , n39839 , n39841 );
xor ( n40500 , n40499 , n40485 );
xor ( n40501 , n40069 , n40071 );
xor ( n40502 , n40501 , n40482 );
not ( n40503 , n40502 );
xor ( n40504 , n40267 , n40269 );
xor ( n40505 , n40504 , n40479 );
xor ( n40506 , n40079 , n40127 );
xor ( n40507 , n40506 , n40261 );
xor ( n40508 , n40081 , n40083 );
xor ( n40509 , n40508 , n40124 );
xor ( n40510 , n40145 , n40255 );
xor ( n40511 , n40510 , n40258 );
and ( n40512 , n40509 , n40511 );
xor ( n40513 , n40130 , n40134 );
xor ( n40514 , n40513 , n40142 );
xor ( n40515 , n40168 , n40249 );
xor ( n40516 , n40515 , n40252 );
and ( n40517 , n40514 , n40516 );
and ( n40518 , n38462 , n35374 );
and ( n40519 , n38003 , n35372 );
nor ( n40520 , n40518 , n40519 );
xnor ( n40521 , n40520 , n34661 );
and ( n40522 , n38979 , n34911 );
and ( n40523 , n38777 , n34909 );
nor ( n40524 , n40522 , n40523 );
xnor ( n40525 , n40524 , n34104 );
and ( n40526 , n40521 , n40525 );
xor ( n40527 , n40335 , n40343 );
xor ( n40528 , n40527 , n40346 );
and ( n40529 , n40525 , n40528 );
and ( n40530 , n40521 , n40528 );
or ( n40531 , n40526 , n40529 , n40530 );
xor ( n40532 , n40304 , n40306 );
xor ( n40533 , n40532 , n40309 );
and ( n40534 , n40531 , n40533 );
xor ( n40535 , n40235 , n40237 );
xor ( n40536 , n40535 , n40240 );
and ( n40537 , n39768 , n33632 );
and ( n40538 , n39759 , n33630 );
nor ( n40539 , n40537 , n40538 );
xnor ( n40540 , n40539 , n28124 );
xor ( n40541 , n40322 , n40323 );
xor ( n40542 , n40541 , n40325 );
and ( n40543 , n40540 , n40542 );
and ( n40544 , n40536 , n40543 );
xor ( n40545 , n40200 , n40213 );
xor ( n40546 , n40545 , n40216 );
xor ( n40547 , n40222 , n40224 );
xor ( n40548 , n40547 , n40227 );
and ( n40549 , n40546 , n40548 );
and ( n40550 , n26678 , n36229 );
and ( n40551 , n26399 , n36690 );
and ( n40552 , n40550 , n40551 );
and ( n40553 , n25959 , n37626 );
and ( n40554 , n40551 , n40553 );
and ( n40555 , n40550 , n40553 );
or ( n40556 , n40552 , n40554 , n40555 );
xor ( n40557 , n40314 , n40315 );
and ( n40558 , n26148 , n37187 );
and ( n40559 , n40557 , n40558 );
and ( n40560 , n25742 , n38204 );
and ( n40561 , n40558 , n40560 );
and ( n40562 , n40557 , n40560 );
or ( n40563 , n40559 , n40561 , n40562 );
and ( n40564 , n40556 , n40563 );
and ( n40565 , n27863 , n27558 );
and ( n40566 , n40563 , n40565 );
and ( n40567 , n40556 , n40565 );
or ( n40568 , n40564 , n40566 , n40567 );
and ( n40569 , n40548 , n40568 );
and ( n40570 , n40546 , n40568 );
or ( n40571 , n40549 , n40569 , n40570 );
and ( n40572 , n40543 , n40571 );
and ( n40573 , n40536 , n40571 );
or ( n40574 , n40544 , n40572 , n40573 );
and ( n40575 , n40534 , n40574 );
and ( n40576 , n26399 , n37187 );
and ( n40577 , n26148 , n37626 );
and ( n40578 , n40576 , n40577 );
and ( n40579 , n25959 , n38204 );
and ( n40580 , n40577 , n40579 );
and ( n40581 , n40576 , n40579 );
or ( n40582 , n40578 , n40580 , n40581 );
xor ( n40583 , n32981 , n33578 );
buf ( n40584 , n40583 );
buf ( n40585 , n40584 );
buf ( n40586 , n40585 );
and ( n40587 , n40586 , n28117 );
and ( n40588 , n40582 , n40587 );
xor ( n40589 , n40550 , n40551 );
xor ( n40590 , n40589 , n40553 );
and ( n40591 , n40587 , n40590 );
and ( n40592 , n40582 , n40590 );
or ( n40593 , n40588 , n40591 , n40592 );
xor ( n40594 , n40329 , n40330 );
xor ( n40595 , n40594 , n40332 );
and ( n40596 , n40593 , n40595 );
xor ( n40597 , n40336 , n40337 );
xor ( n40598 , n40597 , n40340 );
and ( n40599 , n40595 , n40598 );
and ( n40600 , n40593 , n40598 );
or ( n40601 , n40596 , n40599 , n40600 );
xor ( n40602 , n40201 , n40205 );
xor ( n40603 , n40602 , n40210 );
xor ( n40604 , n40316 , n40317 );
xor ( n40605 , n40604 , n40319 );
and ( n40606 , n40603 , n40605 );
xor ( n40607 , n40362 , n40363 );
xor ( n40608 , n40607 , n40365 );
and ( n40609 , n26980 , n35169 );
and ( n40610 , n26782 , n36229 );
and ( n40611 , n40609 , n40610 );
and ( n40612 , n26678 , n36690 );
and ( n40613 , n40610 , n40612 );
and ( n40614 , n40609 , n40612 );
or ( n40615 , n40611 , n40613 , n40614 );
and ( n40616 , n40608 , n40615 );
and ( n40617 , n27591 , n34122 );
and ( n40618 , n27389 , n34817 );
and ( n40619 , n40617 , n40618 );
xor ( n40620 , n33040 , n33576 );
buf ( n40621 , n40620 );
buf ( n40622 , n40621 );
buf ( n40623 , n40622 );
and ( n40624 , n40623 , n28117 );
and ( n40625 , n40618 , n40624 );
and ( n40626 , n40617 , n40624 );
or ( n40627 , n40619 , n40625 , n40626 );
and ( n40628 , n40615 , n40627 );
and ( n40629 , n40608 , n40627 );
or ( n40630 , n40616 , n40628 , n40629 );
and ( n40631 , n40605 , n40630 );
and ( n40632 , n40603 , n40630 );
or ( n40633 , n40606 , n40631 , n40632 );
and ( n40634 , n40601 , n40633 );
and ( n40635 , n27863 , n33739 );
and ( n40636 , n25451 , n39713 );
and ( n40637 , n40635 , n40636 );
and ( n40638 , n25220 , n40196 );
and ( n40639 , n40636 , n40638 );
and ( n40640 , n40635 , n40638 );
or ( n40641 , n40637 , n40639 , n40640 );
buf ( n40642 , n15019 );
buf ( n40643 , n40642 );
and ( n40644 , n24993 , n40643 );
buf ( n40645 , n24731 );
and ( n40646 , n40644 , n40645 );
and ( n40647 , n37159 , n37197 );
and ( n40648 , n37151 , n37194 );
nor ( n40649 , n40647 , n40648 );
xnor ( n40650 , n40649 , n36218 );
and ( n40651 , n40645 , n40650 );
and ( n40652 , n40644 , n40650 );
or ( n40653 , n40646 , n40651 , n40652 );
and ( n40654 , n40641 , n40653 );
and ( n40655 , n38142 , n36910 );
and ( n40656 , n37387 , n36908 );
nor ( n40657 , n40655 , n40656 );
xnor ( n40658 , n40657 , n36221 );
and ( n40659 , n39759 , n34911 );
and ( n40660 , n39500 , n34909 );
nor ( n40661 , n40659 , n40660 );
xnor ( n40662 , n40661 , n34104 );
and ( n40663 , n40658 , n40662 );
and ( n40664 , n40172 , n34352 );
and ( n40665 , n39768 , n34350 );
nor ( n40666 , n40664 , n40665 );
xnor ( n40667 , n40666 , n28532 );
and ( n40668 , n40662 , n40667 );
and ( n40669 , n40658 , n40667 );
or ( n40670 , n40663 , n40668 , n40669 );
and ( n40671 , n40653 , n40670 );
and ( n40672 , n40641 , n40670 );
or ( n40673 , n40654 , n40671 , n40672 );
xor ( n40674 , n40382 , n40383 );
xor ( n40675 , n40674 , n40385 );
xor ( n40676 , n40389 , n40390 );
xor ( n40677 , n40676 , n40395 );
and ( n40678 , n40675 , n40677 );
xor ( n40679 , n40403 , n40407 );
xor ( n40680 , n40679 , n40412 );
and ( n40681 , n40677 , n40680 );
and ( n40682 , n40675 , n40680 );
or ( n40683 , n40678 , n40681 , n40682 );
and ( n40684 , n40673 , n40683 );
xor ( n40685 , n40359 , n40360 );
xor ( n40686 , n40685 , n40368 );
and ( n40687 , n40683 , n40686 );
and ( n40688 , n40673 , n40686 );
or ( n40689 , n40684 , n40687 , n40688 );
and ( n40690 , n40633 , n40689 );
and ( n40691 , n40601 , n40689 );
or ( n40692 , n40634 , n40690 , n40691 );
xor ( n40693 , n40328 , n40349 );
xor ( n40694 , n40693 , n40374 );
and ( n40695 , n40692 , n40694 );
xor ( n40696 , n40448 , n40450 );
xor ( n40697 , n40696 , n40453 );
and ( n40698 , n40694 , n40697 );
and ( n40699 , n40692 , n40697 );
or ( n40700 , n40695 , n40698 , n40699 );
and ( n40701 , n40574 , n40700 );
and ( n40702 , n40534 , n40700 );
or ( n40703 , n40575 , n40701 , n40702 );
and ( n40704 , n40516 , n40703 );
and ( n40705 , n40514 , n40703 );
or ( n40706 , n40517 , n40704 , n40705 );
and ( n40707 , n40511 , n40706 );
and ( n40708 , n40509 , n40706 );
or ( n40709 , n40512 , n40707 , n40708 );
and ( n40710 , n40507 , n40709 );
xor ( n40711 , n40274 , n40276 );
xor ( n40712 , n40711 , n40470 );
and ( n40713 , n40709 , n40712 );
and ( n40714 , n40507 , n40712 );
or ( n40715 , n40710 , n40713 , n40714 );
xor ( n40716 , n40272 , n40473 );
xor ( n40717 , n40716 , n40476 );
and ( n40718 , n40715 , n40717 );
xor ( n40719 , n40292 , n40294 );
xor ( n40720 , n40719 , n40296 );
xor ( n40721 , n40300 , n40312 );
xor ( n40722 , n40721 , n40377 );
and ( n40723 , n40720 , n40722 );
xor ( n40724 , n40456 , n40458 );
xor ( n40725 , n40724 , n40461 );
and ( n40726 , n40722 , n40725 );
and ( n40727 , n40720 , n40725 );
or ( n40728 , n40723 , n40726 , n40727 );
xor ( n40729 , n40281 , n40283 );
xor ( n40730 , n40729 , n40286 );
and ( n40731 , n40728 , n40730 );
xor ( n40732 , n40299 , n40380 );
xor ( n40733 , n40732 , n40464 );
and ( n40734 , n40730 , n40733 );
and ( n40735 , n40728 , n40733 );
or ( n40736 , n40731 , n40734 , n40735 );
xor ( n40737 , n40279 , n40289 );
xor ( n40738 , n40737 , n40467 );
and ( n40739 , n40736 , n40738 );
xor ( n40740 , n40531 , n40533 );
xor ( n40741 , n40352 , n40354 );
xor ( n40742 , n40741 , n40371 );
xor ( n40743 , n40418 , n40442 );
xor ( n40744 , n40743 , n40445 );
and ( n40745 , n40742 , n40744 );
xor ( n40746 , n40521 , n40525 );
xor ( n40747 , n40746 , n40528 );
and ( n40748 , n40744 , n40747 );
and ( n40749 , n40742 , n40747 );
or ( n40750 , n40745 , n40748 , n40749 );
and ( n40751 , n40740 , n40750 );
xor ( n40752 , n40540 , n40542 );
and ( n40753 , n28129 , n27246 );
and ( n40754 , n27962 , n27558 );
and ( n40755 , n40753 , n40754 );
xor ( n40756 , n40557 , n40558 );
xor ( n40757 , n40756 , n40560 );
and ( n40758 , n40754 , n40757 );
and ( n40759 , n40753 , n40757 );
or ( n40760 , n40755 , n40758 , n40759 );
and ( n40761 , n39759 , n34352 );
and ( n40762 , n39500 , n34350 );
nor ( n40763 , n40761 , n40762 );
xnor ( n40764 , n40763 , n28532 );
and ( n40765 , n40760 , n40764 );
and ( n40766 , n40172 , n33632 );
and ( n40767 , n39768 , n33630 );
nor ( n40768 , n40766 , n40767 );
xnor ( n40769 , n40768 , n28124 );
and ( n40770 , n40764 , n40769 );
and ( n40771 , n40760 , n40769 );
or ( n40772 , n40765 , n40770 , n40771 );
and ( n40773 , n40752 , n40772 );
xor ( n40774 , n40388 , n40398 );
xor ( n40775 , n40774 , n40415 );
xor ( n40776 , n40434 , n40436 );
xor ( n40777 , n40776 , n40439 );
and ( n40778 , n40775 , n40777 );
xor ( n40779 , n40556 , n40563 );
xor ( n40780 , n40779 , n40565 );
and ( n40781 , n40777 , n40780 );
and ( n40782 , n40775 , n40780 );
or ( n40783 , n40778 , n40781 , n40782 );
and ( n40784 , n40772 , n40783 );
and ( n40785 , n40752 , n40783 );
or ( n40786 , n40773 , n40784 , n40785 );
and ( n40787 , n40750 , n40786 );
and ( n40788 , n40740 , n40786 );
or ( n40789 , n40751 , n40787 , n40788 );
xor ( n40790 , n40422 , n40426 );
xor ( n40791 , n40790 , n40431 );
and ( n40792 , n25451 , n40196 );
and ( n40793 , n25220 , n40643 );
and ( n40794 , n40792 , n40793 );
and ( n40795 , n25742 , n38737 );
and ( n40796 , n40794 , n40795 );
and ( n40797 , n25623 , n39261 );
and ( n40798 , n40795 , n40797 );
and ( n40799 , n40794 , n40797 );
or ( n40800 , n40796 , n40798 , n40799 );
and ( n40801 , n40791 , n40800 );
and ( n40802 , n40586 , n33632 );
and ( n40803 , n40178 , n33630 );
nor ( n40804 , n40802 , n40803 );
xnor ( n40805 , n40804 , n28124 );
xor ( n40806 , n40617 , n40618 );
xor ( n40807 , n40806 , n40624 );
and ( n40808 , n40805 , n40807 );
and ( n40809 , n27962 , n33739 );
and ( n40810 , n26933 , n36229 );
and ( n40811 , n40809 , n40810 );
and ( n40812 , n26782 , n36690 );
and ( n40813 , n40810 , n40812 );
and ( n40814 , n40809 , n40812 );
or ( n40815 , n40811 , n40813 , n40814 );
and ( n40816 , n40807 , n40815 );
and ( n40817 , n40805 , n40815 );
or ( n40818 , n40808 , n40816 , n40817 );
and ( n40819 , n40800 , n40818 );
and ( n40820 , n40791 , n40818 );
or ( n40821 , n40801 , n40819 , n40820 );
and ( n40822 , n26399 , n37626 );
and ( n40823 , n26148 , n38204 );
and ( n40824 , n40822 , n40823 );
and ( n40825 , n25742 , n39261 );
and ( n40826 , n40823 , n40825 );
and ( n40827 , n40822 , n40825 );
or ( n40828 , n40824 , n40826 , n40827 );
and ( n40829 , n25623 , n39713 );
and ( n40830 , n37387 , n37197 );
and ( n40831 , n37159 , n37194 );
nor ( n40832 , n40830 , n40831 );
xnor ( n40833 , n40832 , n36218 );
and ( n40834 , n40829 , n40833 );
and ( n40835 , n38359 , n36910 );
and ( n40836 , n38142 , n36908 );
nor ( n40837 , n40835 , n40836 );
xnor ( n40838 , n40837 , n36221 );
and ( n40839 , n40833 , n40838 );
and ( n40840 , n40829 , n40838 );
or ( n40841 , n40834 , n40839 , n40840 );
and ( n40842 , n40828 , n40841 );
and ( n40843 , n38462 , n36367 );
and ( n40844 , n38003 , n36365 );
nor ( n40845 , n40843 , n40844 );
xnor ( n40846 , n40845 , n35608 );
and ( n40847 , n38979 , n35911 );
and ( n40848 , n38777 , n35909 );
nor ( n40849 , n40847 , n40848 );
xnor ( n40850 , n40849 , n35161 );
and ( n40851 , n40846 , n40850 );
and ( n40852 , n39500 , n35374 );
and ( n40853 , n39200 , n35372 );
nor ( n40854 , n40852 , n40853 );
xnor ( n40855 , n40854 , n34661 );
and ( n40856 , n40850 , n40855 );
and ( n40857 , n40846 , n40855 );
or ( n40858 , n40851 , n40856 , n40857 );
and ( n40859 , n40841 , n40858 );
and ( n40860 , n40828 , n40858 );
or ( n40861 , n40842 , n40859 , n40860 );
xor ( n40862 , n40635 , n40636 );
xor ( n40863 , n40862 , n40638 );
xor ( n40864 , n40644 , n40645 );
xor ( n40865 , n40864 , n40650 );
and ( n40866 , n40863 , n40865 );
xor ( n40867 , n40658 , n40662 );
xor ( n40868 , n40867 , n40667 );
and ( n40869 , n40865 , n40868 );
and ( n40870 , n40863 , n40868 );
or ( n40871 , n40866 , n40869 , n40870 );
and ( n40872 , n40861 , n40871 );
xor ( n40873 , n40608 , n40615 );
xor ( n40874 , n40873 , n40627 );
and ( n40875 , n40871 , n40874 );
and ( n40876 , n40861 , n40874 );
or ( n40877 , n40872 , n40875 , n40876 );
and ( n40878 , n40821 , n40877 );
xor ( n40879 , n40603 , n40605 );
xor ( n40880 , n40879 , n40630 );
and ( n40881 , n40877 , n40880 );
and ( n40882 , n40821 , n40880 );
or ( n40883 , n40878 , n40881 , n40882 );
xor ( n40884 , n40546 , n40548 );
xor ( n40885 , n40884 , n40568 );
and ( n40886 , n40883 , n40885 );
xor ( n40887 , n40601 , n40633 );
xor ( n40888 , n40887 , n40689 );
and ( n40889 , n40885 , n40888 );
and ( n40890 , n40883 , n40888 );
or ( n40891 , n40886 , n40889 , n40890 );
xor ( n40892 , n40536 , n40543 );
xor ( n40893 , n40892 , n40571 );
and ( n40894 , n40891 , n40893 );
xor ( n40895 , n40692 , n40694 );
xor ( n40896 , n40895 , n40697 );
and ( n40897 , n40893 , n40896 );
and ( n40898 , n40891 , n40896 );
or ( n40899 , n40894 , n40897 , n40898 );
and ( n40900 , n40789 , n40899 );
xor ( n40901 , n40534 , n40574 );
xor ( n40902 , n40901 , n40700 );
and ( n40903 , n40899 , n40902 );
and ( n40904 , n40789 , n40902 );
or ( n40905 , n40900 , n40903 , n40904 );
xor ( n40906 , n40514 , n40516 );
xor ( n40907 , n40906 , n40703 );
and ( n40908 , n40905 , n40907 );
xor ( n40909 , n40728 , n40730 );
xor ( n40910 , n40909 , n40733 );
and ( n40911 , n40907 , n40910 );
and ( n40912 , n40905 , n40910 );
or ( n40913 , n40908 , n40911 , n40912 );
and ( n40914 , n40738 , n40913 );
and ( n40915 , n40736 , n40913 );
or ( n40916 , n40739 , n40914 , n40915 );
xor ( n40917 , n40507 , n40709 );
xor ( n40918 , n40917 , n40712 );
and ( n40919 , n40916 , n40918 );
xor ( n40920 , n40509 , n40511 );
xor ( n40921 , n40920 , n40706 );
xor ( n40922 , n40736 , n40738 );
xor ( n40923 , n40922 , n40913 );
and ( n40924 , n40921 , n40923 );
xor ( n40925 , n40720 , n40722 );
xor ( n40926 , n40925 , n40725 );
and ( n40927 , n39768 , n34352 );
and ( n40928 , n39759 , n34350 );
nor ( n40929 , n40927 , n40928 );
xnor ( n40930 , n40929 , n28532 );
xor ( n40931 , n40582 , n40587 );
xor ( n40932 , n40931 , n40590 );
and ( n40933 , n40930 , n40932 );
xor ( n40934 , n40753 , n40754 );
xor ( n40935 , n40934 , n40757 );
and ( n40936 , n40932 , n40935 );
and ( n40937 , n40930 , n40935 );
or ( n40938 , n40933 , n40936 , n40937 );
and ( n40939 , n37159 , n36910 );
and ( n40940 , n37151 , n36908 );
nor ( n40941 , n40939 , n40940 );
xnor ( n40942 , n40941 , n36221 );
and ( n40943 , n40938 , n40942 );
and ( n40944 , n38142 , n36367 );
and ( n40945 , n37387 , n36365 );
nor ( n40946 , n40944 , n40945 );
xnor ( n40947 , n40946 , n35608 );
and ( n40948 , n40942 , n40947 );
and ( n40949 , n40938 , n40947 );
or ( n40950 , n40943 , n40948 , n40949 );
and ( n40951 , n38003 , n35911 );
and ( n40952 , n38359 , n35909 );
nor ( n40953 , n40951 , n40952 );
xnor ( n40954 , n40953 , n35161 );
xor ( n40955 , n40760 , n40764 );
xor ( n40956 , n40955 , n40769 );
and ( n40957 , n40954 , n40956 );
xor ( n40958 , n40593 , n40595 );
xor ( n40959 , n40958 , n40598 );
and ( n40960 , n40956 , n40959 );
and ( n40961 , n40954 , n40959 );
or ( n40962 , n40957 , n40960 , n40961 );
and ( n40963 , n40950 , n40962 );
xor ( n40964 , n40673 , n40683 );
xor ( n40965 , n40964 , n40686 );
xor ( n40966 , n40641 , n40653 );
xor ( n40967 , n40966 , n40670 );
xor ( n40968 , n40675 , n40677 );
xor ( n40969 , n40968 , n40680 );
and ( n40970 , n40967 , n40969 );
xor ( n40971 , n40792 , n40793 );
and ( n40972 , n26678 , n37187 );
and ( n40973 , n40971 , n40972 );
and ( n40974 , n25959 , n38737 );
and ( n40975 , n40972 , n40974 );
and ( n40976 , n40971 , n40974 );
or ( n40977 , n40973 , n40975 , n40976 );
and ( n40978 , n28129 , n27558 );
and ( n40979 , n40977 , n40978 );
xor ( n40980 , n40576 , n40577 );
xor ( n40981 , n40980 , n40579 );
and ( n40982 , n40978 , n40981 );
and ( n40983 , n40977 , n40981 );
or ( n40984 , n40979 , n40982 , n40983 );
and ( n40985 , n40969 , n40984 );
and ( n40986 , n40967 , n40984 );
or ( n40987 , n40970 , n40985 , n40986 );
and ( n40988 , n40965 , n40987 );
and ( n40989 , n27962 , n28209 );
and ( n40990 , n26933 , n35544 );
and ( n40991 , n40989 , n40990 );
xor ( n40992 , n40794 , n40795 );
xor ( n40993 , n40992 , n40797 );
and ( n40994 , n40990 , n40993 );
and ( n40995 , n40989 , n40993 );
or ( n40996 , n40991 , n40994 , n40995 );
and ( n40997 , n39768 , n34911 );
and ( n40998 , n39759 , n34909 );
nor ( n40999 , n40997 , n40998 );
xnor ( n41000 , n40999 , n34104 );
and ( n41001 , n40623 , n33632 );
and ( n41002 , n40586 , n33630 );
nor ( n41003 , n41001 , n41002 );
xnor ( n41004 , n41003 , n28124 );
and ( n41005 , n41000 , n41004 );
and ( n41006 , n28129 , n33739 );
and ( n41007 , n27962 , n34122 );
and ( n41008 , n41006 , n41007 );
xor ( n41009 , n33096 , n33574 );
buf ( n41010 , n41009 );
buf ( n41011 , n41010 );
buf ( n41012 , n41011 );
and ( n41013 , n41012 , n33632 );
and ( n41014 , n40623 , n33630 );
nor ( n41015 , n41013 , n41014 );
xnor ( n41016 , n41015 , n28124 );
and ( n41017 , n41007 , n41016 );
and ( n41018 , n41006 , n41016 );
or ( n41019 , n41008 , n41017 , n41018 );
and ( n41020 , n41004 , n41019 );
and ( n41021 , n41000 , n41019 );
or ( n41022 , n41005 , n41020 , n41021 );
and ( n41023 , n27863 , n34817 );
and ( n41024 , n27389 , n35544 );
or ( n41025 , n41023 , n41024 );
and ( n41026 , n26980 , n36229 );
and ( n41027 , n26933 , n36690 );
and ( n41028 , n41026 , n41027 );
and ( n41029 , n26678 , n37626 );
and ( n41030 , n41027 , n41029 );
and ( n41031 , n41026 , n41029 );
or ( n41032 , n41028 , n41030 , n41031 );
and ( n41033 , n41025 , n41032 );
and ( n41034 , n25623 , n40196 );
and ( n41035 , n25451 , n40643 );
and ( n41036 , n41034 , n41035 );
buf ( n41037 , n15236 );
buf ( n41038 , n41037 );
and ( n41039 , n25220 , n41038 );
and ( n41040 , n41035 , n41039 );
and ( n41041 , n41034 , n41039 );
or ( n41042 , n41036 , n41040 , n41041 );
and ( n41043 , n41032 , n41042 );
and ( n41044 , n41025 , n41042 );
or ( n41045 , n41033 , n41043 , n41044 );
and ( n41046 , n41022 , n41045 );
buf ( n41047 , n24993 );
and ( n41048 , n38142 , n37197 );
and ( n41049 , n37387 , n37194 );
nor ( n41050 , n41048 , n41049 );
xnor ( n41051 , n41050 , n36218 );
and ( n41052 , n41047 , n41051 );
and ( n41053 , n38003 , n36910 );
and ( n41054 , n38359 , n36908 );
nor ( n41055 , n41053 , n41054 );
xnor ( n41056 , n41055 , n36221 );
and ( n41057 , n41051 , n41056 );
and ( n41058 , n41047 , n41056 );
or ( n41059 , n41052 , n41057 , n41058 );
and ( n41060 , n38777 , n36367 );
and ( n41061 , n38462 , n36365 );
nor ( n41062 , n41060 , n41061 );
xnor ( n41063 , n41062 , n35608 );
and ( n41064 , n39200 , n35911 );
and ( n41065 , n38979 , n35909 );
nor ( n41066 , n41064 , n41065 );
xnor ( n41067 , n41066 , n35161 );
and ( n41068 , n41063 , n41067 );
and ( n41069 , n39759 , n35374 );
and ( n41070 , n39500 , n35372 );
nor ( n41071 , n41069 , n41070 );
xnor ( n41072 , n41071 , n34661 );
and ( n41073 , n41067 , n41072 );
and ( n41074 , n41063 , n41072 );
or ( n41075 , n41068 , n41073 , n41074 );
and ( n41076 , n41059 , n41075 );
xor ( n41077 , n40809 , n40810 );
xor ( n41078 , n41077 , n40812 );
and ( n41079 , n41075 , n41078 );
and ( n41080 , n41059 , n41078 );
or ( n41081 , n41076 , n41079 , n41080 );
and ( n41082 , n41045 , n41081 );
and ( n41083 , n41022 , n41081 );
or ( n41084 , n41046 , n41082 , n41083 );
and ( n41085 , n40996 , n41084 );
xor ( n41086 , n40822 , n40823 );
xor ( n41087 , n41086 , n40825 );
xor ( n41088 , n40829 , n40833 );
xor ( n41089 , n41088 , n40838 );
and ( n41090 , n41087 , n41089 );
xor ( n41091 , n40846 , n40850 );
xor ( n41092 , n41091 , n40855 );
and ( n41093 , n41089 , n41092 );
and ( n41094 , n41087 , n41092 );
or ( n41095 , n41090 , n41093 , n41094 );
xor ( n41096 , n40805 , n40807 );
xor ( n41097 , n41096 , n40815 );
and ( n41098 , n41095 , n41097 );
xor ( n41099 , n40828 , n40841 );
xor ( n41100 , n41099 , n40858 );
and ( n41101 , n41097 , n41100 );
and ( n41102 , n41095 , n41100 );
or ( n41103 , n41098 , n41101 , n41102 );
and ( n41104 , n41084 , n41103 );
and ( n41105 , n40996 , n41103 );
or ( n41106 , n41085 , n41104 , n41105 );
and ( n41107 , n40987 , n41106 );
and ( n41108 , n40965 , n41106 );
or ( n41109 , n40988 , n41107 , n41108 );
and ( n41110 , n40962 , n41109 );
and ( n41111 , n40950 , n41109 );
or ( n41112 , n40963 , n41110 , n41111 );
xor ( n41113 , n40742 , n40744 );
xor ( n41114 , n41113 , n40747 );
xor ( n41115 , n40752 , n40772 );
xor ( n41116 , n41115 , n40783 );
and ( n41117 , n41114 , n41116 );
xor ( n41118 , n40883 , n40885 );
xor ( n41119 , n41118 , n40888 );
and ( n41120 , n41116 , n41119 );
and ( n41121 , n41114 , n41119 );
or ( n41122 , n41117 , n41120 , n41121 );
and ( n41123 , n41112 , n41122 );
xor ( n41124 , n40740 , n40750 );
xor ( n41125 , n41124 , n40786 );
and ( n41126 , n41122 , n41125 );
and ( n41127 , n41112 , n41125 );
or ( n41128 , n41123 , n41126 , n41127 );
and ( n41129 , n40926 , n41128 );
xor ( n41130 , n40789 , n40899 );
xor ( n41131 , n41130 , n40902 );
and ( n41132 , n41128 , n41131 );
and ( n41133 , n40926 , n41131 );
or ( n41134 , n41129 , n41132 , n41133 );
xor ( n41135 , n40905 , n40907 );
xor ( n41136 , n41135 , n40910 );
and ( n41137 , n41134 , n41136 );
xor ( n41138 , n40891 , n40893 );
xor ( n41139 , n41138 , n40896 );
xor ( n41140 , n40775 , n40777 );
xor ( n41141 , n41140 , n40780 );
xor ( n41142 , n40821 , n40877 );
xor ( n41143 , n41142 , n40880 );
and ( n41144 , n41141 , n41143 );
xor ( n41145 , n40938 , n40942 );
xor ( n41146 , n41145 , n40947 );
and ( n41147 , n41143 , n41146 );
and ( n41148 , n41141 , n41146 );
or ( n41149 , n41144 , n41147 , n41148 );
xor ( n41150 , n40954 , n40956 );
xor ( n41151 , n41150 , n40959 );
xor ( n41152 , n40791 , n40800 );
xor ( n41153 , n41152 , n40818 );
xor ( n41154 , n40861 , n40871 );
xor ( n41155 , n41154 , n40874 );
and ( n41156 , n41153 , n41155 );
xor ( n41157 , n40930 , n40932 );
xor ( n41158 , n41157 , n40935 );
and ( n41159 , n41155 , n41158 );
and ( n41160 , n41153 , n41158 );
or ( n41161 , n41156 , n41159 , n41160 );
and ( n41162 , n41151 , n41161 );
and ( n41163 , n26782 , n37187 );
and ( n41164 , n26399 , n38204 );
and ( n41165 , n41163 , n41164 );
and ( n41166 , n26148 , n38737 );
and ( n41167 , n41164 , n41166 );
and ( n41168 , n41163 , n41166 );
or ( n41169 , n41165 , n41167 , n41168 );
and ( n41170 , n27863 , n34122 );
and ( n41171 , n41169 , n41170 );
and ( n41172 , n27591 , n34817 );
and ( n41173 , n41170 , n41172 );
and ( n41174 , n41169 , n41172 );
or ( n41175 , n41171 , n41173 , n41174 );
and ( n41176 , n25623 , n40643 );
and ( n41177 , n25451 , n41038 );
and ( n41178 , n41176 , n41177 );
and ( n41179 , n25959 , n39261 );
and ( n41180 , n41178 , n41179 );
and ( n41181 , n25742 , n39713 );
and ( n41182 , n41179 , n41181 );
and ( n41183 , n41178 , n41181 );
or ( n41184 , n41180 , n41182 , n41183 );
and ( n41185 , n28129 , n28209 );
and ( n41186 , n41184 , n41185 );
and ( n41187 , n27389 , n35169 );
and ( n41188 , n41185 , n41187 );
and ( n41189 , n41184 , n41187 );
or ( n41190 , n41186 , n41188 , n41189 );
and ( n41191 , n41175 , n41190 );
xor ( n41192 , n40609 , n40610 );
xor ( n41193 , n41192 , n40612 );
and ( n41194 , n41190 , n41193 );
and ( n41195 , n41175 , n41193 );
or ( n41196 , n41191 , n41194 , n41195 );
and ( n41197 , n38777 , n35911 );
and ( n41198 , n38462 , n35909 );
nor ( n41199 , n41197 , n41198 );
xnor ( n41200 , n41199 , n35161 );
and ( n41201 , n39200 , n35374 );
and ( n41202 , n38979 , n35372 );
nor ( n41203 , n41201 , n41202 );
xnor ( n41204 , n41203 , n34661 );
and ( n41205 , n41200 , n41204 );
xor ( n41206 , n40977 , n40978 );
xor ( n41207 , n41206 , n40981 );
and ( n41208 , n41204 , n41207 );
and ( n41209 , n41200 , n41207 );
or ( n41210 , n41205 , n41208 , n41209 );
and ( n41211 , n41196 , n41210 );
xor ( n41212 , n40863 , n40865 );
xor ( n41213 , n41212 , n40868 );
xor ( n41214 , n40989 , n40990 );
xor ( n41215 , n41214 , n40993 );
and ( n41216 , n41213 , n41215 );
and ( n41217 , n26980 , n35544 );
and ( n41218 , n41012 , n28117 );
and ( n41219 , n41217 , n41218 );
xor ( n41220 , n40971 , n40972 );
xor ( n41221 , n41220 , n40974 );
and ( n41222 , n41218 , n41221 );
and ( n41223 , n41217 , n41221 );
or ( n41224 , n41219 , n41222 , n41223 );
and ( n41225 , n41215 , n41224 );
and ( n41226 , n41213 , n41224 );
or ( n41227 , n41216 , n41225 , n41226 );
and ( n41228 , n41210 , n41227 );
and ( n41229 , n41196 , n41227 );
or ( n41230 , n41211 , n41228 , n41229 );
and ( n41231 , n41161 , n41230 );
and ( n41232 , n41151 , n41230 );
or ( n41233 , n41162 , n41231 , n41232 );
and ( n41234 , n41149 , n41233 );
xor ( n41235 , n40950 , n40962 );
xor ( n41236 , n41235 , n41109 );
and ( n41237 , n41233 , n41236 );
and ( n41238 , n41149 , n41236 );
or ( n41239 , n41234 , n41237 , n41238 );
and ( n41240 , n41139 , n41239 );
xor ( n41241 , n41112 , n41122 );
xor ( n41242 , n41241 , n41125 );
and ( n41243 , n41239 , n41242 );
and ( n41244 , n41139 , n41242 );
or ( n41245 , n41240 , n41243 , n41244 );
xor ( n41246 , n40926 , n41128 );
xor ( n41247 , n41246 , n41131 );
and ( n41248 , n41245 , n41247 );
xor ( n41249 , n41114 , n41116 );
xor ( n41250 , n41249 , n41119 );
and ( n41251 , n40172 , n34911 );
and ( n41252 , n39768 , n34909 );
nor ( n41253 , n41251 , n41252 );
xnor ( n41254 , n41253 , n34104 );
and ( n41255 , n40586 , n34352 );
and ( n41256 , n40178 , n34350 );
nor ( n41257 , n41255 , n41256 );
xnor ( n41258 , n41257 , n28532 );
and ( n41259 , n41254 , n41258 );
xor ( n41260 , n41163 , n41164 );
xor ( n41261 , n41260 , n41166 );
and ( n41262 , n41258 , n41261 );
and ( n41263 , n41254 , n41261 );
or ( n41264 , n41259 , n41262 , n41263 );
xor ( n41265 , n41006 , n41007 );
xor ( n41266 , n41265 , n41016 );
xnor ( n41267 , n41023 , n41024 );
and ( n41268 , n41266 , n41267 );
and ( n41269 , n27389 , n36229 );
and ( n41270 , n26980 , n36690 );
and ( n41271 , n41269 , n41270 );
and ( n41272 , n26782 , n37626 );
and ( n41273 , n41270 , n41272 );
and ( n41274 , n41269 , n41272 );
or ( n41275 , n41271 , n41273 , n41274 );
and ( n41276 , n41267 , n41275 );
and ( n41277 , n41266 , n41275 );
or ( n41278 , n41268 , n41276 , n41277 );
and ( n41279 , n41264 , n41278 );
and ( n41280 , n28129 , n34122 );
and ( n41281 , n26933 , n37187 );
and ( n41282 , n41280 , n41281 );
and ( n41283 , n26678 , n38204 );
and ( n41284 , n41281 , n41283 );
and ( n41285 , n41280 , n41283 );
or ( n41286 , n41282 , n41284 , n41285 );
and ( n41287 , n25959 , n39713 );
and ( n41288 , n25742 , n40196 );
and ( n41289 , n41287 , n41288 );
and ( n41290 , n38359 , n37197 );
and ( n41291 , n38142 , n37194 );
nor ( n41292 , n41290 , n41291 );
xnor ( n41293 , n41292 , n36218 );
and ( n41294 , n41288 , n41293 );
and ( n41295 , n41287 , n41293 );
or ( n41296 , n41289 , n41294 , n41295 );
and ( n41297 , n41286 , n41296 );
and ( n41298 , n38462 , n36910 );
and ( n41299 , n38003 , n36908 );
nor ( n41300 , n41298 , n41299 );
xnor ( n41301 , n41300 , n36221 );
and ( n41302 , n39500 , n35911 );
and ( n41303 , n39200 , n35909 );
nor ( n41304 , n41302 , n41303 );
xnor ( n41305 , n41304 , n35161 );
and ( n41306 , n41301 , n41305 );
and ( n41307 , n39768 , n35374 );
and ( n41308 , n39759 , n35372 );
nor ( n41309 , n41307 , n41308 );
xnor ( n41310 , n41309 , n34661 );
and ( n41311 , n41305 , n41310 );
and ( n41312 , n41301 , n41310 );
or ( n41313 , n41306 , n41311 , n41312 );
and ( n41314 , n41296 , n41313 );
and ( n41315 , n41286 , n41313 );
or ( n41316 , n41297 , n41314 , n41315 );
and ( n41317 , n41278 , n41316 );
and ( n41318 , n41264 , n41316 );
or ( n41319 , n41279 , n41317 , n41318 );
xor ( n41320 , n41026 , n41027 );
xor ( n41321 , n41320 , n41029 );
xor ( n41322 , n41034 , n41035 );
xor ( n41323 , n41322 , n41039 );
and ( n41324 , n41321 , n41323 );
xor ( n41325 , n41047 , n41051 );
xor ( n41326 , n41325 , n41056 );
and ( n41327 , n41323 , n41326 );
and ( n41328 , n41321 , n41326 );
or ( n41329 , n41324 , n41327 , n41328 );
xor ( n41330 , n41000 , n41004 );
xor ( n41331 , n41330 , n41019 );
and ( n41332 , n41329 , n41331 );
xor ( n41333 , n41025 , n41032 );
xor ( n41334 , n41333 , n41042 );
and ( n41335 , n41331 , n41334 );
and ( n41336 , n41329 , n41334 );
or ( n41337 , n41332 , n41335 , n41336 );
and ( n41338 , n41319 , n41337 );
xor ( n41339 , n41022 , n41045 );
xor ( n41340 , n41339 , n41081 );
and ( n41341 , n41337 , n41340 );
and ( n41342 , n41319 , n41340 );
or ( n41343 , n41338 , n41341 , n41342 );
xor ( n41344 , n40967 , n40969 );
xor ( n41345 , n41344 , n40984 );
and ( n41346 , n41343 , n41345 );
xor ( n41347 , n40996 , n41084 );
xor ( n41348 , n41347 , n41103 );
and ( n41349 , n41345 , n41348 );
and ( n41350 , n41343 , n41348 );
or ( n41351 , n41346 , n41349 , n41350 );
xor ( n41352 , n40965 , n40987 );
xor ( n41353 , n41352 , n41106 );
and ( n41354 , n41351 , n41353 );
and ( n41355 , n40178 , n34352 );
and ( n41356 , n40172 , n34350 );
nor ( n41357 , n41355 , n41356 );
xnor ( n41358 , n41357 , n28532 );
xor ( n41359 , n41169 , n41170 );
xor ( n41360 , n41359 , n41172 );
and ( n41361 , n41358 , n41360 );
xor ( n41362 , n41184 , n41185 );
xor ( n41363 , n41362 , n41187 );
and ( n41364 , n41360 , n41363 );
and ( n41365 , n41358 , n41363 );
or ( n41366 , n41361 , n41364 , n41365 );
and ( n41367 , n38003 , n36367 );
and ( n41368 , n38359 , n36365 );
nor ( n41369 , n41367 , n41368 );
xnor ( n41370 , n41369 , n35608 );
and ( n41371 , n41366 , n41370 );
xor ( n41372 , n41095 , n41097 );
xor ( n41373 , n41372 , n41100 );
xor ( n41374 , n41175 , n41190 );
xor ( n41375 , n41374 , n41193 );
and ( n41376 , n41373 , n41375 );
xor ( n41377 , n41200 , n41204 );
xor ( n41378 , n41377 , n41207 );
and ( n41379 , n41375 , n41378 );
and ( n41380 , n41373 , n41378 );
or ( n41381 , n41376 , n41379 , n41380 );
and ( n41382 , n41371 , n41381 );
xor ( n41383 , n41059 , n41075 );
xor ( n41384 , n41383 , n41078 );
xor ( n41385 , n41087 , n41089 );
xor ( n41386 , n41385 , n41092 );
and ( n41387 , n41384 , n41386 );
xor ( n41388 , n41217 , n41218 );
xor ( n41389 , n41388 , n41221 );
and ( n41390 , n41386 , n41389 );
and ( n41391 , n41384 , n41389 );
or ( n41392 , n41387 , n41390 , n41391 );
xor ( n41393 , n41176 , n41177 );
and ( n41394 , n26399 , n38737 );
and ( n41395 , n41393 , n41394 );
and ( n41396 , n26148 , n39261 );
and ( n41397 , n41394 , n41396 );
and ( n41398 , n41393 , n41396 );
or ( n41399 , n41395 , n41397 , n41398 );
and ( n41400 , n27591 , n35169 );
and ( n41401 , n41399 , n41400 );
xor ( n41402 , n33097 , n33573 );
buf ( n41403 , n41402 );
buf ( n41404 , n41403 );
buf ( n41405 , n41404 );
and ( n41406 , n41405 , n28117 );
and ( n41407 , n41400 , n41406 );
and ( n41408 , n41399 , n41406 );
or ( n41409 , n41401 , n41407 , n41408 );
xor ( n41410 , n41063 , n41067 );
xor ( n41411 , n41410 , n41072 );
xor ( n41412 , n41178 , n41179 );
xor ( n41413 , n41412 , n41181 );
and ( n41414 , n41411 , n41413 );
and ( n41415 , n40623 , n34352 );
and ( n41416 , n40586 , n34350 );
nor ( n41417 , n41415 , n41416 );
xnor ( n41418 , n41417 , n28532 );
xor ( n41419 , n41269 , n41270 );
xor ( n41420 , n41419 , n41272 );
and ( n41421 , n41418 , n41420 );
and ( n41422 , n27863 , n35544 );
and ( n41423 , n27591 , n36229 );
and ( n41424 , n41422 , n41423 );
and ( n41425 , n27389 , n36690 );
and ( n41426 , n41423 , n41425 );
and ( n41427 , n41422 , n41425 );
or ( n41428 , n41424 , n41426 , n41427 );
and ( n41429 , n41420 , n41428 );
and ( n41430 , n41418 , n41428 );
or ( n41431 , n41421 , n41429 , n41430 );
and ( n41432 , n41413 , n41431 );
and ( n41433 , n41411 , n41431 );
or ( n41434 , n41414 , n41432 , n41433 );
and ( n41435 , n41409 , n41434 );
and ( n41436 , n26980 , n37187 );
and ( n41437 , n26933 , n37626 );
and ( n41438 , n41436 , n41437 );
and ( n41439 , n25742 , n40643 );
and ( n41440 , n41437 , n41439 );
and ( n41441 , n41436 , n41439 );
or ( n41442 , n41438 , n41440 , n41441 );
and ( n41443 , n25623 , n41038 );
buf ( n41444 , n15630 );
buf ( n41445 , n41444 );
and ( n41446 , n25451 , n41445 );
and ( n41447 , n41443 , n41446 );
buf ( n41448 , n25220 );
and ( n41449 , n41446 , n41448 );
and ( n41450 , n41443 , n41448 );
or ( n41451 , n41447 , n41449 , n41450 );
and ( n41452 , n41442 , n41451 );
and ( n41453 , n38003 , n37197 );
and ( n41454 , n38359 , n37194 );
nor ( n41455 , n41453 , n41454 );
xnor ( n41456 , n41455 , n36218 );
and ( n41457 , n38777 , n36910 );
and ( n41458 , n38462 , n36908 );
nor ( n41459 , n41457 , n41458 );
xnor ( n41460 , n41459 , n36221 );
and ( n41461 , n41456 , n41460 );
and ( n41462 , n39200 , n36367 );
and ( n41463 , n38979 , n36365 );
nor ( n41464 , n41462 , n41463 );
xnor ( n41465 , n41464 , n35608 );
and ( n41466 , n41460 , n41465 );
and ( n41467 , n41456 , n41465 );
or ( n41468 , n41461 , n41466 , n41467 );
and ( n41469 , n41451 , n41468 );
and ( n41470 , n41442 , n41468 );
or ( n41471 , n41452 , n41469 , n41470 );
xor ( n41472 , n41280 , n41281 );
xor ( n41473 , n41472 , n41283 );
xor ( n41474 , n41287 , n41288 );
xor ( n41475 , n41474 , n41293 );
and ( n41476 , n41473 , n41475 );
xor ( n41477 , n41301 , n41305 );
xor ( n41478 , n41477 , n41310 );
and ( n41479 , n41475 , n41478 );
and ( n41480 , n41473 , n41478 );
or ( n41481 , n41476 , n41479 , n41480 );
and ( n41482 , n41471 , n41481 );
xor ( n41483 , n41254 , n41258 );
xor ( n41484 , n41483 , n41261 );
and ( n41485 , n41481 , n41484 );
and ( n41486 , n41471 , n41484 );
or ( n41487 , n41482 , n41485 , n41486 );
and ( n41488 , n41434 , n41487 );
and ( n41489 , n41409 , n41487 );
or ( n41490 , n41435 , n41488 , n41489 );
and ( n41491 , n41392 , n41490 );
xor ( n41492 , n41266 , n41267 );
xor ( n41493 , n41492 , n41275 );
xor ( n41494 , n41286 , n41296 );
xor ( n41495 , n41494 , n41313 );
and ( n41496 , n41493 , n41495 );
xor ( n41497 , n41321 , n41323 );
xor ( n41498 , n41497 , n41326 );
and ( n41499 , n41495 , n41498 );
and ( n41500 , n41493 , n41498 );
or ( n41501 , n41496 , n41499 , n41500 );
xor ( n41502 , n41264 , n41278 );
xor ( n41503 , n41502 , n41316 );
and ( n41504 , n41501 , n41503 );
xor ( n41505 , n41329 , n41331 );
xor ( n41506 , n41505 , n41334 );
and ( n41507 , n41503 , n41506 );
and ( n41508 , n41501 , n41506 );
or ( n41509 , n41504 , n41507 , n41508 );
and ( n41510 , n41490 , n41509 );
and ( n41511 , n41392 , n41509 );
or ( n41512 , n41491 , n41510 , n41511 );
and ( n41513 , n41381 , n41512 );
and ( n41514 , n41371 , n41512 );
or ( n41515 , n41382 , n41513 , n41514 );
and ( n41516 , n41353 , n41515 );
and ( n41517 , n41351 , n41515 );
or ( n41518 , n41354 , n41516 , n41517 );
and ( n41519 , n41250 , n41518 );
xor ( n41520 , n41153 , n41155 );
xor ( n41521 , n41520 , n41158 );
xor ( n41522 , n41196 , n41210 );
xor ( n41523 , n41522 , n41227 );
and ( n41524 , n41521 , n41523 );
xor ( n41525 , n41343 , n41345 );
xor ( n41526 , n41525 , n41348 );
and ( n41527 , n41523 , n41526 );
and ( n41528 , n41521 , n41526 );
or ( n41529 , n41524 , n41527 , n41528 );
xor ( n41530 , n41141 , n41143 );
xor ( n41531 , n41530 , n41146 );
and ( n41532 , n41529 , n41531 );
xor ( n41533 , n41151 , n41161 );
xor ( n41534 , n41533 , n41230 );
and ( n41535 , n41531 , n41534 );
and ( n41536 , n41529 , n41534 );
or ( n41537 , n41532 , n41535 , n41536 );
and ( n41538 , n41518 , n41537 );
and ( n41539 , n41250 , n41537 );
or ( n41540 , n41519 , n41538 , n41539 );
xor ( n41541 , n41139 , n41239 );
xor ( n41542 , n41541 , n41242 );
and ( n41543 , n41540 , n41542 );
xor ( n41544 , n41149 , n41233 );
xor ( n41545 , n41544 , n41236 );
xor ( n41546 , n41213 , n41215 );
xor ( n41547 , n41546 , n41224 );
xor ( n41548 , n41319 , n41337 );
xor ( n41549 , n41548 , n41340 );
and ( n41550 , n41547 , n41549 );
xor ( n41551 , n41366 , n41370 );
and ( n41552 , n41549 , n41551 );
and ( n41553 , n41547 , n41551 );
or ( n41554 , n41550 , n41552 , n41553 );
xor ( n41555 , n41358 , n41360 );
xor ( n41556 , n41555 , n41363 );
and ( n41557 , n26782 , n38204 );
and ( n41558 , n26678 , n38737 );
and ( n41559 , n41557 , n41558 );
and ( n41560 , n26399 , n39261 );
and ( n41561 , n41558 , n41560 );
and ( n41562 , n41557 , n41560 );
or ( n41563 , n41559 , n41561 , n41562 );
and ( n41564 , n27962 , n34817 );
and ( n41565 , n41563 , n41564 );
and ( n41566 , n41405 , n33632 );
and ( n41567 , n41012 , n33630 );
nor ( n41568 , n41566 , n41567 );
xnor ( n41569 , n41568 , n28124 );
and ( n41570 , n41564 , n41569 );
and ( n41571 , n41563 , n41569 );
or ( n41572 , n41565 , n41570 , n41571 );
and ( n41573 , n27863 , n35169 );
and ( n41574 , n27591 , n35544 );
and ( n41575 , n41573 , n41574 );
xor ( n41576 , n41393 , n41394 );
xor ( n41577 , n41576 , n41396 );
and ( n41578 , n41574 , n41577 );
and ( n41579 , n41573 , n41577 );
or ( n41580 , n41575 , n41578 , n41579 );
and ( n41581 , n41572 , n41580 );
xor ( n41582 , n41399 , n41400 );
xor ( n41583 , n41582 , n41406 );
and ( n41584 , n41580 , n41583 );
and ( n41585 , n41572 , n41583 );
or ( n41586 , n41581 , n41584 , n41585 );
and ( n41587 , n41556 , n41586 );
and ( n41588 , n28129 , n34817 );
and ( n41589 , n41012 , n34352 );
and ( n41590 , n40623 , n34350 );
nor ( n41591 , n41589 , n41590 );
xnor ( n41592 , n41591 , n28532 );
and ( n41593 , n41588 , n41592 );
xor ( n41594 , n41557 , n41558 );
xor ( n41595 , n41594 , n41560 );
and ( n41596 , n41592 , n41595 );
and ( n41597 , n41588 , n41595 );
or ( n41598 , n41593 , n41596 , n41597 );
and ( n41599 , n40178 , n34911 );
and ( n41600 , n40172 , n34909 );
nor ( n41601 , n41599 , n41600 );
xnor ( n41602 , n41601 , n34104 );
and ( n41603 , n41598 , n41602 );
xor ( n41604 , n41563 , n41564 );
xor ( n41605 , n41604 , n41569 );
and ( n41606 , n41602 , n41605 );
and ( n41607 , n41598 , n41605 );
or ( n41608 , n41603 , n41606 , n41607 );
and ( n41609 , n25742 , n41038 );
and ( n41610 , n25623 , n41445 );
and ( n41611 , n41609 , n41610 );
and ( n41612 , n26148 , n39713 );
and ( n41613 , n41611 , n41612 );
and ( n41614 , n25959 , n40196 );
and ( n41615 , n41612 , n41614 );
and ( n41616 , n41611 , n41614 );
or ( n41617 , n41613 , n41615 , n41616 );
xor ( n41618 , n33153 , n33571 );
buf ( n41619 , n41618 );
buf ( n41620 , n41619 );
buf ( n41621 , n41620 );
and ( n41622 , n41621 , n28117 );
and ( n41623 , n41617 , n41622 );
and ( n41624 , n41608 , n41623 );
and ( n41625 , n26782 , n38737 );
and ( n41626 , n26678 , n39261 );
and ( n41627 , n41625 , n41626 );
xor ( n41628 , n33252 , n33567 );
buf ( n41629 , n41628 );
buf ( n41630 , n41629 );
buf ( n41631 , n41630 );
and ( n41632 , n41631 , n28117 );
and ( n41633 , n41626 , n41632 );
and ( n41634 , n41625 , n41632 );
or ( n41635 , n41627 , n41633 , n41634 );
and ( n41636 , n27962 , n35169 );
and ( n41637 , n41635 , n41636 );
and ( n41638 , n41621 , n33632 );
and ( n41639 , n41405 , n33630 );
nor ( n41640 , n41638 , n41639 );
xnor ( n41641 , n41640 , n28124 );
and ( n41642 , n41636 , n41641 );
and ( n41643 , n41635 , n41641 );
or ( n41644 , n41637 , n41642 , n41643 );
and ( n41645 , n39759 , n35911 );
and ( n41646 , n39500 , n35909 );
nor ( n41647 , n41645 , n41646 );
xnor ( n41648 , n41647 , n35161 );
xor ( n41649 , n33200 , n33569 );
buf ( n41650 , n41649 );
buf ( n41651 , n41650 );
buf ( n41652 , n41651 );
and ( n41653 , n41652 , n28117 );
and ( n41654 , n41648 , n41653 );
and ( n41655 , n27389 , n37187 );
and ( n41656 , n26933 , n38204 );
and ( n41657 , n41655 , n41656 );
and ( n41658 , n41653 , n41657 );
and ( n41659 , n41648 , n41657 );
or ( n41660 , n41654 , n41658 , n41659 );
and ( n41661 , n41644 , n41660 );
and ( n41662 , n28129 , n35169 );
and ( n41663 , n27863 , n36229 );
and ( n41664 , n41662 , n41663 );
and ( n41665 , n26399 , n39713 );
and ( n41666 , n41663 , n41665 );
and ( n41667 , n41662 , n41665 );
or ( n41668 , n41664 , n41666 , n41667 );
and ( n41669 , n26148 , n40196 );
and ( n41670 , n25959 , n40643 );
and ( n41671 , n41669 , n41670 );
and ( n41672 , n38462 , n37197 );
and ( n41673 , n38003 , n37194 );
nor ( n41674 , n41672 , n41673 );
xnor ( n41675 , n41674 , n36218 );
and ( n41676 , n41670 , n41675 );
and ( n41677 , n41669 , n41675 );
or ( n41678 , n41671 , n41676 , n41677 );
and ( n41679 , n41668 , n41678 );
and ( n41680 , n38979 , n36910 );
and ( n41681 , n38777 , n36908 );
nor ( n41682 , n41680 , n41681 );
xnor ( n41683 , n41682 , n36221 );
and ( n41684 , n39500 , n36367 );
and ( n41685 , n39200 , n36365 );
nor ( n41686 , n41684 , n41685 );
xnor ( n41687 , n41686 , n35608 );
and ( n41688 , n41683 , n41687 );
and ( n41689 , n40178 , n35374 );
and ( n41690 , n40172 , n35372 );
nor ( n41691 , n41689 , n41690 );
xnor ( n41692 , n41691 , n34661 );
and ( n41693 , n41687 , n41692 );
and ( n41694 , n41683 , n41692 );
or ( n41695 , n41688 , n41693 , n41694 );
and ( n41696 , n41678 , n41695 );
and ( n41697 , n41668 , n41695 );
or ( n41698 , n41679 , n41696 , n41697 );
and ( n41699 , n41660 , n41698 );
and ( n41700 , n41644 , n41698 );
or ( n41701 , n41661 , n41699 , n41700 );
and ( n41702 , n41623 , n41701 );
and ( n41703 , n41608 , n41701 );
or ( n41704 , n41624 , n41702 , n41703 );
and ( n41705 , n41586 , n41704 );
and ( n41706 , n41556 , n41704 );
or ( n41707 , n41587 , n41705 , n41706 );
xor ( n41708 , n41422 , n41423 );
xor ( n41709 , n41708 , n41425 );
xor ( n41710 , n41436 , n41437 );
xor ( n41711 , n41710 , n41439 );
and ( n41712 , n41709 , n41711 );
xor ( n41713 , n41443 , n41446 );
xor ( n41714 , n41713 , n41448 );
and ( n41715 , n41711 , n41714 );
and ( n41716 , n41709 , n41714 );
or ( n41717 , n41712 , n41715 , n41716 );
xor ( n41718 , n41418 , n41420 );
xor ( n41719 , n41718 , n41428 );
and ( n41720 , n41717 , n41719 );
xor ( n41721 , n41442 , n41451 );
xor ( n41722 , n41721 , n41468 );
and ( n41723 , n41719 , n41722 );
and ( n41724 , n41717 , n41722 );
or ( n41725 , n41720 , n41723 , n41724 );
xor ( n41726 , n41411 , n41413 );
xor ( n41727 , n41726 , n41431 );
and ( n41728 , n41725 , n41727 );
xor ( n41729 , n41471 , n41481 );
xor ( n41730 , n41729 , n41484 );
and ( n41731 , n41727 , n41730 );
and ( n41732 , n41725 , n41730 );
or ( n41733 , n41728 , n41731 , n41732 );
xor ( n41734 , n41384 , n41386 );
xor ( n41735 , n41734 , n41389 );
and ( n41736 , n41733 , n41735 );
xor ( n41737 , n41409 , n41434 );
xor ( n41738 , n41737 , n41487 );
and ( n41739 , n41735 , n41738 );
and ( n41740 , n41733 , n41738 );
or ( n41741 , n41736 , n41739 , n41740 );
and ( n41742 , n41707 , n41741 );
xor ( n41743 , n41373 , n41375 );
xor ( n41744 , n41743 , n41378 );
and ( n41745 , n41741 , n41744 );
and ( n41746 , n41707 , n41744 );
or ( n41747 , n41742 , n41745 , n41746 );
and ( n41748 , n41554 , n41747 );
xor ( n41749 , n41371 , n41381 );
xor ( n41750 , n41749 , n41512 );
and ( n41751 , n41747 , n41750 );
and ( n41752 , n41554 , n41750 );
or ( n41753 , n41748 , n41751 , n41752 );
xor ( n41754 , n41351 , n41353 );
xor ( n41755 , n41754 , n41515 );
and ( n41756 , n41753 , n41755 );
xor ( n41757 , n41529 , n41531 );
xor ( n41758 , n41757 , n41534 );
and ( n41759 , n41755 , n41758 );
and ( n41760 , n41753 , n41758 );
or ( n41761 , n41756 , n41759 , n41760 );
and ( n41762 , n41545 , n41761 );
xor ( n41763 , n41250 , n41518 );
xor ( n41764 , n41763 , n41537 );
and ( n41765 , n41761 , n41764 );
and ( n41766 , n41545 , n41764 );
or ( n41767 , n41762 , n41765 , n41766 );
and ( n41768 , n41542 , n41767 );
and ( n41769 , n41540 , n41767 );
or ( n41770 , n41543 , n41768 , n41769 );
and ( n41771 , n41247 , n41770 );
and ( n41772 , n41245 , n41770 );
or ( n41773 , n41248 , n41771 , n41772 );
and ( n41774 , n41136 , n41773 );
and ( n41775 , n41134 , n41773 );
or ( n41776 , n41137 , n41774 , n41775 );
and ( n41777 , n40923 , n41776 );
and ( n41778 , n40921 , n41776 );
or ( n41779 , n40924 , n41777 , n41778 );
and ( n41780 , n40918 , n41779 );
and ( n41781 , n40916 , n41779 );
or ( n41782 , n40919 , n41780 , n41781 );
and ( n41783 , n40717 , n41782 );
and ( n41784 , n40715 , n41782 );
or ( n41785 , n40718 , n41783 , n41784 );
and ( n41786 , n40505 , n41785 );
xor ( n41787 , n40505 , n41785 );
xor ( n41788 , n40715 , n40717 );
xor ( n41789 , n41788 , n41782 );
not ( n41790 , n41789 );
xor ( n41791 , n40916 , n40918 );
xor ( n41792 , n41791 , n41779 );
not ( n41793 , n41792 );
xor ( n41794 , n40921 , n40923 );
xor ( n41795 , n41794 , n41776 );
not ( n41796 , n41795 );
xor ( n41797 , n41134 , n41136 );
xor ( n41798 , n41797 , n41773 );
xor ( n41799 , n41245 , n41247 );
xor ( n41800 , n41799 , n41770 );
xor ( n41801 , n41540 , n41542 );
xor ( n41802 , n41801 , n41767 );
xor ( n41803 , n41545 , n41761 );
xor ( n41804 , n41803 , n41764 );
xor ( n41805 , n41521 , n41523 );
xor ( n41806 , n41805 , n41526 );
xor ( n41807 , n41392 , n41490 );
xor ( n41808 , n41807 , n41509 );
xor ( n41809 , n41501 , n41503 );
xor ( n41810 , n41809 , n41506 );
xor ( n41811 , n41493 , n41495 );
xor ( n41812 , n41811 , n41498 );
xor ( n41813 , n41572 , n41580 );
xor ( n41814 , n41813 , n41583 );
and ( n41815 , n41812 , n41814 );
and ( n41816 , n27962 , n35544 );
and ( n41817 , n41405 , n34352 );
and ( n41818 , n41012 , n34350 );
nor ( n41819 , n41817 , n41818 );
xnor ( n41820 , n41819 , n28532 );
and ( n41821 , n41816 , n41820 );
xor ( n41822 , n41625 , n41626 );
xor ( n41823 , n41822 , n41632 );
and ( n41824 , n41820 , n41823 );
and ( n41825 , n41816 , n41823 );
or ( n41826 , n41821 , n41824 , n41825 );
and ( n41827 , n40172 , n35374 );
and ( n41828 , n39768 , n35372 );
nor ( n41829 , n41827 , n41828 );
xnor ( n41830 , n41829 , n34661 );
and ( n41831 , n41826 , n41830 );
xor ( n41832 , n41635 , n41636 );
xor ( n41833 , n41832 , n41641 );
and ( n41834 , n41830 , n41833 );
and ( n41835 , n41826 , n41833 );
or ( n41836 , n41831 , n41834 , n41835 );
and ( n41837 , n38979 , n36367 );
and ( n41838 , n38777 , n36365 );
nor ( n41839 , n41837 , n41838 );
xnor ( n41840 , n41839 , n35608 );
and ( n41841 , n41836 , n41840 );
xor ( n41842 , n41598 , n41602 );
xor ( n41843 , n41842 , n41605 );
and ( n41844 , n41840 , n41843 );
and ( n41845 , n41836 , n41843 );
or ( n41846 , n41841 , n41844 , n41845 );
and ( n41847 , n41814 , n41846 );
and ( n41848 , n41812 , n41846 );
or ( n41849 , n41815 , n41847 , n41848 );
and ( n41850 , n41810 , n41849 );
xor ( n41851 , n41473 , n41475 );
xor ( n41852 , n41851 , n41478 );
xor ( n41853 , n41573 , n41574 );
xor ( n41854 , n41853 , n41577 );
and ( n41855 , n41852 , n41854 );
xor ( n41856 , n41617 , n41622 );
and ( n41857 , n41854 , n41856 );
and ( n41858 , n41852 , n41856 );
or ( n41859 , n41855 , n41857 , n41858 );
xor ( n41860 , n41456 , n41460 );
xor ( n41861 , n41860 , n41465 );
xor ( n41862 , n41611 , n41612 );
xor ( n41863 , n41862 , n41614 );
and ( n41864 , n41861 , n41863 );
xor ( n41865 , n41588 , n41592 );
xor ( n41866 , n41865 , n41595 );
and ( n41867 , n41863 , n41866 );
and ( n41868 , n41861 , n41866 );
or ( n41869 , n41864 , n41867 , n41868 );
and ( n41870 , n40623 , n34911 );
and ( n41871 , n40586 , n34909 );
nor ( n41872 , n41870 , n41871 );
xnor ( n41873 , n41872 , n34104 );
and ( n41874 , n41652 , n33632 );
and ( n41875 , n41621 , n33630 );
nor ( n41876 , n41874 , n41875 );
xnor ( n41877 , n41876 , n28124 );
and ( n41878 , n41873 , n41877 );
xor ( n41879 , n41609 , n41610 );
and ( n41880 , n41877 , n41879 );
and ( n41881 , n41873 , n41879 );
or ( n41882 , n41878 , n41880 , n41881 );
xor ( n41883 , n41655 , n41656 );
and ( n41884 , n26782 , n39261 );
and ( n41885 , n26678 , n39713 );
and ( n41886 , n41884 , n41885 );
xor ( n41887 , n33290 , n33565 );
buf ( n41888 , n41887 );
buf ( n41889 , n41888 );
buf ( n41890 , n41889 );
and ( n41891 , n41890 , n28117 );
and ( n41892 , n41885 , n41891 );
and ( n41893 , n41884 , n41891 );
or ( n41894 , n41886 , n41892 , n41893 );
and ( n41895 , n41883 , n41894 );
and ( n41896 , n26933 , n38737 );
and ( n41897 , n25959 , n41038 );
and ( n41898 , n41896 , n41897 );
and ( n41899 , n25742 , n41445 );
and ( n41900 , n41897 , n41899 );
and ( n41901 , n41896 , n41899 );
or ( n41902 , n41898 , n41900 , n41901 );
and ( n41903 , n41894 , n41902 );
and ( n41904 , n41883 , n41902 );
or ( n41905 , n41895 , n41903 , n41904 );
and ( n41906 , n41882 , n41905 );
buf ( n41907 , n15810 );
buf ( n41908 , n41907 );
and ( n41909 , n25623 , n41908 );
buf ( n41910 , n25451 );
and ( n41911 , n41909 , n41910 );
and ( n41912 , n38777 , n37197 );
and ( n41913 , n38462 , n37194 );
nor ( n41914 , n41912 , n41913 );
xnor ( n41915 , n41914 , n36218 );
and ( n41916 , n41910 , n41915 );
and ( n41917 , n41909 , n41915 );
or ( n41918 , n41911 , n41916 , n41917 );
and ( n41919 , n39200 , n36910 );
and ( n41920 , n38979 , n36908 );
nor ( n41921 , n41919 , n41920 );
xnor ( n41922 , n41921 , n36221 );
and ( n41923 , n39759 , n36367 );
and ( n41924 , n39500 , n36365 );
nor ( n41925 , n41923 , n41924 );
xnor ( n41926 , n41925 , n35608 );
and ( n41927 , n41922 , n41926 );
and ( n41928 , n40172 , n35911 );
and ( n41929 , n39768 , n35909 );
nor ( n41930 , n41928 , n41929 );
xnor ( n41931 , n41930 , n35161 );
and ( n41932 , n41926 , n41931 );
and ( n41933 , n41922 , n41931 );
or ( n41934 , n41927 , n41932 , n41933 );
and ( n41935 , n41918 , n41934 );
xor ( n41936 , n41662 , n41663 );
xor ( n41937 , n41936 , n41665 );
and ( n41938 , n41934 , n41937 );
and ( n41939 , n41918 , n41937 );
or ( n41940 , n41935 , n41938 , n41939 );
and ( n41941 , n41905 , n41940 );
and ( n41942 , n41882 , n41940 );
or ( n41943 , n41906 , n41941 , n41942 );
and ( n41944 , n41869 , n41943 );
xor ( n41945 , n41648 , n41653 );
xor ( n41946 , n41945 , n41657 );
xor ( n41947 , n41668 , n41678 );
xor ( n41948 , n41947 , n41695 );
and ( n41949 , n41946 , n41948 );
xor ( n41950 , n41709 , n41711 );
xor ( n41951 , n41950 , n41714 );
and ( n41952 , n41948 , n41951 );
and ( n41953 , n41946 , n41951 );
or ( n41954 , n41949 , n41952 , n41953 );
and ( n41955 , n41943 , n41954 );
and ( n41956 , n41869 , n41954 );
or ( n41957 , n41944 , n41955 , n41956 );
and ( n41958 , n41859 , n41957 );
xor ( n41959 , n41608 , n41623 );
xor ( n41960 , n41959 , n41701 );
and ( n41961 , n41957 , n41960 );
and ( n41962 , n41859 , n41960 );
or ( n41963 , n41958 , n41961 , n41962 );
and ( n41964 , n41849 , n41963 );
and ( n41965 , n41810 , n41963 );
or ( n41966 , n41850 , n41964 , n41965 );
and ( n41967 , n41808 , n41966 );
xor ( n41968 , n41547 , n41549 );
xor ( n41969 , n41968 , n41551 );
and ( n41970 , n41966 , n41969 );
and ( n41971 , n41808 , n41969 );
or ( n41972 , n41967 , n41970 , n41971 );
and ( n41973 , n41806 , n41972 );
xor ( n41974 , n41554 , n41747 );
xor ( n41975 , n41974 , n41750 );
and ( n41976 , n41972 , n41975 );
and ( n41977 , n41806 , n41975 );
or ( n41978 , n41973 , n41976 , n41977 );
xor ( n41979 , n41753 , n41755 );
xor ( n41980 , n41979 , n41758 );
and ( n41981 , n41978 , n41980 );
xor ( n41982 , n41707 , n41741 );
xor ( n41983 , n41982 , n41744 );
xor ( n41984 , n41556 , n41586 );
xor ( n41985 , n41984 , n41704 );
xor ( n41986 , n41733 , n41735 );
xor ( n41987 , n41986 , n41738 );
and ( n41988 , n41985 , n41987 );
xor ( n41989 , n41725 , n41727 );
xor ( n41990 , n41989 , n41730 );
xor ( n41991 , n41644 , n41660 );
xor ( n41992 , n41991 , n41698 );
xor ( n41993 , n41717 , n41719 );
xor ( n41994 , n41993 , n41722 );
and ( n41995 , n41992 , n41994 );
xor ( n41996 , n41836 , n41840 );
xor ( n41997 , n41996 , n41843 );
and ( n41998 , n41994 , n41997 );
and ( n41999 , n41992 , n41997 );
or ( n42000 , n41995 , n41998 , n41999 );
and ( n42001 , n41990 , n42000 );
and ( n42002 , n25959 , n41445 );
and ( n42003 , n25742 , n41908 );
and ( n42004 , n42002 , n42003 );
and ( n42005 , n26399 , n40196 );
and ( n42006 , n42004 , n42005 );
and ( n42007 , n26148 , n40643 );
and ( n42008 , n42005 , n42007 );
and ( n42009 , n42004 , n42007 );
or ( n42010 , n42006 , n42008 , n42009 );
and ( n42011 , n27591 , n36690 );
and ( n42012 , n42010 , n42011 );
and ( n42013 , n26980 , n37626 );
and ( n42014 , n42011 , n42013 );
and ( n42015 , n42010 , n42013 );
or ( n42016 , n42012 , n42014 , n42015 );
and ( n42017 , n40586 , n34911 );
and ( n42018 , n40178 , n34909 );
nor ( n42019 , n42017 , n42018 );
xnor ( n42020 , n42019 , n34104 );
or ( n42021 , n42016 , n42020 );
xor ( n42022 , n41669 , n41670 );
xor ( n42023 , n42022 , n41675 );
xor ( n42024 , n41683 , n41687 );
xor ( n42025 , n42024 , n41692 );
and ( n42026 , n42023 , n42025 );
xor ( n42027 , n41816 , n41820 );
xor ( n42028 , n42027 , n41823 );
and ( n42029 , n42025 , n42028 );
and ( n42030 , n42023 , n42028 );
or ( n42031 , n42026 , n42029 , n42030 );
and ( n42032 , n41012 , n34911 );
and ( n42033 , n40623 , n34909 );
nor ( n42034 , n42032 , n42033 );
xnor ( n42035 , n42034 , n34104 );
and ( n42036 , n41621 , n34352 );
and ( n42037 , n41405 , n34350 );
nor ( n42038 , n42036 , n42037 );
xnor ( n42039 , n42038 , n28532 );
and ( n42040 , n42035 , n42039 );
and ( n42041 , n27863 , n37187 );
and ( n42042 , n27389 , n38204 );
and ( n42043 , n42041 , n42042 );
and ( n42044 , n26933 , n39261 );
and ( n42045 , n42042 , n42044 );
and ( n42046 , n42041 , n42044 );
or ( n42047 , n42043 , n42045 , n42046 );
and ( n42048 , n42039 , n42047 );
and ( n42049 , n42035 , n42047 );
or ( n42050 , n42040 , n42048 , n42049 );
and ( n42051 , n26399 , n40643 );
and ( n42052 , n26148 , n41038 );
and ( n42053 , n42051 , n42052 );
and ( n42054 , n38979 , n37197 );
and ( n42055 , n38777 , n37194 );
nor ( n42056 , n42054 , n42055 );
xnor ( n42057 , n42056 , n36218 );
and ( n42058 , n42052 , n42057 );
and ( n42059 , n42051 , n42057 );
or ( n42060 , n42053 , n42058 , n42059 );
and ( n42061 , n39500 , n36910 );
and ( n42062 , n39200 , n36908 );
nor ( n42063 , n42061 , n42062 );
xnor ( n42064 , n42063 , n36221 );
and ( n42065 , n39768 , n36367 );
and ( n42066 , n39759 , n36365 );
nor ( n42067 , n42065 , n42066 );
xnor ( n42068 , n42067 , n35608 );
and ( n42069 , n42064 , n42068 );
and ( n42070 , n40178 , n35911 );
and ( n42071 , n40172 , n35909 );
nor ( n42072 , n42070 , n42071 );
xnor ( n42073 , n42072 , n35161 );
and ( n42074 , n42068 , n42073 );
and ( n42075 , n42064 , n42073 );
or ( n42076 , n42069 , n42074 , n42075 );
and ( n42077 , n42060 , n42076 );
xor ( n42078 , n41896 , n41897 );
xor ( n42079 , n42078 , n41899 );
and ( n42080 , n42076 , n42079 );
and ( n42081 , n42060 , n42079 );
or ( n42082 , n42077 , n42080 , n42081 );
and ( n42083 , n42050 , n42082 );
xor ( n42084 , n41873 , n41877 );
xor ( n42085 , n42084 , n41879 );
and ( n42086 , n42082 , n42085 );
and ( n42087 , n42050 , n42085 );
or ( n42088 , n42083 , n42086 , n42087 );
and ( n42089 , n42031 , n42088 );
xor ( n42090 , n41861 , n41863 );
xor ( n42091 , n42090 , n41866 );
and ( n42092 , n42088 , n42091 );
and ( n42093 , n42031 , n42091 );
or ( n42094 , n42089 , n42092 , n42093 );
and ( n42095 , n42021 , n42094 );
xor ( n42096 , n41852 , n41854 );
xor ( n42097 , n42096 , n41856 );
and ( n42098 , n42094 , n42097 );
and ( n42099 , n42021 , n42097 );
or ( n42100 , n42095 , n42098 , n42099 );
and ( n42101 , n42000 , n42100 );
and ( n42102 , n41990 , n42100 );
or ( n42103 , n42001 , n42101 , n42102 );
and ( n42104 , n41987 , n42103 );
and ( n42105 , n41985 , n42103 );
or ( n42106 , n41988 , n42104 , n42105 );
and ( n42107 , n41983 , n42106 );
xor ( n42108 , n41808 , n41966 );
xor ( n42109 , n42108 , n41969 );
and ( n42110 , n42106 , n42109 );
and ( n42111 , n41983 , n42109 );
or ( n42112 , n42107 , n42110 , n42111 );
xor ( n42113 , n41806 , n41972 );
xor ( n42114 , n42113 , n41975 );
and ( n42115 , n42112 , n42114 );
xor ( n42116 , n41810 , n41849 );
xor ( n42117 , n42116 , n41963 );
xor ( n42118 , n41812 , n41814 );
xor ( n42119 , n42118 , n41846 );
xor ( n42120 , n41859 , n41957 );
xor ( n42121 , n42120 , n41960 );
and ( n42122 , n42119 , n42121 );
xor ( n42123 , n41869 , n41943 );
xor ( n42124 , n42123 , n41954 );
xor ( n42125 , n41882 , n41905 );
xor ( n42126 , n42125 , n41940 );
xor ( n42127 , n41946 , n41948 );
xor ( n42128 , n42127 , n41951 );
and ( n42129 , n42126 , n42128 );
xnor ( n42130 , n42016 , n42020 );
and ( n42131 , n42128 , n42130 );
and ( n42132 , n42126 , n42130 );
or ( n42133 , n42129 , n42131 , n42132 );
and ( n42134 , n42124 , n42133 );
and ( n42135 , n27962 , n36229 );
and ( n42136 , n27863 , n36690 );
and ( n42137 , n42135 , n42136 );
xor ( n42138 , n41884 , n41885 );
xor ( n42139 , n42138 , n41891 );
and ( n42140 , n42136 , n42139 );
and ( n42141 , n42135 , n42139 );
or ( n42142 , n42137 , n42140 , n42141 );
xor ( n42143 , n42010 , n42011 );
xor ( n42144 , n42143 , n42013 );
and ( n42145 , n42142 , n42144 );
xor ( n42146 , n41883 , n41894 );
xor ( n42147 , n42146 , n41902 );
xor ( n42148 , n41918 , n41934 );
xor ( n42149 , n42148 , n41937 );
and ( n42150 , n42147 , n42149 );
xor ( n42151 , n42002 , n42003 );
and ( n42152 , n26678 , n40196 );
and ( n42153 , n42151 , n42152 );
xor ( n42154 , n33327 , n33563 );
buf ( n42155 , n42154 );
buf ( n42156 , n42155 );
buf ( n42157 , n42156 );
and ( n42158 , n42157 , n28117 );
and ( n42159 , n42152 , n42158 );
and ( n42160 , n42151 , n42158 );
or ( n42161 , n42153 , n42159 , n42160 );
and ( n42162 , n27591 , n37187 );
and ( n42163 , n42161 , n42162 );
and ( n42164 , n27389 , n37626 );
and ( n42165 , n42162 , n42164 );
and ( n42166 , n42161 , n42164 );
or ( n42167 , n42163 , n42165 , n42166 );
and ( n42168 , n42149 , n42167 );
and ( n42169 , n42147 , n42167 );
or ( n42170 , n42150 , n42168 , n42169 );
and ( n42171 , n42145 , n42170 );
and ( n42172 , n26980 , n38204 );
and ( n42173 , n41631 , n33632 );
and ( n42174 , n41652 , n33630 );
nor ( n42175 , n42173 , n42174 );
xnor ( n42176 , n42175 , n28124 );
and ( n42177 , n42172 , n42176 );
xor ( n42178 , n42004 , n42005 );
xor ( n42179 , n42178 , n42007 );
and ( n42180 , n42176 , n42179 );
and ( n42181 , n42172 , n42179 );
or ( n42182 , n42177 , n42180 , n42181 );
xor ( n42183 , n41909 , n41910 );
xor ( n42184 , n42183 , n41915 );
xor ( n42185 , n41922 , n41926 );
xor ( n42186 , n42185 , n41931 );
and ( n42187 , n42184 , n42186 );
xor ( n42188 , n42135 , n42136 );
xor ( n42189 , n42188 , n42139 );
and ( n42190 , n42186 , n42189 );
and ( n42191 , n42184 , n42189 );
or ( n42192 , n42187 , n42190 , n42191 );
and ( n42193 , n42182 , n42192 );
and ( n42194 , n26399 , n41038 );
and ( n42195 , n26148 , n41445 );
and ( n42196 , n42194 , n42195 );
and ( n42197 , n25959 , n41908 );
and ( n42198 , n42195 , n42197 );
and ( n42199 , n42194 , n42197 );
or ( n42200 , n42196 , n42198 , n42199 );
and ( n42201 , n26980 , n38737 );
and ( n42202 , n42200 , n42201 );
and ( n42203 , n26782 , n39713 );
and ( n42204 , n42201 , n42203 );
and ( n42205 , n42200 , n42203 );
or ( n42206 , n42202 , n42204 , n42205 );
and ( n42207 , n40623 , n35374 );
and ( n42208 , n40586 , n35372 );
nor ( n42209 , n42207 , n42208 );
xnor ( n42210 , n42209 , n34661 );
xor ( n42211 , n42041 , n42042 );
xor ( n42212 , n42211 , n42044 );
and ( n42213 , n42210 , n42212 );
and ( n42214 , n42206 , n42213 );
and ( n42215 , n41405 , n34911 );
and ( n42216 , n41012 , n34909 );
nor ( n42217 , n42215 , n42216 );
xnor ( n42218 , n42217 , n34104 );
and ( n42219 , n41890 , n33632 );
and ( n42220 , n41631 , n33630 );
nor ( n42221 , n42219 , n42220 );
xnor ( n42222 , n42221 , n28124 );
and ( n42223 , n42218 , n42222 );
and ( n42224 , n28129 , n36690 );
and ( n42225 , n27863 , n37626 );
and ( n42226 , n42224 , n42225 );
and ( n42227 , n27389 , n38737 );
and ( n42228 , n42225 , n42227 );
and ( n42229 , n42224 , n42227 );
or ( n42230 , n42226 , n42228 , n42229 );
and ( n42231 , n42222 , n42230 );
and ( n42232 , n42218 , n42230 );
or ( n42233 , n42223 , n42231 , n42232 );
and ( n42234 , n42213 , n42233 );
and ( n42235 , n42206 , n42233 );
or ( n42236 , n42214 , n42234 , n42235 );
and ( n42237 , n42192 , n42236 );
and ( n42238 , n42182 , n42236 );
or ( n42239 , n42193 , n42237 , n42238 );
and ( n42240 , n42170 , n42239 );
and ( n42241 , n42145 , n42239 );
or ( n42242 , n42171 , n42240 , n42241 );
and ( n42243 , n42133 , n42242 );
and ( n42244 , n42124 , n42242 );
or ( n42245 , n42134 , n42243 , n42244 );
and ( n42246 , n42121 , n42245 );
and ( n42247 , n42119 , n42245 );
or ( n42248 , n42122 , n42246 , n42247 );
and ( n42249 , n42117 , n42248 );
xor ( n42250 , n41985 , n41987 );
xor ( n42251 , n42250 , n42103 );
and ( n42252 , n42248 , n42251 );
and ( n42253 , n42117 , n42251 );
or ( n42254 , n42249 , n42252 , n42253 );
xor ( n42255 , n41983 , n42106 );
xor ( n42256 , n42255 , n42109 );
and ( n42257 , n42254 , n42256 );
xor ( n42258 , n41990 , n42000 );
xor ( n42259 , n42258 , n42100 );
xor ( n42260 , n41992 , n41994 );
xor ( n42261 , n42260 , n41997 );
xor ( n42262 , n42021 , n42094 );
xor ( n42263 , n42262 , n42097 );
and ( n42264 , n42261 , n42263 );
and ( n42265 , n26933 , n39713 );
and ( n42266 , n26782 , n40196 );
and ( n42267 , n42265 , n42266 );
and ( n42268 , n26678 , n40643 );
and ( n42269 , n42266 , n42268 );
and ( n42270 , n42265 , n42268 );
or ( n42271 , n42267 , n42269 , n42270 );
and ( n42272 , n28129 , n36229 );
and ( n42273 , n42271 , n42272 );
and ( n42274 , n27591 , n37626 );
and ( n42275 , n42272 , n42274 );
and ( n42276 , n42271 , n42274 );
or ( n42277 , n42273 , n42275 , n42276 );
and ( n42278 , n27962 , n36690 );
and ( n42279 , n41652 , n34352 );
and ( n42280 , n41621 , n34350 );
nor ( n42281 , n42279 , n42280 );
xnor ( n42282 , n42281 , n28532 );
and ( n42283 , n42278 , n42282 );
xor ( n42284 , n42151 , n42152 );
xor ( n42285 , n42284 , n42158 );
and ( n42286 , n42282 , n42285 );
and ( n42287 , n42278 , n42285 );
or ( n42288 , n42283 , n42286 , n42287 );
and ( n42289 , n42277 , n42288 );
and ( n42290 , n40586 , n35374 );
and ( n42291 , n40178 , n35372 );
nor ( n42292 , n42290 , n42291 );
xnor ( n42293 , n42292 , n34661 );
and ( n42294 , n42288 , n42293 );
and ( n42295 , n42277 , n42293 );
or ( n42296 , n42289 , n42294 , n42295 );
and ( n42297 , n28129 , n35544 );
xor ( n42298 , n42161 , n42162 );
xor ( n42299 , n42298 , n42164 );
and ( n42300 , n42297 , n42299 );
xor ( n42301 , n42172 , n42176 );
xor ( n42302 , n42301 , n42179 );
and ( n42303 , n42299 , n42302 );
and ( n42304 , n42297 , n42302 );
or ( n42305 , n42300 , n42303 , n42304 );
and ( n42306 , n42296 , n42305 );
and ( n42307 , n39768 , n35911 );
and ( n42308 , n39759 , n35909 );
nor ( n42309 , n42307 , n42308 );
xnor ( n42310 , n42309 , n35161 );
and ( n42311 , n42305 , n42310 );
and ( n42312 , n42296 , n42310 );
or ( n42313 , n42306 , n42311 , n42312 );
xor ( n42314 , n41826 , n41830 );
xor ( n42315 , n42314 , n41833 );
and ( n42316 , n42313 , n42315 );
and ( n42317 , n42263 , n42316 );
and ( n42318 , n42261 , n42316 );
or ( n42319 , n42264 , n42317 , n42318 );
and ( n42320 , n42259 , n42319 );
and ( n42321 , n26980 , n39261 );
buf ( n42322 , n15972 );
buf ( n42323 , n42322 );
and ( n42324 , n25742 , n42323 );
and ( n42325 , n42321 , n42324 );
buf ( n42326 , n25623 );
and ( n42327 , n42324 , n42326 );
and ( n42328 , n42321 , n42326 );
or ( n42329 , n42325 , n42327 , n42328 );
and ( n42330 , n39200 , n37197 );
and ( n42331 , n38979 , n37194 );
nor ( n42332 , n42330 , n42331 );
xnor ( n42333 , n42332 , n36218 );
and ( n42334 , n39759 , n36910 );
and ( n42335 , n39500 , n36908 );
nor ( n42336 , n42334 , n42335 );
xnor ( n42337 , n42336 , n36221 );
and ( n42338 , n42333 , n42337 );
and ( n42339 , n40172 , n36367 );
and ( n42340 , n39768 , n36365 );
nor ( n42341 , n42339 , n42340 );
xnor ( n42342 , n42341 , n35608 );
and ( n42343 , n42337 , n42342 );
and ( n42344 , n42333 , n42342 );
or ( n42345 , n42338 , n42343 , n42344 );
and ( n42346 , n42329 , n42345 );
and ( n42347 , n40586 , n35911 );
and ( n42348 , n40178 , n35909 );
nor ( n42349 , n42347 , n42348 );
xnor ( n42350 , n42349 , n35161 );
and ( n42351 , n41012 , n35374 );
and ( n42352 , n40623 , n35372 );
nor ( n42353 , n42351 , n42352 );
xnor ( n42354 , n42353 , n34661 );
and ( n42355 , n42350 , n42354 );
and ( n42356 , n41621 , n34911 );
and ( n42357 , n41405 , n34909 );
nor ( n42358 , n42356 , n42357 );
xnor ( n42359 , n42358 , n34104 );
and ( n42360 , n42354 , n42359 );
and ( n42361 , n42350 , n42359 );
or ( n42362 , n42355 , n42360 , n42361 );
and ( n42363 , n42345 , n42362 );
and ( n42364 , n42329 , n42362 );
or ( n42365 , n42346 , n42363 , n42364 );
xor ( n42366 , n42035 , n42039 );
xor ( n42367 , n42366 , n42047 );
and ( n42368 , n42365 , n42367 );
xor ( n42369 , n42060 , n42076 );
xor ( n42370 , n42369 , n42079 );
and ( n42371 , n42367 , n42370 );
and ( n42372 , n42365 , n42370 );
or ( n42373 , n42368 , n42371 , n42372 );
xor ( n42374 , n42023 , n42025 );
xor ( n42375 , n42374 , n42028 );
and ( n42376 , n42373 , n42375 );
xor ( n42377 , n42050 , n42082 );
xor ( n42378 , n42377 , n42085 );
and ( n42379 , n42375 , n42378 );
and ( n42380 , n42373 , n42378 );
or ( n42381 , n42376 , n42379 , n42380 );
xor ( n42382 , n42031 , n42088 );
xor ( n42383 , n42382 , n42091 );
and ( n42384 , n42381 , n42383 );
xor ( n42385 , n42142 , n42144 );
xor ( n42386 , n42051 , n42052 );
xor ( n42387 , n42386 , n42057 );
xor ( n42388 , n42064 , n42068 );
xor ( n42389 , n42388 , n42073 );
and ( n42390 , n42387 , n42389 );
xor ( n42391 , n42200 , n42201 );
xor ( n42392 , n42391 , n42203 );
and ( n42393 , n42389 , n42392 );
and ( n42394 , n42387 , n42392 );
or ( n42395 , n42390 , n42393 , n42394 );
xor ( n42396 , n42271 , n42272 );
xor ( n42397 , n42396 , n42274 );
xor ( n42398 , n42210 , n42212 );
and ( n42399 , n42397 , n42398 );
and ( n42400 , n42157 , n33632 );
and ( n42401 , n41890 , n33630 );
nor ( n42402 , n42400 , n42401 );
xnor ( n42403 , n42402 , n28124 );
xor ( n42404 , n42194 , n42195 );
xor ( n42405 , n42404 , n42197 );
and ( n42406 , n42403 , n42405 );
and ( n42407 , n42398 , n42406 );
and ( n42408 , n42397 , n42406 );
or ( n42409 , n42399 , n42407 , n42408 );
and ( n42410 , n42395 , n42409 );
xor ( n42411 , n33363 , n33561 );
buf ( n42412 , n42411 );
buf ( n42413 , n42412 );
buf ( n42414 , n42413 );
and ( n42415 , n42414 , n28117 );
and ( n42416 , n26148 , n41908 );
and ( n42417 , n25959 , n42323 );
and ( n42418 , n42416 , n42417 );
and ( n42419 , n42415 , n42418 );
and ( n42420 , n28129 , n37187 );
and ( n42421 , n27962 , n37626 );
and ( n42422 , n42420 , n42421 );
and ( n42423 , n26980 , n39713 );
and ( n42424 , n42421 , n42423 );
and ( n42425 , n42420 , n42423 );
or ( n42426 , n42422 , n42424 , n42425 );
and ( n42427 , n42418 , n42426 );
and ( n42428 , n42415 , n42426 );
or ( n42429 , n42419 , n42427 , n42428 );
and ( n42430 , n26678 , n41038 );
and ( n42431 , n26399 , n41445 );
and ( n42432 , n42430 , n42431 );
and ( n42433 , n39500 , n37197 );
and ( n42434 , n39200 , n37194 );
nor ( n42435 , n42433 , n42434 );
xnor ( n42436 , n42435 , n36218 );
and ( n42437 , n42431 , n42436 );
and ( n42438 , n42430 , n42436 );
or ( n42439 , n42432 , n42437 , n42438 );
and ( n42440 , n39768 , n36910 );
and ( n42441 , n39759 , n36908 );
nor ( n42442 , n42440 , n42441 );
xnor ( n42443 , n42442 , n36221 );
and ( n42444 , n40178 , n36367 );
and ( n42445 , n40172 , n36365 );
nor ( n42446 , n42444 , n42445 );
xnor ( n42447 , n42446 , n35608 );
and ( n42448 , n42443 , n42447 );
and ( n42449 , n40623 , n35911 );
and ( n42450 , n40586 , n35909 );
nor ( n42451 , n42449 , n42450 );
xnor ( n42452 , n42451 , n35161 );
and ( n42453 , n42447 , n42452 );
and ( n42454 , n42443 , n42452 );
or ( n42455 , n42448 , n42453 , n42454 );
and ( n42456 , n42439 , n42455 );
and ( n42457 , n41405 , n35374 );
and ( n42458 , n41012 , n35372 );
nor ( n42459 , n42457 , n42458 );
xnor ( n42460 , n42459 , n34661 );
and ( n42461 , n41652 , n34911 );
and ( n42462 , n41621 , n34909 );
nor ( n42463 , n42461 , n42462 );
xnor ( n42464 , n42463 , n34104 );
and ( n42465 , n42460 , n42464 );
and ( n42466 , n41890 , n34352 );
and ( n42467 , n41631 , n34350 );
nor ( n42468 , n42466 , n42467 );
xnor ( n42469 , n42468 , n28532 );
and ( n42470 , n42464 , n42469 );
and ( n42471 , n42460 , n42469 );
or ( n42472 , n42465 , n42470 , n42471 );
and ( n42473 , n42455 , n42472 );
and ( n42474 , n42439 , n42472 );
or ( n42475 , n42456 , n42473 , n42474 );
and ( n42476 , n42429 , n42475 );
xor ( n42477 , n42224 , n42225 );
xor ( n42478 , n42477 , n42227 );
xor ( n42479 , n42321 , n42324 );
xor ( n42480 , n42479 , n42326 );
and ( n42481 , n42478 , n42480 );
xor ( n42482 , n42333 , n42337 );
xor ( n42483 , n42482 , n42342 );
and ( n42484 , n42480 , n42483 );
and ( n42485 , n42478 , n42483 );
or ( n42486 , n42481 , n42484 , n42485 );
and ( n42487 , n42475 , n42486 );
and ( n42488 , n42429 , n42486 );
or ( n42489 , n42476 , n42487 , n42488 );
and ( n42490 , n42409 , n42489 );
and ( n42491 , n42395 , n42489 );
or ( n42492 , n42410 , n42490 , n42491 );
and ( n42493 , n42385 , n42492 );
xor ( n42494 , n42184 , n42186 );
xor ( n42495 , n42494 , n42189 );
xor ( n42496 , n42206 , n42213 );
xor ( n42497 , n42496 , n42233 );
and ( n42498 , n42495 , n42497 );
xor ( n42499 , n42365 , n42367 );
xor ( n42500 , n42499 , n42370 );
and ( n42501 , n42497 , n42500 );
and ( n42502 , n42495 , n42500 );
or ( n42503 , n42498 , n42501 , n42502 );
and ( n42504 , n42492 , n42503 );
and ( n42505 , n42385 , n42503 );
or ( n42506 , n42493 , n42504 , n42505 );
and ( n42507 , n42383 , n42506 );
and ( n42508 , n42381 , n42506 );
or ( n42509 , n42384 , n42507 , n42508 );
xor ( n42510 , n42147 , n42149 );
xor ( n42511 , n42510 , n42167 );
xor ( n42512 , n42182 , n42192 );
xor ( n42513 , n42512 , n42236 );
and ( n42514 , n42511 , n42513 );
xor ( n42515 , n42373 , n42375 );
xor ( n42516 , n42515 , n42378 );
and ( n42517 , n42513 , n42516 );
and ( n42518 , n42511 , n42516 );
or ( n42519 , n42514 , n42517 , n42518 );
xor ( n42520 , n42126 , n42128 );
xor ( n42521 , n42520 , n42130 );
and ( n42522 , n42519 , n42521 );
xor ( n42523 , n42145 , n42170 );
xor ( n42524 , n42523 , n42239 );
and ( n42525 , n42521 , n42524 );
and ( n42526 , n42519 , n42524 );
or ( n42527 , n42522 , n42525 , n42526 );
and ( n42528 , n42509 , n42527 );
xor ( n42529 , n42124 , n42133 );
xor ( n42530 , n42529 , n42242 );
and ( n42531 , n42527 , n42530 );
and ( n42532 , n42509 , n42530 );
or ( n42533 , n42528 , n42531 , n42532 );
and ( n42534 , n42319 , n42533 );
and ( n42535 , n42259 , n42533 );
or ( n42536 , n42320 , n42534 , n42535 );
xor ( n42537 , n42117 , n42248 );
xor ( n42538 , n42537 , n42251 );
and ( n42539 , n42536 , n42538 );
xor ( n42540 , n42119 , n42121 );
xor ( n42541 , n42540 , n42245 );
xor ( n42542 , n42313 , n42315 );
xor ( n42543 , n42296 , n42305 );
xor ( n42544 , n42543 , n42310 );
xor ( n42545 , n42277 , n42288 );
xor ( n42546 , n42545 , n42293 );
xor ( n42547 , n42297 , n42299 );
xor ( n42548 , n42547 , n42302 );
and ( n42549 , n42546 , n42548 );
xor ( n42550 , n42218 , n42222 );
xor ( n42551 , n42550 , n42230 );
xor ( n42552 , n42329 , n42345 );
xor ( n42553 , n42552 , n42362 );
and ( n42554 , n42551 , n42553 );
xor ( n42555 , n42278 , n42282 );
xor ( n42556 , n42555 , n42285 );
and ( n42557 , n42553 , n42556 );
and ( n42558 , n42551 , n42556 );
or ( n42559 , n42554 , n42557 , n42558 );
and ( n42560 , n42548 , n42559 );
and ( n42561 , n42546 , n42559 );
or ( n42562 , n42549 , n42560 , n42561 );
and ( n42563 , n42544 , n42562 );
xor ( n42564 , n42416 , n42417 );
and ( n42565 , n26782 , n40643 );
and ( n42566 , n42564 , n42565 );
xor ( n42567 , n33399 , n33559 );
buf ( n42568 , n42567 );
buf ( n42569 , n42568 );
buf ( n42570 , n42569 );
and ( n42571 , n42570 , n28117 );
and ( n42572 , n42565 , n42571 );
and ( n42573 , n42564 , n42571 );
or ( n42574 , n42566 , n42572 , n42573 );
and ( n42575 , n27591 , n38204 );
and ( n42576 , n42574 , n42575 );
and ( n42577 , n41631 , n34352 );
and ( n42578 , n41652 , n34350 );
nor ( n42579 , n42577 , n42578 );
xnor ( n42580 , n42579 , n28532 );
and ( n42581 , n42575 , n42580 );
and ( n42582 , n42574 , n42580 );
or ( n42583 , n42576 , n42581 , n42582 );
and ( n42584 , n26678 , n41445 );
and ( n42585 , n26399 , n41908 );
and ( n42586 , n42584 , n42585 );
and ( n42587 , n26148 , n42323 );
and ( n42588 , n42585 , n42587 );
and ( n42589 , n42584 , n42587 );
or ( n42590 , n42586 , n42588 , n42589 );
and ( n42591 , n26933 , n40196 );
and ( n42592 , n42590 , n42591 );
and ( n42593 , n42414 , n33632 );
and ( n42594 , n42157 , n33630 );
nor ( n42595 , n42593 , n42594 );
xnor ( n42596 , n42595 , n28124 );
and ( n42597 , n42591 , n42596 );
and ( n42598 , n42590 , n42596 );
or ( n42599 , n42592 , n42597 , n42598 );
and ( n42600 , n27962 , n37187 );
and ( n42601 , n42599 , n42600 );
xor ( n42602 , n42265 , n42266 );
xor ( n42603 , n42602 , n42268 );
and ( n42604 , n42600 , n42603 );
and ( n42605 , n42599 , n42603 );
or ( n42606 , n42601 , n42604 , n42605 );
and ( n42607 , n42583 , n42606 );
xor ( n42608 , n42350 , n42354 );
xor ( n42609 , n42608 , n42359 );
xor ( n42610 , n42403 , n42405 );
and ( n42611 , n42609 , n42610 );
and ( n42612 , n28129 , n37626 );
and ( n42613 , n27962 , n38204 );
and ( n42614 , n42612 , n42613 );
and ( n42615 , n27389 , n39713 );
and ( n42616 , n42613 , n42615 );
and ( n42617 , n42612 , n42615 );
or ( n42618 , n42614 , n42616 , n42617 );
and ( n42619 , n26782 , n41038 );
buf ( n42620 , n16248 );
buf ( n42621 , n42620 );
and ( n42622 , n25959 , n42621 );
and ( n42623 , n42619 , n42622 );
buf ( n42624 , n25742 );
and ( n42625 , n42622 , n42624 );
and ( n42626 , n42619 , n42624 );
or ( n42627 , n42623 , n42625 , n42626 );
and ( n42628 , n42618 , n42627 );
and ( n42629 , n39759 , n37197 );
and ( n42630 , n39500 , n37194 );
nor ( n42631 , n42629 , n42630 );
xnor ( n42632 , n42631 , n36218 );
and ( n42633 , n40172 , n36910 );
and ( n42634 , n39768 , n36908 );
nor ( n42635 , n42633 , n42634 );
xnor ( n42636 , n42635 , n36221 );
and ( n42637 , n42632 , n42636 );
and ( n42638 , n40586 , n36367 );
and ( n42639 , n40178 , n36365 );
nor ( n42640 , n42638 , n42639 );
xnor ( n42641 , n42640 , n35608 );
and ( n42642 , n42636 , n42641 );
and ( n42643 , n42632 , n42641 );
or ( n42644 , n42637 , n42642 , n42643 );
and ( n42645 , n42627 , n42644 );
and ( n42646 , n42618 , n42644 );
or ( n42647 , n42628 , n42645 , n42646 );
and ( n42648 , n42610 , n42647 );
and ( n42649 , n42609 , n42647 );
or ( n42650 , n42611 , n42648 , n42649 );
and ( n42651 , n42606 , n42650 );
and ( n42652 , n42583 , n42650 );
or ( n42653 , n42607 , n42651 , n42652 );
and ( n42654 , n41012 , n35911 );
and ( n42655 , n40623 , n35909 );
nor ( n42656 , n42654 , n42655 );
xnor ( n42657 , n42656 , n35161 );
and ( n42658 , n41621 , n35374 );
and ( n42659 , n41405 , n35372 );
nor ( n42660 , n42658 , n42659 );
xnor ( n42661 , n42660 , n34661 );
and ( n42662 , n42657 , n42661 );
and ( n42663 , n41631 , n34911 );
and ( n42664 , n41652 , n34909 );
nor ( n42665 , n42663 , n42664 );
xnor ( n42666 , n42665 , n34104 );
and ( n42667 , n42661 , n42666 );
and ( n42668 , n42657 , n42666 );
or ( n42669 , n42662 , n42667 , n42668 );
and ( n42670 , n42157 , n34352 );
and ( n42671 , n41890 , n34350 );
nor ( n42672 , n42670 , n42671 );
xnor ( n42673 , n42672 , n28532 );
and ( n42674 , n42570 , n33632 );
and ( n42675 , n42414 , n33630 );
nor ( n42676 , n42674 , n42675 );
xnor ( n42677 , n42676 , n28124 );
and ( n42678 , n42673 , n42677 );
xor ( n42679 , n33426 , n33557 );
buf ( n42680 , n42679 );
buf ( n42681 , n42680 );
buf ( n42682 , n42681 );
and ( n42683 , n42682 , n28117 );
and ( n42684 , n42677 , n42683 );
and ( n42685 , n42673 , n42683 );
or ( n42686 , n42678 , n42684 , n42685 );
and ( n42687 , n42669 , n42686 );
xor ( n42688 , n42420 , n42421 );
xor ( n42689 , n42688 , n42423 );
and ( n42690 , n42686 , n42689 );
and ( n42691 , n42669 , n42689 );
or ( n42692 , n42687 , n42690 , n42691 );
xor ( n42693 , n42430 , n42431 );
xor ( n42694 , n42693 , n42436 );
xor ( n42695 , n42443 , n42447 );
xor ( n42696 , n42695 , n42452 );
and ( n42697 , n42694 , n42696 );
xor ( n42698 , n42460 , n42464 );
xor ( n42699 , n42698 , n42469 );
and ( n42700 , n42696 , n42699 );
and ( n42701 , n42694 , n42699 );
or ( n42702 , n42697 , n42700 , n42701 );
and ( n42703 , n42692 , n42702 );
xor ( n42704 , n42415 , n42418 );
xor ( n42705 , n42704 , n42426 );
and ( n42706 , n42702 , n42705 );
and ( n42707 , n42692 , n42705 );
or ( n42708 , n42703 , n42706 , n42707 );
xor ( n42709 , n42387 , n42389 );
xor ( n42710 , n42709 , n42392 );
and ( n42711 , n42708 , n42710 );
xor ( n42712 , n42397 , n42398 );
xor ( n42713 , n42712 , n42406 );
and ( n42714 , n42710 , n42713 );
and ( n42715 , n42708 , n42713 );
or ( n42716 , n42711 , n42714 , n42715 );
and ( n42717 , n42653 , n42716 );
xor ( n42718 , n42395 , n42409 );
xor ( n42719 , n42718 , n42489 );
and ( n42720 , n42716 , n42719 );
and ( n42721 , n42653 , n42719 );
or ( n42722 , n42717 , n42720 , n42721 );
and ( n42723 , n42562 , n42722 );
and ( n42724 , n42544 , n42722 );
or ( n42725 , n42563 , n42723 , n42724 );
and ( n42726 , n42542 , n42725 );
xor ( n42727 , n42381 , n42383 );
xor ( n42728 , n42727 , n42506 );
and ( n42729 , n42725 , n42728 );
and ( n42730 , n42542 , n42728 );
or ( n42731 , n42726 , n42729 , n42730 );
xor ( n42732 , n42261 , n42263 );
xor ( n42733 , n42732 , n42316 );
and ( n42734 , n42731 , n42733 );
xor ( n42735 , n42509 , n42527 );
xor ( n42736 , n42735 , n42530 );
and ( n42737 , n42733 , n42736 );
and ( n42738 , n42731 , n42736 );
or ( n42739 , n42734 , n42737 , n42738 );
and ( n42740 , n42541 , n42739 );
xor ( n42741 , n42259 , n42319 );
xor ( n42742 , n42741 , n42533 );
and ( n42743 , n42739 , n42742 );
and ( n42744 , n42541 , n42742 );
or ( n42745 , n42740 , n42743 , n42744 );
and ( n42746 , n42538 , n42745 );
and ( n42747 , n42536 , n42745 );
or ( n42748 , n42539 , n42746 , n42747 );
and ( n42749 , n42256 , n42748 );
and ( n42750 , n42254 , n42748 );
or ( n42751 , n42257 , n42749 , n42750 );
and ( n42752 , n42114 , n42751 );
and ( n42753 , n42112 , n42751 );
or ( n42754 , n42115 , n42752 , n42753 );
and ( n42755 , n41980 , n42754 );
and ( n42756 , n41978 , n42754 );
or ( n42757 , n41981 , n42755 , n42756 );
or ( n42758 , n41804 , n42757 );
or ( n42759 , n41802 , n42758 );
or ( n42760 , n41800 , n42759 );
and ( n42761 , n41798 , n42760 );
xor ( n42762 , n41798 , n42760 );
xnor ( n42763 , n41800 , n42759 );
xnor ( n42764 , n41802 , n42758 );
xnor ( n42765 , n41804 , n42757 );
xor ( n42766 , n41978 , n41980 );
xor ( n42767 , n42766 , n42754 );
xor ( n42768 , n42112 , n42114 );
xor ( n42769 , n42768 , n42751 );
not ( n42770 , n42769 );
xor ( n42771 , n42254 , n42256 );
xor ( n42772 , n42771 , n42748 );
not ( n42773 , n42772 );
xor ( n42774 , n42536 , n42538 );
xor ( n42775 , n42774 , n42745 );
not ( n42776 , n42775 );
xor ( n42777 , n42541 , n42739 );
xor ( n42778 , n42777 , n42742 );
xor ( n42779 , n42519 , n42521 );
xor ( n42780 , n42779 , n42524 );
xor ( n42781 , n42385 , n42492 );
xor ( n42782 , n42781 , n42503 );
xor ( n42783 , n42511 , n42513 );
xor ( n42784 , n42783 , n42516 );
and ( n42785 , n42782 , n42784 );
xor ( n42786 , n42495 , n42497 );
xor ( n42787 , n42786 , n42500 );
xor ( n42788 , n42429 , n42475 );
xor ( n42789 , n42788 , n42486 );
xor ( n42790 , n42574 , n42575 );
xor ( n42791 , n42790 , n42580 );
xor ( n42792 , n42599 , n42600 );
xor ( n42793 , n42792 , n42603 );
and ( n42794 , n42791 , n42793 );
and ( n42795 , n42789 , n42794 );
xor ( n42796 , n42439 , n42455 );
xor ( n42797 , n42796 , n42472 );
xor ( n42798 , n42478 , n42480 );
xor ( n42799 , n42798 , n42483 );
and ( n42800 , n42797 , n42799 );
and ( n42801 , n26980 , n40196 );
and ( n42802 , n26933 , n40643 );
and ( n42803 , n42801 , n42802 );
xor ( n42804 , n42584 , n42585 );
xor ( n42805 , n42804 , n42587 );
and ( n42806 , n42802 , n42805 );
and ( n42807 , n42801 , n42805 );
or ( n42808 , n42803 , n42806 , n42807 );
and ( n42809 , n27863 , n38204 );
and ( n42810 , n42808 , n42809 );
xor ( n42811 , n42590 , n42591 );
xor ( n42812 , n42811 , n42596 );
and ( n42813 , n42809 , n42812 );
and ( n42814 , n42808 , n42812 );
or ( n42815 , n42810 , n42813 , n42814 );
and ( n42816 , n42799 , n42815 );
and ( n42817 , n42797 , n42815 );
or ( n42818 , n42800 , n42816 , n42817 );
and ( n42819 , n42794 , n42818 );
and ( n42820 , n42789 , n42818 );
or ( n42821 , n42795 , n42819 , n42820 );
and ( n42822 , n42787 , n42821 );
and ( n42823 , n27591 , n38737 );
and ( n42824 , n27389 , n39261 );
and ( n42825 , n42823 , n42824 );
xor ( n42826 , n42564 , n42565 );
xor ( n42827 , n42826 , n42571 );
and ( n42828 , n42824 , n42827 );
and ( n42829 , n42823 , n42827 );
or ( n42830 , n42825 , n42828 , n42829 );
and ( n42831 , n26148 , n42621 );
xor ( n42832 , n33460 , n33555 );
buf ( n42833 , n42832 );
buf ( n42834 , n42833 );
buf ( n42835 , n42834 );
and ( n42836 , n42835 , n28117 );
and ( n42837 , n42831 , n42836 );
and ( n42838 , n28129 , n38204 );
and ( n42839 , n27863 , n39261 );
and ( n42840 , n42838 , n42839 );
and ( n42841 , n26980 , n40643 );
and ( n42842 , n42839 , n42841 );
and ( n42843 , n42838 , n42841 );
or ( n42844 , n42840 , n42842 , n42843 );
and ( n42845 , n42837 , n42844 );
and ( n42846 , n26933 , n41038 );
and ( n42847 , n26678 , n41908 );
and ( n42848 , n42846 , n42847 );
and ( n42849 , n26399 , n42323 );
and ( n42850 , n42847 , n42849 );
and ( n42851 , n42846 , n42849 );
or ( n42852 , n42848 , n42850 , n42851 );
and ( n42853 , n42844 , n42852 );
and ( n42854 , n42837 , n42852 );
or ( n42855 , n42845 , n42853 , n42854 );
and ( n42856 , n40178 , n36910 );
and ( n42857 , n40172 , n36908 );
nor ( n42858 , n42856 , n42857 );
xnor ( n42859 , n42858 , n36221 );
and ( n42860 , n40623 , n36367 );
and ( n42861 , n40586 , n36365 );
nor ( n42862 , n42860 , n42861 );
xnor ( n42863 , n42862 , n35608 );
and ( n42864 , n42859 , n42863 );
and ( n42865 , n41652 , n35374 );
and ( n42866 , n41621 , n35372 );
nor ( n42867 , n42865 , n42866 );
xnor ( n42868 , n42867 , n34661 );
and ( n42869 , n42863 , n42868 );
and ( n42870 , n42859 , n42868 );
or ( n42871 , n42864 , n42869 , n42870 );
xor ( n42872 , n42612 , n42613 );
xor ( n42873 , n42872 , n42615 );
and ( n42874 , n42871 , n42873 );
xor ( n42875 , n42619 , n42622 );
xor ( n42876 , n42875 , n42624 );
and ( n42877 , n42873 , n42876 );
and ( n42878 , n42871 , n42876 );
or ( n42879 , n42874 , n42877 , n42878 );
and ( n42880 , n42855 , n42879 );
xor ( n42881 , n42632 , n42636 );
xor ( n42882 , n42881 , n42641 );
xor ( n42883 , n42657 , n42661 );
xor ( n42884 , n42883 , n42666 );
and ( n42885 , n42882 , n42884 );
xor ( n42886 , n42673 , n42677 );
xor ( n42887 , n42886 , n42683 );
and ( n42888 , n42884 , n42887 );
and ( n42889 , n42882 , n42887 );
or ( n42890 , n42885 , n42888 , n42889 );
and ( n42891 , n42879 , n42890 );
and ( n42892 , n42855 , n42890 );
or ( n42893 , n42880 , n42891 , n42892 );
and ( n42894 , n42830 , n42893 );
xor ( n42895 , n42618 , n42627 );
xor ( n42896 , n42895 , n42644 );
xor ( n42897 , n42669 , n42686 );
xor ( n42898 , n42897 , n42689 );
and ( n42899 , n42896 , n42898 );
xor ( n42900 , n42694 , n42696 );
xor ( n42901 , n42900 , n42699 );
and ( n42902 , n42898 , n42901 );
and ( n42903 , n42896 , n42901 );
or ( n42904 , n42899 , n42902 , n42903 );
and ( n42905 , n42893 , n42904 );
and ( n42906 , n42830 , n42904 );
or ( n42907 , n42894 , n42905 , n42906 );
xor ( n42908 , n42551 , n42553 );
xor ( n42909 , n42908 , n42556 );
and ( n42910 , n42907 , n42909 );
xor ( n42911 , n42583 , n42606 );
xor ( n42912 , n42911 , n42650 );
and ( n42913 , n42909 , n42912 );
and ( n42914 , n42907 , n42912 );
or ( n42915 , n42910 , n42913 , n42914 );
and ( n42916 , n42821 , n42915 );
and ( n42917 , n42787 , n42915 );
or ( n42918 , n42822 , n42916 , n42917 );
and ( n42919 , n42784 , n42918 );
and ( n42920 , n42782 , n42918 );
or ( n42921 , n42785 , n42919 , n42920 );
and ( n42922 , n42780 , n42921 );
xor ( n42923 , n42542 , n42725 );
xor ( n42924 , n42923 , n42728 );
and ( n42925 , n42921 , n42924 );
and ( n42926 , n42780 , n42924 );
or ( n42927 , n42922 , n42925 , n42926 );
xor ( n42928 , n42731 , n42733 );
xor ( n42929 , n42928 , n42736 );
and ( n42930 , n42927 , n42929 );
xor ( n42931 , n42544 , n42562 );
xor ( n42932 , n42931 , n42722 );
xor ( n42933 , n42546 , n42548 );
xor ( n42934 , n42933 , n42559 );
xor ( n42935 , n42653 , n42716 );
xor ( n42936 , n42935 , n42719 );
and ( n42937 , n42934 , n42936 );
xor ( n42938 , n42708 , n42710 );
xor ( n42939 , n42938 , n42713 );
xor ( n42940 , n42609 , n42610 );
xor ( n42941 , n42940 , n42647 );
xor ( n42942 , n42692 , n42702 );
xor ( n42943 , n42942 , n42705 );
and ( n42944 , n42941 , n42943 );
xor ( n42945 , n42791 , n42793 );
and ( n42946 , n42943 , n42945 );
and ( n42947 , n42941 , n42945 );
or ( n42948 , n42944 , n42946 , n42947 );
and ( n42949 , n42939 , n42948 );
xor ( n42950 , n42808 , n42809 );
xor ( n42951 , n42950 , n42812 );
xor ( n42952 , n42823 , n42824 );
xor ( n42953 , n42952 , n42827 );
and ( n42954 , n42951 , n42953 );
xor ( n42955 , n42831 , n42836 );
and ( n42956 , n26782 , n41445 );
and ( n42957 , n42955 , n42956 );
and ( n42958 , n42682 , n33632 );
and ( n42959 , n42570 , n33630 );
nor ( n42960 , n42958 , n42959 );
xnor ( n42961 , n42960 , n28124 );
and ( n42962 , n42956 , n42961 );
and ( n42963 , n42955 , n42961 );
or ( n42964 , n42957 , n42962 , n42963 );
and ( n42965 , n27863 , n38737 );
and ( n42966 , n42964 , n42965 );
and ( n42967 , n27591 , n39261 );
and ( n42968 , n42965 , n42967 );
and ( n42969 , n42964 , n42967 );
or ( n42970 , n42966 , n42968 , n42969 );
and ( n42971 , n42953 , n42970 );
and ( n42972 , n42951 , n42970 );
or ( n42973 , n42954 , n42971 , n42972 );
xor ( n42974 , n42801 , n42802 );
xor ( n42975 , n42974 , n42805 );
and ( n42976 , n27389 , n40643 );
and ( n42977 , n26980 , n41038 );
and ( n42978 , n42976 , n42977 );
and ( n42979 , n42570 , n34352 );
and ( n42980 , n42414 , n34350 );
nor ( n42981 , n42979 , n42980 );
xnor ( n42982 , n42981 , n28532 );
and ( n42983 , n42977 , n42982 );
and ( n42984 , n42976 , n42982 );
or ( n42985 , n42978 , n42983 , n42984 );
and ( n42986 , n27962 , n38737 );
and ( n42987 , n42985 , n42986 );
and ( n42988 , n41890 , n34911 );
and ( n42989 , n41631 , n34909 );
nor ( n42990 , n42988 , n42989 );
xnor ( n42991 , n42990 , n34104 );
and ( n42992 , n42986 , n42991 );
and ( n42993 , n42985 , n42991 );
or ( n42994 , n42987 , n42992 , n42993 );
and ( n42995 , n42975 , n42994 );
and ( n42996 , n42414 , n34352 );
and ( n42997 , n42157 , n34350 );
nor ( n42998 , n42996 , n42997 );
xnor ( n42999 , n42998 , n28532 );
and ( n43000 , n26782 , n41908 );
and ( n43001 , n26678 , n42323 );
and ( n43002 , n43000 , n43001 );
and ( n43003 , n26399 , n42621 );
and ( n43004 , n43001 , n43003 );
and ( n43005 , n43000 , n43003 );
or ( n43006 , n43002 , n43004 , n43005 );
and ( n43007 , n42999 , n43006 );
buf ( n43008 , n16310 );
buf ( n43009 , n43008 );
and ( n43010 , n26148 , n43009 );
buf ( n43011 , n25959 );
and ( n43012 , n43010 , n43011 );
and ( n43013 , n40172 , n37197 );
and ( n43014 , n39768 , n37194 );
nor ( n43015 , n43013 , n43014 );
xnor ( n43016 , n43015 , n36218 );
and ( n43017 , n43011 , n43016 );
and ( n43018 , n43010 , n43016 );
or ( n43019 , n43012 , n43017 , n43018 );
and ( n43020 , n43006 , n43019 );
and ( n43021 , n42999 , n43019 );
or ( n43022 , n43007 , n43020 , n43021 );
and ( n43023 , n42994 , n43022 );
and ( n43024 , n42975 , n43022 );
or ( n43025 , n42995 , n43023 , n43024 );
and ( n43026 , n40586 , n36910 );
and ( n43027 , n40178 , n36908 );
nor ( n43028 , n43026 , n43027 );
xnor ( n43029 , n43028 , n36221 );
and ( n43030 , n41012 , n36367 );
and ( n43031 , n40623 , n36365 );
nor ( n43032 , n43030 , n43031 );
xnor ( n43033 , n43032 , n35608 );
and ( n43034 , n43029 , n43033 );
and ( n43035 , n41621 , n35911 );
and ( n43036 , n41405 , n35909 );
nor ( n43037 , n43035 , n43036 );
xnor ( n43038 , n43037 , n35161 );
and ( n43039 , n43033 , n43038 );
and ( n43040 , n43029 , n43038 );
or ( n43041 , n43034 , n43039 , n43040 );
xor ( n43042 , n42838 , n42839 );
xor ( n43043 , n43042 , n42841 );
and ( n43044 , n43041 , n43043 );
xor ( n43045 , n42846 , n42847 );
xor ( n43046 , n43045 , n42849 );
and ( n43047 , n43043 , n43046 );
and ( n43048 , n43041 , n43046 );
or ( n43049 , n43044 , n43047 , n43048 );
xor ( n43050 , n42837 , n42844 );
xor ( n43051 , n43050 , n42852 );
and ( n43052 , n43049 , n43051 );
xor ( n43053 , n42871 , n42873 );
xor ( n43054 , n43053 , n42876 );
and ( n43055 , n43051 , n43054 );
and ( n43056 , n43049 , n43054 );
or ( n43057 , n43052 , n43055 , n43056 );
and ( n43058 , n43025 , n43057 );
xor ( n43059 , n42855 , n42879 );
xor ( n43060 , n43059 , n42890 );
and ( n43061 , n43057 , n43060 );
and ( n43062 , n43025 , n43060 );
or ( n43063 , n43058 , n43061 , n43062 );
and ( n43064 , n42973 , n43063 );
xor ( n43065 , n42797 , n42799 );
xor ( n43066 , n43065 , n42815 );
and ( n43067 , n43063 , n43066 );
and ( n43068 , n42973 , n43066 );
or ( n43069 , n43064 , n43067 , n43068 );
and ( n43070 , n42948 , n43069 );
and ( n43071 , n42939 , n43069 );
or ( n43072 , n42949 , n43070 , n43071 );
and ( n43073 , n42936 , n43072 );
and ( n43074 , n42934 , n43072 );
or ( n43075 , n42937 , n43073 , n43074 );
and ( n43076 , n42932 , n43075 );
xor ( n43077 , n42782 , n42784 );
xor ( n43078 , n43077 , n42918 );
and ( n43079 , n43075 , n43078 );
and ( n43080 , n42932 , n43078 );
or ( n43081 , n43076 , n43079 , n43080 );
xor ( n43082 , n42780 , n42921 );
xor ( n43083 , n43082 , n42924 );
and ( n43084 , n43081 , n43083 );
xor ( n43085 , n42787 , n42821 );
xor ( n43086 , n43085 , n42915 );
xor ( n43087 , n42789 , n42794 );
xor ( n43088 , n43087 , n42818 );
xor ( n43089 , n42907 , n42909 );
xor ( n43090 , n43089 , n42912 );
and ( n43091 , n43088 , n43090 );
xor ( n43092 , n42830 , n42893 );
xor ( n43093 , n43092 , n42904 );
xor ( n43094 , n42896 , n42898 );
xor ( n43095 , n43094 , n42901 );
xor ( n43096 , n42882 , n42884 );
xor ( n43097 , n43096 , n42887 );
xor ( n43098 , n42964 , n42965 );
xor ( n43099 , n43098 , n42967 );
and ( n43100 , n43097 , n43099 );
and ( n43101 , n27591 , n39713 );
and ( n43102 , n27389 , n40196 );
and ( n43103 , n43101 , n43102 );
xor ( n43104 , n42955 , n42956 );
xor ( n43105 , n43104 , n42961 );
and ( n43106 , n43102 , n43105 );
and ( n43107 , n43101 , n43105 );
or ( n43108 , n43103 , n43106 , n43107 );
and ( n43109 , n43099 , n43108 );
and ( n43110 , n43097 , n43108 );
or ( n43111 , n43100 , n43109 , n43110 );
and ( n43112 , n43095 , n43111 );
xor ( n43113 , n42859 , n42863 );
xor ( n43114 , n43113 , n42868 );
xor ( n43115 , n42985 , n42986 );
xor ( n43116 , n43115 , n42991 );
and ( n43117 , n43114 , n43116 );
and ( n43118 , n26678 , n42621 );
and ( n43119 , n26399 , n43009 );
and ( n43120 , n43118 , n43119 );
xor ( n43121 , n33478 , n33553 );
buf ( n43122 , n43121 );
buf ( n43123 , n43122 );
buf ( n43124 , n43123 );
and ( n43125 , n43124 , n33632 );
and ( n43126 , n42835 , n33630 );
nor ( n43127 , n43125 , n43126 );
xnor ( n43128 , n43127 , n28124 );
and ( n43129 , n43119 , n43128 );
and ( n43130 , n43118 , n43128 );
or ( n43131 , n43120 , n43129 , n43130 );
and ( n43132 , n26933 , n41445 );
and ( n43133 , n43131 , n43132 );
and ( n43134 , n42835 , n33632 );
and ( n43135 , n42682 , n33630 );
nor ( n43136 , n43134 , n43135 );
xnor ( n43137 , n43136 , n28124 );
and ( n43138 , n43132 , n43137 );
and ( n43139 , n43131 , n43137 );
or ( n43140 , n43133 , n43138 , n43139 );
and ( n43141 , n43116 , n43140 );
and ( n43142 , n43114 , n43140 );
or ( n43143 , n43117 , n43141 , n43142 );
and ( n43144 , n43124 , n28117 );
xor ( n43145 , n42976 , n42977 );
xor ( n43146 , n43145 , n42982 );
and ( n43147 , n43144 , n43146 );
and ( n43148 , n27962 , n39713 );
and ( n43149 , n27591 , n40643 );
and ( n43150 , n43148 , n43149 );
and ( n43151 , n26933 , n41908 );
and ( n43152 , n43149 , n43151 );
and ( n43153 , n43148 , n43151 );
or ( n43154 , n43150 , n43152 , n43153 );
and ( n43155 , n43146 , n43154 );
and ( n43156 , n43144 , n43154 );
or ( n43157 , n43147 , n43155 , n43156 );
and ( n43158 , n40178 , n37197 );
and ( n43159 , n40172 , n37194 );
nor ( n43160 , n43158 , n43159 );
xnor ( n43161 , n43160 , n36218 );
and ( n43162 , n40623 , n36910 );
and ( n43163 , n40586 , n36908 );
nor ( n43164 , n43162 , n43163 );
xnor ( n43165 , n43164 , n36221 );
and ( n43166 , n43161 , n43165 );
and ( n43167 , n41405 , n36367 );
and ( n43168 , n41012 , n36365 );
nor ( n43169 , n43167 , n43168 );
xnor ( n43170 , n43169 , n35608 );
and ( n43171 , n43165 , n43170 );
and ( n43172 , n43161 , n43170 );
or ( n43173 , n43166 , n43171 , n43172 );
xor ( n43174 , n43000 , n43001 );
xor ( n43175 , n43174 , n43003 );
and ( n43176 , n43173 , n43175 );
xor ( n43177 , n43010 , n43011 );
xor ( n43178 , n43177 , n43016 );
and ( n43179 , n43175 , n43178 );
and ( n43180 , n43173 , n43178 );
or ( n43181 , n43176 , n43179 , n43180 );
and ( n43182 , n43157 , n43181 );
xor ( n43183 , n42999 , n43006 );
xor ( n43184 , n43183 , n43019 );
and ( n43185 , n43181 , n43184 );
and ( n43186 , n43157 , n43184 );
or ( n43187 , n43182 , n43185 , n43186 );
and ( n43188 , n43143 , n43187 );
xor ( n43189 , n42975 , n42994 );
xor ( n43190 , n43189 , n43022 );
and ( n43191 , n43187 , n43190 );
and ( n43192 , n43143 , n43190 );
or ( n43193 , n43188 , n43191 , n43192 );
and ( n43194 , n43111 , n43193 );
and ( n43195 , n43095 , n43193 );
or ( n43196 , n43112 , n43194 , n43195 );
and ( n43197 , n43093 , n43196 );
xor ( n43198 , n42941 , n42943 );
xor ( n43199 , n43198 , n42945 );
and ( n43200 , n43196 , n43199 );
and ( n43201 , n43093 , n43199 );
or ( n43202 , n43197 , n43200 , n43201 );
and ( n43203 , n43090 , n43202 );
and ( n43204 , n43088 , n43202 );
or ( n43205 , n43091 , n43203 , n43204 );
and ( n43206 , n43086 , n43205 );
xor ( n43207 , n42934 , n42936 );
xor ( n43208 , n43207 , n43072 );
and ( n43209 , n43205 , n43208 );
and ( n43210 , n43086 , n43208 );
or ( n43211 , n43206 , n43209 , n43210 );
xor ( n43212 , n42932 , n43075 );
xor ( n43213 , n43212 , n43078 );
and ( n43214 , n43211 , n43213 );
xor ( n43215 , n42939 , n42948 );
xor ( n43216 , n43215 , n43069 );
xor ( n43217 , n42973 , n43063 );
xor ( n43218 , n43217 , n43066 );
xor ( n43219 , n42951 , n42953 );
xor ( n43220 , n43219 , n42970 );
xor ( n43221 , n43025 , n43057 );
xor ( n43222 , n43221 , n43060 );
and ( n43223 , n43220 , n43222 );
xor ( n43224 , n43049 , n43051 );
xor ( n43225 , n43224 , n43054 );
and ( n43226 , n26980 , n41445 );
and ( n43227 , n26782 , n42323 );
and ( n43228 , n43226 , n43227 );
and ( n43229 , n42682 , n34352 );
and ( n43230 , n42570 , n34350 );
nor ( n43231 , n43229 , n43230 );
xnor ( n43232 , n43231 , n28532 );
and ( n43233 , n43227 , n43232 );
and ( n43234 , n43226 , n43232 );
or ( n43235 , n43228 , n43233 , n43234 );
and ( n43236 , n27962 , n39261 );
and ( n43237 , n43235 , n43236 );
and ( n43238 , n27863 , n39713 );
and ( n43239 , n43236 , n43238 );
and ( n43240 , n43235 , n43238 );
or ( n43241 , n43237 , n43239 , n43240 );
and ( n43242 , n26782 , n42621 );
and ( n43243 , n26678 , n43009 );
and ( n43244 , n43242 , n43243 );
xor ( n43245 , n33495 , n33551 );
buf ( n43246 , n43245 );
buf ( n43247 , n43246 );
buf ( n43248 , n43247 );
and ( n43249 , n43248 , n33632 );
and ( n43250 , n43124 , n33630 );
nor ( n43251 , n43249 , n43250 );
xnor ( n43252 , n43251 , n28124 );
and ( n43253 , n43243 , n43252 );
and ( n43254 , n43242 , n43252 );
or ( n43255 , n43244 , n43253 , n43254 );
and ( n43256 , n27389 , n41038 );
and ( n43257 , n43255 , n43256 );
xor ( n43258 , n43118 , n43119 );
xor ( n43259 , n43258 , n43128 );
and ( n43260 , n43256 , n43259 );
and ( n43261 , n43255 , n43259 );
or ( n43262 , n43257 , n43260 , n43261 );
and ( n43263 , n28129 , n38737 );
and ( n43264 , n43262 , n43263 );
and ( n43265 , n41631 , n35374 );
and ( n43266 , n41652 , n35372 );
nor ( n43267 , n43265 , n43266 );
xnor ( n43268 , n43267 , n34661 );
and ( n43269 , n43263 , n43268 );
and ( n43270 , n43262 , n43268 );
or ( n43271 , n43264 , n43269 , n43270 );
and ( n43272 , n43241 , n43271 );
and ( n43273 , n41405 , n35911 );
and ( n43274 , n41012 , n35909 );
nor ( n43275 , n43273 , n43274 );
xnor ( n43276 , n43275 , n35161 );
and ( n43277 , n43271 , n43276 );
and ( n43278 , n43241 , n43276 );
or ( n43279 , n43272 , n43277 , n43278 );
and ( n43280 , n43225 , n43279 );
xor ( n43281 , n43041 , n43043 );
xor ( n43282 , n43281 , n43046 );
xor ( n43283 , n43101 , n43102 );
xor ( n43284 , n43283 , n43105 );
and ( n43285 , n43282 , n43284 );
and ( n43286 , n27591 , n40196 );
and ( n43287 , n42157 , n34911 );
and ( n43288 , n41890 , n34909 );
nor ( n43289 , n43287 , n43288 );
xnor ( n43290 , n43289 , n34104 );
and ( n43291 , n43286 , n43290 );
xor ( n43292 , n43131 , n43132 );
xor ( n43293 , n43292 , n43137 );
and ( n43294 , n43290 , n43293 );
and ( n43295 , n43286 , n43293 );
or ( n43296 , n43291 , n43294 , n43295 );
and ( n43297 , n43284 , n43296 );
and ( n43298 , n43282 , n43296 );
or ( n43299 , n43285 , n43297 , n43298 );
and ( n43300 , n43279 , n43299 );
and ( n43301 , n43225 , n43299 );
or ( n43302 , n43280 , n43300 , n43301 );
and ( n43303 , n43222 , n43302 );
and ( n43304 , n43220 , n43302 );
or ( n43305 , n43223 , n43303 , n43304 );
and ( n43306 , n43218 , n43305 );
xor ( n43307 , n43093 , n43196 );
xor ( n43308 , n43307 , n43199 );
and ( n43309 , n43305 , n43308 );
and ( n43310 , n43218 , n43308 );
or ( n43311 , n43306 , n43309 , n43310 );
and ( n43312 , n43216 , n43311 );
xor ( n43313 , n43088 , n43090 );
xor ( n43314 , n43313 , n43202 );
and ( n43315 , n43311 , n43314 );
and ( n43316 , n43216 , n43314 );
or ( n43317 , n43312 , n43315 , n43316 );
xor ( n43318 , n43086 , n43205 );
xor ( n43319 , n43318 , n43208 );
and ( n43320 , n43317 , n43319 );
xor ( n43321 , n43216 , n43311 );
xor ( n43322 , n43321 , n43314 );
xor ( n43323 , n43029 , n43033 );
xor ( n43324 , n43323 , n43038 );
and ( n43325 , n27389 , n41445 );
and ( n43326 , n26980 , n41908 );
and ( n43327 , n43325 , n43326 );
and ( n43328 , n42835 , n34352 );
and ( n43329 , n42682 , n34350 );
nor ( n43330 , n43328 , n43329 );
xnor ( n43331 , n43330 , n28532 );
and ( n43332 , n43326 , n43331 );
and ( n43333 , n43325 , n43331 );
or ( n43334 , n43327 , n43332 , n43333 );
and ( n43335 , n27863 , n40196 );
and ( n43336 , n43334 , n43335 );
and ( n43337 , n42414 , n34911 );
and ( n43338 , n42157 , n34909 );
nor ( n43339 , n43337 , n43338 );
xnor ( n43340 , n43339 , n34104 );
and ( n43341 , n43335 , n43340 );
and ( n43342 , n43334 , n43340 );
or ( n43343 , n43336 , n43341 , n43342 );
and ( n43344 , n43324 , n43343 );
and ( n43345 , n41890 , n35374 );
and ( n43346 , n41631 , n35372 );
nor ( n43347 , n43345 , n43346 );
xnor ( n43348 , n43347 , n34661 );
and ( n43349 , n43248 , n28117 );
and ( n43350 , n43348 , n43349 );
xor ( n43351 , n43226 , n43227 );
xor ( n43352 , n43351 , n43232 );
and ( n43353 , n43349 , n43352 );
and ( n43354 , n43348 , n43352 );
or ( n43355 , n43350 , n43353 , n43354 );
and ( n43356 , n43343 , n43355 );
and ( n43357 , n43324 , n43355 );
or ( n43358 , n43344 , n43356 , n43357 );
buf ( n43359 , n26148 );
xor ( n43360 , n33511 , n33549 );
buf ( n43361 , n43360 );
buf ( n43362 , n43361 );
buf ( n43363 , n43362 );
and ( n43364 , n43363 , n28117 );
and ( n43365 , n43359 , n43364 );
and ( n43366 , n28129 , n39713 );
and ( n43367 , n27591 , n41038 );
and ( n43368 , n43366 , n43367 );
and ( n43369 , n40586 , n37197 );
and ( n43370 , n40178 , n37194 );
nor ( n43371 , n43369 , n43370 );
xnor ( n43372 , n43371 , n36218 );
and ( n43373 , n43367 , n43372 );
and ( n43374 , n43366 , n43372 );
or ( n43375 , n43368 , n43373 , n43374 );
and ( n43376 , n43365 , n43375 );
and ( n43377 , n41012 , n36910 );
and ( n43378 , n40623 , n36908 );
nor ( n43379 , n43377 , n43378 );
xnor ( n43380 , n43379 , n36221 );
and ( n43381 , n41621 , n36367 );
and ( n43382 , n41405 , n36365 );
nor ( n43383 , n43381 , n43382 );
xnor ( n43384 , n43383 , n35608 );
and ( n43385 , n43380 , n43384 );
and ( n43386 , n42157 , n35374 );
and ( n43387 , n41890 , n35372 );
nor ( n43388 , n43386 , n43387 );
xnor ( n43389 , n43388 , n34661 );
and ( n43390 , n43384 , n43389 );
and ( n43391 , n43380 , n43389 );
or ( n43392 , n43385 , n43390 , n43391 );
and ( n43393 , n43375 , n43392 );
and ( n43394 , n43365 , n43392 );
or ( n43395 , n43376 , n43393 , n43394 );
xor ( n43396 , n43144 , n43146 );
xor ( n43397 , n43396 , n43154 );
and ( n43398 , n43395 , n43397 );
xor ( n43399 , n43173 , n43175 );
xor ( n43400 , n43399 , n43178 );
and ( n43401 , n43397 , n43400 );
and ( n43402 , n43395 , n43400 );
or ( n43403 , n43398 , n43401 , n43402 );
and ( n43404 , n43358 , n43403 );
xor ( n43405 , n43114 , n43116 );
xor ( n43406 , n43405 , n43140 );
and ( n43407 , n43403 , n43406 );
and ( n43408 , n43358 , n43406 );
or ( n43409 , n43404 , n43407 , n43408 );
xor ( n43410 , n43097 , n43099 );
xor ( n43411 , n43410 , n43108 );
and ( n43412 , n43409 , n43411 );
xor ( n43413 , n43143 , n43187 );
xor ( n43414 , n43413 , n43190 );
and ( n43415 , n43411 , n43414 );
and ( n43416 , n43409 , n43414 );
or ( n43417 , n43412 , n43415 , n43416 );
xor ( n43418 , n43095 , n43111 );
xor ( n43419 , n43418 , n43193 );
and ( n43420 , n43417 , n43419 );
and ( n43421 , n39768 , n37197 );
and ( n43422 , n39759 , n37194 );
nor ( n43423 , n43421 , n43422 );
xnor ( n43424 , n43423 , n36218 );
xor ( n43425 , n43241 , n43271 );
xor ( n43426 , n43425 , n43276 );
and ( n43427 , n43424 , n43426 );
xor ( n43428 , n43157 , n43181 );
xor ( n43429 , n43428 , n43184 );
xor ( n43430 , n43262 , n43263 );
xor ( n43431 , n43430 , n43268 );
and ( n43432 , n41652 , n35911 );
and ( n43433 , n41621 , n35909 );
nor ( n43434 , n43432 , n43433 );
xnor ( n43435 , n43434 , n35161 );
xor ( n43436 , n43334 , n43335 );
xor ( n43437 , n43436 , n43340 );
and ( n43438 , n43435 , n43437 );
and ( n43439 , n43431 , n43438 );
xor ( n43440 , n43148 , n43149 );
xor ( n43441 , n43440 , n43151 );
xor ( n43442 , n43161 , n43165 );
xor ( n43443 , n43442 , n43170 );
and ( n43444 , n43441 , n43443 );
buf ( n43445 , n16538 );
buf ( n43446 , n43445 );
and ( n43447 , n26399 , n43446 );
xor ( n43448 , n43359 , n43364 );
and ( n43449 , n43447 , n43448 );
and ( n43450 , n43443 , n43449 );
and ( n43451 , n43441 , n43449 );
or ( n43452 , n43444 , n43450 , n43451 );
and ( n43453 , n43438 , n43452 );
and ( n43454 , n43431 , n43452 );
or ( n43455 , n43439 , n43453 , n43454 );
and ( n43456 , n43429 , n43455 );
xor ( n43457 , n43242 , n43243 );
xor ( n43458 , n43457 , n43252 );
xor ( n43459 , n43325 , n43326 );
xor ( n43460 , n43459 , n43331 );
and ( n43461 , n43458 , n43460 );
and ( n43462 , n27962 , n40643 );
and ( n43463 , n27863 , n41038 );
and ( n43464 , n43462 , n43463 );
and ( n43465 , n27591 , n41445 );
and ( n43466 , n43463 , n43465 );
and ( n43467 , n43462 , n43465 );
or ( n43468 , n43464 , n43466 , n43467 );
and ( n43469 , n43460 , n43468 );
and ( n43470 , n43458 , n43468 );
or ( n43471 , n43461 , n43469 , n43470 );
and ( n43472 , n26782 , n43009 );
and ( n43473 , n40623 , n37197 );
and ( n43474 , n40586 , n37194 );
nor ( n43475 , n43473 , n43474 );
xnor ( n43476 , n43475 , n36218 );
and ( n43477 , n43472 , n43476 );
and ( n43478 , n41405 , n36910 );
and ( n43479 , n41012 , n36908 );
nor ( n43480 , n43478 , n43479 );
xnor ( n43481 , n43480 , n36221 );
and ( n43482 , n43476 , n43481 );
and ( n43483 , n43472 , n43481 );
or ( n43484 , n43477 , n43482 , n43483 );
and ( n43485 , n41652 , n36367 );
and ( n43486 , n41621 , n36365 );
nor ( n43487 , n43485 , n43486 );
xnor ( n43488 , n43487 , n35608 );
and ( n43489 , n41890 , n35911 );
and ( n43490 , n41631 , n35909 );
nor ( n43491 , n43489 , n43490 );
xnor ( n43492 , n43491 , n35161 );
and ( n43493 , n43488 , n43492 );
and ( n43494 , n42682 , n34911 );
and ( n43495 , n42570 , n34909 );
nor ( n43496 , n43494 , n43495 );
xnor ( n43497 , n43496 , n34104 );
and ( n43498 , n43492 , n43497 );
and ( n43499 , n43488 , n43497 );
or ( n43500 , n43493 , n43498 , n43499 );
and ( n43501 , n43484 , n43500 );
xor ( n43502 , n43366 , n43367 );
xor ( n43503 , n43502 , n43372 );
and ( n43504 , n43500 , n43503 );
and ( n43505 , n43484 , n43503 );
or ( n43506 , n43501 , n43504 , n43505 );
and ( n43507 , n43471 , n43506 );
xor ( n43508 , n43348 , n43349 );
xor ( n43509 , n43508 , n43352 );
and ( n43510 , n43506 , n43509 );
and ( n43511 , n43471 , n43509 );
or ( n43512 , n43507 , n43510 , n43511 );
xor ( n43513 , n43324 , n43343 );
xor ( n43514 , n43513 , n43355 );
and ( n43515 , n43512 , n43514 );
xor ( n43516 , n43395 , n43397 );
xor ( n43517 , n43516 , n43400 );
and ( n43518 , n43514 , n43517 );
and ( n43519 , n43512 , n43517 );
or ( n43520 , n43515 , n43518 , n43519 );
and ( n43521 , n43455 , n43520 );
and ( n43522 , n43429 , n43520 );
or ( n43523 , n43456 , n43521 , n43522 );
and ( n43524 , n43427 , n43523 );
xor ( n43525 , n43225 , n43279 );
xor ( n43526 , n43525 , n43299 );
and ( n43527 , n43523 , n43526 );
and ( n43528 , n43427 , n43526 );
or ( n43529 , n43524 , n43527 , n43528 );
and ( n43530 , n43419 , n43529 );
and ( n43531 , n43417 , n43529 );
or ( n43532 , n43420 , n43530 , n43531 );
xor ( n43533 , n43218 , n43305 );
xor ( n43534 , n43533 , n43308 );
and ( n43535 , n43532 , n43534 );
xor ( n43536 , n43220 , n43222 );
xor ( n43537 , n43536 , n43302 );
xor ( n43538 , n43409 , n43411 );
xor ( n43539 , n43538 , n43414 );
xor ( n43540 , n43282 , n43284 );
xor ( n43541 , n43540 , n43296 );
xor ( n43542 , n43358 , n43403 );
xor ( n43543 , n43542 , n43406 );
and ( n43544 , n43541 , n43543 );
xor ( n43545 , n43424 , n43426 );
and ( n43546 , n43543 , n43545 );
and ( n43547 , n43541 , n43545 );
or ( n43548 , n43544 , n43546 , n43547 );
and ( n43549 , n43539 , n43548 );
and ( n43550 , n26980 , n42323 );
and ( n43551 , n26933 , n42621 );
and ( n43552 , n43550 , n43551 );
and ( n43553 , n26678 , n43446 );
and ( n43554 , n43363 , n33632 );
and ( n43555 , n43248 , n33630 );
nor ( n43556 , n43554 , n43555 );
xnor ( n43557 , n43556 , n28124 );
xor ( n43558 , n43553 , n43557 );
xor ( n43559 , n33527 , n33547 );
buf ( n43560 , n43559 );
buf ( n43561 , n43560 );
buf ( n43562 , n43561 );
and ( n43563 , n43562 , n28117 );
xor ( n43564 , n43558 , n43563 );
and ( n43565 , n43551 , n43564 );
and ( n43566 , n43550 , n43564 );
or ( n43567 , n43552 , n43565 , n43566 );
and ( n43568 , n27863 , n40643 );
and ( n43569 , n43567 , n43568 );
and ( n43570 , n42570 , n34911 );
and ( n43571 , n42414 , n34909 );
nor ( n43572 , n43570 , n43571 );
xnor ( n43573 , n43572 , n34104 );
and ( n43574 , n43568 , n43573 );
and ( n43575 , n43567 , n43573 );
or ( n43576 , n43569 , n43574 , n43575 );
and ( n43577 , n28129 , n39261 );
and ( n43578 , n43576 , n43577 );
xor ( n43579 , n43255 , n43256 );
xor ( n43580 , n43579 , n43259 );
and ( n43581 , n43577 , n43580 );
and ( n43582 , n43576 , n43580 );
or ( n43583 , n43578 , n43581 , n43582 );
xor ( n43584 , n43235 , n43236 );
xor ( n43585 , n43584 , n43238 );
and ( n43586 , n43583 , n43585 );
xor ( n43587 , n43286 , n43290 );
xor ( n43588 , n43587 , n43293 );
and ( n43589 , n43585 , n43588 );
and ( n43590 , n43583 , n43588 );
or ( n43591 , n43586 , n43589 , n43590 );
xor ( n43592 , n43365 , n43375 );
xor ( n43593 , n43592 , n43392 );
xor ( n43594 , n43435 , n43437 );
and ( n43595 , n43593 , n43594 );
xor ( n43596 , n43447 , n43448 );
and ( n43597 , n43553 , n43557 );
and ( n43598 , n43557 , n43563 );
and ( n43599 , n43553 , n43563 );
or ( n43600 , n43597 , n43598 , n43599 );
and ( n43601 , n43596 , n43600 );
and ( n43602 , n26933 , n42323 );
and ( n43603 , n43600 , n43602 );
and ( n43604 , n43596 , n43602 );
or ( n43605 , n43601 , n43603 , n43604 );
and ( n43606 , n43594 , n43605 );
and ( n43607 , n43593 , n43605 );
or ( n43608 , n43595 , n43606 , n43607 );
xor ( n43609 , n43380 , n43384 );
xor ( n43610 , n43609 , n43389 );
and ( n43611 , n43124 , n34352 );
and ( n43612 , n42835 , n34350 );
nor ( n43613 , n43611 , n43612 );
xnor ( n43614 , n43613 , n28532 );
buf ( n43615 , n26399 );
xor ( n43616 , n33534 , n33545 );
buf ( n43617 , n43616 );
buf ( n43618 , n43617 );
buf ( n43619 , n43618 );
and ( n43620 , n43619 , n28117 );
and ( n43621 , n43615 , n43620 );
and ( n43622 , n43614 , n43621 );
and ( n43623 , n28129 , n40643 );
and ( n43624 , n27962 , n41038 );
and ( n43625 , n43623 , n43624 );
and ( n43626 , n27389 , n42323 );
and ( n43627 , n43624 , n43626 );
and ( n43628 , n43623 , n43626 );
or ( n43629 , n43625 , n43627 , n43628 );
and ( n43630 , n43621 , n43629 );
and ( n43631 , n43614 , n43629 );
or ( n43632 , n43622 , n43630 , n43631 );
and ( n43633 , n43610 , n43632 );
and ( n43634 , n26980 , n42621 );
and ( n43635 , n41012 , n37197 );
and ( n43636 , n40623 , n37194 );
nor ( n43637 , n43635 , n43636 );
xnor ( n43638 , n43637 , n36218 );
and ( n43639 , n43634 , n43638 );
and ( n43640 , n41621 , n36910 );
and ( n43641 , n41405 , n36908 );
nor ( n43642 , n43640 , n43641 );
xnor ( n43643 , n43642 , n36221 );
and ( n43644 , n43638 , n43643 );
and ( n43645 , n43634 , n43643 );
or ( n43646 , n43639 , n43644 , n43645 );
xor ( n43647 , n43462 , n43463 );
xor ( n43648 , n43647 , n43465 );
and ( n43649 , n43646 , n43648 );
xor ( n43650 , n43472 , n43476 );
xor ( n43651 , n43650 , n43481 );
and ( n43652 , n43648 , n43651 );
and ( n43653 , n43646 , n43651 );
or ( n43654 , n43649 , n43652 , n43653 );
and ( n43655 , n43632 , n43654 );
and ( n43656 , n43610 , n43654 );
or ( n43657 , n43633 , n43655 , n43656 );
xor ( n43658 , n43441 , n43443 );
xor ( n43659 , n43658 , n43449 );
and ( n43660 , n43657 , n43659 );
xor ( n43661 , n43471 , n43506 );
xor ( n43662 , n43661 , n43509 );
and ( n43663 , n43659 , n43662 );
and ( n43664 , n43657 , n43662 );
or ( n43665 , n43660 , n43663 , n43664 );
and ( n43666 , n43608 , n43665 );
xor ( n43667 , n43431 , n43438 );
xor ( n43668 , n43667 , n43452 );
and ( n43669 , n43665 , n43668 );
and ( n43670 , n43608 , n43668 );
or ( n43671 , n43666 , n43669 , n43670 );
and ( n43672 , n43591 , n43671 );
xor ( n43673 , n43429 , n43455 );
xor ( n43674 , n43673 , n43520 );
and ( n43675 , n43671 , n43674 );
and ( n43676 , n43591 , n43674 );
or ( n43677 , n43672 , n43675 , n43676 );
and ( n43678 , n43548 , n43677 );
and ( n43679 , n43539 , n43677 );
or ( n43680 , n43549 , n43678 , n43679 );
and ( n43681 , n43537 , n43680 );
xor ( n43682 , n43417 , n43419 );
xor ( n43683 , n43682 , n43529 );
and ( n43684 , n43680 , n43683 );
and ( n43685 , n43537 , n43683 );
or ( n43686 , n43681 , n43684 , n43685 );
and ( n43687 , n43534 , n43686 );
and ( n43688 , n43532 , n43686 );
or ( n43689 , n43535 , n43687 , n43688 );
and ( n43690 , n43322 , n43689 );
xor ( n43691 , n43532 , n43534 );
xor ( n43692 , n43691 , n43686 );
xor ( n43693 , n43427 , n43523 );
xor ( n43694 , n43693 , n43526 );
xor ( n43695 , n43512 , n43514 );
xor ( n43696 , n43695 , n43517 );
xor ( n43697 , n43583 , n43585 );
xor ( n43698 , n43697 , n43588 );
and ( n43699 , n43696 , n43698 );
xor ( n43700 , n43576 , n43577 );
xor ( n43701 , n43700 , n43580 );
and ( n43702 , n27863 , n41445 );
and ( n43703 , n27591 , n41908 );
and ( n43704 , n43702 , n43703 );
and ( n43705 , n42835 , n34911 );
and ( n43706 , n42682 , n34909 );
nor ( n43707 , n43705 , n43706 );
xnor ( n43708 , n43707 , n34104 );
and ( n43709 , n43703 , n43708 );
and ( n43710 , n43702 , n43708 );
or ( n43711 , n43704 , n43709 , n43710 );
and ( n43712 , n28129 , n40196 );
and ( n43713 , n43711 , n43712 );
xor ( n43714 , n43550 , n43551 );
xor ( n43715 , n43714 , n43564 );
and ( n43716 , n43712 , n43715 );
and ( n43717 , n43711 , n43715 );
or ( n43718 , n43713 , n43716 , n43717 );
and ( n43719 , n41631 , n35911 );
and ( n43720 , n41652 , n35909 );
nor ( n43721 , n43719 , n43720 );
xnor ( n43722 , n43721 , n35161 );
and ( n43723 , n43718 , n43722 );
xor ( n43724 , n43567 , n43568 );
xor ( n43725 , n43724 , n43573 );
and ( n43726 , n43722 , n43725 );
and ( n43727 , n43718 , n43725 );
or ( n43728 , n43723 , n43726 , n43727 );
and ( n43729 , n43701 , n43728 );
xor ( n43730 , n43458 , n43460 );
xor ( n43731 , n43730 , n43468 );
xor ( n43732 , n43484 , n43500 );
xor ( n43733 , n43732 , n43503 );
and ( n43734 , n43731 , n43733 );
xor ( n43735 , n43488 , n43492 );
xor ( n43736 , n43735 , n43497 );
buf ( n43737 , n16732 );
buf ( n43738 , n43737 );
and ( n43739 , n26678 , n43738 );
not ( n43740 , n43739 );
xor ( n43741 , n43615 , n43620 );
and ( n43742 , n43740 , n43741 );
and ( n43743 , n43736 , n43742 );
buf ( n43744 , n43739 );
and ( n43745 , n43742 , n43744 );
and ( n43746 , n43736 , n43744 );
or ( n43747 , n43743 , n43745 , n43746 );
and ( n43748 , n43733 , n43747 );
and ( n43749 , n43731 , n43747 );
or ( n43750 , n43734 , n43748 , n43749 );
and ( n43751 , n43728 , n43750 );
and ( n43752 , n43701 , n43750 );
or ( n43753 , n43729 , n43751 , n43752 );
and ( n43754 , n43698 , n43753 );
and ( n43755 , n43696 , n43753 );
or ( n43756 , n43699 , n43754 , n43755 );
xor ( n43757 , n43541 , n43543 );
xor ( n43758 , n43757 , n43545 );
and ( n43759 , n43756 , n43758 );
xor ( n43760 , n43591 , n43671 );
xor ( n43761 , n43760 , n43674 );
and ( n43762 , n43758 , n43761 );
and ( n43763 , n43756 , n43761 );
or ( n43764 , n43759 , n43762 , n43763 );
and ( n43765 , n43694 , n43764 );
xor ( n43766 , n43539 , n43548 );
xor ( n43767 , n43766 , n43677 );
and ( n43768 , n43764 , n43767 );
and ( n43769 , n43694 , n43767 );
or ( n43770 , n43765 , n43768 , n43769 );
xor ( n43771 , n43537 , n43680 );
xor ( n43772 , n43771 , n43683 );
and ( n43773 , n43770 , n43772 );
xor ( n43774 , n43694 , n43764 );
xor ( n43775 , n43774 , n43767 );
xor ( n43776 , n43608 , n43665 );
xor ( n43777 , n43776 , n43668 );
xor ( n43778 , n43593 , n43594 );
xor ( n43779 , n43778 , n43605 );
xor ( n43780 , n43657 , n43659 );
xor ( n43781 , n43780 , n43662 );
and ( n43782 , n43779 , n43781 );
and ( n43783 , n26782 , n43446 );
and ( n43784 , n43248 , n34352 );
and ( n43785 , n43124 , n34350 );
nor ( n43786 , n43784 , n43785 );
xnor ( n43787 , n43786 , n28532 );
and ( n43788 , n43783 , n43787 );
and ( n43789 , n43562 , n33632 );
and ( n43790 , n43363 , n33630 );
nor ( n43791 , n43789 , n43790 );
xnor ( n43792 , n43791 , n28124 );
and ( n43793 , n43787 , n43792 );
and ( n43794 , n43783 , n43792 );
or ( n43795 , n43788 , n43793 , n43794 );
and ( n43796 , n26782 , n43738 );
and ( n43797 , n43619 , n33632 );
and ( n43798 , n43562 , n33630 );
nor ( n43799 , n43797 , n43798 );
xnor ( n43800 , n43799 , n28124 );
and ( n43801 , n43796 , n43800 );
xor ( n43802 , n33540 , n33543 );
buf ( n43803 , n43802 );
buf ( n43804 , n43803 );
buf ( n43805 , n43804 );
and ( n43806 , n43805 , n28117 );
and ( n43807 , n43800 , n43806 );
and ( n43808 , n43796 , n43806 );
or ( n43809 , n43801 , n43807 , n43808 );
and ( n43810 , n26933 , n43009 );
and ( n43811 , n43809 , n43810 );
xor ( n43812 , n43740 , n43741 );
not ( n43813 , n43812 );
and ( n43814 , n43810 , n43813 );
and ( n43815 , n43809 , n43813 );
or ( n43816 , n43811 , n43814 , n43815 );
and ( n43817 , n43795 , n43816 );
and ( n43818 , n27389 , n41908 );
and ( n43819 , n43816 , n43818 );
and ( n43820 , n43795 , n43818 );
or ( n43821 , n43817 , n43819 , n43820 );
and ( n43822 , n27962 , n40196 );
and ( n43823 , n43821 , n43822 );
xor ( n43824 , n43596 , n43600 );
xor ( n43825 , n43824 , n43602 );
and ( n43826 , n43822 , n43825 );
and ( n43827 , n43821 , n43825 );
or ( n43828 , n43823 , n43826 , n43827 );
and ( n43829 , n43781 , n43828 );
and ( n43830 , n43779 , n43828 );
or ( n43831 , n43782 , n43829 , n43830 );
and ( n43832 , n43777 , n43831 );
and ( n43833 , n41631 , n36367 );
and ( n43834 , n41652 , n36365 );
nor ( n43835 , n43833 , n43834 );
xnor ( n43836 , n43835 , n35608 );
and ( n43837 , n42570 , n35374 );
and ( n43838 , n42414 , n35372 );
nor ( n43839 , n43837 , n43838 );
xnor ( n43840 , n43839 , n34661 );
and ( n43841 , n43836 , n43840 );
xor ( n43842 , n43783 , n43787 );
xor ( n43843 , n43842 , n43792 );
and ( n43844 , n43840 , n43843 );
and ( n43845 , n43836 , n43843 );
or ( n43846 , n43841 , n43844 , n43845 );
xor ( n43847 , n43702 , n43703 );
xor ( n43848 , n43847 , n43708 );
and ( n43849 , n27863 , n41908 );
and ( n43850 , n27591 , n42323 );
and ( n43851 , n43849 , n43850 );
and ( n43852 , n43848 , n43851 );
and ( n43853 , n27389 , n42621 );
and ( n43854 , n43124 , n34911 );
and ( n43855 , n42835 , n34909 );
nor ( n43856 , n43854 , n43855 );
xnor ( n43857 , n43856 , n34104 );
and ( n43858 , n43853 , n43857 );
and ( n43859 , n43851 , n43858 );
and ( n43860 , n43848 , n43858 );
or ( n43861 , n43852 , n43859 , n43860 );
and ( n43862 , n43846 , n43861 );
and ( n43863 , n26980 , n43009 );
and ( n43864 , n26933 , n43446 );
and ( n43865 , n43863 , n43864 );
and ( n43866 , n41405 , n37197 );
and ( n43867 , n41012 , n37194 );
nor ( n43868 , n43866 , n43867 );
xnor ( n43869 , n43868 , n36218 );
and ( n43870 , n43864 , n43869 );
and ( n43871 , n43863 , n43869 );
or ( n43872 , n43865 , n43870 , n43871 );
and ( n43873 , n41652 , n36910 );
and ( n43874 , n41621 , n36908 );
nor ( n43875 , n43873 , n43874 );
xnor ( n43876 , n43875 , n36221 );
and ( n43877 , n41890 , n36367 );
and ( n43878 , n41631 , n36365 );
nor ( n43879 , n43877 , n43878 );
xnor ( n43880 , n43879 , n35608 );
and ( n43881 , n43876 , n43880 );
and ( n43882 , n42414 , n35911 );
and ( n43883 , n42157 , n35909 );
nor ( n43884 , n43882 , n43883 );
xnor ( n43885 , n43884 , n35161 );
and ( n43886 , n43880 , n43885 );
and ( n43887 , n43876 , n43885 );
or ( n43888 , n43881 , n43886 , n43887 );
and ( n43889 , n43872 , n43888 );
xor ( n43890 , n43623 , n43624 );
xor ( n43891 , n43890 , n43626 );
and ( n43892 , n43888 , n43891 );
and ( n43893 , n43872 , n43891 );
or ( n43894 , n43889 , n43892 , n43893 );
and ( n43895 , n43861 , n43894 );
and ( n43896 , n43846 , n43894 );
or ( n43897 , n43862 , n43895 , n43896 );
xor ( n43898 , n43610 , n43632 );
xor ( n43899 , n43898 , n43654 );
and ( n43900 , n43897 , n43899 );
xor ( n43901 , n43718 , n43722 );
xor ( n43902 , n43901 , n43725 );
and ( n43903 , n43899 , n43902 );
and ( n43904 , n43897 , n43902 );
or ( n43905 , n43900 , n43903 , n43904 );
xor ( n43906 , n43614 , n43621 );
xor ( n43907 , n43906 , n43629 );
xor ( n43908 , n43646 , n43648 );
xor ( n43909 , n43908 , n43651 );
and ( n43910 , n43907 , n43909 );
xor ( n43911 , n43711 , n43712 );
xor ( n43912 , n43911 , n43715 );
and ( n43913 , n43909 , n43912 );
and ( n43914 , n43907 , n43912 );
or ( n43915 , n43910 , n43913 , n43914 );
buf ( n43916 , n43812 );
xor ( n43917 , n43634 , n43638 );
xor ( n43918 , n43917 , n43643 );
and ( n43919 , n42682 , n35374 );
and ( n43920 , n42570 , n35372 );
nor ( n43921 , n43919 , n43920 );
xnor ( n43922 , n43921 , n34661 );
and ( n43923 , n43363 , n34352 );
and ( n43924 , n43248 , n34350 );
nor ( n43925 , n43923 , n43924 );
xnor ( n43926 , n43925 , n28532 );
and ( n43927 , n43922 , n43926 );
xor ( n43928 , n43796 , n43800 );
xor ( n43929 , n43928 , n43806 );
and ( n43930 , n43926 , n43929 );
and ( n43931 , n43922 , n43929 );
or ( n43932 , n43927 , n43930 , n43931 );
and ( n43933 , n43918 , n43932 );
xor ( n43934 , n43849 , n43850 );
xor ( n43935 , n43853 , n43857 );
and ( n43936 , n43934 , n43935 );
and ( n43937 , n28129 , n41445 );
and ( n43938 , n27962 , n41908 );
and ( n43939 , n43937 , n43938 );
and ( n43940 , n27863 , n42323 );
and ( n43941 , n43938 , n43940 );
and ( n43942 , n43937 , n43940 );
or ( n43943 , n43939 , n43941 , n43942 );
and ( n43944 , n43935 , n43943 );
and ( n43945 , n43934 , n43943 );
or ( n43946 , n43936 , n43944 , n43945 );
and ( n43947 , n43932 , n43946 );
and ( n43948 , n43918 , n43946 );
or ( n43949 , n43933 , n43947 , n43948 );
and ( n43950 , n43916 , n43949 );
and ( n43951 , n27591 , n42621 );
and ( n43952 , n26980 , n43446 );
and ( n43953 , n43951 , n43952 );
and ( n43954 , n26933 , n43738 );
and ( n43955 , n43952 , n43954 );
and ( n43956 , n43951 , n43954 );
or ( n43957 , n43953 , n43955 , n43956 );
buf ( n43958 , n16750 );
buf ( n43959 , n43958 );
and ( n43960 , n26782 , n43959 );
buf ( n43961 , n26678 );
and ( n43962 , n43960 , n43961 );
and ( n43963 , n41621 , n37197 );
and ( n43964 , n41405 , n37194 );
nor ( n43965 , n43963 , n43964 );
xnor ( n43966 , n43965 , n36218 );
and ( n43967 , n43961 , n43966 );
and ( n43968 , n43960 , n43966 );
or ( n43969 , n43962 , n43967 , n43968 );
and ( n43970 , n43957 , n43969 );
and ( n43971 , n41631 , n36910 );
and ( n43972 , n41652 , n36908 );
nor ( n43973 , n43971 , n43972 );
xnor ( n43974 , n43973 , n36221 );
and ( n43975 , n42157 , n36367 );
and ( n43976 , n41890 , n36365 );
nor ( n43977 , n43975 , n43976 );
xnor ( n43978 , n43977 , n35608 );
and ( n43979 , n43974 , n43978 );
and ( n43980 , n42570 , n35911 );
and ( n43981 , n42414 , n35909 );
nor ( n43982 , n43980 , n43981 );
xnor ( n43983 , n43982 , n35161 );
and ( n43984 , n43978 , n43983 );
and ( n43985 , n43974 , n43983 );
or ( n43986 , n43979 , n43984 , n43985 );
and ( n43987 , n43969 , n43986 );
and ( n43988 , n43957 , n43986 );
or ( n43989 , n43970 , n43987 , n43988 );
and ( n43990 , n42835 , n35374 );
and ( n43991 , n42682 , n35372 );
nor ( n43992 , n43990 , n43991 );
xnor ( n43993 , n43992 , n34661 );
and ( n43994 , n43562 , n34352 );
and ( n43995 , n43363 , n34350 );
nor ( n43996 , n43994 , n43995 );
xnor ( n43997 , n43996 , n28532 );
and ( n43998 , n43993 , n43997 );
and ( n43999 , n43805 , n33632 );
and ( n44000 , n43619 , n33630 );
nor ( n44001 , n43999 , n44000 );
xnor ( n44002 , n44001 , n28124 );
and ( n44003 , n43997 , n44002 );
and ( n44004 , n43993 , n44002 );
or ( n44005 , n43998 , n44003 , n44004 );
xor ( n44006 , n43863 , n43864 );
xor ( n44007 , n44006 , n43869 );
and ( n44008 , n44005 , n44007 );
xor ( n44009 , n43876 , n43880 );
xor ( n44010 , n44009 , n43885 );
and ( n44011 , n44007 , n44010 );
and ( n44012 , n44005 , n44010 );
or ( n44013 , n44008 , n44011 , n44012 );
and ( n44014 , n43989 , n44013 );
xor ( n44015 , n43836 , n43840 );
xor ( n44016 , n44015 , n43843 );
and ( n44017 , n44013 , n44016 );
and ( n44018 , n43989 , n44016 );
or ( n44019 , n44014 , n44017 , n44018 );
and ( n44020 , n43949 , n44019 );
and ( n44021 , n43916 , n44019 );
or ( n44022 , n43950 , n44020 , n44021 );
and ( n44023 , n43915 , n44022 );
xor ( n44024 , n43731 , n43733 );
xor ( n44025 , n44024 , n43747 );
and ( n44026 , n44022 , n44025 );
and ( n44027 , n43915 , n44025 );
or ( n44028 , n44023 , n44026 , n44027 );
and ( n44029 , n43905 , n44028 );
xor ( n44030 , n43701 , n43728 );
xor ( n44031 , n44030 , n43750 );
and ( n44032 , n44028 , n44031 );
and ( n44033 , n43905 , n44031 );
or ( n44034 , n44029 , n44032 , n44033 );
and ( n44035 , n43831 , n44034 );
and ( n44036 , n43777 , n44034 );
or ( n44037 , n43832 , n44035 , n44036 );
xor ( n44038 , n43756 , n43758 );
xor ( n44039 , n44038 , n43761 );
and ( n44040 , n44037 , n44039 );
xor ( n44041 , n43696 , n43698 );
xor ( n44042 , n44041 , n43753 );
xor ( n44043 , n43821 , n43822 );
xor ( n44044 , n44043 , n43825 );
and ( n44045 , n42414 , n35374 );
and ( n44046 , n42157 , n35372 );
nor ( n44047 , n44045 , n44046 );
xnor ( n44048 , n44047 , n34661 );
xor ( n44049 , n43795 , n43816 );
xor ( n44050 , n44049 , n43818 );
and ( n44051 , n44048 , n44050 );
and ( n44052 , n44044 , n44051 );
xor ( n44053 , n43736 , n43742 );
xor ( n44054 , n44053 , n43744 );
xor ( n44055 , n43846 , n43861 );
xor ( n44056 , n44055 , n43894 );
and ( n44057 , n44054 , n44056 );
xor ( n44058 , n43848 , n43851 );
xor ( n44059 , n44058 , n43858 );
xor ( n44060 , n43872 , n43888 );
xor ( n44061 , n44060 , n43891 );
and ( n44062 , n44059 , n44061 );
xor ( n44063 , n43809 , n43810 );
xor ( n44064 , n44063 , n43813 );
and ( n44065 , n44061 , n44064 );
and ( n44066 , n44059 , n44064 );
or ( n44067 , n44062 , n44065 , n44066 );
and ( n44068 , n44056 , n44067 );
and ( n44069 , n44054 , n44067 );
or ( n44070 , n44057 , n44068 , n44069 );
and ( n44071 , n44051 , n44070 );
and ( n44072 , n44044 , n44070 );
or ( n44073 , n44052 , n44071 , n44072 );
xor ( n44074 , n33514 , n33542 );
buf ( n44075 , n44074 );
buf ( n44076 , n44075 );
buf ( n44077 , n44076 );
and ( n44078 , n44077 , n28117 );
and ( n44079 , n44077 , n33630 );
not ( n44080 , n44079 );
and ( n44081 , n44080 , n28124 );
and ( n44082 , n44077 , n33632 );
and ( n44083 , n43805 , n33630 );
nor ( n44084 , n44082 , n44083 );
xnor ( n44085 , n44084 , n28124 );
and ( n44086 , n44081 , n44085 );
and ( n44087 , n44078 , n44086 );
and ( n44088 , n28129 , n41908 );
and ( n44089 , n27962 , n42323 );
and ( n44090 , n44088 , n44089 );
and ( n44091 , n27863 , n42621 );
and ( n44092 , n44089 , n44091 );
and ( n44093 , n44088 , n44091 );
or ( n44094 , n44090 , n44092 , n44093 );
and ( n44095 , n44086 , n44094 );
and ( n44096 , n44078 , n44094 );
or ( n44097 , n44087 , n44095 , n44096 );
and ( n44098 , n27591 , n43009 );
and ( n44099 , n27389 , n43446 );
and ( n44100 , n44098 , n44099 );
and ( n44101 , n26980 , n43738 );
and ( n44102 , n44099 , n44101 );
and ( n44103 , n44098 , n44101 );
or ( n44104 , n44100 , n44102 , n44103 );
and ( n44105 , n41652 , n37197 );
and ( n44106 , n41621 , n37194 );
nor ( n44107 , n44105 , n44106 );
xnor ( n44108 , n44107 , n36218 );
and ( n44109 , n41890 , n36910 );
and ( n44110 , n41631 , n36908 );
nor ( n44111 , n44109 , n44110 );
xnor ( n44112 , n44111 , n36221 );
and ( n44113 , n44108 , n44112 );
and ( n44114 , n42414 , n36367 );
and ( n44115 , n42157 , n36365 );
nor ( n44116 , n44114 , n44115 );
xnor ( n44117 , n44116 , n35608 );
and ( n44118 , n44112 , n44117 );
and ( n44119 , n44108 , n44117 );
or ( n44120 , n44113 , n44118 , n44119 );
and ( n44121 , n44104 , n44120 );
and ( n44122 , n42682 , n35911 );
and ( n44123 , n42570 , n35909 );
nor ( n44124 , n44122 , n44123 );
xnor ( n44125 , n44124 , n35161 );
and ( n44126 , n43124 , n35374 );
and ( n44127 , n42835 , n35372 );
nor ( n44128 , n44126 , n44127 );
xnor ( n44129 , n44128 , n34661 );
and ( n44130 , n44125 , n44129 );
and ( n44131 , n43363 , n34911 );
and ( n44132 , n43248 , n34909 );
nor ( n44133 , n44131 , n44132 );
xnor ( n44134 , n44133 , n34104 );
and ( n44135 , n44129 , n44134 );
and ( n44136 , n44125 , n44134 );
or ( n44137 , n44130 , n44135 , n44136 );
and ( n44138 , n44120 , n44137 );
and ( n44139 , n44104 , n44137 );
or ( n44140 , n44121 , n44138 , n44139 );
and ( n44141 , n44097 , n44140 );
xor ( n44142 , n43937 , n43938 );
xor ( n44143 , n44142 , n43940 );
xor ( n44144 , n43951 , n43952 );
xor ( n44145 , n44144 , n43954 );
and ( n44146 , n44143 , n44145 );
xor ( n44147 , n43960 , n43961 );
xor ( n44148 , n44147 , n43966 );
and ( n44149 , n44145 , n44148 );
and ( n44150 , n44143 , n44148 );
or ( n44151 , n44146 , n44149 , n44150 );
and ( n44152 , n44140 , n44151 );
and ( n44153 , n44097 , n44151 );
or ( n44154 , n44141 , n44152 , n44153 );
xor ( n44155 , n43922 , n43926 );
xor ( n44156 , n44155 , n43929 );
xor ( n44157 , n43934 , n43935 );
xor ( n44158 , n44157 , n43943 );
and ( n44159 , n44156 , n44158 );
xor ( n44160 , n43957 , n43969 );
xor ( n44161 , n44160 , n43986 );
and ( n44162 , n44158 , n44161 );
and ( n44163 , n44156 , n44161 );
or ( n44164 , n44159 , n44162 , n44163 );
and ( n44165 , n44154 , n44164 );
xor ( n44166 , n43918 , n43932 );
xor ( n44167 , n44166 , n43946 );
and ( n44168 , n44164 , n44167 );
and ( n44169 , n44154 , n44167 );
or ( n44170 , n44165 , n44168 , n44169 );
xor ( n44171 , n43907 , n43909 );
xor ( n44172 , n44171 , n43912 );
and ( n44173 , n44170 , n44172 );
xor ( n44174 , n43916 , n43949 );
xor ( n44175 , n44174 , n44019 );
and ( n44176 , n44172 , n44175 );
and ( n44177 , n44170 , n44175 );
or ( n44178 , n44173 , n44176 , n44177 );
xor ( n44179 , n43897 , n43899 );
xor ( n44180 , n44179 , n43902 );
and ( n44181 , n44178 , n44180 );
xor ( n44182 , n43915 , n44022 );
xor ( n44183 , n44182 , n44025 );
and ( n44184 , n44180 , n44183 );
and ( n44185 , n44178 , n44183 );
or ( n44186 , n44181 , n44184 , n44185 );
and ( n44187 , n44073 , n44186 );
xor ( n44188 , n43779 , n43781 );
xor ( n44189 , n44188 , n43828 );
and ( n44190 , n44186 , n44189 );
and ( n44191 , n44073 , n44189 );
or ( n44192 , n44187 , n44190 , n44191 );
and ( n44193 , n44042 , n44192 );
xor ( n44194 , n43777 , n43831 );
xor ( n44195 , n44194 , n44034 );
and ( n44196 , n44192 , n44195 );
and ( n44197 , n44042 , n44195 );
or ( n44198 , n44193 , n44196 , n44197 );
and ( n44199 , n44039 , n44198 );
and ( n44200 , n44037 , n44198 );
or ( n44201 , n44040 , n44199 , n44200 );
and ( n44202 , n43775 , n44201 );
xor ( n44203 , n44037 , n44039 );
xor ( n44204 , n44203 , n44198 );
xor ( n44205 , n43905 , n44028 );
xor ( n44206 , n44205 , n44031 );
xor ( n44207 , n44048 , n44050 );
xor ( n44208 , n44081 , n44085 );
and ( n44209 , n26933 , n43959 );
and ( n44210 , n44208 , n44209 );
and ( n44211 , n43619 , n34352 );
and ( n44212 , n43562 , n34350 );
nor ( n44213 , n44211 , n44212 );
xnor ( n44214 , n44213 , n28532 );
and ( n44215 , n44209 , n44214 );
and ( n44216 , n44208 , n44214 );
or ( n44217 , n44210 , n44215 , n44216 );
and ( n44218 , n27389 , n43009 );
and ( n44219 , n44217 , n44218 );
and ( n44220 , n43248 , n34911 );
and ( n44221 , n43124 , n34909 );
nor ( n44222 , n44220 , n44221 );
xnor ( n44223 , n44222 , n34104 );
and ( n44224 , n44218 , n44223 );
and ( n44225 , n44217 , n44223 );
or ( n44226 , n44219 , n44224 , n44225 );
and ( n44227 , n28129 , n41038 );
and ( n44228 , n44226 , n44227 );
and ( n44229 , n27962 , n41445 );
and ( n44230 , n44227 , n44229 );
and ( n44231 , n44226 , n44229 );
or ( n44232 , n44228 , n44230 , n44231 );
and ( n44233 , n42157 , n35911 );
and ( n44234 , n41890 , n35909 );
nor ( n44235 , n44233 , n44234 );
xnor ( n44236 , n44235 , n35161 );
and ( n44237 , n44232 , n44236 );
and ( n44238 , n44207 , n44237 );
xor ( n44239 , n43989 , n44013 );
xor ( n44240 , n44239 , n44016 );
xor ( n44241 , n44005 , n44007 );
xor ( n44242 , n44241 , n44010 );
xor ( n44243 , n43974 , n43978 );
xor ( n44244 , n44243 , n43983 );
xor ( n44245 , n43993 , n43997 );
xor ( n44246 , n44245 , n44002 );
and ( n44247 , n44244 , n44246 );
and ( n44248 , n28129 , n42323 );
and ( n44249 , n27962 , n42621 );
and ( n44250 , n44248 , n44249 );
and ( n44251 , n27863 , n43009 );
and ( n44252 , n44249 , n44251 );
and ( n44253 , n44248 , n44251 );
or ( n44254 , n44250 , n44252 , n44253 );
and ( n44255 , n27389 , n43738 );
and ( n44256 , n26980 , n43959 );
and ( n44257 , n44255 , n44256 );
buf ( n44258 , n16870 );
buf ( n44259 , n44258 );
and ( n44260 , n26933 , n44259 );
and ( n44261 , n44256 , n44260 );
and ( n44262 , n44255 , n44260 );
or ( n44263 , n44257 , n44261 , n44262 );
and ( n44264 , n44254 , n44263 );
buf ( n44265 , n26782 );
and ( n44266 , n41631 , n37197 );
and ( n44267 , n41652 , n37194 );
nor ( n44268 , n44266 , n44267 );
xnor ( n44269 , n44268 , n36218 );
and ( n44270 , n44265 , n44269 );
and ( n44271 , n42157 , n36910 );
and ( n44272 , n41890 , n36908 );
nor ( n44273 , n44271 , n44272 );
xnor ( n44274 , n44273 , n36221 );
and ( n44275 , n44269 , n44274 );
and ( n44276 , n44265 , n44274 );
or ( n44277 , n44270 , n44275 , n44276 );
and ( n44278 , n44263 , n44277 );
and ( n44279 , n44254 , n44277 );
or ( n44280 , n44264 , n44278 , n44279 );
and ( n44281 , n44246 , n44280 );
and ( n44282 , n44244 , n44280 );
or ( n44283 , n44247 , n44281 , n44282 );
and ( n44284 , n44242 , n44283 );
and ( n44285 , n42570 , n36367 );
and ( n44286 , n42414 , n36365 );
nor ( n44287 , n44285 , n44286 );
xnor ( n44288 , n44287 , n35608 );
and ( n44289 , n42835 , n35911 );
and ( n44290 , n42682 , n35909 );
nor ( n44291 , n44289 , n44290 );
xnor ( n44292 , n44291 , n35161 );
and ( n44293 , n44288 , n44292 );
and ( n44294 , n43562 , n34911 );
and ( n44295 , n43363 , n34909 );
nor ( n44296 , n44294 , n44295 );
xnor ( n44297 , n44296 , n34104 );
and ( n44298 , n44292 , n44297 );
and ( n44299 , n44288 , n44297 );
or ( n44300 , n44293 , n44298 , n44299 );
xor ( n44301 , n44088 , n44089 );
xor ( n44302 , n44301 , n44091 );
and ( n44303 , n44300 , n44302 );
xor ( n44304 , n44098 , n44099 );
xor ( n44305 , n44304 , n44101 );
and ( n44306 , n44302 , n44305 );
and ( n44307 , n44300 , n44305 );
or ( n44308 , n44303 , n44306 , n44307 );
xor ( n44309 , n44078 , n44086 );
xor ( n44310 , n44309 , n44094 );
and ( n44311 , n44308 , n44310 );
xor ( n44312 , n44104 , n44120 );
xor ( n44313 , n44312 , n44137 );
and ( n44314 , n44310 , n44313 );
and ( n44315 , n44308 , n44313 );
or ( n44316 , n44311 , n44314 , n44315 );
and ( n44317 , n44283 , n44316 );
and ( n44318 , n44242 , n44316 );
or ( n44319 , n44284 , n44317 , n44318 );
and ( n44320 , n44240 , n44319 );
xor ( n44321 , n44059 , n44061 );
xor ( n44322 , n44321 , n44064 );
and ( n44323 , n44319 , n44322 );
and ( n44324 , n44240 , n44322 );
or ( n44325 , n44320 , n44323 , n44324 );
and ( n44326 , n44237 , n44325 );
and ( n44327 , n44207 , n44325 );
or ( n44328 , n44238 , n44326 , n44327 );
xor ( n44329 , n44044 , n44051 );
xor ( n44330 , n44329 , n44070 );
and ( n44331 , n44328 , n44330 );
xor ( n44332 , n44178 , n44180 );
xor ( n44333 , n44332 , n44183 );
and ( n44334 , n44330 , n44333 );
and ( n44335 , n44328 , n44333 );
or ( n44336 , n44331 , n44334 , n44335 );
and ( n44337 , n44206 , n44336 );
xor ( n44338 , n44073 , n44186 );
xor ( n44339 , n44338 , n44189 );
and ( n44340 , n44336 , n44339 );
and ( n44341 , n44206 , n44339 );
or ( n44342 , n44337 , n44340 , n44341 );
xor ( n44343 , n44042 , n44192 );
xor ( n44344 , n44343 , n44195 );
and ( n44345 , n44342 , n44344 );
xor ( n44346 , n44206 , n44336 );
xor ( n44347 , n44346 , n44339 );
xor ( n44348 , n44054 , n44056 );
xor ( n44349 , n44348 , n44067 );
xor ( n44350 , n44170 , n44172 );
xor ( n44351 , n44350 , n44175 );
and ( n44352 , n44349 , n44351 );
xor ( n44353 , n44154 , n44164 );
xor ( n44354 , n44353 , n44167 );
xor ( n44355 , n44232 , n44236 );
and ( n44356 , n44354 , n44355 );
xor ( n44357 , n44097 , n44140 );
xor ( n44358 , n44357 , n44151 );
xor ( n44359 , n44156 , n44158 );
xor ( n44360 , n44359 , n44161 );
and ( n44361 , n44358 , n44360 );
xor ( n44362 , n44226 , n44227 );
xor ( n44363 , n44362 , n44229 );
and ( n44364 , n44360 , n44363 );
and ( n44365 , n44358 , n44363 );
or ( n44366 , n44361 , n44364 , n44365 );
and ( n44367 , n44355 , n44366 );
and ( n44368 , n44354 , n44366 );
or ( n44369 , n44356 , n44367 , n44368 );
and ( n44370 , n44351 , n44369 );
and ( n44371 , n44349 , n44369 );
or ( n44372 , n44352 , n44370 , n44371 );
xor ( n44373 , n44328 , n44330 );
xor ( n44374 , n44373 , n44333 );
and ( n44375 , n44372 , n44374 );
xor ( n44376 , n44207 , n44237 );
xor ( n44377 , n44376 , n44325 );
xor ( n44378 , n44143 , n44145 );
xor ( n44379 , n44378 , n44148 );
xor ( n44380 , n44217 , n44218 );
xor ( n44381 , n44380 , n44223 );
and ( n44382 , n44379 , n44381 );
xor ( n44383 , n44108 , n44112 );
xor ( n44384 , n44383 , n44117 );
xor ( n44385 , n44125 , n44129 );
xor ( n44386 , n44385 , n44134 );
and ( n44387 , n44384 , n44386 );
xor ( n44388 , n44208 , n44209 );
xor ( n44389 , n44388 , n44214 );
and ( n44390 , n44386 , n44389 );
and ( n44391 , n44384 , n44389 );
or ( n44392 , n44387 , n44390 , n44391 );
and ( n44393 , n44381 , n44392 );
and ( n44394 , n44379 , n44392 );
or ( n44395 , n44382 , n44393 , n44394 );
and ( n44396 , n43805 , n34352 );
and ( n44397 , n43619 , n34350 );
nor ( n44398 , n44396 , n44397 );
xnor ( n44399 , n44398 , n28532 );
and ( n44400 , n44399 , n44079 );
and ( n44401 , n44077 , n34350 );
not ( n44402 , n44401 );
and ( n44403 , n44402 , n28532 );
and ( n44404 , n44077 , n34352 );
and ( n44405 , n43805 , n34350 );
nor ( n44406 , n44404 , n44405 );
xnor ( n44407 , n44406 , n28532 );
and ( n44408 , n44403 , n44407 );
and ( n44409 , n44079 , n44408 );
and ( n44410 , n44399 , n44408 );
or ( n44411 , n44400 , n44409 , n44410 );
and ( n44412 , n27591 , n43738 );
and ( n44413 , n26980 , n44259 );
and ( n44414 , n44412 , n44413 );
and ( n44415 , n41890 , n37197 );
and ( n44416 , n41631 , n37194 );
nor ( n44417 , n44415 , n44416 );
xnor ( n44418 , n44417 , n36218 );
and ( n44419 , n44413 , n44418 );
and ( n44420 , n44412 , n44418 );
or ( n44421 , n44414 , n44419 , n44420 );
xor ( n44422 , n44248 , n44249 );
xor ( n44423 , n44422 , n44251 );
and ( n44424 , n44421 , n44423 );
xor ( n44425 , n44255 , n44256 );
xor ( n44426 , n44425 , n44260 );
and ( n44427 , n44423 , n44426 );
and ( n44428 , n44421 , n44426 );
or ( n44429 , n44424 , n44427 , n44428 );
and ( n44430 , n44411 , n44429 );
xor ( n44431 , n44254 , n44263 );
xor ( n44432 , n44431 , n44277 );
and ( n44433 , n44429 , n44432 );
and ( n44434 , n44411 , n44432 );
or ( n44435 , n44430 , n44433 , n44434 );
xor ( n44436 , n44244 , n44246 );
xor ( n44437 , n44436 , n44280 );
and ( n44438 , n44435 , n44437 );
xor ( n44439 , n44308 , n44310 );
xor ( n44440 , n44439 , n44313 );
and ( n44441 , n44437 , n44440 );
and ( n44442 , n44435 , n44440 );
or ( n44443 , n44438 , n44441 , n44442 );
and ( n44444 , n44395 , n44443 );
xor ( n44445 , n44242 , n44283 );
xor ( n44446 , n44445 , n44316 );
and ( n44447 , n44443 , n44446 );
and ( n44448 , n44395 , n44446 );
or ( n44449 , n44444 , n44447 , n44448 );
xor ( n44450 , n44240 , n44319 );
xor ( n44451 , n44450 , n44322 );
and ( n44452 , n44449 , n44451 );
xor ( n44453 , n44300 , n44302 );
xor ( n44454 , n44453 , n44305 );
xor ( n44455 , n44403 , n44407 );
and ( n44456 , n27389 , n43959 );
and ( n44457 , n44455 , n44456 );
and ( n44458 , n43619 , n34911 );
and ( n44459 , n43562 , n34909 );
nor ( n44460 , n44458 , n44459 );
xnor ( n44461 , n44460 , n34104 );
and ( n44462 , n44456 , n44461 );
and ( n44463 , n44455 , n44461 );
or ( n44464 , n44457 , n44462 , n44463 );
and ( n44465 , n27591 , n43446 );
and ( n44466 , n44464 , n44465 );
and ( n44467 , n43248 , n35374 );
and ( n44468 , n43124 , n35372 );
nor ( n44469 , n44467 , n44468 );
xnor ( n44470 , n44469 , n34661 );
and ( n44471 , n44465 , n44470 );
and ( n44472 , n44464 , n44470 );
or ( n44473 , n44466 , n44471 , n44472 );
and ( n44474 , n44454 , n44473 );
xor ( n44475 , n44265 , n44269 );
xor ( n44476 , n44475 , n44274 );
xor ( n44477 , n44288 , n44292 );
xor ( n44478 , n44477 , n44297 );
and ( n44479 , n44476 , n44478 );
and ( n44480 , n27591 , n43959 );
buf ( n44481 , n16981 );
buf ( n44482 , n44481 );
and ( n44483 , n26980 , n44482 );
and ( n44484 , n44480 , n44483 );
and ( n44485 , n43805 , n34911 );
and ( n44486 , n43619 , n34909 );
nor ( n44487 , n44485 , n44486 );
xnor ( n44488 , n44487 , n34104 );
and ( n44489 , n44483 , n44488 );
and ( n44490 , n44480 , n44488 );
or ( n44491 , n44484 , n44489 , n44490 );
and ( n44492 , n27863 , n43446 );
and ( n44493 , n44491 , n44492 );
and ( n44494 , n43363 , n35374 );
and ( n44495 , n43248 , n35372 );
nor ( n44496 , n44494 , n44495 );
xnor ( n44497 , n44496 , n34661 );
and ( n44498 , n44492 , n44497 );
and ( n44499 , n44491 , n44497 );
or ( n44500 , n44493 , n44498 , n44499 );
and ( n44501 , n44478 , n44500 );
and ( n44502 , n44476 , n44500 );
or ( n44503 , n44479 , n44501 , n44502 );
and ( n44504 , n44473 , n44503 );
and ( n44505 , n44454 , n44503 );
or ( n44506 , n44474 , n44504 , n44505 );
and ( n44507 , n42414 , n36910 );
and ( n44508 , n42157 , n36908 );
nor ( n44509 , n44507 , n44508 );
xnor ( n44510 , n44509 , n36221 );
and ( n44511 , n42682 , n36367 );
and ( n44512 , n42570 , n36365 );
nor ( n44513 , n44511 , n44512 );
xnor ( n44514 , n44513 , n35608 );
and ( n44515 , n44510 , n44514 );
and ( n44516 , n28129 , n43009 );
and ( n44517 , n27863 , n43738 );
and ( n44518 , n44516 , n44517 );
and ( n44519 , n27389 , n44259 );
and ( n44520 , n44517 , n44519 );
and ( n44521 , n44516 , n44519 );
or ( n44522 , n44518 , n44520 , n44521 );
and ( n44523 , n44514 , n44522 );
and ( n44524 , n44510 , n44522 );
or ( n44525 , n44515 , n44523 , n44524 );
xor ( n44526 , n44399 , n44079 );
xor ( n44527 , n44526 , n44408 );
and ( n44528 , n44525 , n44527 );
xor ( n44529 , n44421 , n44423 );
xor ( n44530 , n44529 , n44426 );
and ( n44531 , n44527 , n44530 );
and ( n44532 , n44525 , n44530 );
or ( n44533 , n44528 , n44531 , n44532 );
xor ( n44534 , n44384 , n44386 );
xor ( n44535 , n44534 , n44389 );
and ( n44536 , n44533 , n44535 );
xor ( n44537 , n44411 , n44429 );
xor ( n44538 , n44537 , n44432 );
and ( n44539 , n44535 , n44538 );
and ( n44540 , n44533 , n44538 );
or ( n44541 , n44536 , n44539 , n44540 );
and ( n44542 , n44506 , n44541 );
xor ( n44543 , n44379 , n44381 );
xor ( n44544 , n44543 , n44392 );
and ( n44545 , n44541 , n44544 );
and ( n44546 , n44506 , n44544 );
or ( n44547 , n44542 , n44545 , n44546 );
xor ( n44548 , n44358 , n44360 );
xor ( n44549 , n44548 , n44363 );
and ( n44550 , n44547 , n44549 );
xor ( n44551 , n44395 , n44443 );
xor ( n44552 , n44551 , n44446 );
and ( n44553 , n44549 , n44552 );
and ( n44554 , n44547 , n44552 );
or ( n44555 , n44550 , n44553 , n44554 );
and ( n44556 , n44451 , n44555 );
and ( n44557 , n44449 , n44555 );
or ( n44558 , n44452 , n44556 , n44557 );
and ( n44559 , n44377 , n44558 );
xor ( n44560 , n44349 , n44351 );
xor ( n44561 , n44560 , n44369 );
and ( n44562 , n44558 , n44561 );
and ( n44563 , n44377 , n44561 );
or ( n44564 , n44559 , n44562 , n44563 );
and ( n44565 , n44374 , n44564 );
and ( n44566 , n44372 , n44564 );
or ( n44567 , n44375 , n44565 , n44566 );
and ( n44568 , n44347 , n44567 );
xor ( n44569 , n44372 , n44374 );
xor ( n44570 , n44569 , n44564 );
xor ( n44571 , n44377 , n44558 );
xor ( n44572 , n44571 , n44561 );
xor ( n44573 , n44354 , n44355 );
xor ( n44574 , n44573 , n44366 );
xor ( n44575 , n44449 , n44451 );
xor ( n44576 , n44575 , n44555 );
and ( n44577 , n44574 , n44576 );
xor ( n44578 , n44435 , n44437 );
xor ( n44579 , n44578 , n44440 );
xor ( n44580 , n44464 , n44465 );
xor ( n44581 , n44580 , n44470 );
and ( n44582 , n28129 , n42621 );
xor ( n44583 , n44491 , n44492 );
xor ( n44584 , n44583 , n44497 );
and ( n44585 , n44582 , n44584 );
and ( n44586 , n44581 , n44585 );
buf ( n44587 , n26933 );
and ( n44588 , n42157 , n37197 );
and ( n44589 , n41890 , n37194 );
nor ( n44590 , n44588 , n44589 );
xnor ( n44591 , n44590 , n36218 );
and ( n44592 , n44587 , n44591 );
and ( n44593 , n42570 , n36910 );
and ( n44594 , n42414 , n36908 );
nor ( n44595 , n44593 , n44594 );
xnor ( n44596 , n44595 , n36221 );
and ( n44597 , n44591 , n44596 );
and ( n44598 , n44587 , n44596 );
or ( n44599 , n44592 , n44597 , n44598 );
xor ( n44600 , n44412 , n44413 );
xor ( n44601 , n44600 , n44418 );
and ( n44602 , n44599 , n44601 );
xor ( n44603 , n44455 , n44456 );
xor ( n44604 , n44603 , n44461 );
and ( n44605 , n44601 , n44604 );
and ( n44606 , n44599 , n44604 );
or ( n44607 , n44602 , n44605 , n44606 );
and ( n44608 , n44585 , n44607 );
and ( n44609 , n44581 , n44607 );
or ( n44610 , n44586 , n44608 , n44609 );
and ( n44611 , n43248 , n35911 );
and ( n44612 , n43124 , n35909 );
nor ( n44613 , n44611 , n44612 );
xnor ( n44614 , n44613 , n35161 );
xor ( n44615 , n44480 , n44483 );
xor ( n44616 , n44615 , n44488 );
and ( n44617 , n44614 , n44616 );
and ( n44618 , n44077 , n34909 );
not ( n44619 , n44618 );
and ( n44620 , n44619 , n34104 );
and ( n44621 , n44077 , n34911 );
and ( n44622 , n43805 , n34909 );
nor ( n44623 , n44621 , n44622 );
xnor ( n44624 , n44623 , n34104 );
and ( n44625 , n44620 , n44624 );
and ( n44626 , n44401 , n44625 );
and ( n44627 , n27863 , n43959 );
and ( n44628 , n27591 , n44259 );
and ( n44629 , n44627 , n44628 );
and ( n44630 , n42414 , n37197 );
and ( n44631 , n42157 , n37194 );
nor ( n44632 , n44630 , n44631 );
xnor ( n44633 , n44632 , n36218 );
and ( n44634 , n44628 , n44633 );
and ( n44635 , n44627 , n44633 );
or ( n44636 , n44629 , n44634 , n44635 );
and ( n44637 , n44625 , n44636 );
and ( n44638 , n44401 , n44636 );
or ( n44639 , n44626 , n44637 , n44638 );
and ( n44640 , n44617 , n44639 );
xor ( n44641 , n44510 , n44514 );
xor ( n44642 , n44641 , n44522 );
and ( n44643 , n44639 , n44642 );
and ( n44644 , n44617 , n44642 );
or ( n44645 , n44640 , n44643 , n44644 );
xor ( n44646 , n44476 , n44478 );
xor ( n44647 , n44646 , n44500 );
and ( n44648 , n44645 , n44647 );
xor ( n44649 , n44525 , n44527 );
xor ( n44650 , n44649 , n44530 );
and ( n44651 , n44647 , n44650 );
and ( n44652 , n44645 , n44650 );
or ( n44653 , n44648 , n44651 , n44652 );
and ( n44654 , n44610 , n44653 );
xor ( n44655 , n44454 , n44473 );
xor ( n44656 , n44655 , n44503 );
and ( n44657 , n44653 , n44656 );
and ( n44658 , n44610 , n44656 );
or ( n44659 , n44654 , n44657 , n44658 );
and ( n44660 , n44579 , n44659 );
xor ( n44661 , n44506 , n44541 );
xor ( n44662 , n44661 , n44544 );
and ( n44663 , n44659 , n44662 );
and ( n44664 , n44579 , n44662 );
or ( n44665 , n44660 , n44663 , n44664 );
xor ( n44666 , n44547 , n44549 );
xor ( n44667 , n44666 , n44552 );
and ( n44668 , n44665 , n44667 );
xor ( n44669 , n44533 , n44535 );
xor ( n44670 , n44669 , n44538 );
xor ( n44671 , n44620 , n44624 );
and ( n44672 , n27389 , n44482 );
and ( n44673 , n44671 , n44672 );
and ( n44674 , n43619 , n35374 );
and ( n44675 , n43562 , n35372 );
nor ( n44676 , n44674 , n44675 );
xnor ( n44677 , n44676 , n34661 );
and ( n44678 , n44672 , n44677 );
and ( n44679 , n44671 , n44677 );
or ( n44680 , n44673 , n44678 , n44679 );
and ( n44681 , n27962 , n43446 );
and ( n44682 , n44680 , n44681 );
and ( n44683 , n43562 , n35374 );
and ( n44684 , n43363 , n35372 );
nor ( n44685 , n44683 , n44684 );
xnor ( n44686 , n44685 , n34661 );
and ( n44687 , n44681 , n44686 );
and ( n44688 , n44680 , n44686 );
or ( n44689 , n44682 , n44687 , n44688 );
and ( n44690 , n27962 , n43009 );
and ( n44691 , n44689 , n44690 );
and ( n44692 , n43124 , n35911 );
and ( n44693 , n42835 , n35909 );
nor ( n44694 , n44692 , n44693 );
xnor ( n44695 , n44694 , n35161 );
and ( n44696 , n44690 , n44695 );
and ( n44697 , n44689 , n44695 );
or ( n44698 , n44691 , n44696 , n44697 );
xor ( n44699 , n44582 , n44584 );
xor ( n44700 , n44516 , n44517 );
xor ( n44701 , n44700 , n44519 );
xor ( n44702 , n44587 , n44591 );
xor ( n44703 , n44702 , n44596 );
and ( n44704 , n44701 , n44703 );
xor ( n44705 , n44614 , n44616 );
and ( n44706 , n44703 , n44705 );
and ( n44707 , n44701 , n44705 );
or ( n44708 , n44704 , n44706 , n44707 );
and ( n44709 , n44699 , n44708 );
xor ( n44710 , n44599 , n44601 );
xor ( n44711 , n44710 , n44604 );
and ( n44712 , n44708 , n44711 );
and ( n44713 , n44699 , n44711 );
or ( n44714 , n44709 , n44712 , n44713 );
and ( n44715 , n44698 , n44714 );
xor ( n44716 , n44581 , n44585 );
xor ( n44717 , n44716 , n44607 );
and ( n44718 , n44714 , n44717 );
and ( n44719 , n44698 , n44717 );
or ( n44720 , n44715 , n44718 , n44719 );
and ( n44721 , n44670 , n44720 );
xor ( n44722 , n44610 , n44653 );
xor ( n44723 , n44722 , n44656 );
and ( n44724 , n44720 , n44723 );
and ( n44725 , n44670 , n44723 );
or ( n44726 , n44721 , n44724 , n44725 );
xor ( n44727 , n44579 , n44659 );
xor ( n44728 , n44727 , n44662 );
and ( n44729 , n44726 , n44728 );
xor ( n44730 , n44645 , n44647 );
xor ( n44731 , n44730 , n44650 );
xor ( n44732 , n44617 , n44639 );
xor ( n44733 , n44732 , n44642 );
xor ( n44734 , n44689 , n44690 );
xor ( n44735 , n44734 , n44695 );
and ( n44736 , n44733 , n44735 );
and ( n44737 , n42682 , n36910 );
and ( n44738 , n42570 , n36908 );
nor ( n44739 , n44737 , n44738 );
xnor ( n44740 , n44739 , n36221 );
and ( n44741 , n43124 , n36367 );
and ( n44742 , n42835 , n36365 );
nor ( n44743 , n44741 , n44742 );
xnor ( n44744 , n44743 , n35608 );
and ( n44745 , n44740 , n44744 );
buf ( n44746 , n26980 );
and ( n44747 , n44746 , n44618 );
and ( n44748 , n44744 , n44747 );
and ( n44749 , n44740 , n44747 );
or ( n44750 , n44745 , n44748 , n44749 );
xor ( n44751 , n44401 , n44625 );
xor ( n44752 , n44751 , n44636 );
and ( n44753 , n44750 , n44752 );
and ( n44754 , n44077 , n35372 );
not ( n44755 , n44754 );
and ( n44756 , n44755 , n34661 );
and ( n44757 , n44077 , n35374 );
and ( n44758 , n43805 , n35372 );
nor ( n44759 , n44757 , n44758 );
xnor ( n44760 , n44759 , n34661 );
and ( n44761 , n44756 , n44760 );
and ( n44762 , n27591 , n44482 );
and ( n44763 , n44761 , n44762 );
and ( n44764 , n43805 , n35374 );
and ( n44765 , n43619 , n35372 );
nor ( n44766 , n44764 , n44765 );
xnor ( n44767 , n44766 , n34661 );
and ( n44768 , n44762 , n44767 );
and ( n44769 , n44761 , n44767 );
or ( n44770 , n44763 , n44768 , n44769 );
and ( n44771 , n27962 , n43738 );
and ( n44772 , n44770 , n44771 );
and ( n44773 , n43363 , n35911 );
and ( n44774 , n43248 , n35909 );
nor ( n44775 , n44773 , n44774 );
xnor ( n44776 , n44775 , n35161 );
and ( n44777 , n44771 , n44776 );
and ( n44778 , n44770 , n44776 );
or ( n44779 , n44772 , n44777 , n44778 );
and ( n44780 , n44752 , n44779 );
and ( n44781 , n44750 , n44779 );
or ( n44782 , n44753 , n44780 , n44781 );
and ( n44783 , n44735 , n44782 );
and ( n44784 , n44733 , n44782 );
or ( n44785 , n44736 , n44783 , n44784 );
and ( n44786 , n44731 , n44785 );
xor ( n44787 , n44698 , n44714 );
xor ( n44788 , n44787 , n44717 );
and ( n44789 , n44785 , n44788 );
and ( n44790 , n44731 , n44788 );
or ( n44791 , n44786 , n44789 , n44790 );
xor ( n44792 , n44670 , n44720 );
xor ( n44793 , n44792 , n44723 );
and ( n44794 , n44791 , n44793 );
xor ( n44795 , n44699 , n44708 );
xor ( n44796 , n44795 , n44711 );
and ( n44797 , n27962 , n43959 );
and ( n44798 , n27863 , n44259 );
and ( n44799 , n44797 , n44798 );
buf ( n44800 , n17035 );
buf ( n44801 , n44800 );
and ( n44802 , n27389 , n44801 );
not ( n44803 , n44802 );
xor ( n44804 , n44746 , n44618 );
xor ( n44805 , n44803 , n44804 );
not ( n44806 , n44805 );
and ( n44807 , n44798 , n44806 );
and ( n44808 , n44797 , n44806 );
or ( n44809 , n44799 , n44807 , n44808 );
and ( n44810 , n28129 , n43446 );
and ( n44811 , n44809 , n44810 );
xor ( n44812 , n44671 , n44672 );
xor ( n44813 , n44812 , n44677 );
and ( n44814 , n44810 , n44813 );
and ( n44815 , n44809 , n44813 );
or ( n44816 , n44811 , n44814 , n44815 );
and ( n44817 , n42835 , n36367 );
and ( n44818 , n42682 , n36365 );
nor ( n44819 , n44817 , n44818 );
xnor ( n44820 , n44819 , n35608 );
and ( n44821 , n44816 , n44820 );
xor ( n44822 , n44680 , n44681 );
xor ( n44823 , n44822 , n44686 );
and ( n44824 , n44820 , n44823 );
and ( n44825 , n44816 , n44823 );
or ( n44826 , n44821 , n44824 , n44825 );
and ( n44827 , n44796 , n44826 );
xor ( n44828 , n44627 , n44628 );
xor ( n44829 , n44828 , n44633 );
and ( n44830 , n44803 , n44804 );
and ( n44831 , n44829 , n44830 );
buf ( n44832 , n44802 );
and ( n44833 , n44830 , n44832 );
and ( n44834 , n44829 , n44832 );
or ( n44835 , n44831 , n44833 , n44834 );
xor ( n44836 , n44701 , n44703 );
xor ( n44837 , n44836 , n44705 );
and ( n44838 , n44835 , n44837 );
and ( n44839 , n42570 , n37197 );
and ( n44840 , n42414 , n37194 );
nor ( n44841 , n44839 , n44840 );
xnor ( n44842 , n44841 , n36218 );
and ( n44843 , n42835 , n36910 );
and ( n44844 , n42682 , n36908 );
nor ( n44845 , n44843 , n44844 );
xnor ( n44846 , n44845 , n36221 );
and ( n44847 , n44842 , n44846 );
and ( n44848 , n28129 , n43959 );
and ( n44849 , n42682 , n37197 );
and ( n44850 , n42570 , n37194 );
nor ( n44851 , n44849 , n44850 );
xnor ( n44852 , n44851 , n36218 );
and ( n44853 , n44848 , n44852 );
and ( n44854 , n43124 , n36910 );
and ( n44855 , n42835 , n36908 );
nor ( n44856 , n44854 , n44855 );
xnor ( n44857 , n44856 , n36221 );
and ( n44858 , n44852 , n44857 );
and ( n44859 , n44848 , n44857 );
or ( n44860 , n44853 , n44858 , n44859 );
and ( n44861 , n44846 , n44860 );
and ( n44862 , n44842 , n44860 );
or ( n44863 , n44847 , n44861 , n44862 );
xor ( n44864 , n44740 , n44744 );
xor ( n44865 , n44864 , n44747 );
and ( n44866 , n44863 , n44865 );
xor ( n44867 , n44770 , n44771 );
xor ( n44868 , n44867 , n44776 );
and ( n44869 , n44865 , n44868 );
and ( n44870 , n44863 , n44868 );
or ( n44871 , n44866 , n44869 , n44870 );
and ( n44872 , n44837 , n44871 );
and ( n44873 , n44835 , n44871 );
or ( n44874 , n44838 , n44872 , n44873 );
and ( n44875 , n44826 , n44874 );
and ( n44876 , n44796 , n44874 );
or ( n44877 , n44827 , n44875 , n44876 );
xor ( n44878 , n44731 , n44785 );
xor ( n44879 , n44878 , n44788 );
and ( n44880 , n44877 , n44879 );
xor ( n44881 , n44733 , n44735 );
xor ( n44882 , n44881 , n44782 );
xor ( n44883 , n44756 , n44760 );
and ( n44884 , n27863 , n44482 );
and ( n44885 , n44883 , n44884 );
and ( n44886 , n27591 , n44801 );
and ( n44887 , n44884 , n44886 );
and ( n44888 , n44883 , n44886 );
or ( n44889 , n44885 , n44887 , n44888 );
and ( n44890 , n28129 , n43738 );
and ( n44891 , n44889 , n44890 );
and ( n44892 , n43562 , n35911 );
and ( n44893 , n43363 , n35909 );
nor ( n44894 , n44892 , n44893 );
xnor ( n44895 , n44894 , n35161 );
and ( n44896 , n44890 , n44895 );
and ( n44897 , n44889 , n44895 );
or ( n44898 , n44891 , n44896 , n44897 );
buf ( n44899 , n44805 );
and ( n44900 , n44898 , n44899 );
xor ( n44901 , n44829 , n44830 );
xor ( n44902 , n44901 , n44832 );
and ( n44903 , n44899 , n44902 );
and ( n44904 , n44898 , n44902 );
or ( n44905 , n44900 , n44903 , n44904 );
xor ( n44906 , n44750 , n44752 );
xor ( n44907 , n44906 , n44779 );
and ( n44908 , n44905 , n44907 );
xor ( n44909 , n44816 , n44820 );
xor ( n44910 , n44909 , n44823 );
and ( n44911 , n44907 , n44910 );
and ( n44912 , n44905 , n44910 );
or ( n44913 , n44908 , n44911 , n44912 );
and ( n44914 , n44882 , n44913 );
xor ( n44915 , n44809 , n44810 );
xor ( n44916 , n44915 , n44813 );
and ( n44917 , n44077 , n35909 );
not ( n44918 , n44917 );
and ( n44919 , n44918 , n35161 );
and ( n44920 , n44077 , n35911 );
and ( n44921 , n43805 , n35909 );
nor ( n44922 , n44920 , n44921 );
xnor ( n44923 , n44922 , n35161 );
and ( n44924 , n44919 , n44923 );
and ( n44925 , n27962 , n44482 );
and ( n44926 , n44924 , n44925 );
and ( n44927 , n27863 , n44801 );
and ( n44928 , n44925 , n44927 );
and ( n44929 , n44924 , n44927 );
or ( n44930 , n44926 , n44928 , n44929 );
and ( n44931 , n27962 , n44259 );
and ( n44932 , n44930 , n44931 );
xor ( n44933 , n44883 , n44884 );
xor ( n44934 , n44933 , n44886 );
and ( n44935 , n44931 , n44934 );
and ( n44936 , n44930 , n44934 );
or ( n44937 , n44932 , n44935 , n44936 );
xor ( n44938 , n44761 , n44762 );
xor ( n44939 , n44938 , n44767 );
and ( n44940 , n44937 , n44939 );
and ( n44941 , n44916 , n44940 );
and ( n44942 , n43248 , n36367 );
and ( n44943 , n43124 , n36365 );
nor ( n44944 , n44942 , n44943 );
xnor ( n44945 , n44944 , n35608 );
xor ( n44946 , n44889 , n44890 );
xor ( n44947 , n44946 , n44895 );
and ( n44948 , n44945 , n44947 );
xor ( n44949 , n44797 , n44798 );
xor ( n44950 , n44949 , n44806 );
and ( n44951 , n44947 , n44950 );
and ( n44952 , n44945 , n44950 );
or ( n44953 , n44948 , n44951 , n44952 );
and ( n44954 , n44940 , n44953 );
and ( n44955 , n44916 , n44953 );
or ( n44956 , n44941 , n44954 , n44955 );
and ( n44957 , n43363 , n36367 );
and ( n44958 , n43248 , n36365 );
nor ( n44959 , n44957 , n44958 );
xnor ( n44960 , n44959 , n35608 );
and ( n44961 , n43619 , n35911 );
and ( n44962 , n43562 , n35909 );
nor ( n44963 , n44961 , n44962 );
xnor ( n44964 , n44963 , n35161 );
and ( n44965 , n44960 , n44964 );
buf ( n44966 , n27389 );
or ( n44967 , n44966 , n44754 );
and ( n44968 , n44964 , n44967 );
and ( n44969 , n44960 , n44967 );
or ( n44970 , n44965 , n44968 , n44969 );
xor ( n44971 , n44842 , n44846 );
xor ( n44972 , n44971 , n44860 );
and ( n44973 , n44970 , n44972 );
and ( n44974 , n28129 , n44259 );
buf ( n44975 , n17176 );
buf ( n44976 , n44975 );
and ( n44977 , n27591 , n44976 );
and ( n44978 , n44974 , n44977 );
and ( n44979 , n43248 , n36910 );
and ( n44980 , n43124 , n36908 );
nor ( n44981 , n44979 , n44980 );
xnor ( n44982 , n44981 , n36221 );
and ( n44983 , n44977 , n44982 );
and ( n44984 , n44974 , n44982 );
or ( n44985 , n44978 , n44983 , n44984 );
xor ( n44986 , n44848 , n44852 );
xor ( n44987 , n44986 , n44857 );
and ( n44988 , n44985 , n44987 );
and ( n44989 , n43562 , n36367 );
and ( n44990 , n43363 , n36365 );
nor ( n44991 , n44989 , n44990 );
xnor ( n44992 , n44991 , n35608 );
and ( n44993 , n43805 , n35911 );
and ( n44994 , n43619 , n35909 );
nor ( n44995 , n44993 , n44994 );
xnor ( n44996 , n44995 , n35161 );
and ( n44997 , n44992 , n44996 );
xnor ( n44998 , n44966 , n44754 );
and ( n44999 , n44996 , n44998 );
and ( n45000 , n44992 , n44998 );
or ( n45001 , n44997 , n44999 , n45000 );
and ( n45002 , n44987 , n45001 );
and ( n45003 , n44985 , n45001 );
or ( n45004 , n44988 , n45002 , n45003 );
and ( n45005 , n44972 , n45004 );
and ( n45006 , n44970 , n45004 );
or ( n45007 , n44973 , n45005 , n45006 );
xor ( n45008 , n44863 , n44865 );
xor ( n45009 , n45008 , n44868 );
and ( n45010 , n45007 , n45009 );
xor ( n45011 , n44898 , n44899 );
xor ( n45012 , n45011 , n44902 );
and ( n45013 , n45009 , n45012 );
and ( n45014 , n45007 , n45012 );
or ( n45015 , n45010 , n45013 , n45014 );
and ( n45016 , n44956 , n45015 );
xor ( n45017 , n44835 , n44837 );
xor ( n45018 , n45017 , n44871 );
and ( n45019 , n45015 , n45018 );
and ( n45020 , n44956 , n45018 );
or ( n45021 , n45016 , n45019 , n45020 );
and ( n45022 , n44913 , n45021 );
and ( n45023 , n44882 , n45021 );
or ( n45024 , n44914 , n45022 , n45023 );
and ( n45025 , n44879 , n45024 );
and ( n45026 , n44877 , n45024 );
or ( n45027 , n44880 , n45025 , n45026 );
and ( n45028 , n44793 , n45027 );
and ( n45029 , n44791 , n45027 );
or ( n45030 , n44794 , n45028 , n45029 );
and ( n45031 , n44728 , n45030 );
and ( n45032 , n44726 , n45030 );
or ( n45033 , n44729 , n45031 , n45032 );
and ( n45034 , n44667 , n45033 );
and ( n45035 , n44665 , n45033 );
or ( n45036 , n44668 , n45034 , n45035 );
and ( n45037 , n44576 , n45036 );
and ( n45038 , n44574 , n45036 );
or ( n45039 , n44577 , n45037 , n45038 );
and ( n45040 , n44572 , n45039 );
xor ( n45041 , n44574 , n44576 );
xor ( n45042 , n45041 , n45036 );
xor ( n45043 , n44665 , n44667 );
xor ( n45044 , n45043 , n45033 );
xor ( n45045 , n44726 , n44728 );
xor ( n45046 , n45045 , n45030 );
xor ( n45047 , n44791 , n44793 );
xor ( n45048 , n45047 , n45027 );
xor ( n45049 , n44796 , n44826 );
xor ( n45050 , n45049 , n44874 );
xor ( n45051 , n44937 , n44939 );
xor ( n45052 , n44945 , n44947 );
xor ( n45053 , n45052 , n44950 );
and ( n45054 , n45051 , n45053 );
xor ( n45055 , n44960 , n44964 );
xor ( n45056 , n45055 , n44967 );
xor ( n45057 , n44930 , n44931 );
xor ( n45058 , n45057 , n44934 );
and ( n45059 , n45056 , n45058 );
xor ( n45060 , n44974 , n44977 );
xor ( n45061 , n45060 , n44982 );
xor ( n45062 , n44924 , n44925 );
xor ( n45063 , n45062 , n44927 );
and ( n45064 , n45061 , n45063 );
xor ( n45065 , n44919 , n44923 );
and ( n45066 , n28129 , n44482 );
and ( n45067 , n45065 , n45066 );
and ( n45068 , n43619 , n36367 );
and ( n45069 , n43562 , n36365 );
nor ( n45070 , n45068 , n45069 );
xnor ( n45071 , n45070 , n35608 );
and ( n45072 , n45066 , n45071 );
and ( n45073 , n45065 , n45071 );
or ( n45074 , n45067 , n45072 , n45073 );
and ( n45075 , n45063 , n45074 );
and ( n45076 , n45061 , n45074 );
or ( n45077 , n45064 , n45075 , n45076 );
and ( n45078 , n45058 , n45077 );
and ( n45079 , n45056 , n45077 );
or ( n45080 , n45059 , n45078 , n45079 );
and ( n45081 , n45053 , n45080 );
and ( n45082 , n45051 , n45080 );
or ( n45083 , n45054 , n45081 , n45082 );
xor ( n45084 , n44916 , n44940 );
xor ( n45085 , n45084 , n44953 );
and ( n45086 , n45083 , n45085 );
xor ( n45087 , n45007 , n45009 );
xor ( n45088 , n45087 , n45012 );
and ( n45089 , n45085 , n45088 );
and ( n45090 , n45083 , n45088 );
or ( n45091 , n45086 , n45089 , n45090 );
xor ( n45092 , n44905 , n44907 );
xor ( n45093 , n45092 , n44910 );
and ( n45094 , n45091 , n45093 );
xor ( n45095 , n44956 , n45015 );
xor ( n45096 , n45095 , n45018 );
and ( n45097 , n45093 , n45096 );
and ( n45098 , n45091 , n45096 );
or ( n45099 , n45094 , n45097 , n45098 );
and ( n45100 , n45050 , n45099 );
xor ( n45101 , n44882 , n44913 );
xor ( n45102 , n45101 , n45021 );
and ( n45103 , n45099 , n45102 );
and ( n45104 , n45050 , n45102 );
or ( n45105 , n45100 , n45103 , n45104 );
xor ( n45106 , n44877 , n44879 );
xor ( n45107 , n45106 , n45024 );
and ( n45108 , n45105 , n45107 );
xor ( n45109 , n45050 , n45099 );
xor ( n45110 , n45109 , n45102 );
xor ( n45111 , n45091 , n45093 );
xor ( n45112 , n45111 , n45096 );
xor ( n45113 , n44970 , n44972 );
xor ( n45114 , n45113 , n45004 );
xor ( n45115 , n44985 , n44987 );
xor ( n45116 , n45115 , n45001 );
and ( n45117 , n43124 , n37197 );
and ( n45118 , n42835 , n37194 );
nor ( n45119 , n45117 , n45118 );
xnor ( n45120 , n45119 , n36218 );
and ( n45121 , n43363 , n36910 );
and ( n45122 , n43248 , n36908 );
nor ( n45123 , n45121 , n45122 );
xnor ( n45124 , n45123 , n36221 );
and ( n45125 , n45120 , n45124 );
xor ( n45126 , n45065 , n45066 );
xor ( n45127 , n45126 , n45071 );
and ( n45128 , n45124 , n45127 );
and ( n45129 , n45120 , n45127 );
or ( n45130 , n45125 , n45128 , n45129 );
and ( n45131 , n42835 , n37197 );
and ( n45132 , n42682 , n37194 );
nor ( n45133 , n45131 , n45132 );
xnor ( n45134 , n45133 , n36218 );
or ( n45135 , n45130 , n45134 );
and ( n45136 , n45116 , n45135 );
and ( n45137 , n27962 , n44801 );
and ( n45138 , n27863 , n44976 );
and ( n45139 , n45137 , n45138 );
buf ( n45140 , n27591 );
and ( n45141 , n45140 , n44917 );
and ( n45142 , n45138 , n45141 );
and ( n45143 , n45137 , n45141 );
or ( n45144 , n45139 , n45142 , n45143 );
xor ( n45145 , n44992 , n44996 );
xor ( n45146 , n45145 , n44998 );
and ( n45147 , n45144 , n45146 );
buf ( n45148 , n17217 );
buf ( n45149 , n45148 );
and ( n45150 , n27863 , n45149 );
and ( n45151 , n43248 , n37197 );
and ( n45152 , n43124 , n37194 );
nor ( n45153 , n45151 , n45152 );
xnor ( n45154 , n45153 , n36218 );
and ( n45155 , n45150 , n45154 );
and ( n45156 , n43562 , n36910 );
and ( n45157 , n43363 , n36908 );
nor ( n45158 , n45156 , n45157 );
xnor ( n45159 , n45158 , n36221 );
and ( n45160 , n45154 , n45159 );
and ( n45161 , n45150 , n45159 );
or ( n45162 , n45155 , n45160 , n45161 );
and ( n45163 , n27962 , n45149 );
and ( n45164 , n44077 , n36365 );
not ( n45165 , n45164 );
and ( n45166 , n45165 , n35608 );
and ( n45167 , n45163 , n45166 );
and ( n45168 , n28129 , n44801 );
and ( n45169 , n45167 , n45168 );
and ( n45170 , n27962 , n44976 );
and ( n45171 , n45168 , n45170 );
and ( n45172 , n45167 , n45170 );
or ( n45173 , n45169 , n45171 , n45172 );
and ( n45174 , n45162 , n45173 );
and ( n45175 , n43805 , n36367 );
and ( n45176 , n43619 , n36365 );
nor ( n45177 , n45175 , n45176 );
xnor ( n45178 , n45177 , n35608 );
xor ( n45179 , n45140 , n44917 );
and ( n45180 , n45178 , n45179 );
and ( n45181 , n28129 , n44976 );
and ( n45182 , n43363 , n37197 );
and ( n45183 , n43248 , n37194 );
nor ( n45184 , n45182 , n45183 );
xnor ( n45185 , n45184 , n36218 );
and ( n45186 , n45181 , n45185 );
and ( n45187 , n43619 , n36910 );
and ( n45188 , n43562 , n36908 );
nor ( n45189 , n45187 , n45188 );
xnor ( n45190 , n45189 , n36221 );
and ( n45191 , n45185 , n45190 );
and ( n45192 , n45181 , n45190 );
or ( n45193 , n45186 , n45191 , n45192 );
and ( n45194 , n45179 , n45193 );
and ( n45195 , n45178 , n45193 );
or ( n45196 , n45180 , n45194 , n45195 );
and ( n45197 , n45173 , n45196 );
and ( n45198 , n45162 , n45196 );
or ( n45199 , n45174 , n45197 , n45198 );
and ( n45200 , n45146 , n45199 );
and ( n45201 , n45144 , n45199 );
or ( n45202 , n45147 , n45200 , n45201 );
and ( n45203 , n45135 , n45202 );
and ( n45204 , n45116 , n45202 );
or ( n45205 , n45136 , n45203 , n45204 );
and ( n45206 , n45114 , n45205 );
xor ( n45207 , n45051 , n45053 );
xor ( n45208 , n45207 , n45080 );
and ( n45209 , n45205 , n45208 );
and ( n45210 , n45114 , n45208 );
or ( n45211 , n45206 , n45209 , n45210 );
xor ( n45212 , n45083 , n45085 );
xor ( n45213 , n45212 , n45088 );
and ( n45214 , n45211 , n45213 );
xor ( n45215 , n45056 , n45058 );
xor ( n45216 , n45215 , n45077 );
xor ( n45217 , n45061 , n45063 );
xor ( n45218 , n45217 , n45074 );
xnor ( n45219 , n45130 , n45134 );
and ( n45220 , n45218 , n45219 );
xor ( n45221 , n45137 , n45138 );
xor ( n45222 , n45221 , n45141 );
xor ( n45223 , n45120 , n45124 );
xor ( n45224 , n45223 , n45127 );
and ( n45225 , n45222 , n45224 );
xor ( n45226 , n45150 , n45154 );
xor ( n45227 , n45226 , n45159 );
xor ( n45228 , n45167 , n45168 );
xor ( n45229 , n45228 , n45170 );
and ( n45230 , n45227 , n45229 );
xor ( n45231 , n45163 , n45166 );
buf ( n45232 , n27863 );
and ( n45233 , n45232 , n45164 );
and ( n45234 , n45231 , n45233 );
and ( n45235 , n44077 , n36367 );
and ( n45236 , n43805 , n36365 );
nor ( n45237 , n45235 , n45236 );
xnor ( n45238 , n45237 , n35608 );
and ( n45239 , n45233 , n45238 );
and ( n45240 , n45231 , n45238 );
or ( n45241 , n45234 , n45239 , n45240 );
and ( n45242 , n45229 , n45241 );
and ( n45243 , n45227 , n45241 );
or ( n45244 , n45230 , n45242 , n45243 );
and ( n45245 , n45224 , n45244 );
and ( n45246 , n45222 , n45244 );
or ( n45247 , n45225 , n45245 , n45246 );
and ( n45248 , n45219 , n45247 );
and ( n45249 , n45218 , n45247 );
or ( n45250 , n45220 , n45248 , n45249 );
and ( n45251 , n45216 , n45250 );
xor ( n45252 , n45116 , n45135 );
xor ( n45253 , n45252 , n45202 );
and ( n45254 , n45250 , n45253 );
and ( n45255 , n45216 , n45253 );
or ( n45256 , n45251 , n45254 , n45255 );
xor ( n45257 , n45114 , n45205 );
xor ( n45258 , n45257 , n45208 );
and ( n45259 , n45256 , n45258 );
xor ( n45260 , n45144 , n45146 );
xor ( n45261 , n45260 , n45199 );
xor ( n45262 , n45162 , n45173 );
xor ( n45263 , n45262 , n45196 );
xor ( n45264 , n45178 , n45179 );
xor ( n45265 , n45264 , n45193 );
and ( n45266 , n28129 , n45149 );
buf ( n45267 , n17247 );
buf ( n45268 , n45267 );
and ( n45269 , n27962 , n45268 );
and ( n45270 , n45266 , n45269 );
and ( n45271 , n43562 , n37197 );
and ( n45272 , n43363 , n37194 );
nor ( n45273 , n45271 , n45272 );
xnor ( n45274 , n45273 , n36218 );
and ( n45275 , n45269 , n45274 );
and ( n45276 , n45266 , n45274 );
or ( n45277 , n45270 , n45275 , n45276 );
xor ( n45278 , n45181 , n45185 );
xor ( n45279 , n45278 , n45190 );
and ( n45280 , n45277 , n45279 );
xor ( n45281 , n45231 , n45233 );
xor ( n45282 , n45281 , n45238 );
and ( n45283 , n45279 , n45282 );
and ( n45284 , n45277 , n45282 );
or ( n45285 , n45280 , n45283 , n45284 );
and ( n45286 , n45265 , n45285 );
xor ( n45287 , n45227 , n45229 );
xor ( n45288 , n45287 , n45241 );
and ( n45289 , n45285 , n45288 );
and ( n45290 , n45265 , n45288 );
or ( n45291 , n45286 , n45289 , n45290 );
and ( n45292 , n45263 , n45291 );
xor ( n45293 , n45222 , n45224 );
xor ( n45294 , n45293 , n45244 );
and ( n45295 , n45291 , n45294 );
and ( n45296 , n45263 , n45294 );
or ( n45297 , n45292 , n45295 , n45296 );
and ( n45298 , n45261 , n45297 );
xor ( n45299 , n45218 , n45219 );
xor ( n45300 , n45299 , n45247 );
and ( n45301 , n45297 , n45300 );
and ( n45302 , n45261 , n45300 );
or ( n45303 , n45298 , n45301 , n45302 );
xor ( n45304 , n45216 , n45250 );
xor ( n45305 , n45304 , n45253 );
or ( n45306 , n45303 , n45305 );
and ( n45307 , n45258 , n45306 );
and ( n45308 , n45256 , n45306 );
or ( n45309 , n45259 , n45307 , n45308 );
and ( n45310 , n45213 , n45309 );
and ( n45311 , n45211 , n45309 );
or ( n45312 , n45214 , n45310 , n45311 );
or ( n45313 , n45112 , n45312 );
or ( n45314 , n45110 , n45313 );
and ( n45315 , n45107 , n45314 );
and ( n45316 , n45105 , n45314 );
or ( n45317 , n45108 , n45315 , n45316 );
or ( n45318 , n45048 , n45317 );
or ( n45319 , n45046 , n45318 );
or ( n45320 , n45044 , n45319 );
or ( n45321 , n45042 , n45320 );
and ( n45322 , n45039 , n45321 );
and ( n45323 , n44572 , n45321 );
or ( n45324 , n45040 , n45322 , n45323 );
or ( n45325 , n44570 , n45324 );
and ( n45326 , n44567 , n45325 );
and ( n45327 , n44347 , n45325 );
or ( n45328 , n44568 , n45326 , n45327 );
and ( n45329 , n44344 , n45328 );
and ( n45330 , n44342 , n45328 );
or ( n45331 , n44345 , n45329 , n45330 );
or ( n45332 , n44204 , n45331 );
and ( n45333 , n44201 , n45332 );
and ( n45334 , n43775 , n45332 );
or ( n45335 , n44202 , n45333 , n45334 );
and ( n45336 , n43772 , n45335 );
and ( n45337 , n43770 , n45335 );
or ( n45338 , n43773 , n45336 , n45337 );
or ( n45339 , n43692 , n45338 );
and ( n45340 , n43689 , n45339 );
and ( n45341 , n43322 , n45339 );
or ( n45342 , n43690 , n45340 , n45341 );
and ( n45343 , n43319 , n45342 );
and ( n45344 , n43317 , n45342 );
or ( n45345 , n43320 , n45343 , n45344 );
and ( n45346 , n43213 , n45345 );
and ( n45347 , n43211 , n45345 );
or ( n45348 , n43214 , n45346 , n45347 );
and ( n45349 , n43083 , n45348 );
and ( n45350 , n43081 , n45348 );
or ( n45351 , n43084 , n45349 , n45350 );
and ( n45352 , n42929 , n45351 );
and ( n45353 , n42927 , n45351 );
or ( n45354 , n42930 , n45352 , n45353 );
and ( n45355 , n42778 , n45354 );
xor ( n45356 , n42778 , n45354 );
xor ( n45357 , n42927 , n42929 );
xor ( n45358 , n45357 , n45351 );
not ( n45359 , n45358 );
xor ( n45360 , n43081 , n43083 );
xor ( n45361 , n45360 , n45348 );
xor ( n45362 , n43211 , n43213 );
xor ( n45363 , n45362 , n45345 );
not ( n45364 , n45363 );
xor ( n45365 , n43317 , n43319 );
xor ( n45366 , n45365 , n45342 );
not ( n45367 , n45366 );
xor ( n45368 , n43322 , n43689 );
xor ( n45369 , n45368 , n45339 );
not ( n45370 , n45369 );
xnor ( n45371 , n43692 , n45338 );
xor ( n45372 , n43770 , n43772 );
xor ( n45373 , n45372 , n45335 );
not ( n45374 , n45373 );
xor ( n45375 , n43775 , n44201 );
xor ( n45376 , n45375 , n45332 );
not ( n45377 , n45376 );
xnor ( n45378 , n44204 , n45331 );
xor ( n45379 , n44342 , n44344 );
xor ( n45380 , n45379 , n45328 );
not ( n45381 , n45380 );
xor ( n45382 , n44347 , n44567 );
xor ( n45383 , n45382 , n45325 );
not ( n45384 , n45383 );
xnor ( n45385 , n44570 , n45324 );
xor ( n45386 , n44572 , n45039 );
xor ( n45387 , n45386 , n45321 );
xnor ( n45388 , n45042 , n45320 );
xnor ( n45389 , n45044 , n45319 );
xnor ( n45390 , n45046 , n45318 );
xnor ( n45391 , n45048 , n45317 );
xor ( n45392 , n45105 , n45107 );
xor ( n45393 , n45392 , n45314 );
not ( n45394 , n45393 );
xnor ( n45395 , n45110 , n45313 );
xnor ( n45396 , n45112 , n45312 );
xor ( n45397 , n45211 , n45213 );
xor ( n45398 , n45397 , n45309 );
xor ( n45399 , n45256 , n45258 );
xor ( n45400 , n45399 , n45306 );
not ( n45401 , n45400 );
xnor ( n45402 , n45303 , n45305 );
xor ( n45403 , n45261 , n45297 );
xor ( n45404 , n45403 , n45300 );
xor ( n45405 , n45263 , n45291 );
xor ( n45406 , n45405 , n45294 );
and ( n45407 , n43805 , n36910 );
and ( n45408 , n43619 , n36908 );
nor ( n45409 , n45407 , n45408 );
xnor ( n45410 , n45409 , n36221 );
xor ( n45411 , n45232 , n45164 );
and ( n45412 , n45410 , n45411 );
and ( n45413 , n28129 , n45268 );
and ( n45414 , n43619 , n37197 );
and ( n45415 , n43562 , n37194 );
nor ( n45416 , n45414 , n45415 );
xnor ( n45417 , n45416 , n36218 );
and ( n45418 , n45413 , n45417 );
and ( n45419 , n44077 , n36910 );
and ( n45420 , n43805 , n36908 );
nor ( n45421 , n45419 , n45420 );
xnor ( n45422 , n45421 , n36221 );
and ( n45423 , n45417 , n45422 );
and ( n45424 , n45413 , n45422 );
or ( n45425 , n45418 , n45423 , n45424 );
and ( n45426 , n45411 , n45425 );
and ( n45427 , n45410 , n45425 );
or ( n45428 , n45412 , n45426 , n45427 );
xor ( n45429 , n45266 , n45269 );
xor ( n45430 , n45429 , n45274 );
and ( n45431 , n44077 , n36908 );
not ( n45432 , n45431 );
and ( n45433 , n45432 , n36221 );
buf ( n45434 , n27962 );
and ( n45435 , n45434 , n45431 );
and ( n45436 , n45433 , n45435 );
xor ( n45437 , n45413 , n45417 );
xor ( n45438 , n45437 , n45422 );
and ( n45439 , n45435 , n45438 );
and ( n45440 , n45433 , n45438 );
or ( n45441 , n45436 , n45439 , n45440 );
and ( n45442 , n45430 , n45441 );
xor ( n45443 , n45410 , n45411 );
xor ( n45444 , n45443 , n45425 );
and ( n45445 , n45441 , n45444 );
and ( n45446 , n45430 , n45444 );
or ( n45447 , n45442 , n45445 , n45446 );
and ( n45448 , n45428 , n45447 );
xor ( n45449 , n45277 , n45279 );
xor ( n45450 , n45449 , n45282 );
and ( n45451 , n45447 , n45450 );
and ( n45452 , n45428 , n45450 );
or ( n45453 , n45448 , n45451 , n45452 );
xor ( n45454 , n45265 , n45285 );
xor ( n45455 , n45454 , n45288 );
and ( n45456 , n45453 , n45455 );
xor ( n45457 , n45453 , n45455 );
xor ( n45458 , n45428 , n45447 );
xor ( n45459 , n45458 , n45450 );
xor ( n45460 , n45430 , n45441 );
xor ( n45461 , n45460 , n45444 );
buf ( n45462 , n17268 );
buf ( n45463 , n45462 );
and ( n45464 , n28129 , n45463 );
and ( n45465 , n43805 , n37197 );
and ( n45466 , n43619 , n37194 );
nor ( n45467 , n45465 , n45466 );
xnor ( n45468 , n45467 , n36218 );
and ( n45469 , n45464 , n45468 );
xor ( n45470 , n45434 , n45431 );
and ( n45471 , n45468 , n45470 );
and ( n45472 , n45464 , n45470 );
or ( n45473 , n45469 , n45471 , n45472 );
xor ( n45474 , n45433 , n45435 );
xor ( n45475 , n45474 , n45438 );
and ( n45476 , n45473 , n45475 );
xor ( n45477 , n45473 , n45475 );
xor ( n45478 , n45464 , n45468 );
xor ( n45479 , n45478 , n45470 );
and ( n45480 , n44077 , n37197 );
and ( n45481 , n43805 , n37194 );
nor ( n45482 , n45480 , n45481 );
xnor ( n45483 , n45482 , n36218 );
and ( n45484 , n44077 , n37194 );
not ( n45485 , n45484 );
and ( n45486 , n45485 , n36218 );
and ( n45487 , n45483 , n45486 );
xor ( n45488 , n45483 , n45486 );
buf ( n45489 , n28129 );
and ( n45490 , n45489 , n45484 );
and ( n45491 , n45488 , n45490 );
or ( n45492 , n45487 , n45491 );
and ( n45493 , n45479 , n45492 );
and ( n45494 , n45477 , n45493 );
or ( n45495 , n45476 , n45494 );
and ( n45496 , n45461 , n45495 );
and ( n45497 , n45459 , n45496 );
and ( n45498 , n45457 , n45497 );
or ( n45499 , n45456 , n45498 );
and ( n45500 , n45406 , n45499 );
and ( n45501 , n45404 , n45500 );
and ( n45502 , n45402 , n45501 );
and ( n45503 , n45401 , n45502 );
or ( n45504 , n45400 , n45503 );
and ( n45505 , n45398 , n45504 );
and ( n45506 , n45396 , n45505 );
and ( n45507 , n45395 , n45506 );
and ( n45508 , n45394 , n45507 );
or ( n45509 , n45393 , n45508 );
and ( n45510 , n45391 , n45509 );
and ( n45511 , n45390 , n45510 );
and ( n45512 , n45389 , n45511 );
and ( n45513 , n45388 , n45512 );
and ( n45514 , n45387 , n45513 );
and ( n45515 , n45385 , n45514 );
and ( n45516 , n45384 , n45515 );
or ( n45517 , n45383 , n45516 );
and ( n45518 , n45381 , n45517 );
or ( n45519 , n45380 , n45518 );
and ( n45520 , n45378 , n45519 );
and ( n45521 , n45377 , n45520 );
or ( n45522 , n45376 , n45521 );
and ( n45523 , n45374 , n45522 );
or ( n45524 , n45373 , n45523 );
and ( n45525 , n45371 , n45524 );
and ( n45526 , n45370 , n45525 );
or ( n45527 , n45369 , n45526 );
and ( n45528 , n45367 , n45527 );
or ( n45529 , n45366 , n45528 );
and ( n45530 , n45364 , n45529 );
or ( n45531 , n45363 , n45530 );
and ( n45532 , n45361 , n45531 );
and ( n45533 , n45359 , n45532 );
or ( n45534 , n45358 , n45533 );
and ( n45535 , n45356 , n45534 );
or ( n45536 , n45355 , n45535 );
and ( n45537 , n42776 , n45536 );
or ( n45538 , n42775 , n45537 );
and ( n45539 , n42773 , n45538 );
or ( n45540 , n42772 , n45539 );
and ( n45541 , n42770 , n45540 );
or ( n45542 , n42769 , n45541 );
and ( n45543 , n42767 , n45542 );
and ( n45544 , n42765 , n45543 );
and ( n45545 , n42764 , n45544 );
and ( n45546 , n42763 , n45545 );
and ( n45547 , n42762 , n45546 );
or ( n45548 , n42761 , n45547 );
and ( n45549 , n41796 , n45548 );
or ( n45550 , n41795 , n45549 );
and ( n45551 , n41793 , n45550 );
or ( n45552 , n41792 , n45551 );
and ( n45553 , n41790 , n45552 );
or ( n45554 , n41789 , n45553 );
and ( n45555 , n41787 , n45554 );
or ( n45556 , n41786 , n45555 );
and ( n45557 , n40503 , n45556 );
or ( n45558 , n40502 , n45557 );
and ( n45559 , n40500 , n45558 );
and ( n45560 , n40498 , n45559 );
and ( n45561 , n40497 , n45560 );
or ( n45562 , n40496 , n45561 );
and ( n45563 , n40494 , n45562 );
or ( n45564 , n40493 , n45563 );
and ( n45565 , n39418 , n45564 );
or ( n45566 , n39417 , n45565 );
and ( n45567 , n39415 , n45566 );
or ( n45568 , n39414 , n45567 );
and ( n45569 , n39412 , n45568 );
and ( n45570 , n39410 , n45569 );
and ( n45571 , n39408 , n45570 );
and ( n45572 , n39406 , n45571 );
and ( n45573 , n39404 , n45572 );
or ( n45574 , n39403 , n45573 );
and ( n45575 , n39401 , n45574 );
and ( n45576 , n39400 , n45575 );
or ( n45577 , n39399 , n45576 );
and ( n45578 , n39397 , n45577 );
or ( n45579 , n39396 , n45578 );
and ( n45580 , n39394 , n45579 );
or ( n45581 , n39393 , n45580 );
and ( n45582 , n39391 , n45581 );
and ( n45583 , n39390 , n45582 );
or ( n45584 , n39389 , n45583 );
and ( n45585 , n39387 , n45584 );
and ( n45586 , n39385 , n45585 );
or ( n45587 , n39384 , n45586 );
and ( n45588 , n35500 , n45587 );
or ( n45589 , n35499 , n45588 );
and ( n45590 , n35248 , n45589 );
and ( n45591 , n35246 , n45590 );
and ( n45592 , n35244 , n45591 );
and ( n45593 , n35242 , n45592 );
or ( n45594 , n35241 , n45593 );
and ( n45595 , n34206 , n45594 );
or ( n45596 , n34205 , n45595 );
and ( n45597 , n34203 , n45596 );
and ( n45598 , n34202 , n45597 );
and ( n45599 , n34201 , n45598 );
or ( n45600 , n34200 , n45599 );
and ( n45601 , n28436 , n45600 );
or ( n45602 , n28435 , n45601 );
and ( n45603 , n28433 , n45602 );
and ( n45604 , n28432 , n45603 );
and ( n45605 , n28430 , n45604 );
or ( n45606 , n28429 , n45605 );
and ( n45607 , n27474 , n45606 );
or ( n45608 , n27473 , n45607 );
and ( n45609 , n26756 , n45608 );
or ( n45610 , n26755 , n45609 );
and ( n45611 , n26635 , n45610 );
or ( n45612 , n26634 , n45611 );
and ( n45613 , n26632 , n45612 );
and ( n45614 , n26630 , n45613 );
or ( n45615 , n26629 , n45614 );
and ( n45616 , n26627 , n45615 );
or ( n45617 , n26626 , n45616 );
and ( n45618 , n26010 , n45617 );
or ( n45619 , n26009 , n45618 );
and ( n45620 , n26007 , n45619 );
or ( n45621 , n26006 , n45620 );
and ( n45622 , n25436 , n45621 );
or ( n45623 , n25435 , n45622 );
and ( n45624 , n25181 , n45623 );
and ( n45625 , n25180 , n45624 );
and ( n45626 , n25179 , n45625 );
or ( n45627 , n25178 , n45626 );
and ( n45628 , n25176 , n45627 );
or ( n45629 , n25175 , n45628 );
and ( n45630 , n25173 , n45629 );
and ( n45631 , n25172 , n45630 );
and ( n45632 , n25171 , n45631 );
and ( n45633 , n25170 , n45632 );
and ( n45634 , n25169 , n45633 );
and ( n45635 , n25168 , n45634 );
and ( n45636 , n25167 , n45635 );
and ( n45637 , n25166 , n45636 );
and ( n45638 , n25165 , n45637 );
and ( n45639 , n25164 , n45638 );
and ( n45640 , n25163 , n45639 );
and ( n45641 , n25162 , n45640 );
and ( n45642 , n25161 , n45641 );
and ( n45643 , n25160 , n45642 );
and ( n45644 , n25159 , n45643 );
and ( n45645 , n25158 , n45644 );
and ( n45646 , n25157 , n45645 );
and ( n45647 , n25156 , n45646 );
and ( n45648 , n25155 , n45647 );
and ( n45649 , n25154 , n45648 );
and ( n45650 , n25153 , n45649 );
and ( n45651 , n25152 , n45650 );
and ( n45652 , n25151 , n45651 );
and ( n45653 , n25150 , n45652 );
and ( n45654 , n25149 , n45653 );
and ( n45655 , n25148 , n45654 );
and ( n45656 , n25147 , n45655 );
and ( n45657 , n25146 , n45656 );
and ( n45658 , n25145 , n45657 );
and ( n45659 , n25144 , n45658 );
and ( n45660 , n25143 , n45659 );
and ( n45661 , n25142 , n45660 );
or ( n45662 , n25141 , n45661 );
and ( n45663 , n24269 , n45662 );
and ( n45664 , n24268 , n45663 );
and ( n45665 , n24267 , n45664 );
xor ( n45666 , n24266 , n45665 );
buf ( n45667 , n45666 );
buf ( n45668 , n45667 );
buf ( n45669 , n45668 );
xor ( n45670 , n20873 , n45669 );
and ( n45671 , n20868 , n45670 );
buf ( n45672 , n45671 );
and ( n45673 , n20871 , n20872 );
and ( n45674 , n20872 , n45669 );
and ( n45675 , n20871 , n45669 );
or ( n45676 , n45673 , n45674 , n45675 );
buf ( n45677 , n45676 );
not ( n45678 , n20860 );
and ( n45679 , n20855 , n20846 );
xor ( n45680 , n45678 , n45679 );
and ( n45681 , n20878 , n20881 );
and ( n45682 , n20881 , n20980 );
and ( n45683 , n20878 , n20980 );
or ( n45684 , n45681 , n45682 , n45683 );
or ( n45685 , n20981 , n24265 );
xnor ( n45686 , n45684 , n45685 );
and ( n45687 , n24266 , n45665 );
xor ( n45688 , n45686 , n45687 );
buf ( n45689 , n45688 );
buf ( n45690 , n45689 );
buf ( n45691 , n45690 );
xor ( n45692 , n45680 , n45691 );
xor ( n45693 , n45677 , n45692 );
xor ( n45694 , n45672 , n45693 );
xor ( n45695 , n24267 , n45664 );
buf ( n45696 , n45695 );
buf ( n45697 , n45696 );
buf ( n45698 , n45697 );
xor ( n45699 , n20834 , n20836 );
xor ( n45700 , n20836 , n20838 );
not ( n45701 , n45700 );
and ( n45702 , n45699 , n45701 );
and ( n45703 , n20855 , n45702 );
not ( n45704 , n45703 );
xnor ( n45705 , n45704 , n20841 );
and ( n45706 , n20864 , n20852 );
and ( n45707 , n20844 , n20850 );
nor ( n45708 , n45706 , n45707 );
xnor ( n45709 , n45708 , n20860 );
and ( n45710 , n45705 , n45709 );
buf ( n45711 , n20708 );
buf ( n45712 , n45711 );
and ( n45713 , n45712 , n20846 );
and ( n45714 , n45709 , n45713 );
and ( n45715 , n45705 , n45713 );
or ( n45716 , n45710 , n45714 , n45715 );
and ( n45717 , n45698 , n45716 );
buf ( n45718 , n45717 );
buf ( n45719 , n20868 );
xor ( n45720 , n45719 , n45670 );
and ( n45721 , n45718 , n45720 );
xor ( n45722 , n20842 , n20861 );
xor ( n45723 , n45722 , n20865 );
xor ( n45724 , n24268 , n45663 );
buf ( n45725 , n45724 );
buf ( n45726 , n45725 );
buf ( n45727 , n45726 );
buf ( n45728 , n17455 );
buf ( n45729 , n45728 );
buf ( n45730 , n17457 );
buf ( n45731 , n45730 );
and ( n45732 , n45729 , n45731 );
not ( n45733 , n45732 );
and ( n45734 , n20838 , n45733 );
not ( n45735 , n45734 );
and ( n45736 , n20844 , n45702 );
and ( n45737 , n20855 , n45700 );
nor ( n45738 , n45736 , n45737 );
xnor ( n45739 , n45738 , n20841 );
and ( n45740 , n45735 , n45739 );
and ( n45741 , n45712 , n20852 );
and ( n45742 , n20864 , n20850 );
nor ( n45743 , n45741 , n45742 );
xnor ( n45744 , n45743 , n20860 );
and ( n45745 , n45739 , n45744 );
and ( n45746 , n45735 , n45744 );
or ( n45747 , n45740 , n45745 , n45746 );
and ( n45748 , n45727 , n45747 );
buf ( n45749 , n45748 );
and ( n45750 , n45723 , n45749 );
buf ( n45751 , n45698 );
xor ( n45752 , n45751 , n45716 );
and ( n45753 , n45749 , n45752 );
and ( n45754 , n45723 , n45752 );
or ( n45755 , n45750 , n45753 , n45754 );
and ( n45756 , n45720 , n45755 );
and ( n45757 , n45718 , n45755 );
or ( n45758 , n45721 , n45756 , n45757 );
xor ( n45759 , n45694 , n45758 );
xor ( n45760 , n45718 , n45720 );
xor ( n45761 , n45760 , n45755 );
buf ( n45762 , n20708 );
buf ( n45763 , n45762 );
and ( n45764 , n45763 , n20846 );
xor ( n45765 , n24269 , n45662 );
buf ( n45766 , n45765 );
buf ( n45767 , n45766 );
buf ( n45768 , n45767 );
and ( n45769 , n45764 , n45768 );
buf ( n45770 , n45769 );
xor ( n45771 , n45705 , n45709 );
xor ( n45772 , n45771 , n45713 );
and ( n45773 , n45770 , n45772 );
xor ( n45774 , n20838 , n45729 );
xor ( n45775 , n45729 , n45731 );
not ( n45776 , n45775 );
and ( n45777 , n45774 , n45776 );
and ( n45778 , n20855 , n45777 );
not ( n45779 , n45778 );
xnor ( n45780 , n45779 , n45734 );
and ( n45781 , n20864 , n45702 );
and ( n45782 , n20844 , n45700 );
nor ( n45783 , n45781 , n45782 );
xnor ( n45784 , n45783 , n20841 );
and ( n45785 , n45780 , n45784 );
and ( n45786 , n45763 , n20852 );
and ( n45787 , n45712 , n20850 );
nor ( n45788 , n45786 , n45787 );
xnor ( n45789 , n45788 , n20860 );
and ( n45790 , n45784 , n45789 );
and ( n45791 , n45780 , n45789 );
or ( n45792 , n45785 , n45790 , n45791 );
buf ( n45793 , n20708 );
buf ( n45794 , n45793 );
and ( n45795 , n45794 , n20846 );
xor ( n45796 , n25142 , n45660 );
buf ( n45797 , n45796 );
buf ( n45798 , n45797 );
buf ( n45799 , n45798 );
and ( n45800 , n45795 , n45799 );
buf ( n45801 , n45800 );
and ( n45802 , n45792 , n45801 );
xor ( n45803 , n45735 , n45739 );
xor ( n45804 , n45803 , n45744 );
and ( n45805 , n45801 , n45804 );
and ( n45806 , n45792 , n45804 );
or ( n45807 , n45802 , n45805 , n45806 );
and ( n45808 , n45772 , n45807 );
and ( n45809 , n45770 , n45807 );
or ( n45810 , n45773 , n45808 , n45809 );
xor ( n45811 , n45723 , n45749 );
xor ( n45812 , n45811 , n45752 );
and ( n45813 , n45810 , n45812 );
buf ( n45814 , n45727 );
xor ( n45815 , n45814 , n45747 );
xor ( n45816 , n45764 , n45768 );
buf ( n45817 , n45816 );
buf ( n45818 , n17459 );
buf ( n45819 , n45818 );
buf ( n45820 , n17461 );
buf ( n45821 , n45820 );
and ( n45822 , n45819 , n45821 );
not ( n45823 , n45822 );
and ( n45824 , n45731 , n45823 );
not ( n45825 , n45824 );
and ( n45826 , n20844 , n45777 );
and ( n45827 , n20855 , n45775 );
nor ( n45828 , n45826 , n45827 );
xnor ( n45829 , n45828 , n45734 );
and ( n45830 , n45825 , n45829 );
and ( n45831 , n45712 , n45702 );
and ( n45832 , n20864 , n45700 );
nor ( n45833 , n45831 , n45832 );
xnor ( n45834 , n45833 , n20841 );
and ( n45835 , n45829 , n45834 );
and ( n45836 , n45825 , n45834 );
or ( n45837 , n45830 , n45835 , n45836 );
and ( n45838 , n45794 , n20852 );
and ( n45839 , n45763 , n20850 );
nor ( n45840 , n45838 , n45839 );
xnor ( n45841 , n45840 , n20860 );
buf ( n45842 , n20708 );
buf ( n45843 , n45842 );
and ( n45844 , n45843 , n20846 );
and ( n45845 , n45841 , n45844 );
xor ( n45846 , n25143 , n45659 );
buf ( n45847 , n45846 );
buf ( n45848 , n45847 );
buf ( n45849 , n45848 );
and ( n45850 , n45844 , n45849 );
and ( n45851 , n45841 , n45849 );
or ( n45852 , n45845 , n45850 , n45851 );
and ( n45853 , n45837 , n45852 );
xor ( n45854 , n45780 , n45784 );
xor ( n45855 , n45854 , n45789 );
and ( n45856 , n45852 , n45855 );
and ( n45857 , n45837 , n45855 );
or ( n45858 , n45853 , n45856 , n45857 );
and ( n45859 , n45817 , n45858 );
xor ( n45860 , n45792 , n45801 );
xor ( n45861 , n45860 , n45804 );
and ( n45862 , n45858 , n45861 );
and ( n45863 , n45817 , n45861 );
or ( n45864 , n45859 , n45862 , n45863 );
and ( n45865 , n45815 , n45864 );
xor ( n45866 , n45770 , n45772 );
xor ( n45867 , n45866 , n45807 );
and ( n45868 , n45864 , n45867 );
and ( n45869 , n45815 , n45867 );
or ( n45870 , n45865 , n45868 , n45869 );
and ( n45871 , n45812 , n45870 );
and ( n45872 , n45810 , n45870 );
or ( n45873 , n45813 , n45871 , n45872 );
or ( n45874 , n45761 , n45873 );
xor ( n45875 , n45759 , n45874 );
xnor ( n45876 , n45761 , n45873 );
xor ( n45877 , n45810 , n45812 );
xor ( n45878 , n45877 , n45870 );
xor ( n45879 , n45815 , n45864 );
xor ( n45880 , n45879 , n45867 );
xor ( n45881 , n45795 , n45799 );
buf ( n45882 , n45881 );
xor ( n45883 , n45731 , n45819 );
xor ( n45884 , n45819 , n45821 );
not ( n45885 , n45884 );
and ( n45886 , n45883 , n45885 );
and ( n45887 , n20855 , n45886 );
not ( n45888 , n45887 );
xnor ( n45889 , n45888 , n45824 );
and ( n45890 , n20864 , n45777 );
and ( n45891 , n20844 , n45775 );
nor ( n45892 , n45890 , n45891 );
xnor ( n45893 , n45892 , n45734 );
and ( n45894 , n45889 , n45893 );
and ( n45895 , n45763 , n45702 );
and ( n45896 , n45712 , n45700 );
nor ( n45897 , n45895 , n45896 );
xnor ( n45898 , n45897 , n20841 );
and ( n45899 , n45893 , n45898 );
and ( n45900 , n45889 , n45898 );
or ( n45901 , n45894 , n45899 , n45900 );
and ( n45902 , n45843 , n20852 );
and ( n45903 , n45794 , n20850 );
nor ( n45904 , n45902 , n45903 );
xnor ( n45905 , n45904 , n20860 );
buf ( n45906 , n20708 );
buf ( n45907 , n45906 );
and ( n45908 , n45907 , n20846 );
and ( n45909 , n45905 , n45908 );
xor ( n45910 , n25144 , n45658 );
buf ( n45911 , n45910 );
buf ( n45912 , n45911 );
buf ( n45913 , n45912 );
and ( n45914 , n45908 , n45913 );
and ( n45915 , n45905 , n45913 );
or ( n45916 , n45909 , n45914 , n45915 );
and ( n45917 , n45901 , n45916 );
buf ( n45918 , n45917 );
and ( n45919 , n45882 , n45918 );
xor ( n45920 , n45837 , n45852 );
xor ( n45921 , n45920 , n45855 );
and ( n45922 , n45918 , n45921 );
and ( n45923 , n45882 , n45921 );
or ( n45924 , n45919 , n45922 , n45923 );
xor ( n45925 , n45817 , n45858 );
xor ( n45926 , n45925 , n45861 );
and ( n45927 , n45924 , n45926 );
xor ( n45928 , n45825 , n45829 );
xor ( n45929 , n45928 , n45834 );
xor ( n45930 , n45841 , n45844 );
xor ( n45931 , n45930 , n45849 );
and ( n45932 , n45929 , n45931 );
buf ( n45933 , n17463 );
buf ( n45934 , n45933 );
buf ( n45935 , n17465 );
buf ( n45936 , n45935 );
and ( n45937 , n45934 , n45936 );
not ( n45938 , n45937 );
and ( n45939 , n45821 , n45938 );
not ( n45940 , n45939 );
and ( n45941 , n20844 , n45886 );
and ( n45942 , n20855 , n45884 );
nor ( n45943 , n45941 , n45942 );
xnor ( n45944 , n45943 , n45824 );
and ( n45945 , n45940 , n45944 );
and ( n45946 , n45712 , n45777 );
and ( n45947 , n20864 , n45775 );
nor ( n45948 , n45946 , n45947 );
xnor ( n45949 , n45948 , n45734 );
and ( n45950 , n45944 , n45949 );
and ( n45951 , n45940 , n45949 );
or ( n45952 , n45945 , n45950 , n45951 );
and ( n45953 , n45794 , n45702 );
and ( n45954 , n45763 , n45700 );
nor ( n45955 , n45953 , n45954 );
xnor ( n45956 , n45955 , n20841 );
and ( n45957 , n45907 , n20852 );
and ( n45958 , n45843 , n20850 );
nor ( n45959 , n45957 , n45958 );
xnor ( n45960 , n45959 , n20860 );
and ( n45961 , n45956 , n45960 );
buf ( n45962 , n20708 );
buf ( n45963 , n45962 );
and ( n45964 , n45963 , n20846 );
and ( n45965 , n45960 , n45964 );
and ( n45966 , n45956 , n45964 );
or ( n45967 , n45961 , n45965 , n45966 );
and ( n45968 , n45952 , n45967 );
buf ( n45969 , n45968 );
and ( n45970 , n45931 , n45969 );
and ( n45971 , n45929 , n45969 );
or ( n45972 , n45932 , n45970 , n45971 );
xor ( n45973 , n45882 , n45918 );
xor ( n45974 , n45973 , n45921 );
and ( n45975 , n45972 , n45974 );
buf ( n45976 , n45901 );
xor ( n45977 , n45976 , n45916 );
xor ( n45978 , n45889 , n45893 );
xor ( n45979 , n45978 , n45898 );
xor ( n45980 , n45905 , n45908 );
xor ( n45981 , n45980 , n45913 );
and ( n45982 , n45979 , n45981 );
xor ( n45983 , n25145 , n45657 );
buf ( n45984 , n45983 );
buf ( n45985 , n45984 );
buf ( n45986 , n45985 );
xor ( n45987 , n45821 , n45934 );
xor ( n45988 , n45934 , n45936 );
not ( n45989 , n45988 );
and ( n45990 , n45987 , n45989 );
and ( n45991 , n20855 , n45990 );
not ( n45992 , n45991 );
xnor ( n45993 , n45992 , n45939 );
and ( n45994 , n20864 , n45886 );
and ( n45995 , n20844 , n45884 );
nor ( n45996 , n45994 , n45995 );
xnor ( n45997 , n45996 , n45824 );
and ( n45998 , n45993 , n45997 );
and ( n45999 , n45763 , n45777 );
and ( n46000 , n45712 , n45775 );
nor ( n46001 , n45999 , n46000 );
xnor ( n46002 , n46001 , n45734 );
and ( n46003 , n45997 , n46002 );
and ( n46004 , n45993 , n46002 );
or ( n46005 , n45998 , n46003 , n46004 );
and ( n46006 , n45986 , n46005 );
buf ( n46007 , n46006 );
and ( n46008 , n45981 , n46007 );
and ( n46009 , n45979 , n46007 );
or ( n46010 , n45982 , n46008 , n46009 );
and ( n46011 , n45977 , n46010 );
xor ( n46012 , n45929 , n45931 );
xor ( n46013 , n46012 , n45969 );
and ( n46014 , n46010 , n46013 );
and ( n46015 , n45977 , n46013 );
or ( n46016 , n46011 , n46014 , n46015 );
and ( n46017 , n45974 , n46016 );
and ( n46018 , n45972 , n46016 );
or ( n46019 , n45975 , n46017 , n46018 );
and ( n46020 , n45926 , n46019 );
and ( n46021 , n45924 , n46019 );
or ( n46022 , n45927 , n46020 , n46021 );
or ( n46023 , n45880 , n46022 );
and ( n46024 , n45878 , n46023 );
xor ( n46025 , n45878 , n46023 );
xnor ( n46026 , n45880 , n46022 );
xor ( n46027 , n45924 , n45926 );
xor ( n46028 , n46027 , n46019 );
xor ( n46029 , n45972 , n45974 );
xor ( n46030 , n46029 , n46016 );
and ( n46031 , n45843 , n45702 );
and ( n46032 , n45794 , n45700 );
nor ( n46033 , n46031 , n46032 );
xnor ( n46034 , n46033 , n20841 );
and ( n46035 , n45963 , n20852 );
and ( n46036 , n45907 , n20850 );
nor ( n46037 , n46035 , n46036 );
xnor ( n46038 , n46037 , n20860 );
and ( n46039 , n46034 , n46038 );
buf ( n46040 , n20708 );
buf ( n46041 , n46040 );
and ( n46042 , n46041 , n20846 );
and ( n46043 , n46038 , n46042 );
and ( n46044 , n46034 , n46042 );
or ( n46045 , n46039 , n46043 , n46044 );
xor ( n46046 , n45940 , n45944 );
xor ( n46047 , n46046 , n45949 );
and ( n46048 , n46045 , n46047 );
xor ( n46049 , n45956 , n45960 );
xor ( n46050 , n46049 , n45964 );
and ( n46051 , n46047 , n46050 );
and ( n46052 , n46045 , n46050 );
or ( n46053 , n46048 , n46051 , n46052 );
buf ( n46054 , n45952 );
xor ( n46055 , n46054 , n45967 );
and ( n46056 , n46053 , n46055 );
xor ( n46057 , n25146 , n45656 );
buf ( n46058 , n46057 );
buf ( n46059 , n46058 );
buf ( n46060 , n46059 );
buf ( n46061 , n17467 );
buf ( n46062 , n46061 );
buf ( n46063 , n17469 );
buf ( n46064 , n46063 );
and ( n46065 , n46062 , n46064 );
not ( n46066 , n46065 );
and ( n46067 , n45936 , n46066 );
not ( n46068 , n46067 );
and ( n46069 , n20844 , n45990 );
and ( n46070 , n20855 , n45988 );
nor ( n46071 , n46069 , n46070 );
xnor ( n46072 , n46071 , n45939 );
and ( n46073 , n46068 , n46072 );
and ( n46074 , n45712 , n45886 );
and ( n46075 , n20864 , n45884 );
nor ( n46076 , n46074 , n46075 );
xnor ( n46077 , n46076 , n45824 );
and ( n46078 , n46072 , n46077 );
and ( n46079 , n46068 , n46077 );
or ( n46080 , n46073 , n46078 , n46079 );
and ( n46081 , n46060 , n46080 );
buf ( n46082 , n46081 );
and ( n46083 , n45794 , n45777 );
and ( n46084 , n45763 , n45775 );
nor ( n46085 , n46083 , n46084 );
xnor ( n46086 , n46085 , n45734 );
and ( n46087 , n45907 , n45702 );
and ( n46088 , n45843 , n45700 );
nor ( n46089 , n46087 , n46088 );
xnor ( n46090 , n46089 , n20841 );
and ( n46091 , n46086 , n46090 );
and ( n46092 , n46041 , n20852 );
and ( n46093 , n45963 , n20850 );
nor ( n46094 , n46092 , n46093 );
xnor ( n46095 , n46094 , n20860 );
and ( n46096 , n46090 , n46095 );
and ( n46097 , n46086 , n46095 );
or ( n46098 , n46091 , n46096 , n46097 );
buf ( n46099 , n20710 );
buf ( n46100 , n46099 );
and ( n46101 , n46100 , n20846 );
xor ( n46102 , n25147 , n45655 );
buf ( n46103 , n46102 );
buf ( n46104 , n46103 );
buf ( n46105 , n46104 );
and ( n46106 , n46101 , n46105 );
buf ( n46107 , n46106 );
and ( n46108 , n46098 , n46107 );
xor ( n46109 , n45993 , n45997 );
xor ( n46110 , n46109 , n46002 );
and ( n46111 , n46107 , n46110 );
and ( n46112 , n46098 , n46110 );
or ( n46113 , n46108 , n46111 , n46112 );
and ( n46114 , n46082 , n46113 );
buf ( n46115 , n45986 );
xor ( n46116 , n46115 , n46005 );
and ( n46117 , n46113 , n46116 );
and ( n46118 , n46082 , n46116 );
or ( n46119 , n46114 , n46117 , n46118 );
and ( n46120 , n46055 , n46119 );
and ( n46121 , n46053 , n46119 );
or ( n46122 , n46056 , n46120 , n46121 );
xor ( n46123 , n45977 , n46010 );
xor ( n46124 , n46123 , n46013 );
and ( n46125 , n46122 , n46124 );
xor ( n46126 , n45979 , n45981 );
xor ( n46127 , n46126 , n46007 );
xor ( n46128 , n46045 , n46047 );
xor ( n46129 , n46128 , n46050 );
xor ( n46130 , n46034 , n46038 );
xor ( n46131 , n46130 , n46042 );
xor ( n46132 , n45936 , n46062 );
xor ( n46133 , n46062 , n46064 );
not ( n46134 , n46133 );
and ( n46135 , n46132 , n46134 );
and ( n46136 , n20855 , n46135 );
not ( n46137 , n46136 );
xnor ( n46138 , n46137 , n46067 );
and ( n46139 , n20864 , n45990 );
and ( n46140 , n20844 , n45988 );
nor ( n46141 , n46139 , n46140 );
xnor ( n46142 , n46141 , n45939 );
and ( n46143 , n46138 , n46142 );
and ( n46144 , n45763 , n45886 );
and ( n46145 , n45712 , n45884 );
nor ( n46146 , n46144 , n46145 );
xnor ( n46147 , n46146 , n45824 );
and ( n46148 , n46142 , n46147 );
and ( n46149 , n46138 , n46147 );
or ( n46150 , n46143 , n46148 , n46149 );
and ( n46151 , n45843 , n45777 );
and ( n46152 , n45794 , n45775 );
nor ( n46153 , n46151 , n46152 );
xnor ( n46154 , n46153 , n45734 );
and ( n46155 , n45963 , n45702 );
and ( n46156 , n45907 , n45700 );
nor ( n46157 , n46155 , n46156 );
xnor ( n46158 , n46157 , n20841 );
and ( n46159 , n46154 , n46158 );
and ( n46160 , n46100 , n20852 );
and ( n46161 , n46041 , n20850 );
nor ( n46162 , n46160 , n46161 );
xnor ( n46163 , n46162 , n20860 );
and ( n46164 , n46158 , n46163 );
and ( n46165 , n46154 , n46163 );
or ( n46166 , n46159 , n46164 , n46165 );
and ( n46167 , n46150 , n46166 );
buf ( n46168 , n20712 );
buf ( n46169 , n46168 );
and ( n46170 , n46169 , n20846 );
xor ( n46171 , n25148 , n45654 );
buf ( n46172 , n46171 );
buf ( n46173 , n46172 );
buf ( n46174 , n46173 );
and ( n46175 , n46170 , n46174 );
buf ( n46176 , n46175 );
and ( n46177 , n46166 , n46176 );
and ( n46178 , n46150 , n46176 );
or ( n46179 , n46167 , n46177 , n46178 );
and ( n46180 , n46131 , n46179 );
xor ( n46181 , n46068 , n46072 );
xor ( n46182 , n46181 , n46077 );
xor ( n46183 , n46086 , n46090 );
xor ( n46184 , n46183 , n46095 );
and ( n46185 , n46182 , n46184 );
xor ( n46186 , n46101 , n46105 );
buf ( n46187 , n46186 );
and ( n46188 , n46184 , n46187 );
and ( n46189 , n46182 , n46187 );
or ( n46190 , n46185 , n46188 , n46189 );
and ( n46191 , n46179 , n46190 );
and ( n46192 , n46131 , n46190 );
or ( n46193 , n46180 , n46191 , n46192 );
and ( n46194 , n46129 , n46193 );
xor ( n46195 , n46082 , n46113 );
xor ( n46196 , n46195 , n46116 );
and ( n46197 , n46193 , n46196 );
and ( n46198 , n46129 , n46196 );
or ( n46199 , n46194 , n46197 , n46198 );
and ( n46200 , n46127 , n46199 );
xor ( n46201 , n46053 , n46055 );
xor ( n46202 , n46201 , n46119 );
and ( n46203 , n46199 , n46202 );
and ( n46204 , n46127 , n46202 );
or ( n46205 , n46200 , n46203 , n46204 );
and ( n46206 , n46124 , n46205 );
and ( n46207 , n46122 , n46205 );
or ( n46208 , n46125 , n46206 , n46207 );
or ( n46209 , n46030 , n46208 );
and ( n46210 , n46028 , n46209 );
xor ( n46211 , n46028 , n46209 );
xnor ( n46212 , n46030 , n46208 );
xor ( n46213 , n46122 , n46124 );
xor ( n46214 , n46213 , n46205 );
xor ( n46215 , n46127 , n46199 );
xor ( n46216 , n46215 , n46202 );
buf ( n46217 , n46060 );
xor ( n46218 , n46217 , n46080 );
xor ( n46219 , n46098 , n46107 );
xor ( n46220 , n46219 , n46110 );
and ( n46221 , n46218 , n46220 );
buf ( n46222 , n17471 );
buf ( n46223 , n46222 );
buf ( n46224 , n17473 );
buf ( n46225 , n46224 );
and ( n46226 , n46223 , n46225 );
not ( n46227 , n46226 );
and ( n46228 , n46064 , n46227 );
not ( n46229 , n46228 );
and ( n46230 , n20844 , n46135 );
and ( n46231 , n20855 , n46133 );
nor ( n46232 , n46230 , n46231 );
xnor ( n46233 , n46232 , n46067 );
and ( n46234 , n46229 , n46233 );
and ( n46235 , n45712 , n45990 );
and ( n46236 , n20864 , n45988 );
nor ( n46237 , n46235 , n46236 );
xnor ( n46238 , n46237 , n45939 );
and ( n46239 , n46233 , n46238 );
and ( n46240 , n46229 , n46238 );
or ( n46241 , n46234 , n46239 , n46240 );
and ( n46242 , n45794 , n45886 );
and ( n46243 , n45763 , n45884 );
nor ( n46244 , n46242 , n46243 );
xnor ( n46245 , n46244 , n45824 );
and ( n46246 , n45907 , n45777 );
and ( n46247 , n45843 , n45775 );
nor ( n46248 , n46246 , n46247 );
xnor ( n46249 , n46248 , n45734 );
and ( n46250 , n46245 , n46249 );
and ( n46251 , n46041 , n45702 );
and ( n46252 , n45963 , n45700 );
nor ( n46253 , n46251 , n46252 );
xnor ( n46254 , n46253 , n20841 );
and ( n46255 , n46249 , n46254 );
and ( n46256 , n46245 , n46254 );
or ( n46257 , n46250 , n46255 , n46256 );
and ( n46258 , n46241 , n46257 );
and ( n46259 , n46169 , n20852 );
and ( n46260 , n46100 , n20850 );
nor ( n46261 , n46259 , n46260 );
xnor ( n46262 , n46261 , n20860 );
buf ( n46263 , n20714 );
buf ( n46264 , n46263 );
and ( n46265 , n46264 , n20846 );
and ( n46266 , n46262 , n46265 );
xor ( n46267 , n25149 , n45653 );
buf ( n46268 , n46267 );
buf ( n46269 , n46268 );
buf ( n46270 , n46269 );
and ( n46271 , n46265 , n46270 );
and ( n46272 , n46262 , n46270 );
or ( n46273 , n46266 , n46271 , n46272 );
and ( n46274 , n46257 , n46273 );
and ( n46275 , n46241 , n46273 );
or ( n46276 , n46258 , n46274 , n46275 );
xor ( n46277 , n46138 , n46142 );
xor ( n46278 , n46277 , n46147 );
xor ( n46279 , n46154 , n46158 );
xor ( n46280 , n46279 , n46163 );
and ( n46281 , n46278 , n46280 );
xor ( n46282 , n46170 , n46174 );
buf ( n46283 , n46282 );
and ( n46284 , n46280 , n46283 );
and ( n46285 , n46278 , n46283 );
or ( n46286 , n46281 , n46284 , n46285 );
and ( n46287 , n46276 , n46286 );
xor ( n46288 , n46150 , n46166 );
xor ( n46289 , n46288 , n46176 );
and ( n46290 , n46286 , n46289 );
and ( n46291 , n46276 , n46289 );
or ( n46292 , n46287 , n46290 , n46291 );
and ( n46293 , n46220 , n46292 );
and ( n46294 , n46218 , n46292 );
or ( n46295 , n46221 , n46293 , n46294 );
xor ( n46296 , n46129 , n46193 );
xor ( n46297 , n46296 , n46196 );
and ( n46298 , n46295 , n46297 );
xor ( n46299 , n46131 , n46179 );
xor ( n46300 , n46299 , n46190 );
xor ( n46301 , n46182 , n46184 );
xor ( n46302 , n46301 , n46187 );
xor ( n46303 , n46064 , n46223 );
xor ( n46304 , n46223 , n46225 );
not ( n46305 , n46304 );
and ( n46306 , n46303 , n46305 );
and ( n46307 , n20855 , n46306 );
not ( n46308 , n46307 );
xnor ( n46309 , n46308 , n46228 );
and ( n46310 , n20864 , n46135 );
and ( n46311 , n20844 , n46133 );
nor ( n46312 , n46310 , n46311 );
xnor ( n46313 , n46312 , n46067 );
and ( n46314 , n46309 , n46313 );
and ( n46315 , n45763 , n45990 );
and ( n46316 , n45712 , n45988 );
nor ( n46317 , n46315 , n46316 );
xnor ( n46318 , n46317 , n45939 );
and ( n46319 , n46313 , n46318 );
and ( n46320 , n46309 , n46318 );
or ( n46321 , n46314 , n46319 , n46320 );
and ( n46322 , n45843 , n45886 );
and ( n46323 , n45794 , n45884 );
nor ( n46324 , n46322 , n46323 );
xnor ( n46325 , n46324 , n45824 );
and ( n46326 , n45963 , n45777 );
and ( n46327 , n45907 , n45775 );
nor ( n46328 , n46326 , n46327 );
xnor ( n46329 , n46328 , n45734 );
and ( n46330 , n46325 , n46329 );
and ( n46331 , n46100 , n45702 );
and ( n46332 , n46041 , n45700 );
nor ( n46333 , n46331 , n46332 );
xnor ( n46334 , n46333 , n20841 );
and ( n46335 , n46329 , n46334 );
and ( n46336 , n46325 , n46334 );
or ( n46337 , n46330 , n46335 , n46336 );
and ( n46338 , n46321 , n46337 );
buf ( n46339 , n46338 );
and ( n46340 , n46264 , n20852 );
and ( n46341 , n46169 , n20850 );
nor ( n46342 , n46340 , n46341 );
xnor ( n46343 , n46342 , n20860 );
buf ( n46344 , n20716 );
buf ( n46345 , n46344 );
and ( n46346 , n46345 , n20846 );
and ( n46347 , n46343 , n46346 );
xor ( n46348 , n25150 , n45652 );
buf ( n46349 , n46348 );
buf ( n46350 , n46349 );
buf ( n46351 , n46350 );
and ( n46352 , n46346 , n46351 );
and ( n46353 , n46343 , n46351 );
or ( n46354 , n46347 , n46352 , n46353 );
xor ( n46355 , n46229 , n46233 );
xor ( n46356 , n46355 , n46238 );
and ( n46357 , n46354 , n46356 );
xor ( n46358 , n46245 , n46249 );
xor ( n46359 , n46358 , n46254 );
and ( n46360 , n46356 , n46359 );
and ( n46361 , n46354 , n46359 );
or ( n46362 , n46357 , n46360 , n46361 );
and ( n46363 , n46339 , n46362 );
xor ( n46364 , n46241 , n46257 );
xor ( n46365 , n46364 , n46273 );
and ( n46366 , n46362 , n46365 );
and ( n46367 , n46339 , n46365 );
or ( n46368 , n46363 , n46366 , n46367 );
and ( n46369 , n46302 , n46368 );
xor ( n46370 , n46276 , n46286 );
xor ( n46371 , n46370 , n46289 );
and ( n46372 , n46368 , n46371 );
and ( n46373 , n46302 , n46371 );
or ( n46374 , n46369 , n46372 , n46373 );
and ( n46375 , n46300 , n46374 );
xor ( n46376 , n46218 , n46220 );
xor ( n46377 , n46376 , n46292 );
and ( n46378 , n46374 , n46377 );
and ( n46379 , n46300 , n46377 );
or ( n46380 , n46375 , n46378 , n46379 );
and ( n46381 , n46297 , n46380 );
and ( n46382 , n46295 , n46380 );
or ( n46383 , n46298 , n46381 , n46382 );
or ( n46384 , n46216 , n46383 );
and ( n46385 , n46214 , n46384 );
xor ( n46386 , n46214 , n46384 );
xnor ( n46387 , n46216 , n46383 );
xor ( n46388 , n46295 , n46297 );
xor ( n46389 , n46388 , n46380 );
xor ( n46390 , n46300 , n46374 );
xor ( n46391 , n46390 , n46377 );
xor ( n46392 , n46278 , n46280 );
xor ( n46393 , n46392 , n46283 );
xor ( n46394 , n46262 , n46265 );
xor ( n46395 , n46394 , n46270 );
buf ( n46396 , n17475 );
buf ( n46397 , n46396 );
buf ( n46398 , n17477 );
buf ( n46399 , n46398 );
and ( n46400 , n46397 , n46399 );
not ( n46401 , n46400 );
and ( n46402 , n46225 , n46401 );
not ( n46403 , n46402 );
and ( n46404 , n20844 , n46306 );
and ( n46405 , n20855 , n46304 );
nor ( n46406 , n46404 , n46405 );
xnor ( n46407 , n46406 , n46228 );
and ( n46408 , n46403 , n46407 );
and ( n46409 , n45712 , n46135 );
and ( n46410 , n20864 , n46133 );
nor ( n46411 , n46409 , n46410 );
xnor ( n46412 , n46411 , n46067 );
and ( n46413 , n46407 , n46412 );
and ( n46414 , n46403 , n46412 );
or ( n46415 , n46408 , n46413 , n46414 );
and ( n46416 , n45794 , n45990 );
and ( n46417 , n45763 , n45988 );
nor ( n46418 , n46416 , n46417 );
xnor ( n46419 , n46418 , n45939 );
and ( n46420 , n45907 , n45886 );
and ( n46421 , n45843 , n45884 );
nor ( n46422 , n46420 , n46421 );
xnor ( n46423 , n46422 , n45824 );
and ( n46424 , n46419 , n46423 );
and ( n46425 , n46041 , n45777 );
and ( n46426 , n45963 , n45775 );
nor ( n46427 , n46425 , n46426 );
xnor ( n46428 , n46427 , n45734 );
and ( n46429 , n46423 , n46428 );
and ( n46430 , n46419 , n46428 );
or ( n46431 , n46424 , n46429 , n46430 );
and ( n46432 , n46415 , n46431 );
buf ( n46433 , n46432 );
and ( n46434 , n46395 , n46433 );
and ( n46435 , n46169 , n45702 );
and ( n46436 , n46100 , n45700 );
nor ( n46437 , n46435 , n46436 );
xnor ( n46438 , n46437 , n20841 );
and ( n46439 , n46345 , n20852 );
and ( n46440 , n46264 , n20850 );
nor ( n46441 , n46439 , n46440 );
xnor ( n46442 , n46441 , n20860 );
and ( n46443 , n46438 , n46442 );
buf ( n46444 , n20718 );
buf ( n46445 , n46444 );
and ( n46446 , n46445 , n20846 );
and ( n46447 , n46442 , n46446 );
and ( n46448 , n46438 , n46446 );
or ( n46449 , n46443 , n46447 , n46448 );
xor ( n46450 , n46309 , n46313 );
xor ( n46451 , n46450 , n46318 );
and ( n46452 , n46449 , n46451 );
xor ( n46453 , n46325 , n46329 );
xor ( n46454 , n46453 , n46334 );
and ( n46455 , n46451 , n46454 );
and ( n46456 , n46449 , n46454 );
or ( n46457 , n46452 , n46455 , n46456 );
and ( n46458 , n46433 , n46457 );
and ( n46459 , n46395 , n46457 );
or ( n46460 , n46434 , n46458 , n46459 );
and ( n46461 , n46393 , n46460 );
xor ( n46462 , n46339 , n46362 );
xor ( n46463 , n46462 , n46365 );
and ( n46464 , n46460 , n46463 );
and ( n46465 , n46393 , n46463 );
or ( n46466 , n46461 , n46464 , n46465 );
xor ( n46467 , n46302 , n46368 );
xor ( n46468 , n46467 , n46371 );
and ( n46469 , n46466 , n46468 );
buf ( n46470 , n46321 );
xor ( n46471 , n46470 , n46337 );
xor ( n46472 , n46354 , n46356 );
xor ( n46473 , n46472 , n46359 );
and ( n46474 , n46471 , n46473 );
xor ( n46475 , n46343 , n46346 );
xor ( n46476 , n46475 , n46351 );
xor ( n46477 , n25151 , n45651 );
buf ( n46478 , n46477 );
buf ( n46479 , n46478 );
buf ( n46480 , n46479 );
and ( n46481 , n46264 , n45702 );
and ( n46482 , n46169 , n45700 );
nor ( n46483 , n46481 , n46482 );
xnor ( n46484 , n46483 , n20841 );
and ( n46485 , n46445 , n20852 );
and ( n46486 , n46345 , n20850 );
nor ( n46487 , n46485 , n46486 );
xnor ( n46488 , n46487 , n20860 );
and ( n46489 , n46484 , n46488 );
and ( n46490 , n46480 , n46489 );
buf ( n46491 , n46490 );
and ( n46492 , n46476 , n46491 );
xor ( n46493 , n46225 , n46397 );
xor ( n46494 , n46397 , n46399 );
not ( n46495 , n46494 );
and ( n46496 , n46493 , n46495 );
and ( n46497 , n20855 , n46496 );
not ( n46498 , n46497 );
xnor ( n46499 , n46498 , n46402 );
and ( n46500 , n20864 , n46306 );
and ( n46501 , n20844 , n46304 );
nor ( n46502 , n46500 , n46501 );
xnor ( n46503 , n46502 , n46228 );
and ( n46504 , n46499 , n46503 );
and ( n46505 , n45763 , n46135 );
and ( n46506 , n45712 , n46133 );
nor ( n46507 , n46505 , n46506 );
xnor ( n46508 , n46507 , n46067 );
and ( n46509 , n46503 , n46508 );
and ( n46510 , n46499 , n46508 );
or ( n46511 , n46504 , n46509 , n46510 );
and ( n46512 , n45843 , n45990 );
and ( n46513 , n45794 , n45988 );
nor ( n46514 , n46512 , n46513 );
xnor ( n46515 , n46514 , n45939 );
and ( n46516 , n45963 , n45886 );
and ( n46517 , n45907 , n45884 );
nor ( n46518 , n46516 , n46517 );
xnor ( n46519 , n46518 , n45824 );
and ( n46520 , n46515 , n46519 );
and ( n46521 , n46100 , n45777 );
and ( n46522 , n46041 , n45775 );
nor ( n46523 , n46521 , n46522 );
xnor ( n46524 , n46523 , n45734 );
and ( n46525 , n46519 , n46524 );
and ( n46526 , n46515 , n46524 );
or ( n46527 , n46520 , n46525 , n46526 );
and ( n46528 , n46511 , n46527 );
buf ( n46529 , n20720 );
buf ( n46530 , n46529 );
and ( n46531 , n46530 , n20846 );
xor ( n46532 , n25152 , n45650 );
buf ( n46533 , n46532 );
buf ( n46534 , n46533 );
buf ( n46535 , n46534 );
and ( n46536 , n46531 , n46535 );
buf ( n46537 , n46536 );
and ( n46538 , n46527 , n46537 );
and ( n46539 , n46511 , n46537 );
or ( n46540 , n46528 , n46538 , n46539 );
and ( n46541 , n46491 , n46540 );
and ( n46542 , n46476 , n46540 );
or ( n46543 , n46492 , n46541 , n46542 );
and ( n46544 , n46473 , n46543 );
and ( n46545 , n46471 , n46543 );
or ( n46546 , n46474 , n46544 , n46545 );
xor ( n46547 , n46393 , n46460 );
xor ( n46548 , n46547 , n46463 );
and ( n46549 , n46546 , n46548 );
xor ( n46550 , n46403 , n46407 );
xor ( n46551 , n46550 , n46412 );
xor ( n46552 , n46419 , n46423 );
xor ( n46553 , n46552 , n46428 );
and ( n46554 , n46551 , n46553 );
xor ( n46555 , n46438 , n46442 );
xor ( n46556 , n46555 , n46446 );
and ( n46557 , n46553 , n46556 );
and ( n46558 , n46551 , n46556 );
or ( n46559 , n46554 , n46557 , n46558 );
buf ( n46560 , n46415 );
xor ( n46561 , n46560 , n46431 );
and ( n46562 , n46559 , n46561 );
xor ( n46563 , n46449 , n46451 );
xor ( n46564 , n46563 , n46454 );
and ( n46565 , n46561 , n46564 );
and ( n46566 , n46559 , n46564 );
or ( n46567 , n46562 , n46565 , n46566 );
xor ( n46568 , n46395 , n46433 );
xor ( n46569 , n46568 , n46457 );
and ( n46570 , n46567 , n46569 );
xor ( n46571 , n46484 , n46488 );
and ( n46572 , n46530 , n20852 );
and ( n46573 , n46445 , n20850 );
nor ( n46574 , n46572 , n46573 );
xnor ( n46575 , n46574 , n20860 );
buf ( n46576 , n20722 );
buf ( n46577 , n46576 );
and ( n46578 , n46577 , n20846 );
and ( n46579 , n46575 , n46578 );
and ( n46580 , n46571 , n46579 );
buf ( n46581 , n17479 );
buf ( n46582 , n46581 );
buf ( n46583 , n17481 );
buf ( n46584 , n46583 );
and ( n46585 , n46582 , n46584 );
not ( n46586 , n46585 );
and ( n46587 , n46399 , n46586 );
not ( n46588 , n46587 );
and ( n46589 , n20844 , n46496 );
and ( n46590 , n20855 , n46494 );
nor ( n46591 , n46589 , n46590 );
xnor ( n46592 , n46591 , n46402 );
and ( n46593 , n46588 , n46592 );
and ( n46594 , n45712 , n46306 );
and ( n46595 , n20864 , n46304 );
nor ( n46596 , n46594 , n46595 );
xnor ( n46597 , n46596 , n46228 );
and ( n46598 , n46592 , n46597 );
and ( n46599 , n46588 , n46597 );
or ( n46600 , n46593 , n46598 , n46599 );
and ( n46601 , n46579 , n46600 );
and ( n46602 , n46571 , n46600 );
or ( n46603 , n46580 , n46601 , n46602 );
and ( n46604 , n45794 , n46135 );
and ( n46605 , n45763 , n46133 );
nor ( n46606 , n46604 , n46605 );
xnor ( n46607 , n46606 , n46067 );
and ( n46608 , n45907 , n45990 );
and ( n46609 , n45843 , n45988 );
nor ( n46610 , n46608 , n46609 );
xnor ( n46611 , n46610 , n45939 );
and ( n46612 , n46607 , n46611 );
and ( n46613 , n46041 , n45886 );
and ( n46614 , n45963 , n45884 );
nor ( n46615 , n46613 , n46614 );
xnor ( n46616 , n46615 , n45824 );
and ( n46617 , n46611 , n46616 );
and ( n46618 , n46607 , n46616 );
or ( n46619 , n46612 , n46617 , n46618 );
and ( n46620 , n46169 , n45777 );
and ( n46621 , n46100 , n45775 );
nor ( n46622 , n46620 , n46621 );
xnor ( n46623 , n46622 , n45734 );
and ( n46624 , n46345 , n45702 );
and ( n46625 , n46264 , n45700 );
nor ( n46626 , n46624 , n46625 );
xnor ( n46627 , n46626 , n20841 );
and ( n46628 , n46623 , n46627 );
xor ( n46629 , n25153 , n45649 );
buf ( n46630 , n46629 );
buf ( n46631 , n46630 );
buf ( n46632 , n46631 );
and ( n46633 , n46627 , n46632 );
and ( n46634 , n46623 , n46632 );
or ( n46635 , n46628 , n46633 , n46634 );
and ( n46636 , n46619 , n46635 );
xor ( n46637 , n46499 , n46503 );
xor ( n46638 , n46637 , n46508 );
and ( n46639 , n46635 , n46638 );
and ( n46640 , n46619 , n46638 );
or ( n46641 , n46636 , n46639 , n46640 );
and ( n46642 , n46603 , n46641 );
buf ( n46643 , n46480 );
xor ( n46644 , n46643 , n46489 );
and ( n46645 , n46641 , n46644 );
and ( n46646 , n46603 , n46644 );
or ( n46647 , n46642 , n46645 , n46646 );
xor ( n46648 , n46476 , n46491 );
xor ( n46649 , n46648 , n46540 );
and ( n46650 , n46647 , n46649 );
xor ( n46651 , n46559 , n46561 );
xor ( n46652 , n46651 , n46564 );
and ( n46653 , n46649 , n46652 );
and ( n46654 , n46647 , n46652 );
or ( n46655 , n46650 , n46653 , n46654 );
and ( n46656 , n46569 , n46655 );
and ( n46657 , n46567 , n46655 );
or ( n46658 , n46570 , n46656 , n46657 );
and ( n46659 , n46548 , n46658 );
and ( n46660 , n46546 , n46658 );
or ( n46661 , n46549 , n46659 , n46660 );
and ( n46662 , n46468 , n46661 );
and ( n46663 , n46466 , n46661 );
or ( n46664 , n46469 , n46662 , n46663 );
or ( n46665 , n46391 , n46664 );
and ( n46666 , n46389 , n46665 );
xor ( n46667 , n46389 , n46665 );
xnor ( n46668 , n46391 , n46664 );
xor ( n46669 , n46466 , n46468 );
xor ( n46670 , n46669 , n46661 );
xor ( n46671 , n46546 , n46548 );
xor ( n46672 , n46671 , n46658 );
xor ( n46673 , n46471 , n46473 );
xor ( n46674 , n46673 , n46543 );
xor ( n46675 , n46567 , n46569 );
xor ( n46676 , n46675 , n46655 );
and ( n46677 , n46674 , n46676 );
xor ( n46678 , n46511 , n46527 );
xor ( n46679 , n46678 , n46537 );
xor ( n46680 , n46551 , n46553 );
xor ( n46681 , n46680 , n46556 );
and ( n46682 , n46679 , n46681 );
xor ( n46683 , n46515 , n46519 );
xor ( n46684 , n46683 , n46524 );
xor ( n46685 , n46531 , n46535 );
buf ( n46686 , n46685 );
and ( n46687 , n46684 , n46686 );
xor ( n46688 , n46575 , n46578 );
and ( n46689 , n46445 , n45702 );
and ( n46690 , n46345 , n45700 );
nor ( n46691 , n46689 , n46690 );
xnor ( n46692 , n46691 , n20841 );
and ( n46693 , n46577 , n20852 );
and ( n46694 , n46530 , n20850 );
nor ( n46695 , n46693 , n46694 );
xnor ( n46696 , n46695 , n20860 );
and ( n46697 , n46692 , n46696 );
and ( n46698 , n46688 , n46697 );
buf ( n46699 , n46698 );
and ( n46700 , n46686 , n46699 );
and ( n46701 , n46684 , n46699 );
or ( n46702 , n46687 , n46700 , n46701 );
and ( n46703 , n46681 , n46702 );
and ( n46704 , n46679 , n46702 );
or ( n46705 , n46682 , n46703 , n46704 );
xor ( n46706 , n46647 , n46649 );
xor ( n46707 , n46706 , n46652 );
and ( n46708 , n46705 , n46707 );
xor ( n46709 , n46399 , n46582 );
xor ( n46710 , n46582 , n46584 );
not ( n46711 , n46710 );
and ( n46712 , n46709 , n46711 );
and ( n46713 , n20855 , n46712 );
not ( n46714 , n46713 );
xnor ( n46715 , n46714 , n46587 );
and ( n46716 , n20864 , n46496 );
and ( n46717 , n20844 , n46494 );
nor ( n46718 , n46716 , n46717 );
xnor ( n46719 , n46718 , n46402 );
and ( n46720 , n46715 , n46719 );
and ( n46721 , n45763 , n46306 );
and ( n46722 , n45712 , n46304 );
nor ( n46723 , n46721 , n46722 );
xnor ( n46724 , n46723 , n46228 );
and ( n46725 , n46719 , n46724 );
and ( n46726 , n46715 , n46724 );
or ( n46727 , n46720 , n46725 , n46726 );
and ( n46728 , n45843 , n46135 );
and ( n46729 , n45794 , n46133 );
nor ( n46730 , n46728 , n46729 );
xnor ( n46731 , n46730 , n46067 );
and ( n46732 , n45963 , n45990 );
and ( n46733 , n45907 , n45988 );
nor ( n46734 , n46732 , n46733 );
xnor ( n46735 , n46734 , n45939 );
and ( n46736 , n46731 , n46735 );
and ( n46737 , n46100 , n45886 );
and ( n46738 , n46041 , n45884 );
nor ( n46739 , n46737 , n46738 );
xnor ( n46740 , n46739 , n45824 );
and ( n46741 , n46735 , n46740 );
and ( n46742 , n46731 , n46740 );
or ( n46743 , n46736 , n46741 , n46742 );
and ( n46744 , n46727 , n46743 );
and ( n46745 , n46264 , n45777 );
and ( n46746 , n46169 , n45775 );
nor ( n46747 , n46745 , n46746 );
xnor ( n46748 , n46747 , n45734 );
buf ( n46749 , n20724 );
buf ( n46750 , n46749 );
and ( n46751 , n46750 , n20846 );
and ( n46752 , n46748 , n46751 );
xor ( n46753 , n25154 , n45648 );
buf ( n46754 , n46753 );
buf ( n46755 , n46754 );
buf ( n46756 , n46755 );
and ( n46757 , n46751 , n46756 );
and ( n46758 , n46748 , n46756 );
or ( n46759 , n46752 , n46757 , n46758 );
and ( n46760 , n46743 , n46759 );
and ( n46761 , n46727 , n46759 );
or ( n46762 , n46744 , n46760 , n46761 );
xor ( n46763 , n46588 , n46592 );
xor ( n46764 , n46763 , n46597 );
xor ( n46765 , n46607 , n46611 );
xor ( n46766 , n46765 , n46616 );
and ( n46767 , n46764 , n46766 );
xor ( n46768 , n46623 , n46627 );
xor ( n46769 , n46768 , n46632 );
and ( n46770 , n46766 , n46769 );
and ( n46771 , n46764 , n46769 );
or ( n46772 , n46767 , n46770 , n46771 );
and ( n46773 , n46762 , n46772 );
xor ( n46774 , n46571 , n46579 );
xor ( n46775 , n46774 , n46600 );
and ( n46776 , n46772 , n46775 );
and ( n46777 , n46762 , n46775 );
or ( n46778 , n46773 , n46776 , n46777 );
xor ( n46779 , n46603 , n46641 );
xor ( n46780 , n46779 , n46644 );
and ( n46781 , n46778 , n46780 );
xor ( n46782 , n46619 , n46635 );
xor ( n46783 , n46782 , n46638 );
xor ( n46784 , n46692 , n46696 );
and ( n46785 , n46530 , n45702 );
and ( n46786 , n46445 , n45700 );
nor ( n46787 , n46785 , n46786 );
xnor ( n46788 , n46787 , n20841 );
and ( n46789 , n46750 , n20852 );
and ( n46790 , n46577 , n20850 );
nor ( n46791 , n46789 , n46790 );
xnor ( n46792 , n46791 , n20860 );
or ( n46793 , n46788 , n46792 );
and ( n46794 , n46784 , n46793 );
buf ( n46795 , n46794 );
buf ( n46796 , n17483 );
buf ( n46797 , n46796 );
buf ( n46798 , n17485 );
buf ( n46799 , n46798 );
and ( n46800 , n46797 , n46799 );
not ( n46801 , n46800 );
and ( n46802 , n46584 , n46801 );
not ( n46803 , n46802 );
and ( n46804 , n20844 , n46712 );
and ( n46805 , n20855 , n46710 );
nor ( n46806 , n46804 , n46805 );
xnor ( n46807 , n46806 , n46587 );
and ( n46808 , n46803 , n46807 );
and ( n46809 , n45712 , n46496 );
and ( n46810 , n20864 , n46494 );
nor ( n46811 , n46809 , n46810 );
xnor ( n46812 , n46811 , n46402 );
and ( n46813 , n46807 , n46812 );
and ( n46814 , n46803 , n46812 );
or ( n46815 , n46808 , n46813 , n46814 );
and ( n46816 , n45794 , n46306 );
and ( n46817 , n45763 , n46304 );
nor ( n46818 , n46816 , n46817 );
xnor ( n46819 , n46818 , n46228 );
and ( n46820 , n45907 , n46135 );
and ( n46821 , n45843 , n46133 );
nor ( n46822 , n46820 , n46821 );
xnor ( n46823 , n46822 , n46067 );
and ( n46824 , n46819 , n46823 );
and ( n46825 , n46041 , n45990 );
and ( n46826 , n45963 , n45988 );
nor ( n46827 , n46825 , n46826 );
xnor ( n46828 , n46827 , n45939 );
and ( n46829 , n46823 , n46828 );
and ( n46830 , n46819 , n46828 );
or ( n46831 , n46824 , n46829 , n46830 );
and ( n46832 , n46815 , n46831 );
and ( n46833 , n46169 , n45886 );
and ( n46834 , n46100 , n45884 );
nor ( n46835 , n46833 , n46834 );
xnor ( n46836 , n46835 , n45824 );
and ( n46837 , n46345 , n45777 );
and ( n46838 , n46264 , n45775 );
nor ( n46839 , n46837 , n46838 );
xnor ( n46840 , n46839 , n45734 );
and ( n46841 , n46836 , n46840 );
buf ( n46842 , n20726 );
buf ( n46843 , n46842 );
and ( n46844 , n46843 , n20846 );
and ( n46845 , n46840 , n46844 );
and ( n46846 , n46836 , n46844 );
or ( n46847 , n46841 , n46845 , n46846 );
and ( n46848 , n46831 , n46847 );
and ( n46849 , n46815 , n46847 );
or ( n46850 , n46832 , n46848 , n46849 );
and ( n46851 , n46795 , n46850 );
xor ( n46852 , n46715 , n46719 );
xor ( n46853 , n46852 , n46724 );
xor ( n46854 , n46731 , n46735 );
xor ( n46855 , n46854 , n46740 );
and ( n46856 , n46853 , n46855 );
xor ( n46857 , n46748 , n46751 );
xor ( n46858 , n46857 , n46756 );
and ( n46859 , n46855 , n46858 );
and ( n46860 , n46853 , n46858 );
or ( n46861 , n46856 , n46859 , n46860 );
and ( n46862 , n46850 , n46861 );
and ( n46863 , n46795 , n46861 );
or ( n46864 , n46851 , n46862 , n46863 );
and ( n46865 , n46783 , n46864 );
buf ( n46866 , n46688 );
xor ( n46867 , n46866 , n46697 );
xor ( n46868 , n46727 , n46743 );
xor ( n46869 , n46868 , n46759 );
and ( n46870 , n46867 , n46869 );
xor ( n46871 , n46764 , n46766 );
xor ( n46872 , n46871 , n46769 );
and ( n46873 , n46869 , n46872 );
and ( n46874 , n46867 , n46872 );
or ( n46875 , n46870 , n46873 , n46874 );
and ( n46876 , n46864 , n46875 );
and ( n46877 , n46783 , n46875 );
or ( n46878 , n46865 , n46876 , n46877 );
and ( n46879 , n46780 , n46878 );
and ( n46880 , n46778 , n46878 );
or ( n46881 , n46781 , n46879 , n46880 );
and ( n46882 , n46707 , n46881 );
and ( n46883 , n46705 , n46881 );
or ( n46884 , n46708 , n46882 , n46883 );
and ( n46885 , n46676 , n46884 );
and ( n46886 , n46674 , n46884 );
or ( n46887 , n46677 , n46885 , n46886 );
or ( n46888 , n46672 , n46887 );
and ( n46889 , n46670 , n46888 );
xor ( n46890 , n46670 , n46888 );
xnor ( n46891 , n46672 , n46887 );
xor ( n46892 , n46674 , n46676 );
xor ( n46893 , n46892 , n46884 );
xor ( n46894 , n46679 , n46681 );
xor ( n46895 , n46894 , n46702 );
xor ( n46896 , n46684 , n46686 );
xor ( n46897 , n46896 , n46699 );
xor ( n46898 , n46762 , n46772 );
xor ( n46899 , n46898 , n46775 );
and ( n46900 , n46897 , n46899 );
xor ( n46901 , n25155 , n45647 );
buf ( n46902 , n46901 );
buf ( n46903 , n46902 );
buf ( n46904 , n46903 );
xnor ( n46905 , n46788 , n46792 );
and ( n46906 , n46904 , n46905 );
buf ( n46907 , n46906 );
xor ( n46908 , n46584 , n46797 );
xor ( n46909 , n46797 , n46799 );
not ( n46910 , n46909 );
and ( n46911 , n46908 , n46910 );
and ( n46912 , n20855 , n46911 );
not ( n46913 , n46912 );
xnor ( n46914 , n46913 , n46802 );
and ( n46915 , n20864 , n46712 );
and ( n46916 , n20844 , n46710 );
nor ( n46917 , n46915 , n46916 );
xnor ( n46918 , n46917 , n46587 );
and ( n46919 , n46914 , n46918 );
and ( n46920 , n45763 , n46496 );
and ( n46921 , n45712 , n46494 );
nor ( n46922 , n46920 , n46921 );
xnor ( n46923 , n46922 , n46402 );
and ( n46924 , n46918 , n46923 );
and ( n46925 , n46914 , n46923 );
or ( n46926 , n46919 , n46924 , n46925 );
and ( n46927 , n45843 , n46306 );
and ( n46928 , n45794 , n46304 );
nor ( n46929 , n46927 , n46928 );
xnor ( n46930 , n46929 , n46228 );
and ( n46931 , n45963 , n46135 );
and ( n46932 , n45907 , n46133 );
nor ( n46933 , n46931 , n46932 );
xnor ( n46934 , n46933 , n46067 );
and ( n46935 , n46930 , n46934 );
and ( n46936 , n46100 , n45990 );
and ( n46937 , n46041 , n45988 );
nor ( n46938 , n46936 , n46937 );
xnor ( n46939 , n46938 , n45939 );
and ( n46940 , n46934 , n46939 );
and ( n46941 , n46930 , n46939 );
or ( n46942 , n46935 , n46940 , n46941 );
and ( n46943 , n46926 , n46942 );
and ( n46944 , n46264 , n45886 );
and ( n46945 , n46169 , n45884 );
nor ( n46946 , n46944 , n46945 );
xnor ( n46947 , n46946 , n45824 );
and ( n46948 , n46445 , n45777 );
and ( n46949 , n46345 , n45775 );
nor ( n46950 , n46948 , n46949 );
xnor ( n46951 , n46950 , n45734 );
and ( n46952 , n46947 , n46951 );
and ( n46953 , n46577 , n45702 );
and ( n46954 , n46530 , n45700 );
nor ( n46955 , n46953 , n46954 );
xnor ( n46956 , n46955 , n20841 );
and ( n46957 , n46951 , n46956 );
and ( n46958 , n46947 , n46956 );
or ( n46959 , n46952 , n46957 , n46958 );
and ( n46960 , n46942 , n46959 );
and ( n46961 , n46926 , n46959 );
or ( n46962 , n46943 , n46960 , n46961 );
and ( n46963 , n46907 , n46962 );
and ( n46964 , n46843 , n20852 );
and ( n46965 , n46750 , n20850 );
nor ( n46966 , n46964 , n46965 );
xnor ( n46967 , n46966 , n20860 );
buf ( n46968 , n20728 );
buf ( n46969 , n46968 );
and ( n46970 , n46969 , n20846 );
and ( n46971 , n46967 , n46970 );
xor ( n46972 , n25156 , n45646 );
buf ( n46973 , n46972 );
buf ( n46974 , n46973 );
buf ( n46975 , n46974 );
and ( n46976 , n46970 , n46975 );
and ( n46977 , n46967 , n46975 );
or ( n46978 , n46971 , n46976 , n46977 );
xor ( n46979 , n46803 , n46807 );
xor ( n46980 , n46979 , n46812 );
and ( n46981 , n46978 , n46980 );
xor ( n46982 , n46819 , n46823 );
xor ( n46983 , n46982 , n46828 );
and ( n46984 , n46980 , n46983 );
and ( n46985 , n46978 , n46983 );
or ( n46986 , n46981 , n46984 , n46985 );
and ( n46987 , n46962 , n46986 );
and ( n46988 , n46907 , n46986 );
or ( n46989 , n46963 , n46987 , n46988 );
buf ( n46990 , n46784 );
xor ( n46991 , n46990 , n46793 );
xor ( n46992 , n46815 , n46831 );
xor ( n46993 , n46992 , n46847 );
and ( n46994 , n46991 , n46993 );
xor ( n46995 , n46853 , n46855 );
xor ( n46996 , n46995 , n46858 );
and ( n46997 , n46993 , n46996 );
and ( n46998 , n46991 , n46996 );
or ( n46999 , n46994 , n46997 , n46998 );
and ( n47000 , n46989 , n46999 );
xor ( n47001 , n46795 , n46850 );
xor ( n47002 , n47001 , n46861 );
and ( n47003 , n46999 , n47002 );
and ( n47004 , n46989 , n47002 );
or ( n47005 , n47000 , n47003 , n47004 );
and ( n47006 , n46899 , n47005 );
and ( n47007 , n46897 , n47005 );
or ( n47008 , n46900 , n47006 , n47007 );
and ( n47009 , n46895 , n47008 );
xor ( n47010 , n46778 , n46780 );
xor ( n47011 , n47010 , n46878 );
and ( n47012 , n47008 , n47011 );
and ( n47013 , n46895 , n47011 );
or ( n47014 , n47009 , n47012 , n47013 );
xor ( n47015 , n46705 , n46707 );
xor ( n47016 , n47015 , n46881 );
and ( n47017 , n47014 , n47016 );
xor ( n47018 , n46783 , n46864 );
xor ( n47019 , n47018 , n46875 );
xor ( n47020 , n46867 , n46869 );
xor ( n47021 , n47020 , n46872 );
xor ( n47022 , n46836 , n46840 );
xor ( n47023 , n47022 , n46844 );
and ( n47024 , n46345 , n45886 );
and ( n47025 , n46264 , n45884 );
nor ( n47026 , n47024 , n47025 );
xnor ( n47027 , n47026 , n45824 );
and ( n47028 , n46530 , n45777 );
and ( n47029 , n46445 , n45775 );
nor ( n47030 , n47028 , n47029 );
xnor ( n47031 , n47030 , n45734 );
or ( n47032 , n47027 , n47031 );
buf ( n47033 , n17487 );
buf ( n47034 , n47033 );
buf ( n47035 , n17489 );
buf ( n47036 , n47035 );
and ( n47037 , n47034 , n47036 );
not ( n47038 , n47037 );
and ( n47039 , n46799 , n47038 );
not ( n47040 , n47039 );
and ( n47041 , n20844 , n46911 );
and ( n47042 , n20855 , n46909 );
nor ( n47043 , n47041 , n47042 );
xnor ( n47044 , n47043 , n46802 );
and ( n47045 , n47040 , n47044 );
and ( n47046 , n45712 , n46712 );
and ( n47047 , n20864 , n46710 );
nor ( n47048 , n47046 , n47047 );
xnor ( n47049 , n47048 , n46587 );
and ( n47050 , n47044 , n47049 );
and ( n47051 , n47040 , n47049 );
or ( n47052 , n47045 , n47050 , n47051 );
and ( n47053 , n47032 , n47052 );
buf ( n47054 , n47053 );
and ( n47055 , n47023 , n47054 );
and ( n47056 , n45794 , n46496 );
and ( n47057 , n45763 , n46494 );
nor ( n47058 , n47056 , n47057 );
xnor ( n47059 , n47058 , n46402 );
and ( n47060 , n45907 , n46306 );
and ( n47061 , n45843 , n46304 );
nor ( n47062 , n47060 , n47061 );
xnor ( n47063 , n47062 , n46228 );
and ( n47064 , n47059 , n47063 );
and ( n47065 , n46041 , n46135 );
and ( n47066 , n45963 , n46133 );
nor ( n47067 , n47065 , n47066 );
xnor ( n47068 , n47067 , n46067 );
and ( n47069 , n47063 , n47068 );
and ( n47070 , n47059 , n47068 );
or ( n47071 , n47064 , n47069 , n47070 );
and ( n47072 , n46169 , n45990 );
and ( n47073 , n46100 , n45988 );
nor ( n47074 , n47072 , n47073 );
xnor ( n47075 , n47074 , n45939 );
and ( n47076 , n46750 , n45702 );
and ( n47077 , n46577 , n45700 );
nor ( n47078 , n47076 , n47077 );
xnor ( n47079 , n47078 , n20841 );
and ( n47080 , n47075 , n47079 );
and ( n47081 , n46969 , n20852 );
and ( n47082 , n46843 , n20850 );
nor ( n47083 , n47081 , n47082 );
xnor ( n47084 , n47083 , n20860 );
and ( n47085 , n47079 , n47084 );
and ( n47086 , n47075 , n47084 );
or ( n47087 , n47080 , n47085 , n47086 );
and ( n47088 , n47071 , n47087 );
buf ( n47089 , n20730 );
buf ( n47090 , n47089 );
and ( n47091 , n47090 , n20846 );
xor ( n47092 , n25157 , n45645 );
buf ( n47093 , n47092 );
buf ( n47094 , n47093 );
buf ( n47095 , n47094 );
and ( n47096 , n47091 , n47095 );
buf ( n47097 , n47096 );
and ( n47098 , n47087 , n47097 );
and ( n47099 , n47071 , n47097 );
or ( n47100 , n47088 , n47098 , n47099 );
and ( n47101 , n47054 , n47100 );
and ( n47102 , n47023 , n47100 );
or ( n47103 , n47055 , n47101 , n47102 );
xor ( n47104 , n46914 , n46918 );
xor ( n47105 , n47104 , n46923 );
xor ( n47106 , n46930 , n46934 );
xor ( n47107 , n47106 , n46939 );
and ( n47108 , n47105 , n47107 );
xor ( n47109 , n46947 , n46951 );
xor ( n47110 , n47109 , n46956 );
and ( n47111 , n47107 , n47110 );
and ( n47112 , n47105 , n47110 );
or ( n47113 , n47108 , n47111 , n47112 );
buf ( n47114 , n46904 );
xor ( n47115 , n47114 , n46905 );
and ( n47116 , n47113 , n47115 );
xor ( n47117 , n46926 , n46942 );
xor ( n47118 , n47117 , n46959 );
and ( n47119 , n47115 , n47118 );
and ( n47120 , n47113 , n47118 );
or ( n47121 , n47116 , n47119 , n47120 );
and ( n47122 , n47103 , n47121 );
xor ( n47123 , n46907 , n46962 );
xor ( n47124 , n47123 , n46986 );
and ( n47125 , n47121 , n47124 );
and ( n47126 , n47103 , n47124 );
or ( n47127 , n47122 , n47125 , n47126 );
and ( n47128 , n47021 , n47127 );
xor ( n47129 , n46989 , n46999 );
xor ( n47130 , n47129 , n47002 );
and ( n47131 , n47127 , n47130 );
and ( n47132 , n47021 , n47130 );
or ( n47133 , n47128 , n47131 , n47132 );
and ( n47134 , n47019 , n47133 );
xor ( n47135 , n46897 , n46899 );
xor ( n47136 , n47135 , n47005 );
and ( n47137 , n47133 , n47136 );
and ( n47138 , n47019 , n47136 );
or ( n47139 , n47134 , n47137 , n47138 );
xor ( n47140 , n46895 , n47008 );
xor ( n47141 , n47140 , n47011 );
and ( n47142 , n47139 , n47141 );
xor ( n47143 , n47019 , n47133 );
xor ( n47144 , n47143 , n47136 );
xor ( n47145 , n46991 , n46993 );
xor ( n47146 , n47145 , n46996 );
xor ( n47147 , n46978 , n46980 );
xor ( n47148 , n47147 , n46983 );
xor ( n47149 , n46967 , n46970 );
xor ( n47150 , n47149 , n46975 );
xnor ( n47151 , n47027 , n47031 );
and ( n47152 , n46264 , n45990 );
and ( n47153 , n46169 , n45988 );
nor ( n47154 , n47152 , n47153 );
xnor ( n47155 , n47154 , n45939 );
and ( n47156 , n46843 , n45702 );
and ( n47157 , n46750 , n45700 );
nor ( n47158 , n47156 , n47157 );
xnor ( n47159 , n47158 , n20841 );
or ( n47160 , n47155 , n47159 );
and ( n47161 , n47151 , n47160 );
and ( n47162 , n46577 , n45777 );
and ( n47163 , n46530 , n45775 );
nor ( n47164 , n47162 , n47163 );
xnor ( n47165 , n47164 , n45734 );
and ( n47166 , n47090 , n20852 );
and ( n47167 , n46969 , n20850 );
nor ( n47168 , n47166 , n47167 );
xnor ( n47169 , n47168 , n20860 );
and ( n47170 , n47165 , n47169 );
and ( n47171 , n47160 , n47170 );
and ( n47172 , n47151 , n47170 );
or ( n47173 , n47161 , n47171 , n47172 );
and ( n47174 , n47150 , n47173 );
xor ( n47175 , n46799 , n47034 );
xor ( n47176 , n47034 , n47036 );
not ( n47177 , n47176 );
and ( n47178 , n47175 , n47177 );
and ( n47179 , n20855 , n47178 );
not ( n47180 , n47179 );
xnor ( n47181 , n47180 , n47039 );
and ( n47182 , n20864 , n46911 );
and ( n47183 , n20844 , n46909 );
nor ( n47184 , n47182 , n47183 );
xnor ( n47185 , n47184 , n46802 );
and ( n47186 , n47181 , n47185 );
and ( n47187 , n45763 , n46712 );
and ( n47188 , n45712 , n46710 );
nor ( n47189 , n47187 , n47188 );
xnor ( n47190 , n47189 , n46587 );
and ( n47191 , n47185 , n47190 );
and ( n47192 , n47181 , n47190 );
or ( n47193 , n47186 , n47191 , n47192 );
and ( n47194 , n45843 , n46496 );
and ( n47195 , n45794 , n46494 );
nor ( n47196 , n47194 , n47195 );
xnor ( n47197 , n47196 , n46402 );
and ( n47198 , n45963 , n46306 );
and ( n47199 , n45907 , n46304 );
nor ( n47200 , n47198 , n47199 );
xnor ( n47201 , n47200 , n46228 );
and ( n47202 , n47197 , n47201 );
and ( n47203 , n46100 , n46135 );
and ( n47204 , n46041 , n46133 );
nor ( n47205 , n47203 , n47204 );
xnor ( n47206 , n47205 , n46067 );
and ( n47207 , n47201 , n47206 );
and ( n47208 , n47197 , n47206 );
or ( n47209 , n47202 , n47207 , n47208 );
and ( n47210 , n47193 , n47209 );
and ( n47211 , n46445 , n45886 );
and ( n47212 , n46345 , n45884 );
nor ( n47213 , n47211 , n47212 );
xnor ( n47214 , n47213 , n45824 );
buf ( n47215 , n20732 );
buf ( n47216 , n47215 );
and ( n47217 , n47216 , n20846 );
and ( n47218 , n47214 , n47217 );
xor ( n47219 , n25158 , n45644 );
buf ( n47220 , n47219 );
buf ( n47221 , n47220 );
buf ( n47222 , n47221 );
and ( n47223 , n47217 , n47222 );
and ( n47224 , n47214 , n47222 );
or ( n47225 , n47218 , n47223 , n47224 );
and ( n47226 , n47209 , n47225 );
and ( n47227 , n47193 , n47225 );
or ( n47228 , n47210 , n47226 , n47227 );
and ( n47229 , n47173 , n47228 );
and ( n47230 , n47150 , n47228 );
or ( n47231 , n47174 , n47229 , n47230 );
and ( n47232 , n47148 , n47231 );
xor ( n47233 , n47040 , n47044 );
xor ( n47234 , n47233 , n47049 );
xor ( n47235 , n47059 , n47063 );
xor ( n47236 , n47235 , n47068 );
and ( n47237 , n47234 , n47236 );
xor ( n47238 , n47075 , n47079 );
xor ( n47239 , n47238 , n47084 );
and ( n47240 , n47236 , n47239 );
and ( n47241 , n47234 , n47239 );
or ( n47242 , n47237 , n47240 , n47241 );
buf ( n47243 , n47032 );
xor ( n47244 , n47243 , n47052 );
and ( n47245 , n47242 , n47244 );
xor ( n47246 , n47071 , n47087 );
xor ( n47247 , n47246 , n47097 );
and ( n47248 , n47244 , n47247 );
and ( n47249 , n47242 , n47247 );
or ( n47250 , n47245 , n47248 , n47249 );
and ( n47251 , n47231 , n47250 );
and ( n47252 , n47148 , n47250 );
or ( n47253 , n47232 , n47251 , n47252 );
and ( n47254 , n47146 , n47253 );
xor ( n47255 , n47103 , n47121 );
xor ( n47256 , n47255 , n47124 );
and ( n47257 , n47253 , n47256 );
and ( n47258 , n47146 , n47256 );
or ( n47259 , n47254 , n47257 , n47258 );
xor ( n47260 , n47021 , n47127 );
xor ( n47261 , n47260 , n47130 );
and ( n47262 , n47259 , n47261 );
xor ( n47263 , n47023 , n47054 );
xor ( n47264 , n47263 , n47100 );
xor ( n47265 , n47113 , n47115 );
xor ( n47266 , n47265 , n47118 );
and ( n47267 , n47264 , n47266 );
xor ( n47268 , n47105 , n47107 );
xor ( n47269 , n47268 , n47110 );
xor ( n47270 , n47091 , n47095 );
buf ( n47271 , n47270 );
xnor ( n47272 , n47155 , n47159 );
xor ( n47273 , n47165 , n47169 );
and ( n47274 , n47272 , n47273 );
buf ( n47275 , n47274 );
and ( n47276 , n47271 , n47275 );
and ( n47277 , n46530 , n45886 );
and ( n47278 , n46445 , n45884 );
nor ( n47279 , n47277 , n47278 );
xnor ( n47280 , n47279 , n45824 );
and ( n47281 , n46750 , n45777 );
and ( n47282 , n46577 , n45775 );
nor ( n47283 , n47281 , n47282 );
xnor ( n47284 , n47283 , n45734 );
and ( n47285 , n47280 , n47284 );
and ( n47286 , n46969 , n45702 );
and ( n47287 , n46843 , n45700 );
nor ( n47288 , n47286 , n47287 );
xnor ( n47289 , n47288 , n20841 );
and ( n47290 , n47284 , n47289 );
and ( n47291 , n47280 , n47289 );
or ( n47292 , n47285 , n47290 , n47291 );
and ( n47293 , n46345 , n45990 );
and ( n47294 , n46264 , n45988 );
nor ( n47295 , n47293 , n47294 );
xnor ( n47296 , n47295 , n45939 );
and ( n47297 , n47216 , n20852 );
and ( n47298 , n47090 , n20850 );
nor ( n47299 , n47297 , n47298 );
xnor ( n47300 , n47299 , n20860 );
or ( n47301 , n47296 , n47300 );
and ( n47302 , n47292 , n47301 );
buf ( n47303 , n17491 );
buf ( n47304 , n47303 );
buf ( n47305 , n17493 );
buf ( n47306 , n47305 );
and ( n47307 , n47304 , n47306 );
not ( n47308 , n47307 );
and ( n47309 , n47036 , n47308 );
not ( n47310 , n47309 );
and ( n47311 , n20844 , n47178 );
and ( n47312 , n20855 , n47176 );
nor ( n47313 , n47311 , n47312 );
xnor ( n47314 , n47313 , n47039 );
and ( n47315 , n47310 , n47314 );
and ( n47316 , n45712 , n46911 );
and ( n47317 , n20864 , n46909 );
nor ( n47318 , n47316 , n47317 );
xnor ( n47319 , n47318 , n46802 );
and ( n47320 , n47314 , n47319 );
and ( n47321 , n47310 , n47319 );
or ( n47322 , n47315 , n47320 , n47321 );
and ( n47323 , n47301 , n47322 );
and ( n47324 , n47292 , n47322 );
or ( n47325 , n47302 , n47323 , n47324 );
and ( n47326 , n47275 , n47325 );
and ( n47327 , n47271 , n47325 );
or ( n47328 , n47276 , n47326 , n47327 );
and ( n47329 , n47269 , n47328 );
and ( n47330 , n45794 , n46712 );
and ( n47331 , n45763 , n46710 );
nor ( n47332 , n47330 , n47331 );
xnor ( n47333 , n47332 , n46587 );
and ( n47334 , n45907 , n46496 );
and ( n47335 , n45843 , n46494 );
nor ( n47336 , n47334 , n47335 );
xnor ( n47337 , n47336 , n46402 );
and ( n47338 , n47333 , n47337 );
and ( n47339 , n46041 , n46306 );
and ( n47340 , n45963 , n46304 );
nor ( n47341 , n47339 , n47340 );
xnor ( n47342 , n47341 , n46228 );
and ( n47343 , n47337 , n47342 );
and ( n47344 , n47333 , n47342 );
or ( n47345 , n47338 , n47343 , n47344 );
and ( n47346 , n46169 , n46135 );
and ( n47347 , n46100 , n46133 );
nor ( n47348 , n47346 , n47347 );
xnor ( n47349 , n47348 , n46067 );
buf ( n47350 , n20734 );
buf ( n47351 , n47350 );
and ( n47352 , n47351 , n20846 );
and ( n47353 , n47349 , n47352 );
xor ( n47354 , n25159 , n45643 );
buf ( n47355 , n47354 );
buf ( n47356 , n47355 );
buf ( n47357 , n47356 );
and ( n47358 , n47352 , n47357 );
and ( n47359 , n47349 , n47357 );
or ( n47360 , n47353 , n47358 , n47359 );
and ( n47361 , n47345 , n47360 );
xor ( n47362 , n47181 , n47185 );
xor ( n47363 , n47362 , n47190 );
and ( n47364 , n47360 , n47363 );
and ( n47365 , n47345 , n47363 );
or ( n47366 , n47361 , n47364 , n47365 );
xor ( n47367 , n47151 , n47160 );
xor ( n47368 , n47367 , n47170 );
and ( n47369 , n47366 , n47368 );
xor ( n47370 , n47193 , n47209 );
xor ( n47371 , n47370 , n47225 );
and ( n47372 , n47368 , n47371 );
and ( n47373 , n47366 , n47371 );
or ( n47374 , n47369 , n47372 , n47373 );
and ( n47375 , n47328 , n47374 );
and ( n47376 , n47269 , n47374 );
or ( n47377 , n47329 , n47375 , n47376 );
and ( n47378 , n47266 , n47377 );
and ( n47379 , n47264 , n47377 );
or ( n47380 , n47267 , n47378 , n47379 );
xor ( n47381 , n47146 , n47253 );
xor ( n47382 , n47381 , n47256 );
and ( n47383 , n47380 , n47382 );
xor ( n47384 , n47148 , n47231 );
xor ( n47385 , n47384 , n47250 );
xor ( n47386 , n47150 , n47173 );
xor ( n47387 , n47386 , n47228 );
xor ( n47388 , n47242 , n47244 );
xor ( n47389 , n47388 , n47247 );
and ( n47390 , n47387 , n47389 );
xor ( n47391 , n47234 , n47236 );
xor ( n47392 , n47391 , n47239 );
xor ( n47393 , n47197 , n47201 );
xor ( n47394 , n47393 , n47206 );
xor ( n47395 , n47214 , n47217 );
xor ( n47396 , n47395 , n47222 );
and ( n47397 , n47394 , n47396 );
xor ( n47398 , n47280 , n47284 );
xor ( n47399 , n47398 , n47289 );
xnor ( n47400 , n47296 , n47300 );
and ( n47401 , n47399 , n47400 );
buf ( n47402 , n47401 );
and ( n47403 , n47396 , n47402 );
and ( n47404 , n47394 , n47402 );
or ( n47405 , n47397 , n47403 , n47404 );
and ( n47406 , n47392 , n47405 );
and ( n47407 , n46445 , n45990 );
and ( n47408 , n46345 , n45988 );
nor ( n47409 , n47407 , n47408 );
xnor ( n47410 , n47409 , n45939 );
and ( n47411 , n47351 , n20852 );
and ( n47412 , n47216 , n20850 );
nor ( n47413 , n47411 , n47412 );
xnor ( n47414 , n47413 , n20860 );
and ( n47415 , n47410 , n47414 );
and ( n47416 , n46577 , n45886 );
and ( n47417 , n46530 , n45884 );
nor ( n47418 , n47416 , n47417 );
xnor ( n47419 , n47418 , n45824 );
and ( n47420 , n46843 , n45777 );
and ( n47421 , n46750 , n45775 );
nor ( n47422 , n47420 , n47421 );
xnor ( n47423 , n47422 , n45734 );
and ( n47424 , n47419 , n47423 );
and ( n47425 , n47415 , n47424 );
xor ( n47426 , n47036 , n47304 );
xor ( n47427 , n47304 , n47306 );
not ( n47428 , n47427 );
and ( n47429 , n47426 , n47428 );
and ( n47430 , n20855 , n47429 );
not ( n47431 , n47430 );
xnor ( n47432 , n47431 , n47309 );
and ( n47433 , n20864 , n47178 );
and ( n47434 , n20844 , n47176 );
nor ( n47435 , n47433 , n47434 );
xnor ( n47436 , n47435 , n47039 );
and ( n47437 , n47432 , n47436 );
and ( n47438 , n45763 , n46911 );
and ( n47439 , n45712 , n46909 );
nor ( n47440 , n47438 , n47439 );
xnor ( n47441 , n47440 , n46802 );
and ( n47442 , n47436 , n47441 );
and ( n47443 , n47432 , n47441 );
or ( n47444 , n47437 , n47442 , n47443 );
and ( n47445 , n47424 , n47444 );
and ( n47446 , n47415 , n47444 );
or ( n47447 , n47425 , n47445 , n47446 );
and ( n47448 , n45843 , n46712 );
and ( n47449 , n45794 , n46710 );
nor ( n47450 , n47448 , n47449 );
xnor ( n47451 , n47450 , n46587 );
and ( n47452 , n45963 , n46496 );
and ( n47453 , n45907 , n46494 );
nor ( n47454 , n47452 , n47453 );
xnor ( n47455 , n47454 , n46402 );
and ( n47456 , n47451 , n47455 );
and ( n47457 , n46100 , n46306 );
and ( n47458 , n46041 , n46304 );
nor ( n47459 , n47457 , n47458 );
xnor ( n47460 , n47459 , n46228 );
and ( n47461 , n47455 , n47460 );
and ( n47462 , n47451 , n47460 );
or ( n47463 , n47456 , n47461 , n47462 );
and ( n47464 , n46264 , n46135 );
and ( n47465 , n46169 , n46133 );
nor ( n47466 , n47464 , n47465 );
xnor ( n47467 , n47466 , n46067 );
and ( n47468 , n47090 , n45702 );
and ( n47469 , n46969 , n45700 );
nor ( n47470 , n47468 , n47469 );
xnor ( n47471 , n47470 , n20841 );
and ( n47472 , n47467 , n47471 );
buf ( n47473 , n20736 );
buf ( n47474 , n47473 );
and ( n47475 , n47474 , n20846 );
and ( n47476 , n47471 , n47475 );
and ( n47477 , n47467 , n47475 );
or ( n47478 , n47472 , n47476 , n47477 );
and ( n47479 , n47463 , n47478 );
xor ( n47480 , n47310 , n47314 );
xor ( n47481 , n47480 , n47319 );
and ( n47482 , n47478 , n47481 );
and ( n47483 , n47463 , n47481 );
or ( n47484 , n47479 , n47482 , n47483 );
and ( n47485 , n47447 , n47484 );
buf ( n47486 , n47272 );
xor ( n47487 , n47486 , n47273 );
and ( n47488 , n47484 , n47487 );
and ( n47489 , n47447 , n47487 );
or ( n47490 , n47485 , n47488 , n47489 );
and ( n47491 , n47405 , n47490 );
and ( n47492 , n47392 , n47490 );
or ( n47493 , n47406 , n47491 , n47492 );
and ( n47494 , n47389 , n47493 );
and ( n47495 , n47387 , n47493 );
or ( n47496 , n47390 , n47494 , n47495 );
and ( n47497 , n47385 , n47496 );
xor ( n47498 , n47264 , n47266 );
xor ( n47499 , n47498 , n47377 );
and ( n47500 , n47496 , n47499 );
and ( n47501 , n47385 , n47499 );
or ( n47502 , n47497 , n47500 , n47501 );
and ( n47503 , n47382 , n47502 );
and ( n47504 , n47380 , n47502 );
or ( n47505 , n47383 , n47503 , n47504 );
and ( n47506 , n47261 , n47505 );
and ( n47507 , n47259 , n47505 );
or ( n47508 , n47262 , n47506 , n47507 );
or ( n47509 , n47144 , n47508 );
and ( n47510 , n47141 , n47509 );
and ( n47511 , n47139 , n47509 );
or ( n47512 , n47142 , n47510 , n47511 );
and ( n47513 , n47016 , n47512 );
and ( n47514 , n47014 , n47512 );
or ( n47515 , n47017 , n47513 , n47514 );
and ( n47516 , n46893 , n47515 );
xor ( n47517 , n46893 , n47515 );
xor ( n47518 , n47014 , n47016 );
xor ( n47519 , n47518 , n47512 );
not ( n47520 , n47519 );
xor ( n47521 , n47139 , n47141 );
xor ( n47522 , n47521 , n47509 );
xnor ( n47523 , n47144 , n47508 );
xor ( n47524 , n47259 , n47261 );
xor ( n47525 , n47524 , n47505 );
xor ( n47526 , n47380 , n47382 );
xor ( n47527 , n47526 , n47502 );
xor ( n47528 , n47269 , n47328 );
xor ( n47529 , n47528 , n47374 );
xor ( n47530 , n47271 , n47275 );
xor ( n47531 , n47530 , n47325 );
xor ( n47532 , n47366 , n47368 );
xor ( n47533 , n47532 , n47371 );
and ( n47534 , n47531 , n47533 );
xor ( n47535 , n47292 , n47301 );
xor ( n47536 , n47535 , n47322 );
xor ( n47537 , n47345 , n47360 );
xor ( n47538 , n47537 , n47363 );
and ( n47539 , n47536 , n47538 );
xor ( n47540 , n47333 , n47337 );
xor ( n47541 , n47540 , n47342 );
xor ( n47542 , n47349 , n47352 );
xor ( n47543 , n47542 , n47357 );
and ( n47544 , n47541 , n47543 );
xor ( n47545 , n25160 , n45642 );
buf ( n47546 , n47545 );
buf ( n47547 , n47546 );
buf ( n47548 , n47547 );
xor ( n47549 , n47410 , n47414 );
and ( n47550 , n47548 , n47549 );
buf ( n47551 , n47550 );
and ( n47552 , n47543 , n47551 );
and ( n47553 , n47541 , n47551 );
or ( n47554 , n47544 , n47552 , n47553 );
and ( n47555 , n47538 , n47554 );
and ( n47556 , n47536 , n47554 );
or ( n47557 , n47539 , n47555 , n47556 );
and ( n47558 , n47533 , n47557 );
and ( n47559 , n47531 , n47557 );
or ( n47560 , n47534 , n47558 , n47559 );
and ( n47561 , n47529 , n47560 );
xor ( n47562 , n47387 , n47389 );
xor ( n47563 , n47562 , n47493 );
and ( n47564 , n47560 , n47563 );
and ( n47565 , n47529 , n47563 );
or ( n47566 , n47561 , n47564 , n47565 );
xor ( n47567 , n47385 , n47496 );
xor ( n47568 , n47567 , n47499 );
and ( n47569 , n47566 , n47568 );
xor ( n47570 , n47419 , n47423 );
and ( n47571 , n46345 , n46135 );
and ( n47572 , n46264 , n46133 );
nor ( n47573 , n47571 , n47572 );
xnor ( n47574 , n47573 , n46067 );
and ( n47575 , n46530 , n45990 );
and ( n47576 , n46445 , n45988 );
nor ( n47577 , n47575 , n47576 );
xnor ( n47578 , n47577 , n45939 );
and ( n47579 , n47574 , n47578 );
and ( n47580 , n47216 , n45702 );
and ( n47581 , n47090 , n45700 );
nor ( n47582 , n47580 , n47581 );
xnor ( n47583 , n47582 , n20841 );
and ( n47584 , n47578 , n47583 );
and ( n47585 , n47574 , n47583 );
or ( n47586 , n47579 , n47584 , n47585 );
and ( n47587 , n47570 , n47586 );
and ( n47588 , n46750 , n45886 );
and ( n47589 , n46577 , n45884 );
nor ( n47590 , n47588 , n47589 );
xnor ( n47591 , n47590 , n45824 );
and ( n47592 , n46969 , n45777 );
and ( n47593 , n46843 , n45775 );
nor ( n47594 , n47592 , n47593 );
xnor ( n47595 , n47594 , n45734 );
and ( n47596 , n47591 , n47595 );
and ( n47597 , n47586 , n47596 );
and ( n47598 , n47570 , n47596 );
or ( n47599 , n47587 , n47597 , n47598 );
buf ( n47600 , n17495 );
buf ( n47601 , n47600 );
buf ( n47602 , n17497 );
buf ( n47603 , n47602 );
and ( n47604 , n47601 , n47603 );
not ( n47605 , n47604 );
and ( n47606 , n47306 , n47605 );
not ( n47607 , n47606 );
and ( n47608 , n20844 , n47429 );
and ( n47609 , n20855 , n47427 );
nor ( n47610 , n47608 , n47609 );
xnor ( n47611 , n47610 , n47309 );
and ( n47612 , n47607 , n47611 );
and ( n47613 , n45712 , n47178 );
and ( n47614 , n20864 , n47176 );
nor ( n47615 , n47613 , n47614 );
xnor ( n47616 , n47615 , n47039 );
and ( n47617 , n47611 , n47616 );
and ( n47618 , n47607 , n47616 );
or ( n47619 , n47612 , n47617 , n47618 );
and ( n47620 , n45794 , n46911 );
and ( n47621 , n45763 , n46909 );
nor ( n47622 , n47620 , n47621 );
xnor ( n47623 , n47622 , n46802 );
and ( n47624 , n45907 , n46712 );
and ( n47625 , n45843 , n46710 );
nor ( n47626 , n47624 , n47625 );
xnor ( n47627 , n47626 , n46587 );
and ( n47628 , n47623 , n47627 );
and ( n47629 , n46041 , n46496 );
and ( n47630 , n45963 , n46494 );
nor ( n47631 , n47629 , n47630 );
xnor ( n47632 , n47631 , n46402 );
and ( n47633 , n47627 , n47632 );
and ( n47634 , n47623 , n47632 );
or ( n47635 , n47628 , n47633 , n47634 );
and ( n47636 , n47619 , n47635 );
and ( n47637 , n46169 , n46306 );
and ( n47638 , n46100 , n46304 );
nor ( n47639 , n47637 , n47638 );
xnor ( n47640 , n47639 , n46228 );
and ( n47641 , n47474 , n20852 );
and ( n47642 , n47351 , n20850 );
nor ( n47643 , n47641 , n47642 );
xnor ( n47644 , n47643 , n20860 );
and ( n47645 , n47640 , n47644 );
buf ( n47646 , n20738 );
buf ( n47647 , n47646 );
and ( n47648 , n47647 , n20846 );
and ( n47649 , n47644 , n47648 );
and ( n47650 , n47640 , n47648 );
or ( n47651 , n47645 , n47649 , n47650 );
and ( n47652 , n47635 , n47651 );
and ( n47653 , n47619 , n47651 );
or ( n47654 , n47636 , n47652 , n47653 );
and ( n47655 , n47599 , n47654 );
xor ( n47656 , n47432 , n47436 );
xor ( n47657 , n47656 , n47441 );
xor ( n47658 , n47451 , n47455 );
xor ( n47659 , n47658 , n47460 );
and ( n47660 , n47657 , n47659 );
xor ( n47661 , n47467 , n47471 );
xor ( n47662 , n47661 , n47475 );
and ( n47663 , n47659 , n47662 );
and ( n47664 , n47657 , n47662 );
or ( n47665 , n47660 , n47663 , n47664 );
and ( n47666 , n47654 , n47665 );
and ( n47667 , n47599 , n47665 );
or ( n47668 , n47655 , n47666 , n47667 );
buf ( n47669 , n47399 );
xor ( n47670 , n47669 , n47400 );
xor ( n47671 , n47415 , n47424 );
xor ( n47672 , n47671 , n47444 );
and ( n47673 , n47670 , n47672 );
xor ( n47674 , n47463 , n47478 );
xor ( n47675 , n47674 , n47481 );
and ( n47676 , n47672 , n47675 );
and ( n47677 , n47670 , n47675 );
or ( n47678 , n47673 , n47676 , n47677 );
and ( n47679 , n47668 , n47678 );
xor ( n47680 , n47394 , n47396 );
xor ( n47681 , n47680 , n47402 );
and ( n47682 , n47678 , n47681 );
and ( n47683 , n47668 , n47681 );
or ( n47684 , n47679 , n47682 , n47683 );
xor ( n47685 , n47392 , n47405 );
xor ( n47686 , n47685 , n47490 );
and ( n47687 , n47684 , n47686 );
xor ( n47688 , n47447 , n47484 );
xor ( n47689 , n47688 , n47487 );
xor ( n47690 , n25161 , n45641 );
buf ( n47691 , n47690 );
buf ( n47692 , n47691 );
buf ( n47693 , n47692 );
xor ( n47694 , n47574 , n47578 );
xor ( n47695 , n47694 , n47583 );
and ( n47696 , n47693 , n47695 );
buf ( n47697 , n47696 );
xor ( n47698 , n47591 , n47595 );
and ( n47699 , n46264 , n46306 );
and ( n47700 , n46169 , n46304 );
nor ( n47701 , n47699 , n47700 );
xnor ( n47702 , n47701 , n46228 );
and ( n47703 , n46843 , n45886 );
and ( n47704 , n46750 , n45884 );
nor ( n47705 , n47703 , n47704 );
xnor ( n47706 , n47705 , n45824 );
and ( n47707 , n47702 , n47706 );
and ( n47708 , n47090 , n45777 );
and ( n47709 , n46969 , n45775 );
nor ( n47710 , n47708 , n47709 );
xnor ( n47711 , n47710 , n45734 );
and ( n47712 , n47706 , n47711 );
and ( n47713 , n47702 , n47711 );
or ( n47714 , n47707 , n47712 , n47713 );
and ( n47715 , n47698 , n47714 );
and ( n47716 , n46445 , n46135 );
and ( n47717 , n46345 , n46133 );
nor ( n47718 , n47716 , n47717 );
xnor ( n47719 , n47718 , n46067 );
not ( n47720 , n47719 );
and ( n47721 , n46577 , n45990 );
and ( n47722 , n46530 , n45988 );
nor ( n47723 , n47721 , n47722 );
xnor ( n47724 , n47723 , n45939 );
and ( n47725 , n47720 , n47724 );
and ( n47726 , n47714 , n47725 );
and ( n47727 , n47698 , n47725 );
or ( n47728 , n47715 , n47726 , n47727 );
and ( n47729 , n47697 , n47728 );
buf ( n47730 , n47719 );
xor ( n47731 , n47306 , n47601 );
xor ( n47732 , n47601 , n47603 );
not ( n47733 , n47732 );
and ( n47734 , n47731 , n47733 );
and ( n47735 , n20855 , n47734 );
not ( n47736 , n47735 );
xnor ( n47737 , n47736 , n47606 );
and ( n47738 , n20864 , n47429 );
and ( n47739 , n20844 , n47427 );
nor ( n47740 , n47738 , n47739 );
xnor ( n47741 , n47740 , n47309 );
and ( n47742 , n47737 , n47741 );
and ( n47743 , n45763 , n47178 );
and ( n47744 , n45712 , n47176 );
nor ( n47745 , n47743 , n47744 );
xnor ( n47746 , n47745 , n47039 );
and ( n47747 , n47741 , n47746 );
and ( n47748 , n47737 , n47746 );
or ( n47749 , n47742 , n47747 , n47748 );
and ( n47750 , n47730 , n47749 );
and ( n47751 , n45843 , n46911 );
and ( n47752 , n45794 , n46909 );
nor ( n47753 , n47751 , n47752 );
xnor ( n47754 , n47753 , n46802 );
and ( n47755 , n45963 , n46712 );
and ( n47756 , n45907 , n46710 );
nor ( n47757 , n47755 , n47756 );
xnor ( n47758 , n47757 , n46587 );
and ( n47759 , n47754 , n47758 );
and ( n47760 , n46100 , n46496 );
and ( n47761 , n46041 , n46494 );
nor ( n47762 , n47760 , n47761 );
xnor ( n47763 , n47762 , n46402 );
and ( n47764 , n47758 , n47763 );
and ( n47765 , n47754 , n47763 );
or ( n47766 , n47759 , n47764 , n47765 );
and ( n47767 , n47749 , n47766 );
and ( n47768 , n47730 , n47766 );
or ( n47769 , n47750 , n47767 , n47768 );
and ( n47770 , n47728 , n47769 );
and ( n47771 , n47697 , n47769 );
or ( n47772 , n47729 , n47770 , n47771 );
and ( n47773 , n47351 , n45702 );
and ( n47774 , n47216 , n45700 );
nor ( n47775 , n47773 , n47774 );
xnor ( n47776 , n47775 , n20841 );
buf ( n47777 , n20740 );
buf ( n47778 , n47777 );
and ( n47779 , n47778 , n20846 );
and ( n47780 , n47776 , n47779 );
xor ( n47781 , n25162 , n45640 );
buf ( n47782 , n47781 );
buf ( n47783 , n47782 );
buf ( n47784 , n47783 );
and ( n47785 , n47779 , n47784 );
and ( n47786 , n47776 , n47784 );
or ( n47787 , n47780 , n47785 , n47786 );
xor ( n47788 , n47607 , n47611 );
xor ( n47789 , n47788 , n47616 );
and ( n47790 , n47787 , n47789 );
xor ( n47791 , n47623 , n47627 );
xor ( n47792 , n47791 , n47632 );
and ( n47793 , n47789 , n47792 );
and ( n47794 , n47787 , n47792 );
or ( n47795 , n47790 , n47793 , n47794 );
buf ( n47796 , n47548 );
xor ( n47797 , n47796 , n47549 );
and ( n47798 , n47795 , n47797 );
xor ( n47799 , n47570 , n47586 );
xor ( n47800 , n47799 , n47596 );
and ( n47801 , n47797 , n47800 );
and ( n47802 , n47795 , n47800 );
or ( n47803 , n47798 , n47801 , n47802 );
and ( n47804 , n47772 , n47803 );
xor ( n47805 , n47541 , n47543 );
xor ( n47806 , n47805 , n47551 );
and ( n47807 , n47803 , n47806 );
and ( n47808 , n47772 , n47806 );
or ( n47809 , n47804 , n47807 , n47808 );
and ( n47810 , n47689 , n47809 );
xor ( n47811 , n47536 , n47538 );
xor ( n47812 , n47811 , n47554 );
and ( n47813 , n47809 , n47812 );
and ( n47814 , n47689 , n47812 );
or ( n47815 , n47810 , n47813 , n47814 );
and ( n47816 , n47686 , n47815 );
and ( n47817 , n47684 , n47815 );
or ( n47818 , n47687 , n47816 , n47817 );
xor ( n47819 , n47529 , n47560 );
xor ( n47820 , n47819 , n47563 );
and ( n47821 , n47818 , n47820 );
xor ( n47822 , n47531 , n47533 );
xor ( n47823 , n47822 , n47557 );
xor ( n47824 , n47668 , n47678 );
xor ( n47825 , n47824 , n47681 );
xor ( n47826 , n47599 , n47654 );
xor ( n47827 , n47826 , n47665 );
xor ( n47828 , n47670 , n47672 );
xor ( n47829 , n47828 , n47675 );
and ( n47830 , n47827 , n47829 );
xor ( n47831 , n47619 , n47635 );
xor ( n47832 , n47831 , n47651 );
xor ( n47833 , n47657 , n47659 );
xor ( n47834 , n47833 , n47662 );
and ( n47835 , n47832 , n47834 );
xor ( n47836 , n47640 , n47644 );
xor ( n47837 , n47836 , n47648 );
and ( n47838 , n47647 , n20852 );
and ( n47839 , n47474 , n20850 );
nor ( n47840 , n47838 , n47839 );
xnor ( n47841 , n47840 , n20860 );
xor ( n47842 , n47720 , n47724 );
or ( n47843 , n47841 , n47842 );
and ( n47844 , n47837 , n47843 );
and ( n47845 , n46345 , n46306 );
and ( n47846 , n46264 , n46304 );
nor ( n47847 , n47845 , n47846 );
xnor ( n47848 , n47847 , n46228 );
and ( n47849 , n46530 , n46135 );
and ( n47850 , n46445 , n46133 );
nor ( n47851 , n47849 , n47850 );
xnor ( n47852 , n47851 , n46067 );
and ( n47853 , n47848 , n47852 );
and ( n47854 , n47216 , n45777 );
and ( n47855 , n47090 , n45775 );
nor ( n47856 , n47854 , n47855 );
xnor ( n47857 , n47856 , n45734 );
and ( n47858 , n47852 , n47857 );
and ( n47859 , n47848 , n47857 );
or ( n47860 , n47853 , n47858 , n47859 );
and ( n47861 , n46750 , n45990 );
and ( n47862 , n46577 , n45988 );
nor ( n47863 , n47861 , n47862 );
xnor ( n47864 , n47863 , n45939 );
and ( n47865 , n46969 , n45886 );
and ( n47866 , n46843 , n45884 );
nor ( n47867 , n47865 , n47866 );
xnor ( n47868 , n47867 , n45824 );
and ( n47869 , n47864 , n47868 );
and ( n47870 , n47474 , n45702 );
and ( n47871 , n47351 , n45700 );
nor ( n47872 , n47870 , n47871 );
xnor ( n47873 , n47872 , n20841 );
and ( n47874 , n47868 , n47873 );
and ( n47875 , n47864 , n47873 );
or ( n47876 , n47869 , n47874 , n47875 );
and ( n47877 , n47860 , n47876 );
buf ( n47878 , n47877 );
and ( n47879 , n47843 , n47878 );
and ( n47880 , n47837 , n47878 );
or ( n47881 , n47844 , n47879 , n47880 );
and ( n47882 , n47834 , n47881 );
and ( n47883 , n47832 , n47881 );
or ( n47884 , n47835 , n47882 , n47883 );
and ( n47885 , n47829 , n47884 );
and ( n47886 , n47827 , n47884 );
or ( n47887 , n47830 , n47885 , n47886 );
and ( n47888 , n47825 , n47887 );
xor ( n47889 , n47689 , n47809 );
xor ( n47890 , n47889 , n47812 );
and ( n47891 , n47887 , n47890 );
and ( n47892 , n47825 , n47890 );
or ( n47893 , n47888 , n47891 , n47892 );
and ( n47894 , n47823 , n47893 );
xor ( n47895 , n47684 , n47686 );
xor ( n47896 , n47895 , n47815 );
and ( n47897 , n47893 , n47896 );
and ( n47898 , n47823 , n47896 );
or ( n47899 , n47894 , n47897 , n47898 );
and ( n47900 , n47820 , n47899 );
and ( n47901 , n47818 , n47899 );
or ( n47902 , n47821 , n47900 , n47901 );
and ( n47903 , n47568 , n47902 );
and ( n47904 , n47566 , n47902 );
or ( n47905 , n47569 , n47903 , n47904 );
and ( n47906 , n47527 , n47905 );
xor ( n47907 , n47527 , n47905 );
xor ( n47908 , n47566 , n47568 );
xor ( n47909 , n47908 , n47902 );
not ( n47910 , n47909 );
xor ( n47911 , n47818 , n47820 );
xor ( n47912 , n47911 , n47899 );
xor ( n47913 , n47823 , n47893 );
xor ( n47914 , n47913 , n47896 );
buf ( n47915 , n17499 );
buf ( n47916 , n47915 );
buf ( n47917 , n17501 );
buf ( n47918 , n47917 );
and ( n47919 , n47916 , n47918 );
not ( n47920 , n47919 );
and ( n47921 , n47603 , n47920 );
not ( n47922 , n47921 );
and ( n47923 , n20844 , n47734 );
and ( n47924 , n20855 , n47732 );
nor ( n47925 , n47923 , n47924 );
xnor ( n47926 , n47925 , n47606 );
and ( n47927 , n47922 , n47926 );
and ( n47928 , n45712 , n47429 );
and ( n47929 , n20864 , n47427 );
nor ( n47930 , n47928 , n47929 );
xnor ( n47931 , n47930 , n47309 );
and ( n47932 , n47926 , n47931 );
and ( n47933 , n47922 , n47931 );
or ( n47934 , n47927 , n47932 , n47933 );
and ( n47935 , n45794 , n47178 );
and ( n47936 , n45763 , n47176 );
nor ( n47937 , n47935 , n47936 );
xnor ( n47938 , n47937 , n47039 );
and ( n47939 , n45907 , n46911 );
and ( n47940 , n45843 , n46909 );
nor ( n47941 , n47939 , n47940 );
xnor ( n47942 , n47941 , n46802 );
and ( n47943 , n47938 , n47942 );
and ( n47944 , n46041 , n46712 );
and ( n47945 , n45963 , n46710 );
nor ( n47946 , n47944 , n47945 );
xnor ( n47947 , n47946 , n46587 );
and ( n47948 , n47942 , n47947 );
and ( n47949 , n47938 , n47947 );
or ( n47950 , n47943 , n47948 , n47949 );
and ( n47951 , n47934 , n47950 );
and ( n47952 , n46169 , n46496 );
and ( n47953 , n46100 , n46494 );
nor ( n47954 , n47952 , n47953 );
xnor ( n47955 , n47954 , n46402 );
and ( n47956 , n47778 , n20852 );
and ( n47957 , n47647 , n20850 );
nor ( n47958 , n47956 , n47957 );
xnor ( n47959 , n47958 , n20860 );
and ( n47960 , n47955 , n47959 );
buf ( n47961 , n20742 );
buf ( n47962 , n47961 );
and ( n47963 , n47962 , n20846 );
and ( n47964 , n47959 , n47963 );
and ( n47965 , n47955 , n47963 );
or ( n47966 , n47960 , n47964 , n47965 );
and ( n47967 , n47950 , n47966 );
and ( n47968 , n47934 , n47966 );
or ( n47969 , n47951 , n47967 , n47968 );
xor ( n47970 , n47737 , n47741 );
xor ( n47971 , n47970 , n47746 );
xor ( n47972 , n47754 , n47758 );
xor ( n47973 , n47972 , n47763 );
and ( n47974 , n47971 , n47973 );
xor ( n47975 , n47776 , n47779 );
xor ( n47976 , n47975 , n47784 );
and ( n47977 , n47973 , n47976 );
and ( n47978 , n47971 , n47976 );
or ( n47979 , n47974 , n47977 , n47978 );
and ( n47980 , n47969 , n47979 );
buf ( n47981 , n47693 );
xor ( n47982 , n47981 , n47695 );
and ( n47983 , n47979 , n47982 );
and ( n47984 , n47969 , n47982 );
or ( n47985 , n47980 , n47983 , n47984 );
xor ( n47986 , n47698 , n47714 );
xor ( n47987 , n47986 , n47725 );
xor ( n47988 , n47730 , n47749 );
xor ( n47989 , n47988 , n47766 );
and ( n47990 , n47987 , n47989 );
xor ( n47991 , n47787 , n47789 );
xor ( n47992 , n47991 , n47792 );
and ( n47993 , n47989 , n47992 );
and ( n47994 , n47987 , n47992 );
or ( n47995 , n47990 , n47993 , n47994 );
and ( n47996 , n47985 , n47995 );
xor ( n47997 , n47697 , n47728 );
xor ( n47998 , n47997 , n47769 );
and ( n47999 , n47995 , n47998 );
and ( n48000 , n47985 , n47998 );
or ( n48001 , n47996 , n47999 , n48000 );
xor ( n48002 , n47772 , n47803 );
xor ( n48003 , n48002 , n47806 );
and ( n48004 , n48001 , n48003 );
xor ( n48005 , n47795 , n47797 );
xor ( n48006 , n48005 , n47800 );
xor ( n48007 , n47702 , n47706 );
xor ( n48008 , n48007 , n47711 );
xnor ( n48009 , n47841 , n47842 );
and ( n48010 , n48008 , n48009 );
xor ( n48011 , n47848 , n47852 );
xor ( n48012 , n48011 , n47857 );
xor ( n48013 , n47864 , n47868 );
xor ( n48014 , n48013 , n47873 );
or ( n48015 , n48012 , n48014 );
xor ( n48016 , n25163 , n45639 );
buf ( n48017 , n48016 );
buf ( n48018 , n48017 );
buf ( n48019 , n48018 );
and ( n48020 , n46445 , n46306 );
and ( n48021 , n46345 , n46304 );
nor ( n48022 , n48020 , n48021 );
xnor ( n48023 , n48022 , n46228 );
and ( n48024 , n46577 , n46135 );
and ( n48025 , n46530 , n46133 );
nor ( n48026 , n48024 , n48025 );
xnor ( n48027 , n48026 , n46067 );
and ( n48028 , n48023 , n48027 );
and ( n48029 , n47351 , n45777 );
and ( n48030 , n47216 , n45775 );
nor ( n48031 , n48029 , n48030 );
xnor ( n48032 , n48031 , n45734 );
and ( n48033 , n48027 , n48032 );
and ( n48034 , n48023 , n48032 );
or ( n48035 , n48028 , n48033 , n48034 );
and ( n48036 , n48019 , n48035 );
buf ( n48037 , n48036 );
and ( n48038 , n48015 , n48037 );
xor ( n48039 , n47603 , n47916 );
xor ( n48040 , n47916 , n47918 );
not ( n48041 , n48040 );
and ( n48042 , n48039 , n48041 );
and ( n48043 , n20855 , n48042 );
not ( n48044 , n48043 );
xnor ( n48045 , n48044 , n47921 );
and ( n48046 , n20864 , n47734 );
and ( n48047 , n20844 , n47732 );
nor ( n48048 , n48046 , n48047 );
xnor ( n48049 , n48048 , n47606 );
and ( n48050 , n48045 , n48049 );
and ( n48051 , n45763 , n47429 );
and ( n48052 , n45712 , n47427 );
nor ( n48053 , n48051 , n48052 );
xnor ( n48054 , n48053 , n47309 );
and ( n48055 , n48049 , n48054 );
and ( n48056 , n48045 , n48054 );
or ( n48057 , n48050 , n48055 , n48056 );
and ( n48058 , n45843 , n47178 );
and ( n48059 , n45794 , n47176 );
nor ( n48060 , n48058 , n48059 );
xnor ( n48061 , n48060 , n47039 );
and ( n48062 , n45963 , n46911 );
and ( n48063 , n45907 , n46909 );
nor ( n48064 , n48062 , n48063 );
xnor ( n48065 , n48064 , n46802 );
and ( n48066 , n48061 , n48065 );
and ( n48067 , n46100 , n46712 );
and ( n48068 , n46041 , n46710 );
nor ( n48069 , n48067 , n48068 );
xnor ( n48070 , n48069 , n46587 );
and ( n48071 , n48065 , n48070 );
and ( n48072 , n48061 , n48070 );
or ( n48073 , n48066 , n48071 , n48072 );
and ( n48074 , n48057 , n48073 );
and ( n48075 , n46264 , n46496 );
and ( n48076 , n46169 , n46494 );
nor ( n48077 , n48075 , n48076 );
xnor ( n48078 , n48077 , n46402 );
and ( n48079 , n46843 , n45990 );
and ( n48080 , n46750 , n45988 );
nor ( n48081 , n48079 , n48080 );
xnor ( n48082 , n48081 , n45939 );
and ( n48083 , n48078 , n48082 );
and ( n48084 , n47090 , n45886 );
and ( n48085 , n46969 , n45884 );
nor ( n48086 , n48084 , n48085 );
xnor ( n48087 , n48086 , n45824 );
and ( n48088 , n48082 , n48087 );
and ( n48089 , n48078 , n48087 );
or ( n48090 , n48083 , n48088 , n48089 );
and ( n48091 , n48073 , n48090 );
and ( n48092 , n48057 , n48090 );
or ( n48093 , n48074 , n48091 , n48092 );
and ( n48094 , n48037 , n48093 );
and ( n48095 , n48015 , n48093 );
or ( n48096 , n48038 , n48094 , n48095 );
and ( n48097 , n48010 , n48096 );
and ( n48098 , n47647 , n45702 );
and ( n48099 , n47474 , n45700 );
nor ( n48100 , n48098 , n48099 );
xnor ( n48101 , n48100 , n20841 );
and ( n48102 , n47962 , n20852 );
and ( n48103 , n47778 , n20850 );
nor ( n48104 , n48102 , n48103 );
xnor ( n48105 , n48104 , n20860 );
and ( n48106 , n48101 , n48105 );
buf ( n48107 , n20744 );
buf ( n48108 , n48107 );
and ( n48109 , n48108 , n20846 );
and ( n48110 , n48105 , n48109 );
and ( n48111 , n48101 , n48109 );
or ( n48112 , n48106 , n48110 , n48111 );
xor ( n48113 , n47922 , n47926 );
xor ( n48114 , n48113 , n47931 );
and ( n48115 , n48112 , n48114 );
xor ( n48116 , n47938 , n47942 );
xor ( n48117 , n48116 , n47947 );
and ( n48118 , n48114 , n48117 );
and ( n48119 , n48112 , n48117 );
or ( n48120 , n48115 , n48118 , n48119 );
buf ( n48121 , n47860 );
xor ( n48122 , n48121 , n47876 );
and ( n48123 , n48120 , n48122 );
xor ( n48124 , n47934 , n47950 );
xor ( n48125 , n48124 , n47966 );
and ( n48126 , n48122 , n48125 );
and ( n48127 , n48120 , n48125 );
or ( n48128 , n48123 , n48126 , n48127 );
and ( n48129 , n48096 , n48128 );
and ( n48130 , n48010 , n48128 );
or ( n48131 , n48097 , n48129 , n48130 );
and ( n48132 , n48006 , n48131 );
xor ( n48133 , n47837 , n47843 );
xor ( n48134 , n48133 , n47878 );
xor ( n48135 , n47969 , n47979 );
xor ( n48136 , n48135 , n47982 );
and ( n48137 , n48134 , n48136 );
xor ( n48138 , n47987 , n47989 );
xor ( n48139 , n48138 , n47992 );
and ( n48140 , n48136 , n48139 );
and ( n48141 , n48134 , n48139 );
or ( n48142 , n48137 , n48140 , n48141 );
and ( n48143 , n48131 , n48142 );
and ( n48144 , n48006 , n48142 );
or ( n48145 , n48132 , n48143 , n48144 );
and ( n48146 , n48003 , n48145 );
and ( n48147 , n48001 , n48145 );
or ( n48148 , n48004 , n48146 , n48147 );
xor ( n48149 , n47825 , n47887 );
xor ( n48150 , n48149 , n47890 );
and ( n48151 , n48148 , n48150 );
xor ( n48152 , n47827 , n47829 );
xor ( n48153 , n48152 , n47884 );
xor ( n48154 , n47832 , n47834 );
xor ( n48155 , n48154 , n47881 );
xor ( n48156 , n47985 , n47995 );
xor ( n48157 , n48156 , n47998 );
and ( n48158 , n48155 , n48157 );
xor ( n48159 , n47971 , n47973 );
xor ( n48160 , n48159 , n47976 );
xor ( n48161 , n48008 , n48009 );
and ( n48162 , n48160 , n48161 );
xor ( n48163 , n47955 , n47959 );
xor ( n48164 , n48163 , n47963 );
xnor ( n48165 , n48012 , n48014 );
and ( n48166 , n48164 , n48165 );
and ( n48167 , n46530 , n46306 );
and ( n48168 , n46445 , n46304 );
nor ( n48169 , n48167 , n48168 );
xnor ( n48170 , n48169 , n46228 );
and ( n48171 , n47474 , n45777 );
and ( n48172 , n47351 , n45775 );
nor ( n48173 , n48171 , n48172 );
xnor ( n48174 , n48173 , n45734 );
and ( n48175 , n48170 , n48174 );
and ( n48176 , n47778 , n45702 );
and ( n48177 , n47647 , n45700 );
nor ( n48178 , n48176 , n48177 );
xnor ( n48179 , n48178 , n20841 );
and ( n48180 , n48174 , n48179 );
and ( n48181 , n48170 , n48179 );
or ( n48182 , n48175 , n48180 , n48181 );
xor ( n48183 , n48023 , n48027 );
xor ( n48184 , n48183 , n48032 );
and ( n48185 , n48182 , n48184 );
and ( n48186 , n48165 , n48185 );
and ( n48187 , n48164 , n48185 );
or ( n48188 , n48166 , n48186 , n48187 );
and ( n48189 , n48161 , n48188 );
and ( n48190 , n48160 , n48188 );
or ( n48191 , n48162 , n48189 , n48190 );
xor ( n48192 , n25164 , n45638 );
buf ( n48193 , n48192 );
buf ( n48194 , n48193 );
buf ( n48195 , n48194 );
and ( n48196 , n46750 , n46135 );
and ( n48197 , n46577 , n46133 );
nor ( n48198 , n48196 , n48197 );
xnor ( n48199 , n48198 , n46067 );
and ( n48200 , n46969 , n45990 );
and ( n48201 , n46843 , n45988 );
nor ( n48202 , n48200 , n48201 );
xnor ( n48203 , n48202 , n45939 );
and ( n48204 , n48199 , n48203 );
and ( n48205 , n47216 , n45886 );
and ( n48206 , n47090 , n45884 );
nor ( n48207 , n48205 , n48206 );
xnor ( n48208 , n48207 , n45824 );
and ( n48209 , n48203 , n48208 );
and ( n48210 , n48199 , n48208 );
or ( n48211 , n48204 , n48209 , n48210 );
and ( n48212 , n48195 , n48211 );
buf ( n48213 , n48212 );
buf ( n48214 , n17503 );
buf ( n48215 , n48214 );
buf ( n48216 , n17505 );
buf ( n48217 , n48216 );
and ( n48218 , n48215 , n48217 );
not ( n48219 , n48218 );
and ( n48220 , n47918 , n48219 );
not ( n48221 , n48220 );
and ( n48222 , n20844 , n48042 );
and ( n48223 , n20855 , n48040 );
nor ( n48224 , n48222 , n48223 );
xnor ( n48225 , n48224 , n47921 );
and ( n48226 , n48221 , n48225 );
and ( n48227 , n45712 , n47734 );
and ( n48228 , n20864 , n47732 );
nor ( n48229 , n48227 , n48228 );
xnor ( n48230 , n48229 , n47606 );
and ( n48231 , n48225 , n48230 );
and ( n48232 , n48221 , n48230 );
or ( n48233 , n48226 , n48231 , n48232 );
and ( n48234 , n45794 , n47429 );
and ( n48235 , n45763 , n47427 );
nor ( n48236 , n48234 , n48235 );
xnor ( n48237 , n48236 , n47309 );
and ( n48238 , n45907 , n47178 );
and ( n48239 , n45843 , n47176 );
nor ( n48240 , n48238 , n48239 );
xnor ( n48241 , n48240 , n47039 );
and ( n48242 , n48237 , n48241 );
and ( n48243 , n46041 , n46911 );
and ( n48244 , n45963 , n46909 );
nor ( n48245 , n48243 , n48244 );
xnor ( n48246 , n48245 , n46802 );
and ( n48247 , n48241 , n48246 );
and ( n48248 , n48237 , n48246 );
or ( n48249 , n48242 , n48247 , n48248 );
and ( n48250 , n48233 , n48249 );
and ( n48251 , n46169 , n46712 );
and ( n48252 , n46100 , n46710 );
nor ( n48253 , n48251 , n48252 );
xnor ( n48254 , n48253 , n46587 );
and ( n48255 , n46345 , n46496 );
and ( n48256 , n46264 , n46494 );
nor ( n48257 , n48255 , n48256 );
xnor ( n48258 , n48257 , n46402 );
and ( n48259 , n48254 , n48258 );
and ( n48260 , n48108 , n20852 );
and ( n48261 , n47962 , n20850 );
nor ( n48262 , n48260 , n48261 );
xnor ( n48263 , n48262 , n20860 );
and ( n48264 , n48258 , n48263 );
and ( n48265 , n48254 , n48263 );
or ( n48266 , n48259 , n48264 , n48265 );
and ( n48267 , n48249 , n48266 );
and ( n48268 , n48233 , n48266 );
or ( n48269 , n48250 , n48267 , n48268 );
and ( n48270 , n48213 , n48269 );
buf ( n48271 , n20746 );
buf ( n48272 , n48271 );
and ( n48273 , n48272 , n20846 );
xor ( n48274 , n25165 , n45637 );
buf ( n48275 , n48274 );
buf ( n48276 , n48275 );
buf ( n48277 , n48276 );
and ( n48278 , n48273 , n48277 );
buf ( n48279 , n48278 );
xor ( n48280 , n48045 , n48049 );
xor ( n48281 , n48280 , n48054 );
and ( n48282 , n48279 , n48281 );
xor ( n48283 , n48061 , n48065 );
xor ( n48284 , n48283 , n48070 );
and ( n48285 , n48281 , n48284 );
and ( n48286 , n48279 , n48284 );
or ( n48287 , n48282 , n48285 , n48286 );
and ( n48288 , n48269 , n48287 );
and ( n48289 , n48213 , n48287 );
or ( n48290 , n48270 , n48288 , n48289 );
buf ( n48291 , n48019 );
xor ( n48292 , n48291 , n48035 );
xor ( n48293 , n48057 , n48073 );
xor ( n48294 , n48293 , n48090 );
and ( n48295 , n48292 , n48294 );
xor ( n48296 , n48112 , n48114 );
xor ( n48297 , n48296 , n48117 );
and ( n48298 , n48294 , n48297 );
and ( n48299 , n48292 , n48297 );
or ( n48300 , n48295 , n48298 , n48299 );
and ( n48301 , n48290 , n48300 );
xor ( n48302 , n48015 , n48037 );
xor ( n48303 , n48302 , n48093 );
and ( n48304 , n48300 , n48303 );
and ( n48305 , n48290 , n48303 );
or ( n48306 , n48301 , n48304 , n48305 );
and ( n48307 , n48191 , n48306 );
xor ( n48308 , n48010 , n48096 );
xor ( n48309 , n48308 , n48128 );
and ( n48310 , n48306 , n48309 );
and ( n48311 , n48191 , n48309 );
or ( n48312 , n48307 , n48310 , n48311 );
and ( n48313 , n48157 , n48312 );
and ( n48314 , n48155 , n48312 );
or ( n48315 , n48158 , n48313 , n48314 );
and ( n48316 , n48153 , n48315 );
xor ( n48317 , n48001 , n48003 );
xor ( n48318 , n48317 , n48145 );
and ( n48319 , n48315 , n48318 );
and ( n48320 , n48153 , n48318 );
or ( n48321 , n48316 , n48319 , n48320 );
and ( n48322 , n48150 , n48321 );
and ( n48323 , n48148 , n48321 );
or ( n48324 , n48151 , n48322 , n48323 );
and ( n48325 , n47914 , n48324 );
xor ( n48326 , n48006 , n48131 );
xor ( n48327 , n48326 , n48142 );
xor ( n48328 , n48134 , n48136 );
xor ( n48329 , n48328 , n48139 );
xor ( n48330 , n48120 , n48122 );
xor ( n48331 , n48330 , n48125 );
xor ( n48332 , n48078 , n48082 );
xor ( n48333 , n48332 , n48087 );
xor ( n48334 , n48101 , n48105 );
xor ( n48335 , n48334 , n48109 );
and ( n48336 , n48333 , n48335 );
xor ( n48337 , n48182 , n48184 );
and ( n48338 , n48335 , n48337 );
and ( n48339 , n48333 , n48337 );
or ( n48340 , n48336 , n48338 , n48339 );
and ( n48341 , n46843 , n46135 );
and ( n48342 , n46750 , n46133 );
nor ( n48343 , n48341 , n48342 );
xnor ( n48344 , n48343 , n46067 );
and ( n48345 , n47090 , n45990 );
and ( n48346 , n46969 , n45988 );
nor ( n48347 , n48345 , n48346 );
xnor ( n48348 , n48347 , n45939 );
and ( n48349 , n48344 , n48348 );
and ( n48350 , n48272 , n20852 );
and ( n48351 , n48108 , n20850 );
nor ( n48352 , n48350 , n48351 );
xnor ( n48353 , n48352 , n20860 );
and ( n48354 , n48348 , n48353 );
and ( n48355 , n48344 , n48353 );
or ( n48356 , n48349 , n48354 , n48355 );
and ( n48357 , n46577 , n46306 );
and ( n48358 , n46530 , n46304 );
nor ( n48359 , n48357 , n48358 );
xnor ( n48360 , n48359 , n46228 );
and ( n48361 , n47351 , n45886 );
and ( n48362 , n47216 , n45884 );
nor ( n48363 , n48361 , n48362 );
xnor ( n48364 , n48363 , n45824 );
and ( n48365 , n48360 , n48364 );
and ( n48366 , n47647 , n45777 );
and ( n48367 , n47474 , n45775 );
nor ( n48368 , n48366 , n48367 );
xnor ( n48369 , n48368 , n45734 );
and ( n48370 , n48364 , n48369 );
and ( n48371 , n48360 , n48369 );
or ( n48372 , n48365 , n48370 , n48371 );
or ( n48373 , n48356 , n48372 );
xor ( n48374 , n48170 , n48174 );
xor ( n48375 , n48374 , n48179 );
xor ( n48376 , n48199 , n48203 );
xor ( n48377 , n48376 , n48208 );
and ( n48378 , n48375 , n48377 );
and ( n48379 , n46264 , n46712 );
and ( n48380 , n46169 , n46710 );
nor ( n48381 , n48379 , n48380 );
xnor ( n48382 , n48381 , n46587 );
buf ( n48383 , n20748 );
buf ( n48384 , n48383 );
and ( n48385 , n48384 , n20846 );
or ( n48386 , n48382 , n48385 );
and ( n48387 , n48377 , n48386 );
and ( n48388 , n48375 , n48386 );
or ( n48389 , n48378 , n48387 , n48388 );
and ( n48390 , n48373 , n48389 );
xor ( n48391 , n47918 , n48215 );
xor ( n48392 , n48215 , n48217 );
not ( n48393 , n48392 );
and ( n48394 , n48391 , n48393 );
and ( n48395 , n20855 , n48394 );
not ( n48396 , n48395 );
xnor ( n48397 , n48396 , n48220 );
and ( n48398 , n20864 , n48042 );
and ( n48399 , n20844 , n48040 );
nor ( n48400 , n48398 , n48399 );
xnor ( n48401 , n48400 , n47921 );
and ( n48402 , n48397 , n48401 );
and ( n48403 , n45763 , n47734 );
and ( n48404 , n45712 , n47732 );
nor ( n48405 , n48403 , n48404 );
xnor ( n48406 , n48405 , n47606 );
and ( n48407 , n48401 , n48406 );
and ( n48408 , n48397 , n48406 );
or ( n48409 , n48402 , n48407 , n48408 );
and ( n48410 , n45843 , n47429 );
and ( n48411 , n45794 , n47427 );
nor ( n48412 , n48410 , n48411 );
xnor ( n48413 , n48412 , n47309 );
and ( n48414 , n45963 , n47178 );
and ( n48415 , n45907 , n47176 );
nor ( n48416 , n48414 , n48415 );
xnor ( n48417 , n48416 , n47039 );
and ( n48418 , n48413 , n48417 );
and ( n48419 , n46100 , n46911 );
and ( n48420 , n46041 , n46909 );
nor ( n48421 , n48419 , n48420 );
xnor ( n48422 , n48421 , n46802 );
and ( n48423 , n48417 , n48422 );
and ( n48424 , n48413 , n48422 );
or ( n48425 , n48418 , n48423 , n48424 );
and ( n48426 , n48409 , n48425 );
and ( n48427 , n46445 , n46496 );
and ( n48428 , n46345 , n46494 );
nor ( n48429 , n48427 , n48428 );
xnor ( n48430 , n48429 , n46402 );
and ( n48431 , n47962 , n45702 );
and ( n48432 , n47778 , n45700 );
nor ( n48433 , n48431 , n48432 );
xnor ( n48434 , n48433 , n20841 );
and ( n48435 , n48430 , n48434 );
xor ( n48436 , n25166 , n45636 );
buf ( n48437 , n48436 );
buf ( n48438 , n48437 );
buf ( n48439 , n48438 );
and ( n48440 , n48434 , n48439 );
and ( n48441 , n48430 , n48439 );
or ( n48442 , n48435 , n48440 , n48441 );
and ( n48443 , n48425 , n48442 );
and ( n48444 , n48409 , n48442 );
or ( n48445 , n48426 , n48443 , n48444 );
and ( n48446 , n48389 , n48445 );
and ( n48447 , n48373 , n48445 );
or ( n48448 , n48390 , n48446 , n48447 );
and ( n48449 , n48340 , n48448 );
xor ( n48450 , n48221 , n48225 );
xor ( n48451 , n48450 , n48230 );
xor ( n48452 , n48237 , n48241 );
xor ( n48453 , n48452 , n48246 );
and ( n48454 , n48451 , n48453 );
xor ( n48455 , n48254 , n48258 );
xor ( n48456 , n48455 , n48263 );
and ( n48457 , n48453 , n48456 );
and ( n48458 , n48451 , n48456 );
or ( n48459 , n48454 , n48457 , n48458 );
buf ( n48460 , n48195 );
xor ( n48461 , n48460 , n48211 );
and ( n48462 , n48459 , n48461 );
xor ( n48463 , n48233 , n48249 );
xor ( n48464 , n48463 , n48266 );
and ( n48465 , n48461 , n48464 );
and ( n48466 , n48459 , n48464 );
or ( n48467 , n48462 , n48465 , n48466 );
and ( n48468 , n48448 , n48467 );
and ( n48469 , n48340 , n48467 );
or ( n48470 , n48449 , n48468 , n48469 );
and ( n48471 , n48331 , n48470 );
xor ( n48472 , n48164 , n48165 );
xor ( n48473 , n48472 , n48185 );
xor ( n48474 , n48213 , n48269 );
xor ( n48475 , n48474 , n48287 );
and ( n48476 , n48473 , n48475 );
xor ( n48477 , n48292 , n48294 );
xor ( n48478 , n48477 , n48297 );
and ( n48479 , n48475 , n48478 );
and ( n48480 , n48473 , n48478 );
or ( n48481 , n48476 , n48479 , n48480 );
and ( n48482 , n48470 , n48481 );
and ( n48483 , n48331 , n48481 );
or ( n48484 , n48471 , n48482 , n48483 );
and ( n48485 , n48329 , n48484 );
xor ( n48486 , n48191 , n48306 );
xor ( n48487 , n48486 , n48309 );
and ( n48488 , n48484 , n48487 );
and ( n48489 , n48329 , n48487 );
or ( n48490 , n48485 , n48488 , n48489 );
and ( n48491 , n48327 , n48490 );
xor ( n48492 , n48155 , n48157 );
xor ( n48493 , n48492 , n48312 );
and ( n48494 , n48490 , n48493 );
and ( n48495 , n48327 , n48493 );
or ( n48496 , n48491 , n48494 , n48495 );
xor ( n48497 , n48153 , n48315 );
xor ( n48498 , n48497 , n48318 );
or ( n48499 , n48496 , n48498 );
xor ( n48500 , n48148 , n48150 );
xor ( n48501 , n48500 , n48321 );
or ( n48502 , n48499 , n48501 );
and ( n48503 , n48324 , n48502 );
and ( n48504 , n47914 , n48502 );
or ( n48505 , n48325 , n48503 , n48504 );
and ( n48506 , n47912 , n48505 );
xor ( n48507 , n47912 , n48505 );
xor ( n48508 , n47914 , n48324 );
xor ( n48509 , n48508 , n48502 );
xnor ( n48510 , n48499 , n48501 );
xnor ( n48511 , n48496 , n48498 );
xor ( n48512 , n48327 , n48490 );
xor ( n48513 , n48512 , n48493 );
xor ( n48514 , n48160 , n48161 );
xor ( n48515 , n48514 , n48188 );
xor ( n48516 , n48290 , n48300 );
xor ( n48517 , n48516 , n48303 );
and ( n48518 , n48515 , n48517 );
xor ( n48519 , n48279 , n48281 );
xor ( n48520 , n48519 , n48284 );
xor ( n48521 , n48273 , n48277 );
buf ( n48522 , n48521 );
xnor ( n48523 , n48356 , n48372 );
and ( n48524 , n48522 , n48523 );
xor ( n48525 , n48344 , n48348 );
xor ( n48526 , n48525 , n48353 );
xor ( n48527 , n48360 , n48364 );
xor ( n48528 , n48527 , n48369 );
and ( n48529 , n48526 , n48528 );
buf ( n48530 , n48529 );
and ( n48531 , n48523 , n48530 );
and ( n48532 , n48522 , n48530 );
or ( n48533 , n48524 , n48531 , n48532 );
and ( n48534 , n48520 , n48533 );
xnor ( n48535 , n48382 , n48385 );
and ( n48536 , n47216 , n45990 );
and ( n48537 , n47090 , n45988 );
nor ( n48538 , n48536 , n48537 );
xnor ( n48539 , n48538 , n45939 );
and ( n48540 , n48108 , n45702 );
and ( n48541 , n47962 , n45700 );
nor ( n48542 , n48540 , n48541 );
xnor ( n48543 , n48542 , n20841 );
and ( n48544 , n48539 , n48543 );
and ( n48545 , n48384 , n20852 );
and ( n48546 , n48272 , n20850 );
nor ( n48547 , n48545 , n48546 );
xnor ( n48548 , n48547 , n20860 );
and ( n48549 , n48543 , n48548 );
and ( n48550 , n48539 , n48548 );
or ( n48551 , n48544 , n48549 , n48550 );
and ( n48552 , n48535 , n48551 );
and ( n48553 , n47474 , n45886 );
and ( n48554 , n47351 , n45884 );
nor ( n48555 , n48553 , n48554 );
xnor ( n48556 , n48555 , n45824 );
and ( n48557 , n47778 , n45777 );
and ( n48558 , n47647 , n45775 );
nor ( n48559 , n48557 , n48558 );
xnor ( n48560 , n48559 , n45734 );
or ( n48561 , n48556 , n48560 );
and ( n48562 , n48551 , n48561 );
and ( n48563 , n48535 , n48561 );
or ( n48564 , n48552 , n48562 , n48563 );
buf ( n48565 , n17507 );
buf ( n48566 , n48565 );
buf ( n48567 , n17509 );
buf ( n48568 , n48567 );
and ( n48569 , n48566 , n48568 );
not ( n48570 , n48569 );
and ( n48571 , n48217 , n48570 );
not ( n48572 , n48571 );
and ( n48573 , n20844 , n48394 );
and ( n48574 , n20855 , n48392 );
nor ( n48575 , n48573 , n48574 );
xnor ( n48576 , n48575 , n48220 );
and ( n48577 , n48572 , n48576 );
and ( n48578 , n45712 , n48042 );
and ( n48579 , n20864 , n48040 );
nor ( n48580 , n48578 , n48579 );
xnor ( n48581 , n48580 , n47921 );
and ( n48582 , n48576 , n48581 );
and ( n48583 , n48572 , n48581 );
or ( n48584 , n48577 , n48582 , n48583 );
and ( n48585 , n45794 , n47734 );
and ( n48586 , n45763 , n47732 );
nor ( n48587 , n48585 , n48586 );
xnor ( n48588 , n48587 , n47606 );
and ( n48589 , n45907 , n47429 );
and ( n48590 , n45843 , n47427 );
nor ( n48591 , n48589 , n48590 );
xnor ( n48592 , n48591 , n47309 );
and ( n48593 , n48588 , n48592 );
and ( n48594 , n46041 , n47178 );
and ( n48595 , n45963 , n47176 );
nor ( n48596 , n48594 , n48595 );
xnor ( n48597 , n48596 , n47039 );
and ( n48598 , n48592 , n48597 );
and ( n48599 , n48588 , n48597 );
or ( n48600 , n48593 , n48598 , n48599 );
and ( n48601 , n48584 , n48600 );
and ( n48602 , n46169 , n46911 );
and ( n48603 , n46100 , n46909 );
nor ( n48604 , n48602 , n48603 );
xnor ( n48605 , n48604 , n46802 );
and ( n48606 , n46345 , n46712 );
and ( n48607 , n46264 , n46710 );
nor ( n48608 , n48606 , n48607 );
xnor ( n48609 , n48608 , n46587 );
and ( n48610 , n48605 , n48609 );
and ( n48611 , n46530 , n46496 );
and ( n48612 , n46445 , n46494 );
nor ( n48613 , n48611 , n48612 );
xnor ( n48614 , n48613 , n46402 );
and ( n48615 , n48609 , n48614 );
and ( n48616 , n48605 , n48614 );
or ( n48617 , n48610 , n48615 , n48616 );
and ( n48618 , n48600 , n48617 );
and ( n48619 , n48584 , n48617 );
or ( n48620 , n48601 , n48618 , n48619 );
and ( n48621 , n48564 , n48620 );
and ( n48622 , n46750 , n46306 );
and ( n48623 , n46577 , n46304 );
nor ( n48624 , n48622 , n48623 );
xnor ( n48625 , n48624 , n46228 );
and ( n48626 , n46969 , n46135 );
and ( n48627 , n46843 , n46133 );
nor ( n48628 , n48626 , n48627 );
xnor ( n48629 , n48628 , n46067 );
and ( n48630 , n48625 , n48629 );
buf ( n48631 , n20750 );
buf ( n48632 , n48631 );
and ( n48633 , n48632 , n20846 );
and ( n48634 , n48629 , n48633 );
and ( n48635 , n48625 , n48633 );
or ( n48636 , n48630 , n48634 , n48635 );
xor ( n48637 , n48397 , n48401 );
xor ( n48638 , n48637 , n48406 );
and ( n48639 , n48636 , n48638 );
xor ( n48640 , n48413 , n48417 );
xor ( n48641 , n48640 , n48422 );
and ( n48642 , n48638 , n48641 );
and ( n48643 , n48636 , n48641 );
or ( n48644 , n48639 , n48642 , n48643 );
and ( n48645 , n48620 , n48644 );
and ( n48646 , n48564 , n48644 );
or ( n48647 , n48621 , n48645 , n48646 );
and ( n48648 , n48533 , n48647 );
and ( n48649 , n48520 , n48647 );
or ( n48650 , n48534 , n48648 , n48649 );
xor ( n48651 , n48375 , n48377 );
xor ( n48652 , n48651 , n48386 );
xor ( n48653 , n48409 , n48425 );
xor ( n48654 , n48653 , n48442 );
and ( n48655 , n48652 , n48654 );
xor ( n48656 , n48451 , n48453 );
xor ( n48657 , n48656 , n48456 );
and ( n48658 , n48654 , n48657 );
and ( n48659 , n48652 , n48657 );
or ( n48660 , n48655 , n48658 , n48659 );
xor ( n48661 , n48333 , n48335 );
xor ( n48662 , n48661 , n48337 );
and ( n48663 , n48660 , n48662 );
xor ( n48664 , n48373 , n48389 );
xor ( n48665 , n48664 , n48445 );
and ( n48666 , n48662 , n48665 );
and ( n48667 , n48660 , n48665 );
or ( n48668 , n48663 , n48666 , n48667 );
and ( n48669 , n48650 , n48668 );
xor ( n48670 , n48340 , n48448 );
xor ( n48671 , n48670 , n48467 );
and ( n48672 , n48668 , n48671 );
and ( n48673 , n48650 , n48671 );
or ( n48674 , n48669 , n48672 , n48673 );
and ( n48675 , n48517 , n48674 );
and ( n48676 , n48515 , n48674 );
or ( n48677 , n48518 , n48675 , n48676 );
xor ( n48678 , n48329 , n48484 );
xor ( n48679 , n48678 , n48487 );
and ( n48680 , n48677 , n48679 );
xor ( n48681 , n48331 , n48470 );
xor ( n48682 , n48681 , n48481 );
xor ( n48683 , n48473 , n48475 );
xor ( n48684 , n48683 , n48478 );
xor ( n48685 , n48459 , n48461 );
xor ( n48686 , n48685 , n48464 );
xor ( n48687 , n48430 , n48434 );
xor ( n48688 , n48687 , n48439 );
xor ( n48689 , n25167 , n45635 );
buf ( n48690 , n48689 );
buf ( n48691 , n48690 );
buf ( n48692 , n48691 );
xor ( n48693 , n48539 , n48543 );
xor ( n48694 , n48693 , n48548 );
and ( n48695 , n48692 , n48694 );
buf ( n48696 , n48695 );
and ( n48697 , n48688 , n48696 );
xnor ( n48698 , n48556 , n48560 );
and ( n48699 , n46264 , n46911 );
and ( n48700 , n46169 , n46909 );
nor ( n48701 , n48699 , n48700 );
xnor ( n48702 , n48701 , n46802 );
and ( n48703 , n46445 , n46712 );
and ( n48704 , n46345 , n46710 );
nor ( n48705 , n48703 , n48704 );
xnor ( n48706 , n48705 , n46587 );
and ( n48707 , n48702 , n48706 );
buf ( n48708 , n20752 );
buf ( n48709 , n48708 );
and ( n48710 , n48709 , n20846 );
and ( n48711 , n48706 , n48710 );
and ( n48712 , n48702 , n48710 );
or ( n48713 , n48707 , n48711 , n48712 );
and ( n48714 , n48698 , n48713 );
and ( n48715 , n47647 , n45886 );
and ( n48716 , n47474 , n45884 );
nor ( n48717 , n48715 , n48716 );
xnor ( n48718 , n48717 , n45824 );
and ( n48719 , n48272 , n45702 );
and ( n48720 , n48108 , n45700 );
nor ( n48721 , n48719 , n48720 );
xnor ( n48722 , n48721 , n20841 );
and ( n48723 , n48718 , n48722 );
and ( n48724 , n48632 , n20852 );
and ( n48725 , n48384 , n20850 );
nor ( n48726 , n48724 , n48725 );
xnor ( n48727 , n48726 , n20860 );
and ( n48728 , n48722 , n48727 );
and ( n48729 , n48718 , n48727 );
or ( n48730 , n48723 , n48728 , n48729 );
and ( n48731 , n48713 , n48730 );
and ( n48732 , n48698 , n48730 );
or ( n48733 , n48714 , n48731 , n48732 );
and ( n48734 , n48696 , n48733 );
and ( n48735 , n48688 , n48733 );
or ( n48736 , n48697 , n48734 , n48735 );
xor ( n48737 , n48217 , n48566 );
xor ( n48738 , n48566 , n48568 );
not ( n48739 , n48738 );
and ( n48740 , n48737 , n48739 );
and ( n48741 , n20855 , n48740 );
not ( n48742 , n48741 );
xnor ( n48743 , n48742 , n48571 );
and ( n48744 , n20864 , n48394 );
and ( n48745 , n20844 , n48392 );
nor ( n48746 , n48744 , n48745 );
xnor ( n48747 , n48746 , n48220 );
and ( n48748 , n48743 , n48747 );
and ( n48749 , n45763 , n48042 );
and ( n48750 , n45712 , n48040 );
nor ( n48751 , n48749 , n48750 );
xnor ( n48752 , n48751 , n47921 );
and ( n48753 , n48747 , n48752 );
and ( n48754 , n48743 , n48752 );
or ( n48755 , n48748 , n48753 , n48754 );
and ( n48756 , n45843 , n47734 );
and ( n48757 , n45794 , n47732 );
nor ( n48758 , n48756 , n48757 );
xnor ( n48759 , n48758 , n47606 );
and ( n48760 , n45963 , n47429 );
and ( n48761 , n45907 , n47427 );
nor ( n48762 , n48760 , n48761 );
xnor ( n48763 , n48762 , n47309 );
and ( n48764 , n48759 , n48763 );
and ( n48765 , n46100 , n47178 );
and ( n48766 , n46041 , n47176 );
nor ( n48767 , n48765 , n48766 );
xnor ( n48768 , n48767 , n47039 );
and ( n48769 , n48763 , n48768 );
and ( n48770 , n48759 , n48768 );
or ( n48771 , n48764 , n48769 , n48770 );
and ( n48772 , n48755 , n48771 );
and ( n48773 , n46577 , n46496 );
and ( n48774 , n46530 , n46494 );
nor ( n48775 , n48773 , n48774 );
xnor ( n48776 , n48775 , n46402 );
and ( n48777 , n46843 , n46306 );
and ( n48778 , n46750 , n46304 );
nor ( n48779 , n48777 , n48778 );
xnor ( n48780 , n48779 , n46228 );
and ( n48781 , n48776 , n48780 );
and ( n48782 , n47090 , n46135 );
and ( n48783 , n46969 , n46133 );
nor ( n48784 , n48782 , n48783 );
xnor ( n48785 , n48784 , n46067 );
and ( n48786 , n48780 , n48785 );
and ( n48787 , n48776 , n48785 );
or ( n48788 , n48781 , n48786 , n48787 );
and ( n48789 , n48771 , n48788 );
and ( n48790 , n48755 , n48788 );
or ( n48791 , n48772 , n48789 , n48790 );
and ( n48792 , n47351 , n45990 );
and ( n48793 , n47216 , n45988 );
nor ( n48794 , n48792 , n48793 );
xnor ( n48795 , n48794 , n45939 );
and ( n48796 , n47962 , n45777 );
and ( n48797 , n47778 , n45775 );
nor ( n48798 , n48796 , n48797 );
xnor ( n48799 , n48798 , n45734 );
and ( n48800 , n48795 , n48799 );
xor ( n48801 , n25168 , n45634 );
buf ( n48802 , n48801 );
buf ( n48803 , n48802 );
buf ( n48804 , n48803 );
and ( n48805 , n48799 , n48804 );
and ( n48806 , n48795 , n48804 );
or ( n48807 , n48800 , n48805 , n48806 );
xor ( n48808 , n48572 , n48576 );
xor ( n48809 , n48808 , n48581 );
and ( n48810 , n48807 , n48809 );
xor ( n48811 , n48588 , n48592 );
xor ( n48812 , n48811 , n48597 );
and ( n48813 , n48809 , n48812 );
and ( n48814 , n48807 , n48812 );
or ( n48815 , n48810 , n48813 , n48814 );
and ( n48816 , n48791 , n48815 );
buf ( n48817 , n48526 );
xor ( n48818 , n48817 , n48528 );
and ( n48819 , n48815 , n48818 );
and ( n48820 , n48791 , n48818 );
or ( n48821 , n48816 , n48819 , n48820 );
and ( n48822 , n48736 , n48821 );
xor ( n48823 , n48535 , n48551 );
xor ( n48824 , n48823 , n48561 );
xor ( n48825 , n48584 , n48600 );
xor ( n48826 , n48825 , n48617 );
and ( n48827 , n48824 , n48826 );
xor ( n48828 , n48636 , n48638 );
xor ( n48829 , n48828 , n48641 );
and ( n48830 , n48826 , n48829 );
and ( n48831 , n48824 , n48829 );
or ( n48832 , n48827 , n48830 , n48831 );
and ( n48833 , n48821 , n48832 );
and ( n48834 , n48736 , n48832 );
or ( n48835 , n48822 , n48833 , n48834 );
and ( n48836 , n48686 , n48835 );
xor ( n48837 , n48522 , n48523 );
xor ( n48838 , n48837 , n48530 );
xor ( n48839 , n48564 , n48620 );
xor ( n48840 , n48839 , n48644 );
and ( n48841 , n48838 , n48840 );
xor ( n48842 , n48652 , n48654 );
xor ( n48843 , n48842 , n48657 );
and ( n48844 , n48840 , n48843 );
and ( n48845 , n48838 , n48843 );
or ( n48846 , n48841 , n48844 , n48845 );
and ( n48847 , n48835 , n48846 );
and ( n48848 , n48686 , n48846 );
or ( n48849 , n48836 , n48847 , n48848 );
and ( n48850 , n48684 , n48849 );
xor ( n48851 , n48650 , n48668 );
xor ( n48852 , n48851 , n48671 );
and ( n48853 , n48849 , n48852 );
and ( n48854 , n48684 , n48852 );
or ( n48855 , n48850 , n48853 , n48854 );
and ( n48856 , n48682 , n48855 );
xor ( n48857 , n48515 , n48517 );
xor ( n48858 , n48857 , n48674 );
and ( n48859 , n48855 , n48858 );
and ( n48860 , n48682 , n48858 );
or ( n48861 , n48856 , n48859 , n48860 );
and ( n48862 , n48679 , n48861 );
and ( n48863 , n48677 , n48861 );
or ( n48864 , n48680 , n48862 , n48863 );
and ( n48865 , n48513 , n48864 );
xor ( n48866 , n48513 , n48864 );
xor ( n48867 , n48677 , n48679 );
xor ( n48868 , n48867 , n48861 );
not ( n48869 , n48868 );
xor ( n48870 , n48682 , n48855 );
xor ( n48871 , n48870 , n48858 );
xor ( n48872 , n48520 , n48533 );
xor ( n48873 , n48872 , n48647 );
xor ( n48874 , n48660 , n48662 );
xor ( n48875 , n48874 , n48665 );
and ( n48876 , n48873 , n48875 );
xor ( n48877 , n48605 , n48609 );
xor ( n48878 , n48877 , n48614 );
xor ( n48879 , n48625 , n48629 );
xor ( n48880 , n48879 , n48633 );
and ( n48881 , n48878 , n48880 );
and ( n48882 , n47474 , n45990 );
and ( n48883 , n47351 , n45988 );
nor ( n48884 , n48882 , n48883 );
xnor ( n48885 , n48884 , n45939 );
and ( n48886 , n48108 , n45777 );
and ( n48887 , n47962 , n45775 );
nor ( n48888 , n48886 , n48887 );
xnor ( n48889 , n48888 , n45734 );
and ( n48890 , n48885 , n48889 );
and ( n48891 , n48384 , n45702 );
and ( n48892 , n48272 , n45700 );
nor ( n48893 , n48891 , n48892 );
xnor ( n48894 , n48893 , n20841 );
and ( n48895 , n48889 , n48894 );
and ( n48896 , n48885 , n48894 );
or ( n48897 , n48890 , n48895 , n48896 );
xor ( n48898 , n48702 , n48706 );
xor ( n48899 , n48898 , n48710 );
and ( n48900 , n48897 , n48899 );
and ( n48901 , n48880 , n48900 );
and ( n48902 , n48878 , n48900 );
or ( n48903 , n48881 , n48901 , n48902 );
xor ( n48904 , n48718 , n48722 );
xor ( n48905 , n48904 , n48727 );
and ( n48906 , n46345 , n46911 );
and ( n48907 , n46264 , n46909 );
nor ( n48908 , n48906 , n48907 );
xnor ( n48909 , n48908 , n46802 );
and ( n48910 , n46530 , n46712 );
and ( n48911 , n46445 , n46710 );
nor ( n48912 , n48910 , n48911 );
xnor ( n48913 , n48912 , n46587 );
and ( n48914 , n48909 , n48913 );
and ( n48915 , n48905 , n48914 );
buf ( n48916 , n48915 );
and ( n48917 , n47778 , n45886 );
and ( n48918 , n47647 , n45884 );
nor ( n48919 , n48917 , n48918 );
xnor ( n48920 , n48919 , n45824 );
and ( n48921 , n48709 , n20852 );
and ( n48922 , n48632 , n20850 );
nor ( n48923 , n48921 , n48922 );
xnor ( n48924 , n48923 , n20860 );
and ( n48925 , n48920 , n48924 );
buf ( n48926 , n17511 );
buf ( n48927 , n48926 );
buf ( n48928 , n17513 );
buf ( n48929 , n48928 );
and ( n48930 , n48927 , n48929 );
not ( n48931 , n48930 );
and ( n48932 , n48568 , n48931 );
not ( n48933 , n48932 );
and ( n48934 , n20844 , n48740 );
and ( n48935 , n20855 , n48738 );
nor ( n48936 , n48934 , n48935 );
xnor ( n48937 , n48936 , n48571 );
and ( n48938 , n48933 , n48937 );
and ( n48939 , n45712 , n48394 );
and ( n48940 , n20864 , n48392 );
nor ( n48941 , n48939 , n48940 );
xnor ( n48942 , n48941 , n48220 );
and ( n48943 , n48937 , n48942 );
and ( n48944 , n48933 , n48942 );
or ( n48945 , n48938 , n48943 , n48944 );
and ( n48946 , n48925 , n48945 );
and ( n48947 , n45794 , n48042 );
and ( n48948 , n45763 , n48040 );
nor ( n48949 , n48947 , n48948 );
xnor ( n48950 , n48949 , n47921 );
and ( n48951 , n45907 , n47734 );
and ( n48952 , n45843 , n47732 );
nor ( n48953 , n48951 , n48952 );
xnor ( n48954 , n48953 , n47606 );
and ( n48955 , n48950 , n48954 );
and ( n48956 , n46041 , n47429 );
and ( n48957 , n45963 , n47427 );
nor ( n48958 , n48956 , n48957 );
xnor ( n48959 , n48958 , n47309 );
and ( n48960 , n48954 , n48959 );
and ( n48961 , n48950 , n48959 );
or ( n48962 , n48955 , n48960 , n48961 );
and ( n48963 , n48945 , n48962 );
and ( n48964 , n48925 , n48962 );
or ( n48965 , n48946 , n48963 , n48964 );
and ( n48966 , n48916 , n48965 );
and ( n48967 , n46169 , n47178 );
and ( n48968 , n46100 , n47176 );
nor ( n48969 , n48967 , n48968 );
xnor ( n48970 , n48969 , n47039 );
and ( n48971 , n46750 , n46496 );
and ( n48972 , n46577 , n46494 );
nor ( n48973 , n48971 , n48972 );
xnor ( n48974 , n48973 , n46402 );
and ( n48975 , n48970 , n48974 );
and ( n48976 , n46969 , n46306 );
and ( n48977 , n46843 , n46304 );
nor ( n48978 , n48976 , n48977 );
xnor ( n48979 , n48978 , n46228 );
and ( n48980 , n48974 , n48979 );
and ( n48981 , n48970 , n48979 );
or ( n48982 , n48975 , n48980 , n48981 );
and ( n48983 , n47216 , n46135 );
and ( n48984 , n47090 , n46133 );
nor ( n48985 , n48983 , n48984 );
xnor ( n48986 , n48985 , n46067 );
buf ( n48987 , n20754 );
buf ( n48988 , n48987 );
and ( n48989 , n48988 , n20846 );
and ( n48990 , n48986 , n48989 );
xor ( n48991 , n25169 , n45633 );
buf ( n48992 , n48991 );
buf ( n48993 , n48992 );
buf ( n48994 , n48993 );
and ( n48995 , n48989 , n48994 );
and ( n48996 , n48986 , n48994 );
or ( n48997 , n48990 , n48995 , n48996 );
and ( n48998 , n48982 , n48997 );
xor ( n48999 , n48743 , n48747 );
xor ( n49000 , n48999 , n48752 );
and ( n49001 , n48997 , n49000 );
and ( n49002 , n48982 , n49000 );
or ( n49003 , n48998 , n49001 , n49002 );
and ( n49004 , n48965 , n49003 );
and ( n49005 , n48916 , n49003 );
or ( n49006 , n48966 , n49004 , n49005 );
and ( n49007 , n48903 , n49006 );
xor ( n49008 , n48759 , n48763 );
xor ( n49009 , n49008 , n48768 );
xor ( n49010 , n48776 , n48780 );
xor ( n49011 , n49010 , n48785 );
and ( n49012 , n49009 , n49011 );
xor ( n49013 , n48795 , n48799 );
xor ( n49014 , n49013 , n48804 );
and ( n49015 , n49011 , n49014 );
and ( n49016 , n49009 , n49014 );
or ( n49017 , n49012 , n49015 , n49016 );
buf ( n49018 , n48692 );
xor ( n49019 , n49018 , n48694 );
and ( n49020 , n49017 , n49019 );
xor ( n49021 , n48698 , n48713 );
xor ( n49022 , n49021 , n48730 );
and ( n49023 , n49019 , n49022 );
and ( n49024 , n49017 , n49022 );
or ( n49025 , n49020 , n49023 , n49024 );
and ( n49026 , n49006 , n49025 );
and ( n49027 , n48903 , n49025 );
or ( n49028 , n49007 , n49026 , n49027 );
xor ( n49029 , n48688 , n48696 );
xor ( n49030 , n49029 , n48733 );
xor ( n49031 , n48791 , n48815 );
xor ( n49032 , n49031 , n48818 );
and ( n49033 , n49030 , n49032 );
xor ( n49034 , n48824 , n48826 );
xor ( n49035 , n49034 , n48829 );
and ( n49036 , n49032 , n49035 );
and ( n49037 , n49030 , n49035 );
or ( n49038 , n49033 , n49036 , n49037 );
and ( n49039 , n49028 , n49038 );
xor ( n49040 , n48736 , n48821 );
xor ( n49041 , n49040 , n48832 );
and ( n49042 , n49038 , n49041 );
and ( n49043 , n49028 , n49041 );
or ( n49044 , n49039 , n49042 , n49043 );
and ( n49045 , n48875 , n49044 );
and ( n49046 , n48873 , n49044 );
or ( n49047 , n48876 , n49045 , n49046 );
xor ( n49048 , n48684 , n48849 );
xor ( n49049 , n49048 , n48852 );
and ( n49050 , n49047 , n49049 );
xor ( n49051 , n48686 , n48835 );
xor ( n49052 , n49051 , n48846 );
xor ( n49053 , n48838 , n48840 );
xor ( n49054 , n49053 , n48843 );
xor ( n49055 , n48755 , n48771 );
xor ( n49056 , n49055 , n48788 );
xor ( n49057 , n48807 , n48809 );
xor ( n49058 , n49057 , n48812 );
and ( n49059 , n49056 , n49058 );
xor ( n49060 , n48897 , n48899 );
xor ( n49061 , n48885 , n48889 );
xor ( n49062 , n49061 , n48894 );
xor ( n49063 , n48909 , n48913 );
and ( n49064 , n49062 , n49063 );
buf ( n49065 , n49064 );
and ( n49066 , n49060 , n49065 );
xor ( n49067 , n48920 , n48924 );
and ( n49068 , n47090 , n46306 );
and ( n49069 , n46969 , n46304 );
nor ( n49070 , n49068 , n49069 );
xnor ( n49071 , n49070 , n46228 );
and ( n49072 , n47351 , n46135 );
and ( n49073 , n47216 , n46133 );
nor ( n49074 , n49072 , n49073 );
xnor ( n49075 , n49074 , n46067 );
and ( n49076 , n49071 , n49075 );
and ( n49077 , n48272 , n45777 );
and ( n49078 , n48108 , n45775 );
nor ( n49079 , n49077 , n49078 );
xnor ( n49080 , n49079 , n45734 );
and ( n49081 , n49075 , n49080 );
and ( n49082 , n49071 , n49080 );
or ( n49083 , n49076 , n49081 , n49082 );
and ( n49084 , n49067 , n49083 );
and ( n49085 , n47647 , n45990 );
and ( n49086 , n47474 , n45988 );
nor ( n49087 , n49085 , n49086 );
xnor ( n49088 , n49087 , n45939 );
and ( n49089 , n47962 , n45886 );
and ( n49090 , n47778 , n45884 );
nor ( n49091 , n49089 , n49090 );
xnor ( n49092 , n49091 , n45824 );
and ( n49093 , n49088 , n49092 );
and ( n49094 , n48988 , n20852 );
and ( n49095 , n48709 , n20850 );
nor ( n49096 , n49094 , n49095 );
xnor ( n49097 , n49096 , n20860 );
and ( n49098 , n49092 , n49097 );
and ( n49099 , n49088 , n49097 );
or ( n49100 , n49093 , n49098 , n49099 );
and ( n49101 , n49083 , n49100 );
and ( n49102 , n49067 , n49100 );
or ( n49103 , n49084 , n49101 , n49102 );
and ( n49104 , n49065 , n49103 );
and ( n49105 , n49060 , n49103 );
or ( n49106 , n49066 , n49104 , n49105 );
and ( n49107 , n49058 , n49106 );
and ( n49108 , n49056 , n49106 );
or ( n49109 , n49059 , n49107 , n49108 );
and ( n49110 , n46264 , n47178 );
and ( n49111 , n46169 , n47176 );
nor ( n49112 , n49110 , n49111 );
xnor ( n49113 , n49112 , n47039 );
buf ( n49114 , n20756 );
buf ( n49115 , n49114 );
and ( n49116 , n49115 , n20846 );
and ( n49117 , n49113 , n49116 );
xor ( n49118 , n48568 , n48927 );
xor ( n49119 , n48927 , n48929 );
not ( n49120 , n49119 );
and ( n49121 , n49118 , n49120 );
and ( n49122 , n20855 , n49121 );
not ( n49123 , n49122 );
xnor ( n49124 , n49123 , n48932 );
and ( n49125 , n20864 , n48740 );
and ( n49126 , n20844 , n48738 );
nor ( n49127 , n49125 , n49126 );
xnor ( n49128 , n49127 , n48571 );
and ( n49129 , n49124 , n49128 );
and ( n49130 , n45763 , n48394 );
and ( n49131 , n45712 , n48392 );
nor ( n49132 , n49130 , n49131 );
xnor ( n49133 , n49132 , n48220 );
and ( n49134 , n49128 , n49133 );
and ( n49135 , n49124 , n49133 );
or ( n49136 , n49129 , n49134 , n49135 );
and ( n49137 , n49117 , n49136 );
and ( n49138 , n45843 , n48042 );
and ( n49139 , n45794 , n48040 );
nor ( n49140 , n49138 , n49139 );
xnor ( n49141 , n49140 , n47921 );
and ( n49142 , n45963 , n47734 );
and ( n49143 , n45907 , n47732 );
nor ( n49144 , n49142 , n49143 );
xnor ( n49145 , n49144 , n47606 );
and ( n49146 , n49141 , n49145 );
and ( n49147 , n46100 , n47429 );
and ( n49148 , n46041 , n47427 );
nor ( n49149 , n49147 , n49148 );
xnor ( n49150 , n49149 , n47309 );
and ( n49151 , n49145 , n49150 );
and ( n49152 , n49141 , n49150 );
or ( n49153 , n49146 , n49151 , n49152 );
and ( n49154 , n49136 , n49153 );
and ( n49155 , n49117 , n49153 );
or ( n49156 , n49137 , n49154 , n49155 );
and ( n49157 , n46445 , n46911 );
and ( n49158 , n46345 , n46909 );
nor ( n49159 , n49157 , n49158 );
xnor ( n49160 , n49159 , n46802 );
and ( n49161 , n46577 , n46712 );
and ( n49162 , n46530 , n46710 );
nor ( n49163 , n49161 , n49162 );
xnor ( n49164 , n49163 , n46587 );
and ( n49165 , n49160 , n49164 );
and ( n49166 , n46843 , n46496 );
and ( n49167 , n46750 , n46494 );
nor ( n49168 , n49166 , n49167 );
xnor ( n49169 , n49168 , n46402 );
and ( n49170 , n49164 , n49169 );
and ( n49171 , n49160 , n49169 );
or ( n49172 , n49165 , n49170 , n49171 );
and ( n49173 , n48632 , n45702 );
and ( n49174 , n48384 , n45700 );
nor ( n49175 , n49173 , n49174 );
xnor ( n49176 , n49175 , n20841 );
xor ( n49177 , n25170 , n45632 );
buf ( n49178 , n49177 );
buf ( n49179 , n49178 );
buf ( n49180 , n49179 );
and ( n49181 , n49176 , n49180 );
buf ( n49182 , n49181 );
and ( n49183 , n49172 , n49182 );
xor ( n49184 , n48933 , n48937 );
xor ( n49185 , n49184 , n48942 );
and ( n49186 , n49182 , n49185 );
and ( n49187 , n49172 , n49185 );
or ( n49188 , n49183 , n49186 , n49187 );
and ( n49189 , n49156 , n49188 );
xor ( n49190 , n48950 , n48954 );
xor ( n49191 , n49190 , n48959 );
xor ( n49192 , n48970 , n48974 );
xor ( n49193 , n49192 , n48979 );
and ( n49194 , n49191 , n49193 );
xor ( n49195 , n48986 , n48989 );
xor ( n49196 , n49195 , n48994 );
and ( n49197 , n49193 , n49196 );
and ( n49198 , n49191 , n49196 );
or ( n49199 , n49194 , n49197 , n49198 );
and ( n49200 , n49188 , n49199 );
and ( n49201 , n49156 , n49199 );
or ( n49202 , n49189 , n49200 , n49201 );
buf ( n49203 , n48905 );
xor ( n49204 , n49203 , n48914 );
xor ( n49205 , n48925 , n48945 );
xor ( n49206 , n49205 , n48962 );
and ( n49207 , n49204 , n49206 );
xor ( n49208 , n48982 , n48997 );
xor ( n49209 , n49208 , n49000 );
and ( n49210 , n49206 , n49209 );
and ( n49211 , n49204 , n49209 );
or ( n49212 , n49207 , n49210 , n49211 );
and ( n49213 , n49202 , n49212 );
xor ( n49214 , n48878 , n48880 );
xor ( n49215 , n49214 , n48900 );
and ( n49216 , n49212 , n49215 );
and ( n49217 , n49202 , n49215 );
or ( n49218 , n49213 , n49216 , n49217 );
and ( n49219 , n49109 , n49218 );
xor ( n49220 , n48903 , n49006 );
xor ( n49221 , n49220 , n49025 );
and ( n49222 , n49218 , n49221 );
and ( n49223 , n49109 , n49221 );
or ( n49224 , n49219 , n49222 , n49223 );
and ( n49225 , n49054 , n49224 );
xor ( n49226 , n49028 , n49038 );
xor ( n49227 , n49226 , n49041 );
and ( n49228 , n49224 , n49227 );
and ( n49229 , n49054 , n49227 );
or ( n49230 , n49225 , n49228 , n49229 );
and ( n49231 , n49052 , n49230 );
xor ( n49232 , n48873 , n48875 );
xor ( n49233 , n49232 , n49044 );
and ( n49234 , n49230 , n49233 );
and ( n49235 , n49052 , n49233 );
or ( n49236 , n49231 , n49234 , n49235 );
and ( n49237 , n49049 , n49236 );
and ( n49238 , n49047 , n49236 );
or ( n49239 , n49050 , n49237 , n49238 );
and ( n49240 , n48871 , n49239 );
xor ( n49241 , n48871 , n49239 );
xor ( n49242 , n49047 , n49049 );
xor ( n49243 , n49242 , n49236 );
not ( n49244 , n49243 );
xor ( n49245 , n49052 , n49230 );
xor ( n49246 , n49245 , n49233 );
xor ( n49247 , n49030 , n49032 );
xor ( n49248 , n49247 , n49035 );
xor ( n49249 , n48916 , n48965 );
xor ( n49250 , n49249 , n49003 );
xor ( n49251 , n49017 , n49019 );
xor ( n49252 , n49251 , n49022 );
and ( n49253 , n49250 , n49252 );
xor ( n49254 , n49009 , n49011 );
xor ( n49255 , n49254 , n49014 );
xor ( n49256 , n49071 , n49075 );
xor ( n49257 , n49256 , n49080 );
xor ( n49258 , n49088 , n49092 );
xor ( n49259 , n49258 , n49097 );
and ( n49260 , n49257 , n49259 );
xor ( n49261 , n49113 , n49116 );
and ( n49262 , n49259 , n49261 );
and ( n49263 , n49257 , n49261 );
or ( n49264 , n49260 , n49262 , n49263 );
and ( n49265 , n47216 , n46306 );
and ( n49266 , n47090 , n46304 );
nor ( n49267 , n49265 , n49266 );
xnor ( n49268 , n49267 , n46228 );
and ( n49269 , n47474 , n46135 );
and ( n49270 , n47351 , n46133 );
nor ( n49271 , n49269 , n49270 );
xnor ( n49272 , n49271 , n46067 );
and ( n49273 , n49268 , n49272 );
and ( n49274 , n47778 , n45990 );
and ( n49275 , n47647 , n45988 );
nor ( n49276 , n49274 , n49275 );
xnor ( n49277 , n49276 , n45939 );
and ( n49278 , n49272 , n49277 );
and ( n49279 , n49268 , n49277 );
or ( n49280 , n49273 , n49278 , n49279 );
and ( n49281 , n46345 , n47178 );
and ( n49282 , n46264 , n47176 );
nor ( n49283 , n49281 , n49282 );
xnor ( n49284 , n49283 , n47039 );
and ( n49285 , n46530 , n46911 );
and ( n49286 , n46445 , n46909 );
nor ( n49287 , n49285 , n49286 );
xnor ( n49288 , n49287 , n46802 );
and ( n49289 , n49284 , n49288 );
and ( n49290 , n49280 , n49289 );
and ( n49291 , n48384 , n45777 );
and ( n49292 , n48272 , n45775 );
nor ( n49293 , n49291 , n49292 );
xnor ( n49294 , n49293 , n45734 );
and ( n49295 , n48709 , n45702 );
and ( n49296 , n48632 , n45700 );
nor ( n49297 , n49295 , n49296 );
xnor ( n49298 , n49297 , n20841 );
and ( n49299 , n49294 , n49298 );
and ( n49300 , n49289 , n49299 );
and ( n49301 , n49280 , n49299 );
or ( n49302 , n49290 , n49300 , n49301 );
and ( n49303 , n49264 , n49302 );
buf ( n49304 , n17515 );
buf ( n49305 , n49304 );
buf ( n49306 , n17517 );
buf ( n49307 , n49306 );
and ( n49308 , n49305 , n49307 );
not ( n49309 , n49308 );
and ( n49310 , n48929 , n49309 );
not ( n49311 , n49310 );
and ( n49312 , n20844 , n49121 );
and ( n49313 , n20855 , n49119 );
nor ( n49314 , n49312 , n49313 );
xnor ( n49315 , n49314 , n48932 );
and ( n49316 , n49311 , n49315 );
and ( n49317 , n45712 , n48740 );
and ( n49318 , n20864 , n48738 );
nor ( n49319 , n49317 , n49318 );
xnor ( n49320 , n49319 , n48571 );
and ( n49321 , n49315 , n49320 );
and ( n49322 , n49311 , n49320 );
or ( n49323 , n49316 , n49321 , n49322 );
and ( n49324 , n45794 , n48394 );
and ( n49325 , n45763 , n48392 );
nor ( n49326 , n49324 , n49325 );
xnor ( n49327 , n49326 , n48220 );
and ( n49328 , n45907 , n48042 );
and ( n49329 , n45843 , n48040 );
nor ( n49330 , n49328 , n49329 );
xnor ( n49331 , n49330 , n47921 );
and ( n49332 , n49327 , n49331 );
and ( n49333 , n46041 , n47734 );
and ( n49334 , n45963 , n47732 );
nor ( n49335 , n49333 , n49334 );
xnor ( n49336 , n49335 , n47606 );
and ( n49337 , n49331 , n49336 );
and ( n49338 , n49327 , n49336 );
or ( n49339 , n49332 , n49337 , n49338 );
and ( n49340 , n49323 , n49339 );
and ( n49341 , n46169 , n47429 );
and ( n49342 , n46100 , n47427 );
nor ( n49343 , n49341 , n49342 );
xnor ( n49344 , n49343 , n47309 );
and ( n49345 , n46750 , n46712 );
and ( n49346 , n46577 , n46710 );
nor ( n49347 , n49345 , n49346 );
xnor ( n49348 , n49347 , n46587 );
and ( n49349 , n49344 , n49348 );
and ( n49350 , n46969 , n46496 );
and ( n49351 , n46843 , n46494 );
nor ( n49352 , n49350 , n49351 );
xnor ( n49353 , n49352 , n46402 );
and ( n49354 , n49348 , n49353 );
and ( n49355 , n49344 , n49353 );
or ( n49356 , n49349 , n49354 , n49355 );
and ( n49357 , n49339 , n49356 );
and ( n49358 , n49323 , n49356 );
or ( n49359 , n49340 , n49357 , n49358 );
and ( n49360 , n49302 , n49359 );
and ( n49361 , n49264 , n49359 );
or ( n49362 , n49303 , n49360 , n49361 );
and ( n49363 , n49255 , n49362 );
and ( n49364 , n48108 , n45886 );
and ( n49365 , n47962 , n45884 );
nor ( n49366 , n49364 , n49365 );
xnor ( n49367 , n49366 , n45824 );
and ( n49368 , n49115 , n20852 );
and ( n49369 , n48988 , n20850 );
nor ( n49370 , n49368 , n49369 );
xnor ( n49371 , n49370 , n20860 );
and ( n49372 , n49367 , n49371 );
buf ( n49373 , n20758 );
buf ( n49374 , n49373 );
and ( n49375 , n49374 , n20846 );
and ( n49376 , n49371 , n49375 );
and ( n49377 , n49367 , n49375 );
or ( n49378 , n49372 , n49376 , n49377 );
xor ( n49379 , n49124 , n49128 );
xor ( n49380 , n49379 , n49133 );
and ( n49381 , n49378 , n49380 );
xor ( n49382 , n49141 , n49145 );
xor ( n49383 , n49382 , n49150 );
and ( n49384 , n49380 , n49383 );
and ( n49385 , n49378 , n49383 );
or ( n49386 , n49381 , n49384 , n49385 );
buf ( n49387 , n49062 );
xor ( n49388 , n49387 , n49063 );
and ( n49389 , n49386 , n49388 );
xor ( n49390 , n49067 , n49083 );
xor ( n49391 , n49390 , n49100 );
and ( n49392 , n49388 , n49391 );
and ( n49393 , n49386 , n49391 );
or ( n49394 , n49389 , n49392 , n49393 );
and ( n49395 , n49362 , n49394 );
and ( n49396 , n49255 , n49394 );
or ( n49397 , n49363 , n49395 , n49396 );
and ( n49398 , n49252 , n49397 );
and ( n49399 , n49250 , n49397 );
or ( n49400 , n49253 , n49398 , n49399 );
and ( n49401 , n49248 , n49400 );
xor ( n49402 , n49117 , n49136 );
xor ( n49403 , n49402 , n49153 );
xor ( n49404 , n49172 , n49182 );
xor ( n49405 , n49404 , n49185 );
and ( n49406 , n49403 , n49405 );
xor ( n49407 , n49191 , n49193 );
xor ( n49408 , n49407 , n49196 );
and ( n49409 , n49405 , n49408 );
and ( n49410 , n49403 , n49408 );
or ( n49411 , n49406 , n49409 , n49410 );
xor ( n49412 , n49060 , n49065 );
xor ( n49413 , n49412 , n49103 );
and ( n49414 , n49411 , n49413 );
xor ( n49415 , n49156 , n49188 );
xor ( n49416 , n49415 , n49199 );
and ( n49417 , n49413 , n49416 );
and ( n49418 , n49411 , n49416 );
or ( n49419 , n49414 , n49417 , n49418 );
xor ( n49420 , n49056 , n49058 );
xor ( n49421 , n49420 , n49106 );
and ( n49422 , n49419 , n49421 );
xor ( n49423 , n49202 , n49212 );
xor ( n49424 , n49423 , n49215 );
and ( n49425 , n49421 , n49424 );
and ( n49426 , n49419 , n49424 );
or ( n49427 , n49422 , n49425 , n49426 );
and ( n49428 , n49400 , n49427 );
and ( n49429 , n49248 , n49427 );
or ( n49430 , n49401 , n49428 , n49429 );
xor ( n49431 , n49054 , n49224 );
xor ( n49432 , n49431 , n49227 );
and ( n49433 , n49430 , n49432 );
xor ( n49434 , n49109 , n49218 );
xor ( n49435 , n49434 , n49221 );
xor ( n49436 , n49204 , n49206 );
xor ( n49437 , n49436 , n49209 );
xor ( n49438 , n49160 , n49164 );
xor ( n49439 , n49438 , n49169 );
xor ( n49440 , n49176 , n49180 );
buf ( n49441 , n49440 );
and ( n49442 , n49439 , n49441 );
and ( n49443 , n47647 , n46135 );
and ( n49444 , n47474 , n46133 );
nor ( n49445 , n49443 , n49444 );
xnor ( n49446 , n49445 , n46067 );
and ( n49447 , n47962 , n45990 );
and ( n49448 , n47778 , n45988 );
nor ( n49449 , n49447 , n49448 );
xnor ( n49450 , n49449 , n45939 );
and ( n49451 , n49446 , n49450 );
and ( n49452 , n49374 , n20852 );
and ( n49453 , n49115 , n20850 );
nor ( n49454 , n49452 , n49453 );
xnor ( n49455 , n49454 , n20860 );
and ( n49456 , n49450 , n49455 );
and ( n49457 , n49446 , n49455 );
or ( n49458 , n49451 , n49456 , n49457 );
and ( n49459 , n47351 , n46306 );
and ( n49460 , n47216 , n46304 );
nor ( n49461 , n49459 , n49460 );
xnor ( n49462 , n49461 , n46228 );
and ( n49463 , n48632 , n45777 );
and ( n49464 , n48384 , n45775 );
nor ( n49465 , n49463 , n49464 );
xnor ( n49466 , n49465 , n45734 );
and ( n49467 , n49462 , n49466 );
and ( n49468 , n48988 , n45702 );
and ( n49469 , n48709 , n45700 );
nor ( n49470 , n49468 , n49469 );
xnor ( n49471 , n49470 , n20841 );
and ( n49472 , n49466 , n49471 );
and ( n49473 , n49462 , n49471 );
or ( n49474 , n49467 , n49472 , n49473 );
and ( n49475 , n49458 , n49474 );
and ( n49476 , n49441 , n49475 );
and ( n49477 , n49439 , n49475 );
or ( n49478 , n49442 , n49476 , n49477 );
xor ( n49479 , n25171 , n45631 );
buf ( n49480 , n49479 );
buf ( n49481 , n49480 );
buf ( n49482 , n49481 );
xor ( n49483 , n49268 , n49272 );
xor ( n49484 , n49483 , n49277 );
and ( n49485 , n49482 , n49484 );
buf ( n49486 , n49485 );
xor ( n49487 , n49284 , n49288 );
xor ( n49488 , n49294 , n49298 );
and ( n49489 , n49487 , n49488 );
and ( n49490 , n46264 , n47429 );
and ( n49491 , n46169 , n47427 );
nor ( n49492 , n49490 , n49491 );
xnor ( n49493 , n49492 , n47309 );
and ( n49494 , n46445 , n47178 );
and ( n49495 , n46345 , n47176 );
nor ( n49496 , n49494 , n49495 );
xnor ( n49497 , n49496 , n47039 );
and ( n49498 , n49493 , n49497 );
and ( n49499 , n46577 , n46911 );
and ( n49500 , n46530 , n46909 );
nor ( n49501 , n49499 , n49500 );
xnor ( n49502 , n49501 , n46802 );
and ( n49503 , n49497 , n49502 );
and ( n49504 , n49493 , n49502 );
or ( n49505 , n49498 , n49503 , n49504 );
and ( n49506 , n49488 , n49505 );
and ( n49507 , n49487 , n49505 );
or ( n49508 , n49489 , n49506 , n49507 );
and ( n49509 , n49486 , n49508 );
xor ( n49510 , n48929 , n49305 );
xor ( n49511 , n49305 , n49307 );
not ( n49512 , n49511 );
and ( n49513 , n49510 , n49512 );
and ( n49514 , n20855 , n49513 );
not ( n49515 , n49514 );
xnor ( n49516 , n49515 , n49310 );
and ( n49517 , n20864 , n49121 );
and ( n49518 , n20844 , n49119 );
nor ( n49519 , n49517 , n49518 );
xnor ( n49520 , n49519 , n48932 );
and ( n49521 , n49516 , n49520 );
and ( n49522 , n45763 , n48740 );
and ( n49523 , n45712 , n48738 );
nor ( n49524 , n49522 , n49523 );
xnor ( n49525 , n49524 , n48571 );
and ( n49526 , n49520 , n49525 );
and ( n49527 , n49516 , n49525 );
or ( n49528 , n49521 , n49526 , n49527 );
and ( n49529 , n45843 , n48394 );
and ( n49530 , n45794 , n48392 );
nor ( n49531 , n49529 , n49530 );
xnor ( n49532 , n49531 , n48220 );
and ( n49533 , n45963 , n48042 );
and ( n49534 , n45907 , n48040 );
nor ( n49535 , n49533 , n49534 );
xnor ( n49536 , n49535 , n47921 );
and ( n49537 , n49532 , n49536 );
and ( n49538 , n46100 , n47734 );
and ( n49539 , n46041 , n47732 );
nor ( n49540 , n49538 , n49539 );
xnor ( n49541 , n49540 , n47606 );
and ( n49542 , n49536 , n49541 );
and ( n49543 , n49532 , n49541 );
or ( n49544 , n49537 , n49542 , n49543 );
and ( n49545 , n49528 , n49544 );
and ( n49546 , n46843 , n46712 );
and ( n49547 , n46750 , n46710 );
nor ( n49548 , n49546 , n49547 );
xnor ( n49549 , n49548 , n46587 );
and ( n49550 , n47090 , n46496 );
and ( n49551 , n46969 , n46494 );
nor ( n49552 , n49550 , n49551 );
xnor ( n49553 , n49552 , n46402 );
and ( n49554 , n49549 , n49553 );
and ( n49555 , n48272 , n45886 );
and ( n49556 , n48108 , n45884 );
nor ( n49557 , n49555 , n49556 );
xnor ( n49558 , n49557 , n45824 );
and ( n49559 , n49553 , n49558 );
and ( n49560 , n49549 , n49558 );
or ( n49561 , n49554 , n49559 , n49560 );
and ( n49562 , n49544 , n49561 );
and ( n49563 , n49528 , n49561 );
or ( n49564 , n49545 , n49562 , n49563 );
and ( n49565 , n49508 , n49564 );
and ( n49566 , n49486 , n49564 );
or ( n49567 , n49509 , n49565 , n49566 );
and ( n49568 , n49478 , n49567 );
buf ( n49569 , n20760 );
buf ( n49570 , n49569 );
and ( n49571 , n49570 , n20846 );
xor ( n49572 , n25172 , n45630 );
buf ( n49573 , n49572 );
buf ( n49574 , n49573 );
buf ( n49575 , n49574 );
and ( n49576 , n49571 , n49575 );
buf ( n49577 , n49576 );
xor ( n49578 , n49311 , n49315 );
xor ( n49579 , n49578 , n49320 );
and ( n49580 , n49577 , n49579 );
xor ( n49581 , n49327 , n49331 );
xor ( n49582 , n49581 , n49336 );
and ( n49583 , n49579 , n49582 );
and ( n49584 , n49577 , n49582 );
or ( n49585 , n49580 , n49583 , n49584 );
xor ( n49586 , n49257 , n49259 );
xor ( n49587 , n49586 , n49261 );
and ( n49588 , n49585 , n49587 );
xor ( n49589 , n49280 , n49289 );
xor ( n49590 , n49589 , n49299 );
and ( n49591 , n49587 , n49590 );
and ( n49592 , n49585 , n49590 );
or ( n49593 , n49588 , n49591 , n49592 );
and ( n49594 , n49567 , n49593 );
and ( n49595 , n49478 , n49593 );
or ( n49596 , n49568 , n49594 , n49595 );
and ( n49597 , n49437 , n49596 );
xor ( n49598 , n49264 , n49302 );
xor ( n49599 , n49598 , n49359 );
xor ( n49600 , n49386 , n49388 );
xor ( n49601 , n49600 , n49391 );
and ( n49602 , n49599 , n49601 );
xor ( n49603 , n49403 , n49405 );
xor ( n49604 , n49603 , n49408 );
and ( n49605 , n49601 , n49604 );
and ( n49606 , n49599 , n49604 );
or ( n49607 , n49602 , n49605 , n49606 );
and ( n49608 , n49596 , n49607 );
and ( n49609 , n49437 , n49607 );
or ( n49610 , n49597 , n49608 , n49609 );
xor ( n49611 , n49250 , n49252 );
xor ( n49612 , n49611 , n49397 );
and ( n49613 , n49610 , n49612 );
xor ( n49614 , n49419 , n49421 );
xor ( n49615 , n49614 , n49424 );
and ( n49616 , n49612 , n49615 );
and ( n49617 , n49610 , n49615 );
or ( n49618 , n49613 , n49616 , n49617 );
and ( n49619 , n49435 , n49618 );
xor ( n49620 , n49248 , n49400 );
xor ( n49621 , n49620 , n49427 );
and ( n49622 , n49618 , n49621 );
and ( n49623 , n49435 , n49621 );
or ( n49624 , n49619 , n49622 , n49623 );
and ( n49625 , n49432 , n49624 );
and ( n49626 , n49430 , n49624 );
or ( n49627 , n49433 , n49625 , n49626 );
and ( n49628 , n49246 , n49627 );
xor ( n49629 , n49246 , n49627 );
xor ( n49630 , n49430 , n49432 );
xor ( n49631 , n49630 , n49624 );
xor ( n49632 , n49435 , n49618 );
xor ( n49633 , n49632 , n49621 );
xor ( n49634 , n49255 , n49362 );
xor ( n49635 , n49634 , n49394 );
xor ( n49636 , n49411 , n49413 );
xor ( n49637 , n49636 , n49416 );
and ( n49638 , n49635 , n49637 );
xor ( n49639 , n49323 , n49339 );
xor ( n49640 , n49639 , n49356 );
xor ( n49641 , n49378 , n49380 );
xor ( n49642 , n49641 , n49383 );
and ( n49643 , n49640 , n49642 );
xor ( n49644 , n49344 , n49348 );
xor ( n49645 , n49644 , n49353 );
xor ( n49646 , n49367 , n49371 );
xor ( n49647 , n49646 , n49375 );
and ( n49648 , n49645 , n49647 );
xor ( n49649 , n49458 , n49474 );
and ( n49650 , n49647 , n49649 );
and ( n49651 , n49645 , n49649 );
or ( n49652 , n49648 , n49650 , n49651 );
and ( n49653 , n49642 , n49652 );
and ( n49654 , n49640 , n49652 );
or ( n49655 , n49643 , n49653 , n49654 );
xor ( n49656 , n49446 , n49450 );
xor ( n49657 , n49656 , n49455 );
xor ( n49658 , n49493 , n49497 );
xor ( n49659 , n49658 , n49502 );
and ( n49660 , n49657 , n49659 );
xor ( n49661 , n49462 , n49466 );
xor ( n49662 , n49661 , n49471 );
and ( n49663 , n49659 , n49662 );
and ( n49664 , n49657 , n49662 );
or ( n49665 , n49660 , n49663 , n49664 );
and ( n49666 , n46530 , n47178 );
and ( n49667 , n46445 , n47176 );
nor ( n49668 , n49666 , n49667 );
xnor ( n49669 , n49668 , n47039 );
and ( n49670 , n46750 , n46911 );
and ( n49671 , n46577 , n46909 );
nor ( n49672 , n49670 , n49671 );
xnor ( n49673 , n49672 , n46802 );
and ( n49674 , n49669 , n49673 );
and ( n49675 , n46969 , n46712 );
and ( n49676 , n46843 , n46710 );
nor ( n49677 , n49675 , n49676 );
xnor ( n49678 , n49677 , n46587 );
and ( n49679 , n49673 , n49678 );
and ( n49680 , n49669 , n49678 );
or ( n49681 , n49674 , n49679 , n49680 );
and ( n49682 , n48108 , n45990 );
and ( n49683 , n47962 , n45988 );
nor ( n49684 , n49682 , n49683 );
xnor ( n49685 , n49684 , n45939 );
and ( n49686 , n49115 , n45702 );
and ( n49687 , n48988 , n45700 );
nor ( n49688 , n49686 , n49687 );
xnor ( n49689 , n49688 , n20841 );
or ( n49690 , n49685 , n49689 );
and ( n49691 , n49681 , n49690 );
and ( n49692 , n47474 , n46306 );
and ( n49693 , n47351 , n46304 );
nor ( n49694 , n49692 , n49693 );
xnor ( n49695 , n49694 , n46228 );
and ( n49696 , n49570 , n20852 );
and ( n49697 , n49374 , n20850 );
nor ( n49698 , n49696 , n49697 );
xnor ( n49699 , n49698 , n20860 );
and ( n49700 , n49695 , n49699 );
and ( n49701 , n49690 , n49700 );
and ( n49702 , n49681 , n49700 );
or ( n49703 , n49691 , n49701 , n49702 );
and ( n49704 , n49665 , n49703 );
buf ( n49705 , n17519 );
buf ( n49706 , n49705 );
buf ( n49707 , n17521 );
buf ( n49708 , n49707 );
and ( n49709 , n49706 , n49708 );
not ( n49710 , n49709 );
and ( n49711 , n49307 , n49710 );
not ( n49712 , n49711 );
and ( n49713 , n20844 , n49513 );
and ( n49714 , n20855 , n49511 );
nor ( n49715 , n49713 , n49714 );
xnor ( n49716 , n49715 , n49310 );
and ( n49717 , n49712 , n49716 );
and ( n49718 , n45712 , n49121 );
and ( n49719 , n20864 , n49119 );
nor ( n49720 , n49718 , n49719 );
xnor ( n49721 , n49720 , n48932 );
and ( n49722 , n49716 , n49721 );
and ( n49723 , n49712 , n49721 );
or ( n49724 , n49717 , n49722 , n49723 );
and ( n49725 , n45794 , n48740 );
and ( n49726 , n45763 , n48738 );
nor ( n49727 , n49725 , n49726 );
xnor ( n49728 , n49727 , n48571 );
and ( n49729 , n45907 , n48394 );
and ( n49730 , n45843 , n48392 );
nor ( n49731 , n49729 , n49730 );
xnor ( n49732 , n49731 , n48220 );
and ( n49733 , n49728 , n49732 );
and ( n49734 , n46041 , n48042 );
and ( n49735 , n45963 , n48040 );
nor ( n49736 , n49734 , n49735 );
xnor ( n49737 , n49736 , n47921 );
and ( n49738 , n49732 , n49737 );
and ( n49739 , n49728 , n49737 );
or ( n49740 , n49733 , n49738 , n49739 );
and ( n49741 , n49724 , n49740 );
and ( n49742 , n46169 , n47734 );
and ( n49743 , n46100 , n47732 );
nor ( n49744 , n49742 , n49743 );
xnor ( n49745 , n49744 , n47606 );
and ( n49746 , n46345 , n47429 );
and ( n49747 , n46264 , n47427 );
nor ( n49748 , n49746 , n49747 );
xnor ( n49749 , n49748 , n47309 );
and ( n49750 , n49745 , n49749 );
and ( n49751 , n47216 , n46496 );
and ( n49752 , n47090 , n46494 );
nor ( n49753 , n49751 , n49752 );
xnor ( n49754 , n49753 , n46402 );
and ( n49755 , n49749 , n49754 );
and ( n49756 , n49745 , n49754 );
or ( n49757 , n49750 , n49755 , n49756 );
and ( n49758 , n49740 , n49757 );
and ( n49759 , n49724 , n49757 );
or ( n49760 , n49741 , n49758 , n49759 );
and ( n49761 , n49703 , n49760 );
and ( n49762 , n49665 , n49760 );
or ( n49763 , n49704 , n49761 , n49762 );
and ( n49764 , n47778 , n46135 );
and ( n49765 , n47647 , n46133 );
nor ( n49766 , n49764 , n49765 );
xnor ( n49767 , n49766 , n46067 );
and ( n49768 , n48384 , n45886 );
and ( n49769 , n48272 , n45884 );
nor ( n49770 , n49768 , n49769 );
xnor ( n49771 , n49770 , n45824 );
and ( n49772 , n49767 , n49771 );
and ( n49773 , n48709 , n45777 );
and ( n49774 , n48632 , n45775 );
nor ( n49775 , n49773 , n49774 );
xnor ( n49776 , n49775 , n45734 );
and ( n49777 , n49771 , n49776 );
and ( n49778 , n49767 , n49776 );
or ( n49779 , n49772 , n49777 , n49778 );
buf ( n49780 , n20762 );
buf ( n49781 , n49780 );
and ( n49782 , n49781 , n20846 );
xor ( n49783 , n25173 , n45629 );
buf ( n49784 , n49783 );
buf ( n49785 , n49784 );
buf ( n49786 , n49785 );
and ( n49787 , n49782 , n49786 );
buf ( n49788 , n49787 );
and ( n49789 , n49779 , n49788 );
xor ( n49790 , n49516 , n49520 );
xor ( n49791 , n49790 , n49525 );
and ( n49792 , n49788 , n49791 );
and ( n49793 , n49779 , n49791 );
or ( n49794 , n49789 , n49792 , n49793 );
xor ( n49795 , n49532 , n49536 );
xor ( n49796 , n49795 , n49541 );
xor ( n49797 , n49549 , n49553 );
xor ( n49798 , n49797 , n49558 );
and ( n49799 , n49796 , n49798 );
xor ( n49800 , n49571 , n49575 );
buf ( n49801 , n49800 );
and ( n49802 , n49798 , n49801 );
and ( n49803 , n49796 , n49801 );
or ( n49804 , n49799 , n49802 , n49803 );
and ( n49805 , n49794 , n49804 );
buf ( n49806 , n49482 );
xor ( n49807 , n49806 , n49484 );
and ( n49808 , n49804 , n49807 );
and ( n49809 , n49794 , n49807 );
or ( n49810 , n49805 , n49808 , n49809 );
and ( n49811 , n49763 , n49810 );
xor ( n49812 , n49487 , n49488 );
xor ( n49813 , n49812 , n49505 );
xor ( n49814 , n49528 , n49544 );
xor ( n49815 , n49814 , n49561 );
and ( n49816 , n49813 , n49815 );
xor ( n49817 , n49577 , n49579 );
xor ( n49818 , n49817 , n49582 );
and ( n49819 , n49815 , n49818 );
and ( n49820 , n49813 , n49818 );
or ( n49821 , n49816 , n49819 , n49820 );
and ( n49822 , n49810 , n49821 );
and ( n49823 , n49763 , n49821 );
or ( n49824 , n49811 , n49822 , n49823 );
and ( n49825 , n49655 , n49824 );
xor ( n49826 , n49439 , n49441 );
xor ( n49827 , n49826 , n49475 );
xor ( n49828 , n49486 , n49508 );
xor ( n49829 , n49828 , n49564 );
and ( n49830 , n49827 , n49829 );
xor ( n49831 , n49585 , n49587 );
xor ( n49832 , n49831 , n49590 );
and ( n49833 , n49829 , n49832 );
and ( n49834 , n49827 , n49832 );
or ( n49835 , n49830 , n49833 , n49834 );
and ( n49836 , n49824 , n49835 );
and ( n49837 , n49655 , n49835 );
or ( n49838 , n49825 , n49836 , n49837 );
and ( n49839 , n49637 , n49838 );
and ( n49840 , n49635 , n49838 );
or ( n49841 , n49638 , n49839 , n49840 );
xor ( n49842 , n49610 , n49612 );
xor ( n49843 , n49842 , n49615 );
and ( n49844 , n49841 , n49843 );
xor ( n49845 , n49437 , n49596 );
xor ( n49846 , n49845 , n49607 );
xor ( n49847 , n49478 , n49567 );
xor ( n49848 , n49847 , n49593 );
xor ( n49849 , n49599 , n49601 );
xor ( n49850 , n49849 , n49604 );
and ( n49851 , n49848 , n49850 );
xor ( n49852 , n49669 , n49673 );
xor ( n49853 , n49852 , n49678 );
xnor ( n49854 , n49685 , n49689 );
and ( n49855 , n49853 , n49854 );
xor ( n49856 , n49695 , n49699 );
and ( n49857 , n49854 , n49856 );
and ( n49858 , n49853 , n49856 );
or ( n49859 , n49855 , n49857 , n49858 );
and ( n49860 , n47962 , n46135 );
and ( n49861 , n47778 , n46133 );
nor ( n49862 , n49860 , n49861 );
xnor ( n49863 , n49862 , n46067 );
and ( n49864 , n48272 , n45990 );
and ( n49865 , n48108 , n45988 );
nor ( n49866 , n49864 , n49865 );
xnor ( n49867 , n49866 , n45939 );
and ( n49868 , n49863 , n49867 );
and ( n49869 , n49781 , n20852 );
and ( n49870 , n49570 , n20850 );
nor ( n49871 , n49869 , n49870 );
xnor ( n49872 , n49871 , n20860 );
and ( n49873 , n49867 , n49872 );
and ( n49874 , n49863 , n49872 );
or ( n49875 , n49868 , n49873 , n49874 );
and ( n49876 , n46577 , n47178 );
and ( n49877 , n46530 , n47176 );
nor ( n49878 , n49876 , n49877 );
xnor ( n49879 , n49878 , n47039 );
and ( n49880 , n46843 , n46911 );
and ( n49881 , n46750 , n46909 );
nor ( n49882 , n49880 , n49881 );
xnor ( n49883 , n49882 , n46802 );
and ( n49884 , n49879 , n49883 );
and ( n49885 , n47090 , n46712 );
and ( n49886 , n46969 , n46710 );
nor ( n49887 , n49885 , n49886 );
xnor ( n49888 , n49887 , n46587 );
and ( n49889 , n49883 , n49888 );
and ( n49890 , n49879 , n49888 );
or ( n49891 , n49884 , n49889 , n49890 );
and ( n49892 , n49875 , n49891 );
xor ( n49893 , n49307 , n49706 );
xor ( n49894 , n49706 , n49708 );
not ( n49895 , n49894 );
and ( n49896 , n49893 , n49895 );
and ( n49897 , n20855 , n49896 );
not ( n49898 , n49897 );
xnor ( n49899 , n49898 , n49711 );
and ( n49900 , n20864 , n49513 );
and ( n49901 , n20844 , n49511 );
nor ( n49902 , n49900 , n49901 );
xnor ( n49903 , n49902 , n49310 );
and ( n49904 , n49899 , n49903 );
and ( n49905 , n45763 , n49121 );
and ( n49906 , n45712 , n49119 );
nor ( n49907 , n49905 , n49906 );
xnor ( n49908 , n49907 , n48932 );
and ( n49909 , n49903 , n49908 );
and ( n49910 , n49899 , n49908 );
or ( n49911 , n49904 , n49909 , n49910 );
and ( n49912 , n49891 , n49911 );
and ( n49913 , n49875 , n49911 );
or ( n49914 , n49892 , n49912 , n49913 );
and ( n49915 , n49859 , n49914 );
and ( n49916 , n45843 , n48740 );
and ( n49917 , n45794 , n48738 );
nor ( n49918 , n49916 , n49917 );
xnor ( n49919 , n49918 , n48571 );
and ( n49920 , n45963 , n48394 );
and ( n49921 , n45907 , n48392 );
nor ( n49922 , n49920 , n49921 );
xnor ( n49923 , n49922 , n48220 );
and ( n49924 , n49919 , n49923 );
and ( n49925 , n46100 , n48042 );
and ( n49926 , n46041 , n48040 );
nor ( n49927 , n49925 , n49926 );
xnor ( n49928 , n49927 , n47921 );
and ( n49929 , n49923 , n49928 );
and ( n49930 , n49919 , n49928 );
or ( n49931 , n49924 , n49929 , n49930 );
and ( n49932 , n46264 , n47734 );
and ( n49933 , n46169 , n47732 );
nor ( n49934 , n49932 , n49933 );
xnor ( n49935 , n49934 , n47606 );
and ( n49936 , n46445 , n47429 );
and ( n49937 , n46345 , n47427 );
nor ( n49938 , n49936 , n49937 );
xnor ( n49939 , n49938 , n47309 );
and ( n49940 , n49935 , n49939 );
and ( n49941 , n47351 , n46496 );
and ( n49942 , n47216 , n46494 );
nor ( n49943 , n49941 , n49942 );
xnor ( n49944 , n49943 , n46402 );
and ( n49945 , n49939 , n49944 );
and ( n49946 , n49935 , n49944 );
or ( n49947 , n49940 , n49945 , n49946 );
and ( n49948 , n49931 , n49947 );
and ( n49949 , n47647 , n46306 );
and ( n49950 , n47474 , n46304 );
nor ( n49951 , n49949 , n49950 );
xnor ( n49952 , n49951 , n46228 );
and ( n49953 , n48632 , n45886 );
and ( n49954 , n48384 , n45884 );
nor ( n49955 , n49953 , n49954 );
xnor ( n49956 , n49955 , n45824 );
and ( n49957 , n49952 , n49956 );
and ( n49958 , n48988 , n45777 );
and ( n49959 , n48709 , n45775 );
nor ( n49960 , n49958 , n49959 );
xnor ( n49961 , n49960 , n45734 );
and ( n49962 , n49956 , n49961 );
and ( n49963 , n49952 , n49961 );
or ( n49964 , n49957 , n49962 , n49963 );
and ( n49965 , n49947 , n49964 );
and ( n49966 , n49931 , n49964 );
or ( n49967 , n49948 , n49965 , n49966 );
and ( n49968 , n49914 , n49967 );
and ( n49969 , n49859 , n49967 );
or ( n49970 , n49915 , n49968 , n49969 );
and ( n49971 , n49374 , n45702 );
and ( n49972 , n49115 , n45700 );
nor ( n49973 , n49971 , n49972 );
xnor ( n49974 , n49973 , n20841 );
buf ( n49975 , n20764 );
buf ( n49976 , n49975 );
and ( n49977 , n49976 , n20846 );
and ( n49978 , n49974 , n49977 );
xor ( n49979 , n25176 , n45627 );
buf ( n49980 , n49979 );
buf ( n49981 , n49980 );
buf ( n49982 , n49981 );
and ( n49983 , n49977 , n49982 );
and ( n49984 , n49974 , n49982 );
or ( n49985 , n49978 , n49983 , n49984 );
xor ( n49986 , n49712 , n49716 );
xor ( n49987 , n49986 , n49721 );
and ( n49988 , n49985 , n49987 );
xor ( n49989 , n49728 , n49732 );
xor ( n49990 , n49989 , n49737 );
and ( n49991 , n49987 , n49990 );
and ( n49992 , n49985 , n49990 );
or ( n49993 , n49988 , n49991 , n49992 );
xor ( n49994 , n49745 , n49749 );
xor ( n49995 , n49994 , n49754 );
xor ( n49996 , n49767 , n49771 );
xor ( n49997 , n49996 , n49776 );
and ( n49998 , n49995 , n49997 );
xor ( n49999 , n49782 , n49786 );
buf ( n50000 , n49999 );
and ( n50001 , n49997 , n50000 );
and ( n50002 , n49995 , n50000 );
or ( n50003 , n49998 , n50001 , n50002 );
and ( n50004 , n49993 , n50003 );
xor ( n50005 , n49657 , n49659 );
xor ( n50006 , n50005 , n49662 );
and ( n50007 , n50003 , n50006 );
and ( n50008 , n49993 , n50006 );
or ( n50009 , n50004 , n50007 , n50008 );
and ( n50010 , n49970 , n50009 );
xor ( n50011 , n49681 , n49690 );
xor ( n50012 , n50011 , n49700 );
xor ( n50013 , n49724 , n49740 );
xor ( n50014 , n50013 , n49757 );
and ( n50015 , n50012 , n50014 );
xor ( n50016 , n49779 , n49788 );
xor ( n50017 , n50016 , n49791 );
and ( n50018 , n50014 , n50017 );
and ( n50019 , n50012 , n50017 );
or ( n50020 , n50015 , n50018 , n50019 );
and ( n50021 , n50009 , n50020 );
and ( n50022 , n49970 , n50020 );
or ( n50023 , n50010 , n50021 , n50022 );
xor ( n50024 , n49645 , n49647 );
xor ( n50025 , n50024 , n49649 );
xor ( n50026 , n49665 , n49703 );
xor ( n50027 , n50026 , n49760 );
and ( n50028 , n50025 , n50027 );
xor ( n50029 , n49794 , n49804 );
xor ( n50030 , n50029 , n49807 );
and ( n50031 , n50027 , n50030 );
and ( n50032 , n50025 , n50030 );
or ( n50033 , n50028 , n50031 , n50032 );
and ( n50034 , n50023 , n50033 );
xor ( n50035 , n49640 , n49642 );
xor ( n50036 , n50035 , n49652 );
and ( n50037 , n50033 , n50036 );
and ( n50038 , n50023 , n50036 );
or ( n50039 , n50034 , n50037 , n50038 );
and ( n50040 , n49850 , n50039 );
and ( n50041 , n49848 , n50039 );
or ( n50042 , n49851 , n50040 , n50041 );
and ( n50043 , n49846 , n50042 );
xor ( n50044 , n49635 , n49637 );
xor ( n50045 , n50044 , n49838 );
and ( n50046 , n50042 , n50045 );
and ( n50047 , n49846 , n50045 );
or ( n50048 , n50043 , n50046 , n50047 );
and ( n50049 , n49843 , n50048 );
and ( n50050 , n49841 , n50048 );
or ( n50051 , n49844 , n50049 , n50050 );
and ( n50052 , n49633 , n50051 );
xor ( n50053 , n49841 , n49843 );
xor ( n50054 , n50053 , n50048 );
xor ( n50055 , n49655 , n49824 );
xor ( n50056 , n50055 , n49835 );
xor ( n50057 , n49763 , n49810 );
xor ( n50058 , n50057 , n49821 );
xor ( n50059 , n49827 , n49829 );
xor ( n50060 , n50059 , n49832 );
and ( n50061 , n50058 , n50060 );
xor ( n50062 , n49813 , n49815 );
xor ( n50063 , n50062 , n49818 );
xor ( n50064 , n49796 , n49798 );
xor ( n50065 , n50064 , n49801 );
xor ( n50066 , n49863 , n49867 );
xor ( n50067 , n50066 , n49872 );
xor ( n50068 , n49879 , n49883 );
xor ( n50069 , n50068 , n49888 );
and ( n50070 , n50067 , n50069 );
buf ( n50071 , n50070 );
and ( n50072 , n47778 , n46306 );
and ( n50073 , n47647 , n46304 );
nor ( n50074 , n50072 , n50073 );
xnor ( n50075 , n50074 , n46228 );
and ( n50076 , n48108 , n46135 );
and ( n50077 , n47962 , n46133 );
nor ( n50078 , n50076 , n50077 );
xnor ( n50079 , n50078 , n46067 );
and ( n50080 , n50075 , n50079 );
and ( n50081 , n48709 , n45886 );
and ( n50082 , n48632 , n45884 );
nor ( n50083 , n50081 , n50082 );
xnor ( n50084 , n50083 , n45824 );
and ( n50085 , n50079 , n50084 );
and ( n50086 , n50075 , n50084 );
or ( n50087 , n50080 , n50085 , n50086 );
and ( n50088 , n48384 , n45990 );
and ( n50089 , n48272 , n45988 );
nor ( n50090 , n50088 , n50089 );
xnor ( n50091 , n50090 , n45939 );
and ( n50092 , n49115 , n45777 );
and ( n50093 , n48988 , n45775 );
nor ( n50094 , n50092 , n50093 );
xnor ( n50095 , n50094 , n45734 );
and ( n50096 , n50091 , n50095 );
and ( n50097 , n49976 , n20852 );
and ( n50098 , n49781 , n20850 );
nor ( n50099 , n50097 , n50098 );
xnor ( n50100 , n50099 , n20860 );
and ( n50101 , n50095 , n50100 );
and ( n50102 , n50091 , n50100 );
or ( n50103 , n50096 , n50101 , n50102 );
and ( n50104 , n50087 , n50103 );
buf ( n50105 , n17523 );
buf ( n50106 , n50105 );
buf ( n50107 , n17525 );
buf ( n50108 , n50107 );
and ( n50109 , n50106 , n50108 );
not ( n50110 , n50109 );
and ( n50111 , n49708 , n50110 );
not ( n50112 , n50111 );
and ( n50113 , n20844 , n49896 );
and ( n50114 , n20855 , n49894 );
nor ( n50115 , n50113 , n50114 );
xnor ( n50116 , n50115 , n49711 );
and ( n50117 , n50112 , n50116 );
and ( n50118 , n45712 , n49513 );
and ( n50119 , n20864 , n49511 );
nor ( n50120 , n50118 , n50119 );
xnor ( n50121 , n50120 , n49310 );
and ( n50122 , n50116 , n50121 );
and ( n50123 , n50112 , n50121 );
or ( n50124 , n50117 , n50122 , n50123 );
and ( n50125 , n50103 , n50124 );
and ( n50126 , n50087 , n50124 );
or ( n50127 , n50104 , n50125 , n50126 );
and ( n50128 , n50071 , n50127 );
and ( n50129 , n45794 , n49121 );
and ( n50130 , n45763 , n49119 );
nor ( n50131 , n50129 , n50130 );
xnor ( n50132 , n50131 , n48932 );
and ( n50133 , n45907 , n48740 );
and ( n50134 , n45843 , n48738 );
nor ( n50135 , n50133 , n50134 );
xnor ( n50136 , n50135 , n48571 );
and ( n50137 , n50132 , n50136 );
and ( n50138 , n46041 , n48394 );
and ( n50139 , n45963 , n48392 );
nor ( n50140 , n50138 , n50139 );
xnor ( n50141 , n50140 , n48220 );
and ( n50142 , n50136 , n50141 );
and ( n50143 , n50132 , n50141 );
or ( n50144 , n50137 , n50142 , n50143 );
and ( n50145 , n46169 , n48042 );
and ( n50146 , n46100 , n48040 );
nor ( n50147 , n50145 , n50146 );
xnor ( n50148 , n50147 , n47921 );
and ( n50149 , n46345 , n47734 );
and ( n50150 , n46264 , n47732 );
nor ( n50151 , n50149 , n50150 );
xnor ( n50152 , n50151 , n47606 );
and ( n50153 , n50148 , n50152 );
and ( n50154 , n46530 , n47429 );
and ( n50155 , n46445 , n47427 );
nor ( n50156 , n50154 , n50155 );
xnor ( n50157 , n50156 , n47309 );
and ( n50158 , n50152 , n50157 );
and ( n50159 , n50148 , n50157 );
or ( n50160 , n50153 , n50158 , n50159 );
and ( n50161 , n50144 , n50160 );
and ( n50162 , n46750 , n47178 );
and ( n50163 , n46577 , n47176 );
nor ( n50164 , n50162 , n50163 );
xnor ( n50165 , n50164 , n47039 );
and ( n50166 , n46969 , n46911 );
and ( n50167 , n46843 , n46909 );
nor ( n50168 , n50166 , n50167 );
xnor ( n50169 , n50168 , n46802 );
and ( n50170 , n50165 , n50169 );
and ( n50171 , n47216 , n46712 );
and ( n50172 , n47090 , n46710 );
nor ( n50173 , n50171 , n50172 );
xnor ( n50174 , n50173 , n46587 );
and ( n50175 , n50169 , n50174 );
and ( n50176 , n50165 , n50174 );
or ( n50177 , n50170 , n50175 , n50176 );
and ( n50178 , n50160 , n50177 );
and ( n50179 , n50144 , n50177 );
or ( n50180 , n50161 , n50178 , n50179 );
and ( n50181 , n50127 , n50180 );
and ( n50182 , n50071 , n50180 );
or ( n50183 , n50128 , n50181 , n50182 );
and ( n50184 , n50065 , n50183 );
and ( n50185 , n47474 , n46496 );
and ( n50186 , n47351 , n46494 );
nor ( n50187 , n50185 , n50186 );
xnor ( n50188 , n50187 , n46402 );
and ( n50189 , n49570 , n45702 );
and ( n50190 , n49374 , n45700 );
nor ( n50191 , n50189 , n50190 );
xnor ( n50192 , n50191 , n20841 );
and ( n50193 , n50188 , n50192 );
buf ( n50194 , n20766 );
buf ( n50195 , n50194 );
and ( n50196 , n50195 , n20846 );
and ( n50197 , n50192 , n50196 );
and ( n50198 , n50188 , n50196 );
or ( n50199 , n50193 , n50197 , n50198 );
xor ( n50200 , n49899 , n49903 );
xor ( n50201 , n50200 , n49908 );
and ( n50202 , n50199 , n50201 );
xor ( n50203 , n49919 , n49923 );
xor ( n50204 , n50203 , n49928 );
and ( n50205 , n50201 , n50204 );
and ( n50206 , n50199 , n50204 );
or ( n50207 , n50202 , n50205 , n50206 );
xor ( n50208 , n49935 , n49939 );
xor ( n50209 , n50208 , n49944 );
xor ( n50210 , n49952 , n49956 );
xor ( n50211 , n50210 , n49961 );
and ( n50212 , n50209 , n50211 );
xor ( n50213 , n49974 , n49977 );
xor ( n50214 , n50213 , n49982 );
and ( n50215 , n50211 , n50214 );
and ( n50216 , n50209 , n50214 );
or ( n50217 , n50212 , n50215 , n50216 );
and ( n50218 , n50207 , n50217 );
xor ( n50219 , n49853 , n49854 );
xor ( n50220 , n50219 , n49856 );
and ( n50221 , n50217 , n50220 );
and ( n50222 , n50207 , n50220 );
or ( n50223 , n50218 , n50221 , n50222 );
and ( n50224 , n50183 , n50223 );
and ( n50225 , n50065 , n50223 );
or ( n50226 , n50184 , n50224 , n50225 );
and ( n50227 , n50063 , n50226 );
xor ( n50228 , n49875 , n49891 );
xor ( n50229 , n50228 , n49911 );
xor ( n50230 , n49931 , n49947 );
xor ( n50231 , n50230 , n49964 );
and ( n50232 , n50229 , n50231 );
xor ( n50233 , n49985 , n49987 );
xor ( n50234 , n50233 , n49990 );
and ( n50235 , n50231 , n50234 );
and ( n50236 , n50229 , n50234 );
or ( n50237 , n50232 , n50235 , n50236 );
xor ( n50238 , n49859 , n49914 );
xor ( n50239 , n50238 , n49967 );
and ( n50240 , n50237 , n50239 );
xor ( n50241 , n49993 , n50003 );
xor ( n50242 , n50241 , n50006 );
and ( n50243 , n50239 , n50242 );
and ( n50244 , n50237 , n50242 );
or ( n50245 , n50240 , n50243 , n50244 );
and ( n50246 , n50226 , n50245 );
and ( n50247 , n50063 , n50245 );
or ( n50248 , n50227 , n50246 , n50247 );
and ( n50249 , n50060 , n50248 );
and ( n50250 , n50058 , n50248 );
or ( n50251 , n50061 , n50249 , n50250 );
and ( n50252 , n50056 , n50251 );
xor ( n50253 , n49848 , n49850 );
xor ( n50254 , n50253 , n50039 );
and ( n50255 , n50251 , n50254 );
and ( n50256 , n50056 , n50254 );
or ( n50257 , n50252 , n50255 , n50256 );
xor ( n50258 , n49846 , n50042 );
xor ( n50259 , n50258 , n50045 );
and ( n50260 , n50257 , n50259 );
xor ( n50261 , n50023 , n50033 );
xor ( n50262 , n50261 , n50036 );
xor ( n50263 , n49970 , n50009 );
xor ( n50264 , n50263 , n50020 );
xor ( n50265 , n50025 , n50027 );
xor ( n50266 , n50265 , n50030 );
and ( n50267 , n50264 , n50266 );
xor ( n50268 , n50012 , n50014 );
xor ( n50269 , n50268 , n50017 );
xor ( n50270 , n49995 , n49997 );
xor ( n50271 , n50270 , n50000 );
xor ( n50272 , n25179 , n45625 );
buf ( n50273 , n50272 );
buf ( n50274 , n50273 );
buf ( n50275 , n50274 );
xor ( n50276 , n50075 , n50079 );
xor ( n50277 , n50276 , n50084 );
and ( n50278 , n50275 , n50277 );
buf ( n50279 , n50278 );
xor ( n50280 , n50091 , n50095 );
xor ( n50281 , n50280 , n50100 );
and ( n50282 , n46264 , n48042 );
and ( n50283 , n46169 , n48040 );
nor ( n50284 , n50282 , n50283 );
xnor ( n50285 , n50284 , n47921 );
and ( n50286 , n46577 , n47429 );
and ( n50287 , n46530 , n47427 );
nor ( n50288 , n50286 , n50287 );
xnor ( n50289 , n50288 , n47309 );
and ( n50290 , n50285 , n50289 );
and ( n50291 , n46843 , n47178 );
and ( n50292 , n46750 , n47176 );
nor ( n50293 , n50291 , n50292 );
xnor ( n50294 , n50293 , n47039 );
and ( n50295 , n50289 , n50294 );
and ( n50296 , n50285 , n50294 );
or ( n50297 , n50290 , n50295 , n50296 );
and ( n50298 , n50281 , n50297 );
and ( n50299 , n47962 , n46306 );
and ( n50300 , n47778 , n46304 );
nor ( n50301 , n50299 , n50300 );
xnor ( n50302 , n50301 , n46228 );
and ( n50303 , n48988 , n45886 );
and ( n50304 , n48709 , n45884 );
nor ( n50305 , n50303 , n50304 );
xnor ( n50306 , n50305 , n45824 );
and ( n50307 , n50302 , n50306 );
and ( n50308 , n49781 , n45702 );
and ( n50309 , n49570 , n45700 );
nor ( n50310 , n50308 , n50309 );
xnor ( n50311 , n50310 , n20841 );
and ( n50312 , n50306 , n50311 );
and ( n50313 , n50302 , n50311 );
or ( n50314 , n50307 , n50312 , n50313 );
and ( n50315 , n50297 , n50314 );
and ( n50316 , n50281 , n50314 );
or ( n50317 , n50298 , n50315 , n50316 );
and ( n50318 , n50279 , n50317 );
and ( n50319 , n48632 , n45990 );
and ( n50320 , n48384 , n45988 );
nor ( n50321 , n50319 , n50320 );
xnor ( n50322 , n50321 , n45939 );
and ( n50323 , n49374 , n45777 );
and ( n50324 , n49115 , n45775 );
nor ( n50325 , n50323 , n50324 );
xnor ( n50326 , n50325 , n45734 );
and ( n50327 , n50322 , n50326 );
and ( n50328 , n50195 , n20852 );
and ( n50329 , n49976 , n20850 );
nor ( n50330 , n50328 , n50329 );
xnor ( n50331 , n50330 , n20860 );
and ( n50332 , n50326 , n50331 );
and ( n50333 , n50322 , n50331 );
or ( n50334 , n50327 , n50332 , n50333 );
xor ( n50335 , n49708 , n50106 );
xor ( n50336 , n50106 , n50108 );
not ( n50337 , n50336 );
and ( n50338 , n50335 , n50337 );
and ( n50339 , n20855 , n50338 );
not ( n50340 , n50339 );
xnor ( n50341 , n50340 , n50111 );
and ( n50342 , n20864 , n49896 );
and ( n50343 , n20844 , n49894 );
nor ( n50344 , n50342 , n50343 );
xnor ( n50345 , n50344 , n49711 );
and ( n50346 , n50341 , n50345 );
and ( n50347 , n45763 , n49513 );
and ( n50348 , n45712 , n49511 );
nor ( n50349 , n50347 , n50348 );
xnor ( n50350 , n50349 , n49310 );
and ( n50351 , n50345 , n50350 );
and ( n50352 , n50341 , n50350 );
or ( n50353 , n50346 , n50351 , n50352 );
and ( n50354 , n50334 , n50353 );
and ( n50355 , n45843 , n49121 );
and ( n50356 , n45794 , n49119 );
nor ( n50357 , n50355 , n50356 );
xnor ( n50358 , n50357 , n48932 );
and ( n50359 , n45963 , n48740 );
and ( n50360 , n45907 , n48738 );
nor ( n50361 , n50359 , n50360 );
xnor ( n50362 , n50361 , n48571 );
and ( n50363 , n50358 , n50362 );
and ( n50364 , n46100 , n48394 );
and ( n50365 , n46041 , n48392 );
nor ( n50366 , n50364 , n50365 );
xnor ( n50367 , n50366 , n48220 );
and ( n50368 , n50362 , n50367 );
and ( n50369 , n50358 , n50367 );
or ( n50370 , n50363 , n50368 , n50369 );
and ( n50371 , n50353 , n50370 );
and ( n50372 , n50334 , n50370 );
or ( n50373 , n50354 , n50371 , n50372 );
and ( n50374 , n50317 , n50373 );
and ( n50375 , n50279 , n50373 );
or ( n50376 , n50318 , n50374 , n50375 );
and ( n50377 , n50271 , n50376 );
and ( n50378 , n46445 , n47734 );
and ( n50379 , n46345 , n47732 );
nor ( n50380 , n50378 , n50379 );
xnor ( n50381 , n50380 , n47606 );
and ( n50382 , n47090 , n46911 );
and ( n50383 , n46969 , n46909 );
nor ( n50384 , n50382 , n50383 );
xnor ( n50385 , n50384 , n46802 );
and ( n50386 , n50381 , n50385 );
and ( n50387 , n47351 , n46712 );
and ( n50388 , n47216 , n46710 );
nor ( n50389 , n50387 , n50388 );
xnor ( n50390 , n50389 , n46587 );
and ( n50391 , n50385 , n50390 );
and ( n50392 , n50381 , n50390 );
or ( n50393 , n50386 , n50391 , n50392 );
and ( n50394 , n47647 , n46496 );
and ( n50395 , n47474 , n46494 );
nor ( n50396 , n50394 , n50395 );
xnor ( n50397 , n50396 , n46402 );
and ( n50398 , n48272 , n46135 );
and ( n50399 , n48108 , n46133 );
nor ( n50400 , n50398 , n50399 );
xnor ( n50401 , n50400 , n46067 );
and ( n50402 , n50397 , n50401 );
buf ( n50403 , n20768 );
buf ( n50404 , n50403 );
and ( n50405 , n50404 , n20846 );
and ( n50406 , n50401 , n50405 );
and ( n50407 , n50397 , n50405 );
or ( n50408 , n50402 , n50406 , n50407 );
and ( n50409 , n50393 , n50408 );
xor ( n50410 , n50112 , n50116 );
xor ( n50411 , n50410 , n50121 );
and ( n50412 , n50408 , n50411 );
and ( n50413 , n50393 , n50411 );
or ( n50414 , n50409 , n50412 , n50413 );
xor ( n50415 , n50132 , n50136 );
xor ( n50416 , n50415 , n50141 );
xor ( n50417 , n50148 , n50152 );
xor ( n50418 , n50417 , n50157 );
and ( n50419 , n50416 , n50418 );
xor ( n50420 , n50165 , n50169 );
xor ( n50421 , n50420 , n50174 );
and ( n50422 , n50418 , n50421 );
and ( n50423 , n50416 , n50421 );
or ( n50424 , n50419 , n50422 , n50423 );
and ( n50425 , n50414 , n50424 );
buf ( n50426 , n50067 );
xor ( n50427 , n50426 , n50069 );
and ( n50428 , n50424 , n50427 );
and ( n50429 , n50414 , n50427 );
or ( n50430 , n50425 , n50428 , n50429 );
and ( n50431 , n50376 , n50430 );
and ( n50432 , n50271 , n50430 );
or ( n50433 , n50377 , n50431 , n50432 );
and ( n50434 , n50269 , n50433 );
xor ( n50435 , n50087 , n50103 );
xor ( n50436 , n50435 , n50124 );
xor ( n50437 , n50144 , n50160 );
xor ( n50438 , n50437 , n50177 );
and ( n50439 , n50436 , n50438 );
xor ( n50440 , n50199 , n50201 );
xor ( n50441 , n50440 , n50204 );
and ( n50442 , n50438 , n50441 );
and ( n50443 , n50436 , n50441 );
or ( n50444 , n50439 , n50442 , n50443 );
xor ( n50445 , n50071 , n50127 );
xor ( n50446 , n50445 , n50180 );
and ( n50447 , n50444 , n50446 );
xor ( n50448 , n50207 , n50217 );
xor ( n50449 , n50448 , n50220 );
and ( n50450 , n50446 , n50449 );
and ( n50451 , n50444 , n50449 );
or ( n50452 , n50447 , n50450 , n50451 );
and ( n50453 , n50433 , n50452 );
and ( n50454 , n50269 , n50452 );
or ( n50455 , n50434 , n50453 , n50454 );
and ( n50456 , n50266 , n50455 );
and ( n50457 , n50264 , n50455 );
or ( n50458 , n50267 , n50456 , n50457 );
and ( n50459 , n50262 , n50458 );
xor ( n50460 , n50058 , n50060 );
xor ( n50461 , n50460 , n50248 );
and ( n50462 , n50458 , n50461 );
and ( n50463 , n50262 , n50461 );
or ( n50464 , n50459 , n50462 , n50463 );
xor ( n50465 , n50056 , n50251 );
xor ( n50466 , n50465 , n50254 );
and ( n50467 , n50464 , n50466 );
xor ( n50468 , n50063 , n50226 );
xor ( n50469 , n50468 , n50245 );
xor ( n50470 , n50065 , n50183 );
xor ( n50471 , n50470 , n50223 );
xor ( n50472 , n50237 , n50239 );
xor ( n50473 , n50472 , n50242 );
and ( n50474 , n50471 , n50473 );
xor ( n50475 , n50229 , n50231 );
xor ( n50476 , n50475 , n50234 );
xor ( n50477 , n50209 , n50211 );
xor ( n50478 , n50477 , n50214 );
xor ( n50479 , n50188 , n50192 );
xor ( n50480 , n50479 , n50196 );
xor ( n50481 , n50302 , n50306 );
xor ( n50482 , n50481 , n50311 );
xor ( n50483 , n50322 , n50326 );
xor ( n50484 , n50483 , n50331 );
and ( n50485 , n50482 , n50484 );
and ( n50486 , n50480 , n50485 );
xor ( n50487 , n25180 , n45624 );
buf ( n50488 , n50487 );
buf ( n50489 , n50488 );
buf ( n50490 , n50489 );
xor ( n50491 , n50285 , n50289 );
xor ( n50492 , n50491 , n50294 );
and ( n50493 , n50490 , n50492 );
buf ( n50494 , n50493 );
and ( n50495 , n50485 , n50494 );
and ( n50496 , n50480 , n50494 );
or ( n50497 , n50486 , n50495 , n50496 );
and ( n50498 , n50478 , n50497 );
and ( n50499 , n46345 , n48042 );
and ( n50500 , n46264 , n48040 );
nor ( n50501 , n50499 , n50500 );
xnor ( n50502 , n50501 , n47921 );
and ( n50503 , n46530 , n47734 );
and ( n50504 , n46445 , n47732 );
nor ( n50505 , n50503 , n50504 );
xnor ( n50506 , n50505 , n47606 );
and ( n50507 , n50502 , n50506 );
and ( n50508 , n46750 , n47429 );
and ( n50509 , n46577 , n47427 );
nor ( n50510 , n50508 , n50509 );
xnor ( n50511 , n50510 , n47309 );
and ( n50512 , n50506 , n50511 );
and ( n50513 , n50502 , n50511 );
or ( n50514 , n50507 , n50512 , n50513 );
and ( n50515 , n49115 , n45886 );
and ( n50516 , n48988 , n45884 );
nor ( n50517 , n50515 , n50516 );
xnor ( n50518 , n50517 , n45824 );
and ( n50519 , n49570 , n45777 );
and ( n50520 , n49374 , n45775 );
nor ( n50521 , n50519 , n50520 );
xnor ( n50522 , n50521 , n45734 );
and ( n50523 , n50518 , n50522 );
and ( n50524 , n50404 , n20852 );
and ( n50525 , n50195 , n20850 );
nor ( n50526 , n50524 , n50525 );
xnor ( n50527 , n50526 , n20860 );
and ( n50528 , n50522 , n50527 );
and ( n50529 , n50518 , n50527 );
or ( n50530 , n50523 , n50528 , n50529 );
and ( n50531 , n50514 , n50530 );
and ( n50532 , n48384 , n46135 );
and ( n50533 , n48272 , n46133 );
nor ( n50534 , n50532 , n50533 );
xnor ( n50535 , n50534 , n46067 );
and ( n50536 , n48709 , n45990 );
and ( n50537 , n48632 , n45988 );
nor ( n50538 , n50536 , n50537 );
xnor ( n50539 , n50538 , n45939 );
and ( n50540 , n50535 , n50539 );
and ( n50541 , n49976 , n45702 );
and ( n50542 , n49781 , n45700 );
nor ( n50543 , n50541 , n50542 );
xnor ( n50544 , n50543 , n20841 );
and ( n50545 , n50539 , n50544 );
and ( n50546 , n50535 , n50544 );
or ( n50547 , n50540 , n50545 , n50546 );
and ( n50548 , n50530 , n50547 );
and ( n50549 , n50514 , n50547 );
or ( n50550 , n50531 , n50548 , n50549 );
buf ( n50551 , n17527 );
buf ( n50552 , n50551 );
buf ( n50553 , n17529 );
buf ( n50554 , n50553 );
and ( n50555 , n50552 , n50554 );
not ( n50556 , n50555 );
and ( n50557 , n50108 , n50556 );
not ( n50558 , n50557 );
and ( n50559 , n20844 , n50338 );
and ( n50560 , n20855 , n50336 );
nor ( n50561 , n50559 , n50560 );
xnor ( n50562 , n50561 , n50111 );
and ( n50563 , n50558 , n50562 );
and ( n50564 , n45712 , n49896 );
and ( n50565 , n20864 , n49894 );
nor ( n50566 , n50564 , n50565 );
xnor ( n50567 , n50566 , n49711 );
and ( n50568 , n50562 , n50567 );
and ( n50569 , n50558 , n50567 );
or ( n50570 , n50563 , n50568 , n50569 );
and ( n50571 , n45794 , n49513 );
and ( n50572 , n45763 , n49511 );
nor ( n50573 , n50571 , n50572 );
xnor ( n50574 , n50573 , n49310 );
and ( n50575 , n45907 , n49121 );
and ( n50576 , n45843 , n49119 );
nor ( n50577 , n50575 , n50576 );
xnor ( n50578 , n50577 , n48932 );
and ( n50579 , n50574 , n50578 );
and ( n50580 , n46041 , n48740 );
and ( n50581 , n45963 , n48738 );
nor ( n50582 , n50580 , n50581 );
xnor ( n50583 , n50582 , n48571 );
and ( n50584 , n50578 , n50583 );
and ( n50585 , n50574 , n50583 );
or ( n50586 , n50579 , n50584 , n50585 );
and ( n50587 , n50570 , n50586 );
and ( n50588 , n46169 , n48394 );
and ( n50589 , n46100 , n48392 );
nor ( n50590 , n50588 , n50589 );
xnor ( n50591 , n50590 , n48220 );
and ( n50592 , n46969 , n47178 );
and ( n50593 , n46843 , n47176 );
nor ( n50594 , n50592 , n50593 );
xnor ( n50595 , n50594 , n47039 );
and ( n50596 , n50591 , n50595 );
and ( n50597 , n47216 , n46911 );
and ( n50598 , n47090 , n46909 );
nor ( n50599 , n50597 , n50598 );
xnor ( n50600 , n50599 , n46802 );
and ( n50601 , n50595 , n50600 );
and ( n50602 , n50591 , n50600 );
or ( n50603 , n50596 , n50601 , n50602 );
and ( n50604 , n50586 , n50603 );
and ( n50605 , n50570 , n50603 );
or ( n50606 , n50587 , n50604 , n50605 );
and ( n50607 , n50550 , n50606 );
and ( n50608 , n47474 , n46712 );
and ( n50609 , n47351 , n46710 );
nor ( n50610 , n50608 , n50609 );
xnor ( n50611 , n50610 , n46587 );
and ( n50612 , n47778 , n46496 );
and ( n50613 , n47647 , n46494 );
nor ( n50614 , n50612 , n50613 );
xnor ( n50615 , n50614 , n46402 );
and ( n50616 , n50611 , n50615 );
and ( n50617 , n48108 , n46306 );
and ( n50618 , n47962 , n46304 );
nor ( n50619 , n50617 , n50618 );
xnor ( n50620 , n50619 , n46228 );
and ( n50621 , n50615 , n50620 );
and ( n50622 , n50611 , n50620 );
or ( n50623 , n50616 , n50621 , n50622 );
buf ( n50624 , n20770 );
buf ( n50625 , n50624 );
and ( n50626 , n50625 , n20846 );
xor ( n50627 , n25181 , n45623 );
buf ( n50628 , n50627 );
buf ( n50629 , n50628 );
buf ( n50630 , n50629 );
and ( n50631 , n50626 , n50630 );
buf ( n50632 , n50631 );
and ( n50633 , n50623 , n50632 );
xor ( n50634 , n50341 , n50345 );
xor ( n50635 , n50634 , n50350 );
and ( n50636 , n50632 , n50635 );
and ( n50637 , n50623 , n50635 );
or ( n50638 , n50633 , n50636 , n50637 );
and ( n50639 , n50606 , n50638 );
and ( n50640 , n50550 , n50638 );
or ( n50641 , n50607 , n50639 , n50640 );
and ( n50642 , n50497 , n50641 );
and ( n50643 , n50478 , n50641 );
or ( n50644 , n50498 , n50642 , n50643 );
and ( n50645 , n50476 , n50644 );
xor ( n50646 , n50358 , n50362 );
xor ( n50647 , n50646 , n50367 );
xor ( n50648 , n50381 , n50385 );
xor ( n50649 , n50648 , n50390 );
and ( n50650 , n50647 , n50649 );
xor ( n50651 , n50397 , n50401 );
xor ( n50652 , n50651 , n50405 );
and ( n50653 , n50649 , n50652 );
and ( n50654 , n50647 , n50652 );
or ( n50655 , n50650 , n50653 , n50654 );
buf ( n50656 , n50275 );
xor ( n50657 , n50656 , n50277 );
and ( n50658 , n50655 , n50657 );
xor ( n50659 , n50281 , n50297 );
xor ( n50660 , n50659 , n50314 );
and ( n50661 , n50657 , n50660 );
and ( n50662 , n50655 , n50660 );
or ( n50663 , n50658 , n50661 , n50662 );
xor ( n50664 , n50334 , n50353 );
xor ( n50665 , n50664 , n50370 );
xor ( n50666 , n50393 , n50408 );
xor ( n50667 , n50666 , n50411 );
and ( n50668 , n50665 , n50667 );
xor ( n50669 , n50416 , n50418 );
xor ( n50670 , n50669 , n50421 );
and ( n50671 , n50667 , n50670 );
and ( n50672 , n50665 , n50670 );
or ( n50673 , n50668 , n50671 , n50672 );
and ( n50674 , n50663 , n50673 );
xor ( n50675 , n50279 , n50317 );
xor ( n50676 , n50675 , n50373 );
and ( n50677 , n50673 , n50676 );
and ( n50678 , n50663 , n50676 );
or ( n50679 , n50674 , n50677 , n50678 );
and ( n50680 , n50644 , n50679 );
and ( n50681 , n50476 , n50679 );
or ( n50682 , n50645 , n50680 , n50681 );
and ( n50683 , n50473 , n50682 );
and ( n50684 , n50471 , n50682 );
or ( n50685 , n50474 , n50683 , n50684 );
and ( n50686 , n50469 , n50685 );
xor ( n50687 , n50264 , n50266 );
xor ( n50688 , n50687 , n50455 );
and ( n50689 , n50685 , n50688 );
and ( n50690 , n50469 , n50688 );
or ( n50691 , n50686 , n50689 , n50690 );
xor ( n50692 , n50262 , n50458 );
xor ( n50693 , n50692 , n50461 );
and ( n50694 , n50691 , n50693 );
xor ( n50695 , n50269 , n50433 );
xor ( n50696 , n50695 , n50452 );
xor ( n50697 , n50271 , n50376 );
xor ( n50698 , n50697 , n50430 );
xor ( n50699 , n50444 , n50446 );
xor ( n50700 , n50699 , n50449 );
and ( n50701 , n50698 , n50700 );
xor ( n50702 , n50414 , n50424 );
xor ( n50703 , n50702 , n50427 );
xor ( n50704 , n50436 , n50438 );
xor ( n50705 , n50704 , n50441 );
and ( n50706 , n50703 , n50705 );
xor ( n50707 , n50482 , n50484 );
xor ( n50708 , n50518 , n50522 );
xor ( n50709 , n50708 , n50527 );
xor ( n50710 , n50535 , n50539 );
xor ( n50711 , n50710 , n50544 );
or ( n50712 , n50709 , n50711 );
and ( n50713 , n50707 , n50712 );
xor ( n50714 , n50502 , n50506 );
xor ( n50715 , n50714 , n50511 );
and ( n50716 , n46264 , n48394 );
and ( n50717 , n46169 , n48392 );
nor ( n50718 , n50716 , n50717 );
xnor ( n50719 , n50718 , n48220 );
and ( n50720 , n47351 , n46911 );
and ( n50721 , n47216 , n46909 );
nor ( n50722 , n50720 , n50721 );
xnor ( n50723 , n50722 , n46802 );
and ( n50724 , n50719 , n50723 );
buf ( n50725 , n20772 );
buf ( n50726 , n50725 );
and ( n50727 , n50726 , n20846 );
and ( n50728 , n50723 , n50727 );
and ( n50729 , n50719 , n50727 );
or ( n50730 , n50724 , n50728 , n50729 );
and ( n50731 , n50715 , n50730 );
and ( n50732 , n49374 , n45886 );
and ( n50733 , n49115 , n45884 );
nor ( n50734 , n50732 , n50733 );
xnor ( n50735 , n50734 , n45824 );
and ( n50736 , n49781 , n45777 );
and ( n50737 , n49570 , n45775 );
nor ( n50738 , n50736 , n50737 );
xnor ( n50739 , n50738 , n45734 );
and ( n50740 , n50735 , n50739 );
and ( n50741 , n50625 , n20852 );
and ( n50742 , n50404 , n20850 );
nor ( n50743 , n50741 , n50742 );
xnor ( n50744 , n50743 , n20860 );
and ( n50745 , n50739 , n50744 );
and ( n50746 , n50735 , n50744 );
or ( n50747 , n50740 , n50745 , n50746 );
and ( n50748 , n50730 , n50747 );
and ( n50749 , n50715 , n50747 );
or ( n50750 , n50731 , n50748 , n50749 );
and ( n50751 , n50712 , n50750 );
and ( n50752 , n50707 , n50750 );
or ( n50753 , n50713 , n50751 , n50752 );
and ( n50754 , n48272 , n46306 );
and ( n50755 , n48108 , n46304 );
nor ( n50756 , n50754 , n50755 );
xnor ( n50757 , n50756 , n46228 );
and ( n50758 , n48632 , n46135 );
and ( n50759 , n48384 , n46133 );
nor ( n50760 , n50758 , n50759 );
xnor ( n50761 , n50760 , n46067 );
and ( n50762 , n50757 , n50761 );
and ( n50763 , n48988 , n45990 );
and ( n50764 , n48709 , n45988 );
nor ( n50765 , n50763 , n50764 );
xnor ( n50766 , n50765 , n45939 );
and ( n50767 , n50761 , n50766 );
and ( n50768 , n50757 , n50766 );
or ( n50769 , n50762 , n50767 , n50768 );
and ( n50770 , n46843 , n47429 );
and ( n50771 , n46750 , n47427 );
nor ( n50772 , n50770 , n50771 );
xnor ( n50773 , n50772 , n47309 );
and ( n50774 , n47090 , n47178 );
and ( n50775 , n46969 , n47176 );
nor ( n50776 , n50774 , n50775 );
xnor ( n50777 , n50776 , n47039 );
or ( n50778 , n50773 , n50777 );
and ( n50779 , n50769 , n50778 );
xor ( n50780 , n50108 , n50552 );
xor ( n50781 , n50552 , n50554 );
not ( n50782 , n50781 );
and ( n50783 , n50780 , n50782 );
and ( n50784 , n20855 , n50783 );
not ( n50785 , n50784 );
xnor ( n50786 , n50785 , n50557 );
and ( n50787 , n20864 , n50338 );
and ( n50788 , n20844 , n50336 );
nor ( n50789 , n50787 , n50788 );
xnor ( n50790 , n50789 , n50111 );
and ( n50791 , n50786 , n50790 );
and ( n50792 , n45763 , n49896 );
and ( n50793 , n45712 , n49894 );
nor ( n50794 , n50792 , n50793 );
xnor ( n50795 , n50794 , n49711 );
and ( n50796 , n50790 , n50795 );
and ( n50797 , n50786 , n50795 );
or ( n50798 , n50791 , n50796 , n50797 );
and ( n50799 , n50778 , n50798 );
and ( n50800 , n50769 , n50798 );
or ( n50801 , n50779 , n50799 , n50800 );
and ( n50802 , n45843 , n49513 );
and ( n50803 , n45794 , n49511 );
nor ( n50804 , n50802 , n50803 );
xnor ( n50805 , n50804 , n49310 );
and ( n50806 , n45963 , n49121 );
and ( n50807 , n45907 , n49119 );
nor ( n50808 , n50806 , n50807 );
xnor ( n50809 , n50808 , n48932 );
and ( n50810 , n50805 , n50809 );
and ( n50811 , n46100 , n48740 );
and ( n50812 , n46041 , n48738 );
nor ( n50813 , n50811 , n50812 );
xnor ( n50814 , n50813 , n48571 );
and ( n50815 , n50809 , n50814 );
and ( n50816 , n50805 , n50814 );
or ( n50817 , n50810 , n50815 , n50816 );
and ( n50818 , n46445 , n48042 );
and ( n50819 , n46345 , n48040 );
nor ( n50820 , n50818 , n50819 );
xnor ( n50821 , n50820 , n47921 );
and ( n50822 , n46577 , n47734 );
and ( n50823 , n46530 , n47732 );
nor ( n50824 , n50822 , n50823 );
xnor ( n50825 , n50824 , n47606 );
and ( n50826 , n50821 , n50825 );
and ( n50827 , n47647 , n46712 );
and ( n50828 , n47474 , n46710 );
nor ( n50829 , n50827 , n50828 );
xnor ( n50830 , n50829 , n46587 );
and ( n50831 , n50825 , n50830 );
and ( n50832 , n50821 , n50830 );
or ( n50833 , n50826 , n50831 , n50832 );
and ( n50834 , n50817 , n50833 );
and ( n50835 , n47962 , n46496 );
and ( n50836 , n47778 , n46494 );
nor ( n50837 , n50835 , n50836 );
xnor ( n50838 , n50837 , n46402 );
and ( n50839 , n50195 , n45702 );
and ( n50840 , n49976 , n45700 );
nor ( n50841 , n50839 , n50840 );
xnor ( n50842 , n50841 , n20841 );
and ( n50843 , n50838 , n50842 );
xor ( n50844 , n25436 , n45621 );
buf ( n50845 , n50844 );
buf ( n50846 , n50845 );
buf ( n50847 , n50846 );
and ( n50848 , n50842 , n50847 );
and ( n50849 , n50838 , n50847 );
or ( n50850 , n50843 , n50848 , n50849 );
and ( n50851 , n50833 , n50850 );
and ( n50852 , n50817 , n50850 );
or ( n50853 , n50834 , n50851 , n50852 );
and ( n50854 , n50801 , n50853 );
xor ( n50855 , n50558 , n50562 );
xor ( n50856 , n50855 , n50567 );
xor ( n50857 , n50574 , n50578 );
xor ( n50858 , n50857 , n50583 );
and ( n50859 , n50856 , n50858 );
xor ( n50860 , n50591 , n50595 );
xor ( n50861 , n50860 , n50600 );
and ( n50862 , n50858 , n50861 );
and ( n50863 , n50856 , n50861 );
or ( n50864 , n50859 , n50862 , n50863 );
and ( n50865 , n50853 , n50864 );
and ( n50866 , n50801 , n50864 );
or ( n50867 , n50854 , n50865 , n50866 );
and ( n50868 , n50753 , n50867 );
buf ( n50869 , n50490 );
xor ( n50870 , n50869 , n50492 );
xor ( n50871 , n50514 , n50530 );
xor ( n50872 , n50871 , n50547 );
and ( n50873 , n50870 , n50872 );
xor ( n50874 , n50570 , n50586 );
xor ( n50875 , n50874 , n50603 );
and ( n50876 , n50872 , n50875 );
and ( n50877 , n50870 , n50875 );
or ( n50878 , n50873 , n50876 , n50877 );
and ( n50879 , n50867 , n50878 );
and ( n50880 , n50753 , n50878 );
or ( n50881 , n50868 , n50879 , n50880 );
and ( n50882 , n50705 , n50881 );
and ( n50883 , n50703 , n50881 );
or ( n50884 , n50706 , n50882 , n50883 );
and ( n50885 , n50700 , n50884 );
and ( n50886 , n50698 , n50884 );
or ( n50887 , n50701 , n50885 , n50886 );
and ( n50888 , n50696 , n50887 );
xor ( n50889 , n50471 , n50473 );
xor ( n50890 , n50889 , n50682 );
and ( n50891 , n50887 , n50890 );
and ( n50892 , n50696 , n50890 );
or ( n50893 , n50888 , n50891 , n50892 );
xor ( n50894 , n50469 , n50685 );
xor ( n50895 , n50894 , n50688 );
and ( n50896 , n50893 , n50895 );
xor ( n50897 , n50480 , n50485 );
xor ( n50898 , n50897 , n50494 );
xor ( n50899 , n50550 , n50606 );
xor ( n50900 , n50899 , n50638 );
and ( n50901 , n50898 , n50900 );
xor ( n50902 , n50655 , n50657 );
xor ( n50903 , n50902 , n50660 );
and ( n50904 , n50900 , n50903 );
and ( n50905 , n50898 , n50903 );
or ( n50906 , n50901 , n50904 , n50905 );
xor ( n50907 , n50478 , n50497 );
xor ( n50908 , n50907 , n50641 );
and ( n50909 , n50906 , n50908 );
xor ( n50910 , n50663 , n50673 );
xor ( n50911 , n50910 , n50676 );
and ( n50912 , n50908 , n50911 );
and ( n50913 , n50906 , n50911 );
or ( n50914 , n50909 , n50912 , n50913 );
xor ( n50915 , n50476 , n50644 );
xor ( n50916 , n50915 , n50679 );
and ( n50917 , n50914 , n50916 );
xor ( n50918 , n50665 , n50667 );
xor ( n50919 , n50918 , n50670 );
xor ( n50920 , n50623 , n50632 );
xor ( n50921 , n50920 , n50635 );
xor ( n50922 , n50647 , n50649 );
xor ( n50923 , n50922 , n50652 );
and ( n50924 , n50921 , n50923 );
xor ( n50925 , n50611 , n50615 );
xor ( n50926 , n50925 , n50620 );
xor ( n50927 , n50626 , n50630 );
buf ( n50928 , n50927 );
and ( n50929 , n50926 , n50928 );
xnor ( n50930 , n50709 , n50711 );
and ( n50931 , n50928 , n50930 );
and ( n50932 , n50926 , n50930 );
or ( n50933 , n50929 , n50931 , n50932 );
and ( n50934 , n50923 , n50933 );
and ( n50935 , n50921 , n50933 );
or ( n50936 , n50924 , n50934 , n50935 );
and ( n50937 , n50919 , n50936 );
xor ( n50938 , n50719 , n50723 );
xor ( n50939 , n50938 , n50727 );
xor ( n50940 , n50735 , n50739 );
xor ( n50941 , n50940 , n50744 );
and ( n50942 , n50939 , n50941 );
buf ( n50943 , n50942 );
xor ( n50944 , n50757 , n50761 );
xor ( n50945 , n50944 , n50766 );
xnor ( n50946 , n50773 , n50777 );
and ( n50947 , n50945 , n50946 );
and ( n50948 , n46345 , n48394 );
and ( n50949 , n46264 , n48392 );
nor ( n50950 , n50948 , n50949 );
xnor ( n50951 , n50950 , n48220 );
and ( n50952 , n46530 , n48042 );
and ( n50953 , n46445 , n48040 );
nor ( n50954 , n50952 , n50953 );
xnor ( n50955 , n50954 , n47921 );
and ( n50956 , n50951 , n50955 );
and ( n50957 , n47474 , n46911 );
and ( n50958 , n47351 , n46909 );
nor ( n50959 , n50957 , n50958 );
xnor ( n50960 , n50959 , n46802 );
and ( n50961 , n50955 , n50960 );
and ( n50962 , n50951 , n50960 );
or ( n50963 , n50956 , n50961 , n50962 );
and ( n50964 , n50946 , n50963 );
and ( n50965 , n50945 , n50963 );
or ( n50966 , n50947 , n50964 , n50965 );
and ( n50967 , n50943 , n50966 );
and ( n50968 , n48709 , n46135 );
and ( n50969 , n48632 , n46133 );
nor ( n50970 , n50968 , n50969 );
xnor ( n50971 , n50970 , n46067 );
and ( n50972 , n49976 , n45777 );
and ( n50973 , n49781 , n45775 );
nor ( n50974 , n50972 , n50973 );
xnor ( n50975 , n50974 , n45734 );
and ( n50976 , n50971 , n50975 );
and ( n50977 , n50404 , n45702 );
and ( n50978 , n50195 , n45700 );
nor ( n50979 , n50977 , n50978 );
xnor ( n50980 , n50979 , n20841 );
and ( n50981 , n50975 , n50980 );
and ( n50982 , n50971 , n50980 );
or ( n50983 , n50976 , n50981 , n50982 );
and ( n50984 , n48384 , n46306 );
and ( n50985 , n48272 , n46304 );
nor ( n50986 , n50984 , n50985 );
xnor ( n50987 , n50986 , n46228 );
and ( n50988 , n49115 , n45990 );
and ( n50989 , n48988 , n45988 );
nor ( n50990 , n50988 , n50989 );
xnor ( n50991 , n50990 , n45939 );
or ( n50992 , n50987 , n50991 );
and ( n50993 , n50983 , n50992 );
buf ( n50994 , n17531 );
buf ( n50995 , n50994 );
buf ( n50996 , n17533 );
buf ( n50997 , n50996 );
and ( n50998 , n50995 , n50997 );
not ( n50999 , n50998 );
and ( n51000 , n50554 , n50999 );
not ( n51001 , n51000 );
and ( n51002 , n20844 , n50783 );
and ( n51003 , n20855 , n50781 );
nor ( n51004 , n51002 , n51003 );
xnor ( n51005 , n51004 , n50557 );
and ( n51006 , n51001 , n51005 );
and ( n51007 , n45712 , n50338 );
and ( n51008 , n20864 , n50336 );
nor ( n51009 , n51007 , n51008 );
xnor ( n51010 , n51009 , n50111 );
and ( n51011 , n51005 , n51010 );
and ( n51012 , n51001 , n51010 );
or ( n51013 , n51006 , n51011 , n51012 );
and ( n51014 , n50992 , n51013 );
and ( n51015 , n50983 , n51013 );
or ( n51016 , n50993 , n51014 , n51015 );
and ( n51017 , n50966 , n51016 );
and ( n51018 , n50943 , n51016 );
or ( n51019 , n50967 , n51017 , n51018 );
and ( n51020 , n45794 , n49896 );
and ( n51021 , n45763 , n49894 );
nor ( n51022 , n51020 , n51021 );
xnor ( n51023 , n51022 , n49711 );
and ( n51024 , n45907 , n49513 );
and ( n51025 , n45843 , n49511 );
nor ( n51026 , n51024 , n51025 );
xnor ( n51027 , n51026 , n49310 );
and ( n51028 , n51023 , n51027 );
and ( n51029 , n46041 , n49121 );
and ( n51030 , n45963 , n49119 );
nor ( n51031 , n51029 , n51030 );
xnor ( n51032 , n51031 , n48932 );
and ( n51033 , n51027 , n51032 );
and ( n51034 , n51023 , n51032 );
or ( n51035 , n51028 , n51033 , n51034 );
and ( n51036 , n46169 , n48740 );
and ( n51037 , n46100 , n48738 );
nor ( n51038 , n51036 , n51037 );
xnor ( n51039 , n51038 , n48571 );
and ( n51040 , n46750 , n47734 );
and ( n51041 , n46577 , n47732 );
nor ( n51042 , n51040 , n51041 );
xnor ( n51043 , n51042 , n47606 );
and ( n51044 , n51039 , n51043 );
and ( n51045 , n46969 , n47429 );
and ( n51046 , n46843 , n47427 );
nor ( n51047 , n51045 , n51046 );
xnor ( n51048 , n51047 , n47309 );
and ( n51049 , n51043 , n51048 );
and ( n51050 , n51039 , n51048 );
or ( n51051 , n51044 , n51049 , n51050 );
and ( n51052 , n51035 , n51051 );
and ( n51053 , n47216 , n47178 );
and ( n51054 , n47090 , n47176 );
nor ( n51055 , n51053 , n51054 );
xnor ( n51056 , n51055 , n47039 );
and ( n51057 , n47778 , n46712 );
and ( n51058 , n47647 , n46710 );
nor ( n51059 , n51057 , n51058 );
xnor ( n51060 , n51059 , n46587 );
and ( n51061 , n51056 , n51060 );
and ( n51062 , n48108 , n46496 );
and ( n51063 , n47962 , n46494 );
nor ( n51064 , n51062 , n51063 );
xnor ( n51065 , n51064 , n46402 );
and ( n51066 , n51060 , n51065 );
and ( n51067 , n51056 , n51065 );
or ( n51068 , n51061 , n51066 , n51067 );
and ( n51069 , n51051 , n51068 );
and ( n51070 , n51035 , n51068 );
or ( n51071 , n51052 , n51069 , n51070 );
and ( n51072 , n50726 , n20852 );
and ( n51073 , n50625 , n20850 );
nor ( n51074 , n51072 , n51073 );
xnor ( n51075 , n51074 , n20860 );
buf ( n51076 , n20774 );
buf ( n51077 , n51076 );
and ( n51078 , n51077 , n20846 );
and ( n51079 , n51075 , n51078 );
xor ( n51080 , n26007 , n45619 );
buf ( n51081 , n51080 );
buf ( n51082 , n51081 );
buf ( n51083 , n51082 );
and ( n51084 , n51078 , n51083 );
and ( n51085 , n51075 , n51083 );
or ( n51086 , n51079 , n51084 , n51085 );
xor ( n51087 , n50786 , n50790 );
xor ( n51088 , n51087 , n50795 );
and ( n51089 , n51086 , n51088 );
xor ( n51090 , n50805 , n50809 );
xor ( n51091 , n51090 , n50814 );
and ( n51092 , n51088 , n51091 );
and ( n51093 , n51086 , n51091 );
or ( n51094 , n51089 , n51092 , n51093 );
and ( n51095 , n51071 , n51094 );
xor ( n51096 , n50715 , n50730 );
xor ( n51097 , n51096 , n50747 );
and ( n51098 , n51094 , n51097 );
and ( n51099 , n51071 , n51097 );
or ( n51100 , n51095 , n51098 , n51099 );
and ( n51101 , n51019 , n51100 );
xor ( n51102 , n50769 , n50778 );
xor ( n51103 , n51102 , n50798 );
xor ( n51104 , n50817 , n50833 );
xor ( n51105 , n51104 , n50850 );
and ( n51106 , n51103 , n51105 );
xor ( n51107 , n50856 , n50858 );
xor ( n51108 , n51107 , n50861 );
and ( n51109 , n51105 , n51108 );
and ( n51110 , n51103 , n51108 );
or ( n51111 , n51106 , n51109 , n51110 );
and ( n51112 , n51100 , n51111 );
and ( n51113 , n51019 , n51111 );
or ( n51114 , n51101 , n51112 , n51113 );
and ( n51115 , n50936 , n51114 );
and ( n51116 , n50919 , n51114 );
or ( n51117 , n50937 , n51115 , n51116 );
xor ( n51118 , n50707 , n50712 );
xor ( n51119 , n51118 , n50750 );
xor ( n51120 , n50801 , n50853 );
xor ( n51121 , n51120 , n50864 );
and ( n51122 , n51119 , n51121 );
xor ( n51123 , n50870 , n50872 );
xor ( n51124 , n51123 , n50875 );
and ( n51125 , n51121 , n51124 );
and ( n51126 , n51119 , n51124 );
or ( n51127 , n51122 , n51125 , n51126 );
xor ( n51128 , n50753 , n50867 );
xor ( n51129 , n51128 , n50878 );
and ( n51130 , n51127 , n51129 );
xor ( n51131 , n50898 , n50900 );
xor ( n51132 , n51131 , n50903 );
and ( n51133 , n51129 , n51132 );
and ( n51134 , n51127 , n51132 );
or ( n51135 , n51130 , n51133 , n51134 );
and ( n51136 , n51117 , n51135 );
xor ( n51137 , n50703 , n50705 );
xor ( n51138 , n51137 , n50881 );
and ( n51139 , n51135 , n51138 );
and ( n51140 , n51117 , n51138 );
or ( n51141 , n51136 , n51139 , n51140 );
and ( n51142 , n50916 , n51141 );
and ( n51143 , n50914 , n51141 );
or ( n51144 , n50917 , n51142 , n51143 );
xor ( n51145 , n50696 , n50887 );
xor ( n51146 , n51145 , n50890 );
and ( n51147 , n51144 , n51146 );
xor ( n51148 , n50698 , n50700 );
xor ( n51149 , n51148 , n50884 );
xor ( n51150 , n50906 , n50908 );
xor ( n51151 , n51150 , n50911 );
xor ( n51152 , n50821 , n50825 );
xor ( n51153 , n51152 , n50830 );
xor ( n51154 , n50838 , n50842 );
xor ( n51155 , n51154 , n50847 );
and ( n51156 , n51153 , n51155 );
and ( n51157 , n46445 , n48394 );
and ( n51158 , n46345 , n48392 );
nor ( n51159 , n51157 , n51158 );
xnor ( n51160 , n51159 , n48220 );
and ( n51161 , n47647 , n46911 );
and ( n51162 , n47474 , n46909 );
nor ( n51163 , n51161 , n51162 );
xnor ( n51164 , n51163 , n46802 );
and ( n51165 , n51160 , n51164 );
and ( n51166 , n47962 , n46712 );
and ( n51167 , n47778 , n46710 );
nor ( n51168 , n51166 , n51167 );
xnor ( n51169 , n51168 , n46587 );
and ( n51170 , n51164 , n51169 );
and ( n51171 , n51160 , n51169 );
or ( n51172 , n51165 , n51170 , n51171 );
and ( n51173 , n49570 , n45886 );
and ( n51174 , n49374 , n45884 );
nor ( n51175 , n51173 , n51174 );
xnor ( n51176 , n51175 , n45824 );
and ( n51177 , n51172 , n51176 );
and ( n51178 , n51155 , n51177 );
and ( n51179 , n51153 , n51177 );
or ( n51180 , n51156 , n51178 , n51179 );
xor ( n51181 , n50951 , n50955 );
xor ( n51182 , n51181 , n50960 );
xor ( n51183 , n50971 , n50975 );
xor ( n51184 , n51183 , n50980 );
and ( n51185 , n51182 , n51184 );
buf ( n51186 , n51185 );
xnor ( n51187 , n50987 , n50991 );
and ( n51188 , n48988 , n46135 );
and ( n51189 , n48709 , n46133 );
nor ( n51190 , n51188 , n51189 );
xnor ( n51191 , n51190 , n46067 );
and ( n51192 , n50195 , n45777 );
and ( n51193 , n49976 , n45775 );
nor ( n51194 , n51192 , n51193 );
xnor ( n51195 , n51194 , n45734 );
and ( n51196 , n51191 , n51195 );
and ( n51197 , n50625 , n45702 );
and ( n51198 , n50404 , n45700 );
nor ( n51199 , n51197 , n51198 );
xnor ( n51200 , n51199 , n20841 );
and ( n51201 , n51195 , n51200 );
and ( n51202 , n51191 , n51200 );
or ( n51203 , n51196 , n51201 , n51202 );
and ( n51204 , n51187 , n51203 );
and ( n51205 , n48632 , n46306 );
and ( n51206 , n48384 , n46304 );
nor ( n51207 , n51205 , n51206 );
xnor ( n51208 , n51207 , n46228 );
and ( n51209 , n49374 , n45990 );
and ( n51210 , n49115 , n45988 );
nor ( n51211 , n51209 , n51210 );
xnor ( n51212 , n51211 , n45939 );
or ( n51213 , n51208 , n51212 );
and ( n51214 , n51203 , n51213 );
and ( n51215 , n51187 , n51213 );
or ( n51216 , n51204 , n51214 , n51215 );
and ( n51217 , n51186 , n51216 );
xor ( n51218 , n50554 , n50995 );
xor ( n51219 , n50995 , n50997 );
not ( n51220 , n51219 );
and ( n51221 , n51218 , n51220 );
and ( n51222 , n20855 , n51221 );
not ( n51223 , n51222 );
xnor ( n51224 , n51223 , n51000 );
and ( n51225 , n20864 , n50783 );
and ( n51226 , n20844 , n50781 );
nor ( n51227 , n51225 , n51226 );
xnor ( n51228 , n51227 , n50557 );
and ( n51229 , n51224 , n51228 );
and ( n51230 , n45763 , n50338 );
and ( n51231 , n45712 , n50336 );
nor ( n51232 , n51230 , n51231 );
xnor ( n51233 , n51232 , n50111 );
and ( n51234 , n51228 , n51233 );
and ( n51235 , n51224 , n51233 );
or ( n51236 , n51229 , n51234 , n51235 );
and ( n51237 , n45843 , n49896 );
and ( n51238 , n45794 , n49894 );
nor ( n51239 , n51237 , n51238 );
xnor ( n51240 , n51239 , n49711 );
and ( n51241 , n45963 , n49513 );
and ( n51242 , n45907 , n49511 );
nor ( n51243 , n51241 , n51242 );
xnor ( n51244 , n51243 , n49310 );
and ( n51245 , n51240 , n51244 );
and ( n51246 , n46100 , n49121 );
and ( n51247 , n46041 , n49119 );
nor ( n51248 , n51246 , n51247 );
xnor ( n51249 , n51248 , n48932 );
and ( n51250 , n51244 , n51249 );
and ( n51251 , n51240 , n51249 );
or ( n51252 , n51245 , n51250 , n51251 );
and ( n51253 , n51236 , n51252 );
and ( n51254 , n46264 , n48740 );
and ( n51255 , n46169 , n48738 );
nor ( n51256 , n51254 , n51255 );
xnor ( n51257 , n51256 , n48571 );
and ( n51258 , n46577 , n48042 );
and ( n51259 , n46530 , n48040 );
nor ( n51260 , n51258 , n51259 );
xnor ( n51261 , n51260 , n47921 );
and ( n51262 , n51257 , n51261 );
and ( n51263 , n46843 , n47734 );
and ( n51264 , n46750 , n47732 );
nor ( n51265 , n51263 , n51264 );
xnor ( n51266 , n51265 , n47606 );
and ( n51267 , n51261 , n51266 );
and ( n51268 , n51257 , n51266 );
or ( n51269 , n51262 , n51267 , n51268 );
and ( n51270 , n51252 , n51269 );
and ( n51271 , n51236 , n51269 );
or ( n51272 , n51253 , n51270 , n51271 );
and ( n51273 , n51216 , n51272 );
and ( n51274 , n51186 , n51272 );
or ( n51275 , n51217 , n51273 , n51274 );
and ( n51276 , n51180 , n51275 );
and ( n51277 , n47090 , n47429 );
and ( n51278 , n46969 , n47427 );
nor ( n51279 , n51277 , n51278 );
xnor ( n51280 , n51279 , n47309 );
and ( n51281 , n47351 , n47178 );
and ( n51282 , n47216 , n47176 );
nor ( n51283 , n51281 , n51282 );
xnor ( n51284 , n51283 , n47039 );
and ( n51285 , n51280 , n51284 );
and ( n51286 , n48272 , n46496 );
and ( n51287 , n48108 , n46494 );
nor ( n51288 , n51286 , n51287 );
xnor ( n51289 , n51288 , n46402 );
and ( n51290 , n51284 , n51289 );
and ( n51291 , n51280 , n51289 );
or ( n51292 , n51285 , n51290 , n51291 );
and ( n51293 , n51077 , n20852 );
and ( n51294 , n50726 , n20850 );
nor ( n51295 , n51293 , n51294 );
xnor ( n51296 , n51295 , n20860 );
buf ( n51297 , n20776 );
buf ( n51298 , n51297 );
and ( n51299 , n51298 , n20846 );
and ( n51300 , n51296 , n51299 );
xor ( n51301 , n26010 , n45617 );
buf ( n51302 , n51301 );
buf ( n51303 , n51302 );
buf ( n51304 , n51303 );
and ( n51305 , n51299 , n51304 );
and ( n51306 , n51296 , n51304 );
or ( n51307 , n51300 , n51305 , n51306 );
and ( n51308 , n51292 , n51307 );
xor ( n51309 , n51001 , n51005 );
xor ( n51310 , n51309 , n51010 );
and ( n51311 , n51307 , n51310 );
and ( n51312 , n51292 , n51310 );
or ( n51313 , n51308 , n51311 , n51312 );
xor ( n51314 , n51023 , n51027 );
xor ( n51315 , n51314 , n51032 );
xor ( n51316 , n51039 , n51043 );
xor ( n51317 , n51316 , n51048 );
and ( n51318 , n51315 , n51317 );
xor ( n51319 , n51056 , n51060 );
xor ( n51320 , n51319 , n51065 );
and ( n51321 , n51317 , n51320 );
and ( n51322 , n51315 , n51320 );
or ( n51323 , n51318 , n51321 , n51322 );
and ( n51324 , n51313 , n51323 );
buf ( n51325 , n50939 );
xor ( n51326 , n51325 , n50941 );
and ( n51327 , n51323 , n51326 );
and ( n51328 , n51313 , n51326 );
or ( n51329 , n51324 , n51327 , n51328 );
and ( n51330 , n51275 , n51329 );
and ( n51331 , n51180 , n51329 );
or ( n51332 , n51276 , n51330 , n51331 );
xor ( n51333 , n50945 , n50946 );
xor ( n51334 , n51333 , n50963 );
xor ( n51335 , n50983 , n50992 );
xor ( n51336 , n51335 , n51013 );
and ( n51337 , n51334 , n51336 );
xor ( n51338 , n51035 , n51051 );
xor ( n51339 , n51338 , n51068 );
and ( n51340 , n51336 , n51339 );
and ( n51341 , n51334 , n51339 );
or ( n51342 , n51337 , n51340 , n51341 );
xor ( n51343 , n50926 , n50928 );
xor ( n51344 , n51343 , n50930 );
and ( n51345 , n51342 , n51344 );
xor ( n51346 , n50943 , n50966 );
xor ( n51347 , n51346 , n51016 );
and ( n51348 , n51344 , n51347 );
and ( n51349 , n51342 , n51347 );
or ( n51350 , n51345 , n51348 , n51349 );
and ( n51351 , n51332 , n51350 );
xor ( n51352 , n50921 , n50923 );
xor ( n51353 , n51352 , n50933 );
and ( n51354 , n51350 , n51353 );
and ( n51355 , n51332 , n51353 );
or ( n51356 , n51351 , n51354 , n51355 );
xor ( n51357 , n50919 , n50936 );
xor ( n51358 , n51357 , n51114 );
and ( n51359 , n51356 , n51358 );
xor ( n51360 , n51127 , n51129 );
xor ( n51361 , n51360 , n51132 );
and ( n51362 , n51358 , n51361 );
and ( n51363 , n51356 , n51361 );
or ( n51364 , n51359 , n51362 , n51363 );
and ( n51365 , n51151 , n51364 );
xor ( n51366 , n51117 , n51135 );
xor ( n51367 , n51366 , n51138 );
and ( n51368 , n51364 , n51367 );
and ( n51369 , n51151 , n51367 );
or ( n51370 , n51365 , n51368 , n51369 );
and ( n51371 , n51149 , n51370 );
xor ( n51372 , n50914 , n50916 );
xor ( n51373 , n51372 , n51141 );
and ( n51374 , n51370 , n51373 );
and ( n51375 , n51149 , n51373 );
or ( n51376 , n51371 , n51374 , n51375 );
and ( n51377 , n51146 , n51376 );
and ( n51378 , n51144 , n51376 );
or ( n51379 , n51147 , n51377 , n51378 );
and ( n51380 , n50895 , n51379 );
and ( n51381 , n50893 , n51379 );
or ( n51382 , n50896 , n51380 , n51381 );
and ( n51383 , n50693 , n51382 );
and ( n51384 , n50691 , n51382 );
or ( n51385 , n50694 , n51383 , n51384 );
and ( n51386 , n50466 , n51385 );
and ( n51387 , n50464 , n51385 );
or ( n51388 , n50467 , n51386 , n51387 );
and ( n51389 , n50259 , n51388 );
and ( n51390 , n50257 , n51388 );
or ( n51391 , n50260 , n51389 , n51390 );
or ( n51392 , n50054 , n51391 );
and ( n51393 , n50051 , n51392 );
and ( n51394 , n49633 , n51392 );
or ( n51395 , n50052 , n51393 , n51394 );
and ( n51396 , n49631 , n51395 );
xor ( n51397 , n49631 , n51395 );
xor ( n51398 , n49633 , n50051 );
xor ( n51399 , n51398 , n51392 );
not ( n51400 , n51399 );
xnor ( n51401 , n50054 , n51391 );
xor ( n51402 , n50257 , n50259 );
xor ( n51403 , n51402 , n51388 );
not ( n51404 , n51403 );
xor ( n51405 , n50464 , n50466 );
xor ( n51406 , n51405 , n51385 );
xor ( n51407 , n50691 , n50693 );
xor ( n51408 , n51407 , n51382 );
not ( n51409 , n51408 );
xor ( n51410 , n50893 , n50895 );
xor ( n51411 , n51410 , n51379 );
xor ( n51412 , n51144 , n51146 );
xor ( n51413 , n51412 , n51376 );
xor ( n51414 , n51149 , n51370 );
xor ( n51415 , n51414 , n51373 );
xor ( n51416 , n51151 , n51364 );
xor ( n51417 , n51416 , n51367 );
xor ( n51418 , n51019 , n51100 );
xor ( n51419 , n51418 , n51111 );
xor ( n51420 , n51119 , n51121 );
xor ( n51421 , n51420 , n51124 );
and ( n51422 , n51419 , n51421 );
xor ( n51423 , n51071 , n51094 );
xor ( n51424 , n51423 , n51097 );
xor ( n51425 , n51103 , n51105 );
xor ( n51426 , n51425 , n51108 );
and ( n51427 , n51424 , n51426 );
xor ( n51428 , n51086 , n51088 );
xor ( n51429 , n51428 , n51091 );
xor ( n51430 , n51075 , n51078 );
xor ( n51431 , n51430 , n51083 );
xor ( n51432 , n51172 , n51176 );
and ( n51433 , n51431 , n51432 );
and ( n51434 , n46750 , n48042 );
and ( n51435 , n46577 , n48040 );
nor ( n51436 , n51434 , n51435 );
xnor ( n51437 , n51436 , n47921 );
and ( n51438 , n47216 , n47429 );
and ( n51439 , n47090 , n47427 );
nor ( n51440 , n51438 , n51439 );
xnor ( n51441 , n51440 , n47309 );
and ( n51442 , n51437 , n51441 );
and ( n51443 , n47474 , n47178 );
and ( n51444 , n47351 , n47176 );
nor ( n51445 , n51443 , n51444 );
xnor ( n51446 , n51445 , n47039 );
and ( n51447 , n51441 , n51446 );
and ( n51448 , n51437 , n51446 );
or ( n51449 , n51442 , n51447 , n51448 );
and ( n51450 , n49781 , n45886 );
and ( n51451 , n49570 , n45884 );
nor ( n51452 , n51450 , n51451 );
xnor ( n51453 , n51452 , n45824 );
or ( n51454 , n51449 , n51453 );
and ( n51455 , n51432 , n51454 );
and ( n51456 , n51431 , n51454 );
or ( n51457 , n51433 , n51455 , n51456 );
and ( n51458 , n51429 , n51457 );
xor ( n51459 , n51191 , n51195 );
xor ( n51460 , n51459 , n51200 );
xor ( n51461 , n51160 , n51164 );
xor ( n51462 , n51461 , n51169 );
and ( n51463 , n51460 , n51462 );
buf ( n51464 , n51463 );
xnor ( n51465 , n51208 , n51212 );
and ( n51466 , n49115 , n46135 );
and ( n51467 , n48988 , n46133 );
nor ( n51468 , n51466 , n51467 );
xnor ( n51469 , n51468 , n46067 );
and ( n51470 , n50404 , n45777 );
and ( n51471 , n50195 , n45775 );
nor ( n51472 , n51470 , n51471 );
xnor ( n51473 , n51472 , n45734 );
and ( n51474 , n51469 , n51473 );
and ( n51475 , n51298 , n20852 );
and ( n51476 , n51077 , n20850 );
nor ( n51477 , n51475 , n51476 );
xnor ( n51478 , n51477 , n20860 );
and ( n51479 , n51473 , n51478 );
and ( n51480 , n51469 , n51478 );
or ( n51481 , n51474 , n51479 , n51480 );
and ( n51482 , n51465 , n51481 );
and ( n51483 , n46345 , n48740 );
and ( n51484 , n46264 , n48738 );
nor ( n51485 , n51483 , n51484 );
xnor ( n51486 , n51485 , n48571 );
and ( n51487 , n46969 , n47734 );
and ( n51488 , n46843 , n47732 );
nor ( n51489 , n51487 , n51488 );
xnor ( n51490 , n51489 , n47606 );
or ( n51491 , n51486 , n51490 );
and ( n51492 , n51481 , n51491 );
and ( n51493 , n51465 , n51491 );
or ( n51494 , n51482 , n51492 , n51493 );
and ( n51495 , n51464 , n51494 );
and ( n51496 , n48709 , n46306 );
and ( n51497 , n48632 , n46304 );
nor ( n51498 , n51496 , n51497 );
xnor ( n51499 , n51498 , n46228 );
and ( n51500 , n49976 , n45886 );
and ( n51501 , n49781 , n45884 );
nor ( n51502 , n51500 , n51501 );
xnor ( n51503 , n51502 , n45824 );
or ( n51504 , n51499 , n51503 );
and ( n51505 , n50726 , n45702 );
and ( n51506 , n50625 , n45700 );
nor ( n51507 , n51505 , n51506 );
xnor ( n51508 , n51507 , n20841 );
buf ( n51509 , n20778 );
buf ( n51510 , n51509 );
and ( n51511 , n51510 , n20846 );
or ( n51512 , n51508 , n51511 );
and ( n51513 , n51504 , n51512 );
buf ( n51514 , n17535 );
buf ( n51515 , n51514 );
buf ( n51516 , n17537 );
buf ( n51517 , n51516 );
and ( n51518 , n51515 , n51517 );
not ( n51519 , n51518 );
and ( n51520 , n50997 , n51519 );
not ( n51521 , n51520 );
and ( n51522 , n20844 , n51221 );
and ( n51523 , n20855 , n51219 );
nor ( n51524 , n51522 , n51523 );
xnor ( n51525 , n51524 , n51000 );
and ( n51526 , n51521 , n51525 );
and ( n51527 , n45712 , n50783 );
and ( n51528 , n20864 , n50781 );
nor ( n51529 , n51527 , n51528 );
xnor ( n51530 , n51529 , n50557 );
and ( n51531 , n51525 , n51530 );
and ( n51532 , n51521 , n51530 );
or ( n51533 , n51526 , n51531 , n51532 );
and ( n51534 , n51512 , n51533 );
and ( n51535 , n51504 , n51533 );
or ( n51536 , n51513 , n51534 , n51535 );
and ( n51537 , n51494 , n51536 );
and ( n51538 , n51464 , n51536 );
or ( n51539 , n51495 , n51537 , n51538 );
and ( n51540 , n51457 , n51539 );
and ( n51541 , n51429 , n51539 );
or ( n51542 , n51458 , n51540 , n51541 );
and ( n51543 , n51426 , n51542 );
and ( n51544 , n51424 , n51542 );
or ( n51545 , n51427 , n51543 , n51544 );
and ( n51546 , n51421 , n51545 );
and ( n51547 , n51419 , n51545 );
or ( n51548 , n51422 , n51546 , n51547 );
xor ( n51549 , n51356 , n51358 );
xor ( n51550 , n51549 , n51361 );
and ( n51551 , n51548 , n51550 );
and ( n51552 , n45794 , n50338 );
and ( n51553 , n45763 , n50336 );
nor ( n51554 , n51552 , n51553 );
xnor ( n51555 , n51554 , n50111 );
and ( n51556 , n45907 , n49896 );
and ( n51557 , n45843 , n49894 );
nor ( n51558 , n51556 , n51557 );
xnor ( n51559 , n51558 , n49711 );
and ( n51560 , n51555 , n51559 );
and ( n51561 , n46041 , n49513 );
and ( n51562 , n45963 , n49511 );
nor ( n51563 , n51561 , n51562 );
xnor ( n51564 , n51563 , n49310 );
and ( n51565 , n51559 , n51564 );
and ( n51566 , n51555 , n51564 );
or ( n51567 , n51560 , n51565 , n51566 );
and ( n51568 , n46169 , n49121 );
and ( n51569 , n46100 , n49119 );
nor ( n51570 , n51568 , n51569 );
xnor ( n51571 , n51570 , n48932 );
and ( n51572 , n46530 , n48394 );
and ( n51573 , n46445 , n48392 );
nor ( n51574 , n51572 , n51573 );
xnor ( n51575 , n51574 , n48220 );
and ( n51576 , n51571 , n51575 );
and ( n51577 , n47778 , n46911 );
and ( n51578 , n47647 , n46909 );
nor ( n51579 , n51577 , n51578 );
xnor ( n51580 , n51579 , n46802 );
and ( n51581 , n51575 , n51580 );
and ( n51582 , n51571 , n51580 );
or ( n51583 , n51576 , n51581 , n51582 );
and ( n51584 , n51567 , n51583 );
and ( n51585 , n48108 , n46712 );
and ( n51586 , n47962 , n46710 );
nor ( n51587 , n51585 , n51586 );
xnor ( n51588 , n51587 , n46587 );
and ( n51589 , n48384 , n46496 );
and ( n51590 , n48272 , n46494 );
nor ( n51591 , n51589 , n51590 );
xnor ( n51592 , n51591 , n46402 );
and ( n51593 , n51588 , n51592 );
and ( n51594 , n49570 , n45990 );
and ( n51595 , n49374 , n45988 );
nor ( n51596 , n51594 , n51595 );
xnor ( n51597 , n51596 , n45939 );
and ( n51598 , n51592 , n51597 );
and ( n51599 , n51588 , n51597 );
or ( n51600 , n51593 , n51598 , n51599 );
and ( n51601 , n51583 , n51600 );
and ( n51602 , n51567 , n51600 );
or ( n51603 , n51584 , n51601 , n51602 );
xor ( n51604 , n51224 , n51228 );
xor ( n51605 , n51604 , n51233 );
xor ( n51606 , n51240 , n51244 );
xor ( n51607 , n51606 , n51249 );
and ( n51608 , n51605 , n51607 );
xor ( n51609 , n51257 , n51261 );
xor ( n51610 , n51609 , n51266 );
and ( n51611 , n51607 , n51610 );
and ( n51612 , n51605 , n51610 );
or ( n51613 , n51608 , n51611 , n51612 );
and ( n51614 , n51603 , n51613 );
buf ( n51615 , n51182 );
xor ( n51616 , n51615 , n51184 );
and ( n51617 , n51613 , n51616 );
and ( n51618 , n51603 , n51616 );
or ( n51619 , n51614 , n51617 , n51618 );
xor ( n51620 , n51187 , n51203 );
xor ( n51621 , n51620 , n51213 );
xor ( n51622 , n51236 , n51252 );
xor ( n51623 , n51622 , n51269 );
and ( n51624 , n51621 , n51623 );
xor ( n51625 , n51292 , n51307 );
xor ( n51626 , n51625 , n51310 );
and ( n51627 , n51623 , n51626 );
and ( n51628 , n51621 , n51626 );
or ( n51629 , n51624 , n51627 , n51628 );
and ( n51630 , n51619 , n51629 );
xor ( n51631 , n51153 , n51155 );
xor ( n51632 , n51631 , n51177 );
and ( n51633 , n51629 , n51632 );
and ( n51634 , n51619 , n51632 );
or ( n51635 , n51630 , n51633 , n51634 );
xor ( n51636 , n51186 , n51216 );
xor ( n51637 , n51636 , n51272 );
xor ( n51638 , n51313 , n51323 );
xor ( n51639 , n51638 , n51326 );
and ( n51640 , n51637 , n51639 );
xor ( n51641 , n51334 , n51336 );
xor ( n51642 , n51641 , n51339 );
and ( n51643 , n51639 , n51642 );
and ( n51644 , n51637 , n51642 );
or ( n51645 , n51640 , n51643 , n51644 );
and ( n51646 , n51635 , n51645 );
xor ( n51647 , n51180 , n51275 );
xor ( n51648 , n51647 , n51329 );
and ( n51649 , n51645 , n51648 );
and ( n51650 , n51635 , n51648 );
or ( n51651 , n51646 , n51649 , n51650 );
xor ( n51652 , n51332 , n51350 );
xor ( n51653 , n51652 , n51353 );
and ( n51654 , n51651 , n51653 );
xor ( n51655 , n51342 , n51344 );
xor ( n51656 , n51655 , n51347 );
xor ( n51657 , n51315 , n51317 );
xor ( n51658 , n51657 , n51320 );
xor ( n51659 , n51280 , n51284 );
xor ( n51660 , n51659 , n51289 );
xor ( n51661 , n51296 , n51299 );
xor ( n51662 , n51661 , n51304 );
and ( n51663 , n51660 , n51662 );
xnor ( n51664 , n51449 , n51453 );
and ( n51665 , n51662 , n51664 );
and ( n51666 , n51660 , n51664 );
or ( n51667 , n51663 , n51665 , n51666 );
and ( n51668 , n51658 , n51667 );
xor ( n51669 , n26627 , n45615 );
buf ( n51670 , n51669 );
buf ( n51671 , n51670 );
buf ( n51672 , n51671 );
xor ( n51673 , n51469 , n51473 );
xor ( n51674 , n51673 , n51478 );
and ( n51675 , n51672 , n51674 );
buf ( n51676 , n51675 );
xor ( n51677 , n51437 , n51441 );
xor ( n51678 , n51677 , n51446 );
xnor ( n51679 , n51486 , n51490 );
and ( n51680 , n51678 , n51679 );
xnor ( n51681 , n51499 , n51503 );
and ( n51682 , n51679 , n51681 );
and ( n51683 , n51678 , n51681 );
or ( n51684 , n51680 , n51682 , n51683 );
and ( n51685 , n51676 , n51684 );
xnor ( n51686 , n51508 , n51511 );
and ( n51687 , n46577 , n48394 );
and ( n51688 , n46530 , n48392 );
nor ( n51689 , n51687 , n51688 );
xnor ( n51690 , n51689 , n48220 );
and ( n51691 , n46843 , n48042 );
and ( n51692 , n46750 , n48040 );
nor ( n51693 , n51691 , n51692 );
xnor ( n51694 , n51693 , n47921 );
and ( n51695 , n51690 , n51694 );
and ( n51696 , n47962 , n46911 );
and ( n51697 , n47778 , n46909 );
nor ( n51698 , n51696 , n51697 );
xnor ( n51699 , n51698 , n46802 );
and ( n51700 , n51694 , n51699 );
and ( n51701 , n51690 , n51699 );
or ( n51702 , n51695 , n51700 , n51701 );
and ( n51703 , n51686 , n51702 );
and ( n51704 , n49374 , n46135 );
and ( n51705 , n49115 , n46133 );
nor ( n51706 , n51704 , n51705 );
xnor ( n51707 , n51706 , n46067 );
and ( n51708 , n50625 , n45777 );
and ( n51709 , n50404 , n45775 );
nor ( n51710 , n51708 , n51709 );
xnor ( n51711 , n51710 , n45734 );
and ( n51712 , n51707 , n51711 );
and ( n51713 , n51077 , n45702 );
and ( n51714 , n50726 , n45700 );
nor ( n51715 , n51713 , n51714 );
xnor ( n51716 , n51715 , n20841 );
and ( n51717 , n51711 , n51716 );
and ( n51718 , n51707 , n51716 );
or ( n51719 , n51712 , n51717 , n51718 );
and ( n51720 , n51702 , n51719 );
and ( n51721 , n51686 , n51719 );
or ( n51722 , n51703 , n51720 , n51721 );
and ( n51723 , n51684 , n51722 );
and ( n51724 , n51676 , n51722 );
or ( n51725 , n51685 , n51723 , n51724 );
and ( n51726 , n51667 , n51725 );
and ( n51727 , n51658 , n51725 );
or ( n51728 , n51668 , n51726 , n51727 );
and ( n51729 , n49781 , n45990 );
and ( n51730 , n49570 , n45988 );
nor ( n51731 , n51729 , n51730 );
xnor ( n51732 , n51731 , n45939 );
buf ( n51733 , n20780 );
buf ( n51734 , n51733 );
and ( n51735 , n51734 , n20846 );
or ( n51736 , n51732 , n51735 );
and ( n51737 , n50195 , n45886 );
and ( n51738 , n49976 , n45884 );
nor ( n51739 , n51737 , n51738 );
xnor ( n51740 , n51739 , n45824 );
and ( n51741 , n51510 , n20852 );
and ( n51742 , n51298 , n20850 );
nor ( n51743 , n51741 , n51742 );
xnor ( n51744 , n51743 , n20860 );
or ( n51745 , n51740 , n51744 );
and ( n51746 , n51736 , n51745 );
xor ( n51747 , n50997 , n51515 );
xor ( n51748 , n51515 , n51517 );
not ( n51749 , n51748 );
and ( n51750 , n51747 , n51749 );
and ( n51751 , n20855 , n51750 );
not ( n51752 , n51751 );
xnor ( n51753 , n51752 , n51520 );
and ( n51754 , n20864 , n51221 );
and ( n51755 , n20844 , n51219 );
nor ( n51756 , n51754 , n51755 );
xnor ( n51757 , n51756 , n51000 );
and ( n51758 , n51753 , n51757 );
and ( n51759 , n45763 , n50783 );
and ( n51760 , n45712 , n50781 );
nor ( n51761 , n51759 , n51760 );
xnor ( n51762 , n51761 , n50557 );
and ( n51763 , n51757 , n51762 );
and ( n51764 , n51753 , n51762 );
or ( n51765 , n51758 , n51763 , n51764 );
and ( n51766 , n51745 , n51765 );
and ( n51767 , n51736 , n51765 );
or ( n51768 , n51746 , n51766 , n51767 );
and ( n51769 , n45843 , n50338 );
and ( n51770 , n45794 , n50336 );
nor ( n51771 , n51769 , n51770 );
xnor ( n51772 , n51771 , n50111 );
and ( n51773 , n45963 , n49896 );
and ( n51774 , n45907 , n49894 );
nor ( n51775 , n51773 , n51774 );
xnor ( n51776 , n51775 , n49711 );
and ( n51777 , n51772 , n51776 );
and ( n51778 , n46100 , n49513 );
and ( n51779 , n46041 , n49511 );
nor ( n51780 , n51778 , n51779 );
xnor ( n51781 , n51780 , n49310 );
and ( n51782 , n51776 , n51781 );
and ( n51783 , n51772 , n51781 );
or ( n51784 , n51777 , n51782 , n51783 );
and ( n51785 , n46264 , n49121 );
and ( n51786 , n46169 , n49119 );
nor ( n51787 , n51785 , n51786 );
xnor ( n51788 , n51787 , n48932 );
and ( n51789 , n46445 , n48740 );
and ( n51790 , n46345 , n48738 );
nor ( n51791 , n51789 , n51790 );
xnor ( n51792 , n51791 , n48571 );
and ( n51793 , n51788 , n51792 );
and ( n51794 , n47090 , n47734 );
and ( n51795 , n46969 , n47732 );
nor ( n51796 , n51794 , n51795 );
xnor ( n51797 , n51796 , n47606 );
and ( n51798 , n51792 , n51797 );
and ( n51799 , n51788 , n51797 );
or ( n51800 , n51793 , n51798 , n51799 );
and ( n51801 , n51784 , n51800 );
and ( n51802 , n47351 , n47429 );
and ( n51803 , n47216 , n47427 );
nor ( n51804 , n51802 , n51803 );
xnor ( n51805 , n51804 , n47309 );
and ( n51806 , n47647 , n47178 );
and ( n51807 , n47474 , n47176 );
nor ( n51808 , n51806 , n51807 );
xnor ( n51809 , n51808 , n47039 );
and ( n51810 , n51805 , n51809 );
and ( n51811 , n48272 , n46712 );
and ( n51812 , n48108 , n46710 );
nor ( n51813 , n51811 , n51812 );
xnor ( n51814 , n51813 , n46587 );
and ( n51815 , n51809 , n51814 );
and ( n51816 , n51805 , n51814 );
or ( n51817 , n51810 , n51815 , n51816 );
and ( n51818 , n51800 , n51817 );
and ( n51819 , n51784 , n51817 );
or ( n51820 , n51801 , n51818 , n51819 );
and ( n51821 , n51768 , n51820 );
and ( n51822 , n48632 , n46496 );
and ( n51823 , n48384 , n46494 );
nor ( n51824 , n51822 , n51823 );
xnor ( n51825 , n51824 , n46402 );
and ( n51826 , n48988 , n46306 );
and ( n51827 , n48709 , n46304 );
nor ( n51828 , n51826 , n51827 );
xnor ( n51829 , n51828 , n46228 );
and ( n51830 , n51825 , n51829 );
xor ( n51831 , n26630 , n45613 );
buf ( n51832 , n51831 );
buf ( n51833 , n51832 );
buf ( n51834 , n51833 );
and ( n51835 , n51829 , n51834 );
and ( n51836 , n51825 , n51834 );
or ( n51837 , n51830 , n51835 , n51836 );
xor ( n51838 , n51521 , n51525 );
xor ( n51839 , n51838 , n51530 );
and ( n51840 , n51837 , n51839 );
xor ( n51841 , n51555 , n51559 );
xor ( n51842 , n51841 , n51564 );
and ( n51843 , n51839 , n51842 );
and ( n51844 , n51837 , n51842 );
or ( n51845 , n51840 , n51843 , n51844 );
and ( n51846 , n51820 , n51845 );
and ( n51847 , n51768 , n51845 );
or ( n51848 , n51821 , n51846 , n51847 );
buf ( n51849 , n51460 );
xor ( n51850 , n51849 , n51462 );
xor ( n51851 , n51465 , n51481 );
xor ( n51852 , n51851 , n51491 );
and ( n51853 , n51850 , n51852 );
xor ( n51854 , n51504 , n51512 );
xor ( n51855 , n51854 , n51533 );
and ( n51856 , n51852 , n51855 );
and ( n51857 , n51850 , n51855 );
or ( n51858 , n51853 , n51856 , n51857 );
and ( n51859 , n51848 , n51858 );
xor ( n51860 , n51431 , n51432 );
xor ( n51861 , n51860 , n51454 );
and ( n51862 , n51858 , n51861 );
and ( n51863 , n51848 , n51861 );
or ( n51864 , n51859 , n51862 , n51863 );
and ( n51865 , n51728 , n51864 );
xor ( n51866 , n51464 , n51494 );
xor ( n51867 , n51866 , n51536 );
xor ( n51868 , n51603 , n51613 );
xor ( n51869 , n51868 , n51616 );
and ( n51870 , n51867 , n51869 );
xor ( n51871 , n51621 , n51623 );
xor ( n51872 , n51871 , n51626 );
and ( n51873 , n51869 , n51872 );
and ( n51874 , n51867 , n51872 );
or ( n51875 , n51870 , n51873 , n51874 );
and ( n51876 , n51864 , n51875 );
and ( n51877 , n51728 , n51875 );
or ( n51878 , n51865 , n51876 , n51877 );
and ( n51879 , n51656 , n51878 );
xor ( n51880 , n51429 , n51457 );
xor ( n51881 , n51880 , n51539 );
xor ( n51882 , n51619 , n51629 );
xor ( n51883 , n51882 , n51632 );
and ( n51884 , n51881 , n51883 );
xor ( n51885 , n51637 , n51639 );
xor ( n51886 , n51885 , n51642 );
and ( n51887 , n51883 , n51886 );
and ( n51888 , n51881 , n51886 );
or ( n51889 , n51884 , n51887 , n51888 );
and ( n51890 , n51878 , n51889 );
and ( n51891 , n51656 , n51889 );
or ( n51892 , n51879 , n51890 , n51891 );
and ( n51893 , n51653 , n51892 );
and ( n51894 , n51651 , n51892 );
or ( n51895 , n51654 , n51893 , n51894 );
and ( n51896 , n51550 , n51895 );
and ( n51897 , n51548 , n51895 );
or ( n51898 , n51551 , n51896 , n51897 );
or ( n51899 , n51417 , n51898 );
or ( n51900 , n51415 , n51899 );
and ( n51901 , n51413 , n51900 );
xor ( n51902 , n51413 , n51900 );
xnor ( n51903 , n51415 , n51899 );
xnor ( n51904 , n51417 , n51898 );
xor ( n51905 , n51419 , n51421 );
xor ( n51906 , n51905 , n51545 );
xor ( n51907 , n51424 , n51426 );
xor ( n51908 , n51907 , n51542 );
xor ( n51909 , n51635 , n51645 );
xor ( n51910 , n51909 , n51648 );
and ( n51911 , n51908 , n51910 );
xor ( n51912 , n51567 , n51583 );
xor ( n51913 , n51912 , n51600 );
xor ( n51914 , n51605 , n51607 );
xor ( n51915 , n51914 , n51610 );
and ( n51916 , n51913 , n51915 );
xor ( n51917 , n51571 , n51575 );
xor ( n51918 , n51917 , n51580 );
xor ( n51919 , n51588 , n51592 );
xor ( n51920 , n51919 , n51597 );
and ( n51921 , n51918 , n51920 );
xor ( n51922 , n51690 , n51694 );
xor ( n51923 , n51922 , n51699 );
xor ( n51924 , n51707 , n51711 );
xor ( n51925 , n51924 , n51716 );
and ( n51926 , n51923 , n51925 );
buf ( n51927 , n51926 );
and ( n51928 , n51920 , n51927 );
and ( n51929 , n51918 , n51927 );
or ( n51930 , n51921 , n51928 , n51929 );
and ( n51931 , n51915 , n51930 );
and ( n51932 , n51913 , n51930 );
or ( n51933 , n51916 , n51931 , n51932 );
xnor ( n51934 , n51732 , n51735 );
xnor ( n51935 , n51740 , n51744 );
and ( n51936 , n51934 , n51935 );
and ( n51937 , n49570 , n46135 );
and ( n51938 , n49374 , n46133 );
nor ( n51939 , n51937 , n51938 );
xnor ( n51940 , n51939 , n46067 );
and ( n51941 , n50726 , n45777 );
and ( n51942 , n50625 , n45775 );
nor ( n51943 , n51941 , n51942 );
xnor ( n51944 , n51943 , n45734 );
and ( n51945 , n51940 , n51944 );
and ( n51946 , n51298 , n45702 );
and ( n51947 , n51077 , n45700 );
nor ( n51948 , n51946 , n51947 );
xnor ( n51949 , n51948 , n20841 );
and ( n51950 , n51944 , n51949 );
and ( n51951 , n51940 , n51949 );
or ( n51952 , n51945 , n51950 , n51951 );
and ( n51953 , n51935 , n51952 );
and ( n51954 , n51934 , n51952 );
or ( n51955 , n51936 , n51953 , n51954 );
and ( n51956 , n49115 , n46306 );
and ( n51957 , n48988 , n46304 );
nor ( n51958 , n51956 , n51957 );
xnor ( n51959 , n51958 , n46228 );
and ( n51960 , n49976 , n45990 );
and ( n51961 , n49781 , n45988 );
nor ( n51962 , n51960 , n51961 );
xnor ( n51963 , n51962 , n45939 );
and ( n51964 , n51959 , n51963 );
and ( n51965 , n50404 , n45886 );
and ( n51966 , n50195 , n45884 );
nor ( n51967 , n51965 , n51966 );
xnor ( n51968 , n51967 , n45824 );
and ( n51969 , n51963 , n51968 );
and ( n51970 , n51959 , n51968 );
or ( n51971 , n51964 , n51969 , n51970 );
and ( n51972 , n46750 , n48394 );
and ( n51973 , n46577 , n48392 );
nor ( n51974 , n51972 , n51973 );
xnor ( n51975 , n51974 , n48220 );
and ( n51976 , n47474 , n47429 );
and ( n51977 , n47351 , n47427 );
nor ( n51978 , n51976 , n51977 );
xnor ( n51979 , n51978 , n47309 );
and ( n51980 , n51975 , n51979 );
and ( n51981 , n48384 , n46712 );
and ( n51982 , n48272 , n46710 );
nor ( n51983 , n51981 , n51982 );
xnor ( n51984 , n51983 , n46587 );
and ( n51985 , n51979 , n51984 );
and ( n51986 , n51975 , n51984 );
or ( n51987 , n51980 , n51985 , n51986 );
and ( n51988 , n51971 , n51987 );
and ( n51989 , n46530 , n48740 );
and ( n51990 , n46445 , n48738 );
nor ( n51991 , n51989 , n51990 );
xnor ( n51992 , n51991 , n48571 );
and ( n51993 , n47216 , n47734 );
and ( n51994 , n47090 , n47732 );
nor ( n51995 , n51993 , n51994 );
xnor ( n51996 , n51995 , n47606 );
or ( n51997 , n51992 , n51996 );
and ( n51998 , n51987 , n51997 );
and ( n51999 , n51971 , n51997 );
or ( n52000 , n51988 , n51998 , n51999 );
and ( n52001 , n51955 , n52000 );
buf ( n52002 , n17539 );
buf ( n52003 , n52002 );
buf ( n52004 , n17541 );
buf ( n52005 , n52004 );
and ( n52006 , n52003 , n52005 );
not ( n52007 , n52006 );
and ( n52008 , n51517 , n52007 );
not ( n52009 , n52008 );
and ( n52010 , n20844 , n51750 );
and ( n52011 , n20855 , n51748 );
nor ( n52012 , n52010 , n52011 );
xnor ( n52013 , n52012 , n51520 );
and ( n52014 , n52009 , n52013 );
and ( n52015 , n45712 , n51221 );
and ( n52016 , n20864 , n51219 );
nor ( n52017 , n52015 , n52016 );
xnor ( n52018 , n52017 , n51000 );
and ( n52019 , n52013 , n52018 );
and ( n52020 , n52009 , n52018 );
or ( n52021 , n52014 , n52019 , n52020 );
and ( n52022 , n45794 , n50783 );
and ( n52023 , n45763 , n50781 );
nor ( n52024 , n52022 , n52023 );
xnor ( n52025 , n52024 , n50557 );
and ( n52026 , n45907 , n50338 );
and ( n52027 , n45843 , n50336 );
nor ( n52028 , n52026 , n52027 );
xnor ( n52029 , n52028 , n50111 );
and ( n52030 , n52025 , n52029 );
and ( n52031 , n46041 , n49896 );
and ( n52032 , n45963 , n49894 );
nor ( n52033 , n52031 , n52032 );
xnor ( n52034 , n52033 , n49711 );
and ( n52035 , n52029 , n52034 );
and ( n52036 , n52025 , n52034 );
or ( n52037 , n52030 , n52035 , n52036 );
and ( n52038 , n52021 , n52037 );
and ( n52039 , n46169 , n49513 );
and ( n52040 , n46100 , n49511 );
nor ( n52041 , n52039 , n52040 );
xnor ( n52042 , n52041 , n49310 );
and ( n52043 , n46345 , n49121 );
and ( n52044 , n46264 , n49119 );
nor ( n52045 , n52043 , n52044 );
xnor ( n52046 , n52045 , n48932 );
and ( n52047 , n52042 , n52046 );
and ( n52048 , n46969 , n48042 );
and ( n52049 , n46843 , n48040 );
nor ( n52050 , n52048 , n52049 );
xnor ( n52051 , n52050 , n47921 );
and ( n52052 , n52046 , n52051 );
and ( n52053 , n52042 , n52051 );
or ( n52054 , n52047 , n52052 , n52053 );
and ( n52055 , n52037 , n52054 );
and ( n52056 , n52021 , n52054 );
or ( n52057 , n52038 , n52055 , n52056 );
and ( n52058 , n52000 , n52057 );
and ( n52059 , n51955 , n52057 );
or ( n52060 , n52001 , n52058 , n52059 );
and ( n52061 , n47778 , n47178 );
and ( n52062 , n47647 , n47176 );
nor ( n52063 , n52061 , n52062 );
xnor ( n52064 , n52063 , n47039 );
and ( n52065 , n48108 , n46911 );
and ( n52066 , n47962 , n46909 );
nor ( n52067 , n52065 , n52066 );
xnor ( n52068 , n52067 , n46802 );
and ( n52069 , n52064 , n52068 );
and ( n52070 , n48709 , n46496 );
and ( n52071 , n48632 , n46494 );
nor ( n52072 , n52070 , n52071 );
xnor ( n52073 , n52072 , n46402 );
and ( n52074 , n52068 , n52073 );
and ( n52075 , n52064 , n52073 );
or ( n52076 , n52069 , n52074 , n52075 );
and ( n52077 , n51734 , n20852 );
and ( n52078 , n51510 , n20850 );
nor ( n52079 , n52077 , n52078 );
xnor ( n52080 , n52079 , n20860 );
buf ( n52081 , n20782 );
buf ( n52082 , n52081 );
and ( n52083 , n52082 , n20846 );
and ( n52084 , n52080 , n52083 );
xor ( n52085 , n26632 , n45612 );
buf ( n52086 , n52085 );
buf ( n52087 , n52086 );
buf ( n52088 , n52087 );
and ( n52089 , n52083 , n52088 );
and ( n52090 , n52080 , n52088 );
or ( n52091 , n52084 , n52089 , n52090 );
and ( n52092 , n52076 , n52091 );
xor ( n52093 , n51753 , n51757 );
xor ( n52094 , n52093 , n51762 );
and ( n52095 , n52091 , n52094 );
and ( n52096 , n52076 , n52094 );
or ( n52097 , n52092 , n52095 , n52096 );
xor ( n52098 , n51772 , n51776 );
xor ( n52099 , n52098 , n51781 );
xor ( n52100 , n51788 , n51792 );
xor ( n52101 , n52100 , n51797 );
and ( n52102 , n52099 , n52101 );
xor ( n52103 , n51805 , n51809 );
xor ( n52104 , n52103 , n51814 );
and ( n52105 , n52101 , n52104 );
and ( n52106 , n52099 , n52104 );
or ( n52107 , n52102 , n52105 , n52106 );
and ( n52108 , n52097 , n52107 );
buf ( n52109 , n51672 );
xor ( n52110 , n52109 , n51674 );
and ( n52111 , n52107 , n52110 );
and ( n52112 , n52097 , n52110 );
or ( n52113 , n52108 , n52111 , n52112 );
and ( n52114 , n52060 , n52113 );
xor ( n52115 , n51678 , n51679 );
xor ( n52116 , n52115 , n51681 );
xor ( n52117 , n51686 , n51702 );
xor ( n52118 , n52117 , n51719 );
and ( n52119 , n52116 , n52118 );
xor ( n52120 , n51736 , n51745 );
xor ( n52121 , n52120 , n51765 );
and ( n52122 , n52118 , n52121 );
and ( n52123 , n52116 , n52121 );
or ( n52124 , n52119 , n52122 , n52123 );
and ( n52125 , n52113 , n52124 );
and ( n52126 , n52060 , n52124 );
or ( n52127 , n52114 , n52125 , n52126 );
and ( n52128 , n51933 , n52127 );
xor ( n52129 , n51660 , n51662 );
xor ( n52130 , n52129 , n51664 );
xor ( n52131 , n51676 , n51684 );
xor ( n52132 , n52131 , n51722 );
and ( n52133 , n52130 , n52132 );
xor ( n52134 , n51768 , n51820 );
xor ( n52135 , n52134 , n51845 );
and ( n52136 , n52132 , n52135 );
and ( n52137 , n52130 , n52135 );
or ( n52138 , n52133 , n52136 , n52137 );
and ( n52139 , n52127 , n52138 );
and ( n52140 , n51933 , n52138 );
or ( n52141 , n52128 , n52139 , n52140 );
xor ( n52142 , n51658 , n51667 );
xor ( n52143 , n52142 , n51725 );
xor ( n52144 , n51848 , n51858 );
xor ( n52145 , n52144 , n51861 );
and ( n52146 , n52143 , n52145 );
xor ( n52147 , n51867 , n51869 );
xor ( n52148 , n52147 , n51872 );
and ( n52149 , n52145 , n52148 );
and ( n52150 , n52143 , n52148 );
or ( n52151 , n52146 , n52149 , n52150 );
and ( n52152 , n52141 , n52151 );
xor ( n52153 , n51728 , n51864 );
xor ( n52154 , n52153 , n51875 );
and ( n52155 , n52151 , n52154 );
and ( n52156 , n52141 , n52154 );
or ( n52157 , n52152 , n52155 , n52156 );
and ( n52158 , n51910 , n52157 );
and ( n52159 , n51908 , n52157 );
or ( n52160 , n51911 , n52158 , n52159 );
and ( n52161 , n51906 , n52160 );
xor ( n52162 , n51651 , n51653 );
xor ( n52163 , n52162 , n51892 );
and ( n52164 , n52160 , n52163 );
and ( n52165 , n51906 , n52163 );
or ( n52166 , n52161 , n52164 , n52165 );
xor ( n52167 , n51548 , n51550 );
xor ( n52168 , n52167 , n51895 );
and ( n52169 , n52166 , n52168 );
xor ( n52170 , n52166 , n52168 );
xor ( n52171 , n51656 , n51878 );
xor ( n52172 , n52171 , n51889 );
xor ( n52173 , n51881 , n51883 );
xor ( n52174 , n52173 , n51886 );
xor ( n52175 , n51850 , n51852 );
xor ( n52176 , n52175 , n51855 );
xor ( n52177 , n51784 , n51800 );
xor ( n52178 , n52177 , n51817 );
xor ( n52179 , n51837 , n51839 );
xor ( n52180 , n52179 , n51842 );
and ( n52181 , n52178 , n52180 );
xor ( n52182 , n51825 , n51829 );
xor ( n52183 , n52182 , n51834 );
xor ( n52184 , n51940 , n51944 );
xor ( n52185 , n52184 , n51949 );
xor ( n52186 , n51959 , n51963 );
xor ( n52187 , n52186 , n51968 );
or ( n52188 , n52185 , n52187 );
and ( n52189 , n52183 , n52188 );
xor ( n52190 , n51975 , n51979 );
xor ( n52191 , n52190 , n51984 );
xnor ( n52192 , n51992 , n51996 );
and ( n52193 , n52191 , n52192 );
buf ( n52194 , n52193 );
and ( n52195 , n52188 , n52194 );
and ( n52196 , n52183 , n52194 );
or ( n52197 , n52189 , n52195 , n52196 );
and ( n52198 , n52180 , n52197 );
and ( n52199 , n52178 , n52197 );
or ( n52200 , n52181 , n52198 , n52199 );
and ( n52201 , n52176 , n52200 );
and ( n52202 , n47090 , n48042 );
and ( n52203 , n46969 , n48040 );
nor ( n52204 , n52202 , n52203 );
xnor ( n52205 , n52204 , n47921 );
and ( n52206 , n48272 , n46911 );
and ( n52207 , n48108 , n46909 );
nor ( n52208 , n52206 , n52207 );
xnor ( n52209 , n52208 , n46802 );
and ( n52210 , n52205 , n52209 );
and ( n52211 , n48632 , n46712 );
and ( n52212 , n48384 , n46710 );
nor ( n52213 , n52211 , n52212 );
xnor ( n52214 , n52213 , n46587 );
and ( n52215 , n52209 , n52214 );
and ( n52216 , n52205 , n52214 );
or ( n52217 , n52210 , n52215 , n52216 );
and ( n52218 , n49374 , n46306 );
and ( n52219 , n49115 , n46304 );
nor ( n52220 , n52218 , n52219 );
xnor ( n52221 , n52220 , n46228 );
and ( n52222 , n50195 , n45990 );
and ( n52223 , n49976 , n45988 );
nor ( n52224 , n52222 , n52223 );
xnor ( n52225 , n52224 , n45939 );
and ( n52226 , n52221 , n52225 );
and ( n52227 , n51510 , n45702 );
and ( n52228 , n51298 , n45700 );
nor ( n52229 , n52227 , n52228 );
xnor ( n52230 , n52229 , n20841 );
and ( n52231 , n52225 , n52230 );
and ( n52232 , n52221 , n52230 );
or ( n52233 , n52226 , n52231 , n52232 );
and ( n52234 , n52217 , n52233 );
and ( n52235 , n46577 , n48740 );
and ( n52236 , n46530 , n48738 );
nor ( n52237 , n52235 , n52236 );
xnor ( n52238 , n52237 , n48571 );
and ( n52239 , n47351 , n47734 );
and ( n52240 , n47216 , n47732 );
nor ( n52241 , n52239 , n52240 );
xnor ( n52242 , n52241 , n47606 );
or ( n52243 , n52238 , n52242 );
and ( n52244 , n52233 , n52243 );
and ( n52245 , n52217 , n52243 );
or ( n52246 , n52234 , n52244 , n52245 );
and ( n52247 , n49781 , n46135 );
and ( n52248 , n49570 , n46133 );
nor ( n52249 , n52247 , n52248 );
xnor ( n52250 , n52249 , n46067 );
and ( n52251 , n51077 , n45777 );
and ( n52252 , n50726 , n45775 );
nor ( n52253 , n52251 , n52252 );
xnor ( n52254 , n52253 , n45734 );
or ( n52255 , n52250 , n52254 );
and ( n52256 , n46843 , n48394 );
and ( n52257 , n46750 , n48392 );
nor ( n52258 , n52256 , n52257 );
xnor ( n52259 , n52258 , n48220 );
and ( n52260 , n47647 , n47429 );
and ( n52261 , n47474 , n47427 );
nor ( n52262 , n52260 , n52261 );
xnor ( n52263 , n52262 , n47309 );
and ( n52264 , n52259 , n52263 );
and ( n52265 , n52255 , n52264 );
xor ( n52266 , n51517 , n52003 );
xor ( n52267 , n52003 , n52005 );
not ( n52268 , n52267 );
and ( n52269 , n52266 , n52268 );
and ( n52270 , n20855 , n52269 );
not ( n52271 , n52270 );
xnor ( n52272 , n52271 , n52008 );
and ( n52273 , n20864 , n51750 );
and ( n52274 , n20844 , n51748 );
nor ( n52275 , n52273 , n52274 );
xnor ( n52276 , n52275 , n51520 );
and ( n52277 , n52272 , n52276 );
and ( n52278 , n45763 , n51221 );
and ( n52279 , n45712 , n51219 );
nor ( n52280 , n52278 , n52279 );
xnor ( n52281 , n52280 , n51000 );
and ( n52282 , n52276 , n52281 );
and ( n52283 , n52272 , n52281 );
or ( n52284 , n52277 , n52282 , n52283 );
and ( n52285 , n52264 , n52284 );
and ( n52286 , n52255 , n52284 );
or ( n52287 , n52265 , n52285 , n52286 );
and ( n52288 , n52246 , n52287 );
and ( n52289 , n45843 , n50783 );
and ( n52290 , n45794 , n50781 );
nor ( n52291 , n52289 , n52290 );
xnor ( n52292 , n52291 , n50557 );
and ( n52293 , n45963 , n50338 );
and ( n52294 , n45907 , n50336 );
nor ( n52295 , n52293 , n52294 );
xnor ( n52296 , n52295 , n50111 );
and ( n52297 , n52292 , n52296 );
and ( n52298 , n46100 , n49896 );
and ( n52299 , n46041 , n49894 );
nor ( n52300 , n52298 , n52299 );
xnor ( n52301 , n52300 , n49711 );
and ( n52302 , n52296 , n52301 );
and ( n52303 , n52292 , n52301 );
or ( n52304 , n52297 , n52302 , n52303 );
and ( n52305 , n46264 , n49513 );
and ( n52306 , n46169 , n49511 );
nor ( n52307 , n52305 , n52306 );
xnor ( n52308 , n52307 , n49310 );
and ( n52309 , n46445 , n49121 );
and ( n52310 , n46345 , n49119 );
nor ( n52311 , n52309 , n52310 );
xnor ( n52312 , n52311 , n48932 );
and ( n52313 , n52308 , n52312 );
and ( n52314 , n47962 , n47178 );
and ( n52315 , n47778 , n47176 );
nor ( n52316 , n52314 , n52315 );
xnor ( n52317 , n52316 , n47039 );
and ( n52318 , n52312 , n52317 );
and ( n52319 , n52308 , n52317 );
or ( n52320 , n52313 , n52318 , n52319 );
and ( n52321 , n52304 , n52320 );
and ( n52322 , n48988 , n46496 );
and ( n52323 , n48709 , n46494 );
nor ( n52324 , n52322 , n52323 );
xnor ( n52325 , n52324 , n46402 );
and ( n52326 , n50625 , n45886 );
and ( n52327 , n50404 , n45884 );
nor ( n52328 , n52326 , n52327 );
xnor ( n52329 , n52328 , n45824 );
and ( n52330 , n52325 , n52329 );
buf ( n52331 , n20784 );
buf ( n52332 , n52331 );
and ( n52333 , n52332 , n20846 );
and ( n52334 , n52329 , n52333 );
and ( n52335 , n52325 , n52333 );
or ( n52336 , n52330 , n52334 , n52335 );
and ( n52337 , n52320 , n52336 );
and ( n52338 , n52304 , n52336 );
or ( n52339 , n52321 , n52337 , n52338 );
and ( n52340 , n52287 , n52339 );
and ( n52341 , n52246 , n52339 );
or ( n52342 , n52288 , n52340 , n52341 );
xor ( n52343 , n52009 , n52013 );
xor ( n52344 , n52343 , n52018 );
xor ( n52345 , n52025 , n52029 );
xor ( n52346 , n52345 , n52034 );
and ( n52347 , n52344 , n52346 );
xor ( n52348 , n52042 , n52046 );
xor ( n52349 , n52348 , n52051 );
and ( n52350 , n52346 , n52349 );
and ( n52351 , n52344 , n52349 );
or ( n52352 , n52347 , n52350 , n52351 );
buf ( n52353 , n51923 );
xor ( n52354 , n52353 , n51925 );
and ( n52355 , n52352 , n52354 );
xor ( n52356 , n51934 , n51935 );
xor ( n52357 , n52356 , n51952 );
and ( n52358 , n52354 , n52357 );
and ( n52359 , n52352 , n52357 );
or ( n52360 , n52355 , n52358 , n52359 );
and ( n52361 , n52342 , n52360 );
xor ( n52362 , n51971 , n51987 );
xor ( n52363 , n52362 , n51997 );
xor ( n52364 , n52021 , n52037 );
xor ( n52365 , n52364 , n52054 );
and ( n52366 , n52363 , n52365 );
xor ( n52367 , n52076 , n52091 );
xor ( n52368 , n52367 , n52094 );
and ( n52369 , n52365 , n52368 );
and ( n52370 , n52363 , n52368 );
or ( n52371 , n52366 , n52369 , n52370 );
and ( n52372 , n52360 , n52371 );
and ( n52373 , n52342 , n52371 );
or ( n52374 , n52361 , n52372 , n52373 );
and ( n52375 , n52200 , n52374 );
and ( n52376 , n52176 , n52374 );
or ( n52377 , n52201 , n52375 , n52376 );
xor ( n52378 , n51918 , n51920 );
xor ( n52379 , n52378 , n51927 );
xor ( n52380 , n51955 , n52000 );
xor ( n52381 , n52380 , n52057 );
and ( n52382 , n52379 , n52381 );
xor ( n52383 , n52097 , n52107 );
xor ( n52384 , n52383 , n52110 );
and ( n52385 , n52381 , n52384 );
and ( n52386 , n52379 , n52384 );
or ( n52387 , n52382 , n52385 , n52386 );
xor ( n52388 , n51913 , n51915 );
xor ( n52389 , n52388 , n51930 );
and ( n52390 , n52387 , n52389 );
xor ( n52391 , n52060 , n52113 );
xor ( n52392 , n52391 , n52124 );
and ( n52393 , n52389 , n52392 );
and ( n52394 , n52387 , n52392 );
or ( n52395 , n52390 , n52393 , n52394 );
and ( n52396 , n52377 , n52395 );
xor ( n52397 , n51933 , n52127 );
xor ( n52398 , n52397 , n52138 );
and ( n52399 , n52395 , n52398 );
and ( n52400 , n52377 , n52398 );
or ( n52401 , n52396 , n52399 , n52400 );
and ( n52402 , n52174 , n52401 );
xor ( n52403 , n52141 , n52151 );
xor ( n52404 , n52403 , n52154 );
and ( n52405 , n52401 , n52404 );
and ( n52406 , n52174 , n52404 );
or ( n52407 , n52402 , n52405 , n52406 );
and ( n52408 , n52172 , n52407 );
xor ( n52409 , n51908 , n51910 );
xor ( n52410 , n52409 , n52157 );
and ( n52411 , n52407 , n52410 );
and ( n52412 , n52172 , n52410 );
or ( n52413 , n52408 , n52411 , n52412 );
xor ( n52414 , n51906 , n52160 );
xor ( n52415 , n52414 , n52163 );
and ( n52416 , n52413 , n52415 );
xor ( n52417 , n52413 , n52415 );
xor ( n52418 , n52172 , n52407 );
xor ( n52419 , n52418 , n52410 );
xor ( n52420 , n52143 , n52145 );
xor ( n52421 , n52420 , n52148 );
xor ( n52422 , n52130 , n52132 );
xor ( n52423 , n52422 , n52135 );
xor ( n52424 , n52116 , n52118 );
xor ( n52425 , n52424 , n52121 );
xor ( n52426 , n52099 , n52101 );
xor ( n52427 , n52426 , n52104 );
xor ( n52428 , n52064 , n52068 );
xor ( n52429 , n52428 , n52073 );
xor ( n52430 , n52080 , n52083 );
xor ( n52431 , n52430 , n52088 );
and ( n52432 , n52429 , n52431 );
xnor ( n52433 , n52185 , n52187 );
and ( n52434 , n52431 , n52433 );
and ( n52435 , n52429 , n52433 );
or ( n52436 , n52432 , n52434 , n52435 );
and ( n52437 , n52427 , n52436 );
and ( n52438 , n46969 , n48394 );
and ( n52439 , n46843 , n48392 );
nor ( n52440 , n52438 , n52439 );
xnor ( n52441 , n52440 , n48220 );
and ( n52442 , n47216 , n48042 );
and ( n52443 , n47090 , n48040 );
nor ( n52444 , n52442 , n52443 );
xnor ( n52445 , n52444 , n47921 );
and ( n52446 , n52441 , n52445 );
and ( n52447 , n48384 , n46911 );
and ( n52448 , n48272 , n46909 );
nor ( n52449 , n52447 , n52448 );
xnor ( n52450 , n52449 , n46802 );
and ( n52451 , n52445 , n52450 );
and ( n52452 , n52441 , n52450 );
or ( n52453 , n52446 , n52451 , n52452 );
and ( n52454 , n52082 , n20852 );
and ( n52455 , n51734 , n20850 );
nor ( n52456 , n52454 , n52455 );
xnor ( n52457 , n52456 , n20860 );
or ( n52458 , n52453 , n52457 );
xor ( n52459 , n26635 , n45610 );
buf ( n52460 , n52459 );
buf ( n52461 , n52460 );
buf ( n52462 , n52461 );
xor ( n52463 , n52205 , n52209 );
xor ( n52464 , n52463 , n52214 );
and ( n52465 , n52462 , n52464 );
buf ( n52466 , n52465 );
and ( n52467 , n52458 , n52466 );
xor ( n52468 , n52221 , n52225 );
xor ( n52469 , n52468 , n52230 );
xnor ( n52470 , n52238 , n52242 );
and ( n52471 , n52469 , n52470 );
xnor ( n52472 , n52250 , n52254 );
and ( n52473 , n52470 , n52472 );
and ( n52474 , n52469 , n52472 );
or ( n52475 , n52471 , n52473 , n52474 );
and ( n52476 , n52466 , n52475 );
and ( n52477 , n52458 , n52475 );
or ( n52478 , n52467 , n52476 , n52477 );
and ( n52479 , n52436 , n52478 );
and ( n52480 , n52427 , n52478 );
or ( n52481 , n52437 , n52479 , n52480 );
and ( n52482 , n52425 , n52481 );
xor ( n52483 , n52259 , n52263 );
and ( n52484 , n49976 , n46135 );
and ( n52485 , n49781 , n46133 );
nor ( n52486 , n52484 , n52485 );
xnor ( n52487 , n52486 , n46067 );
and ( n52488 , n50726 , n45886 );
and ( n52489 , n50625 , n45884 );
nor ( n52490 , n52488 , n52489 );
xnor ( n52491 , n52490 , n45824 );
and ( n52492 , n52487 , n52491 );
and ( n52493 , n51734 , n45702 );
and ( n52494 , n51510 , n45700 );
nor ( n52495 , n52493 , n52494 );
xnor ( n52496 , n52495 , n20841 );
and ( n52497 , n52491 , n52496 );
and ( n52498 , n52487 , n52496 );
or ( n52499 , n52492 , n52497 , n52498 );
and ( n52500 , n52483 , n52499 );
and ( n52501 , n46750 , n48740 );
and ( n52502 , n46577 , n48738 );
nor ( n52503 , n52501 , n52502 );
xnor ( n52504 , n52503 , n48571 );
and ( n52505 , n47474 , n47734 );
and ( n52506 , n47351 , n47732 );
nor ( n52507 , n52505 , n52506 );
xnor ( n52508 , n52507 , n47606 );
or ( n52509 , n52504 , n52508 );
and ( n52510 , n52499 , n52509 );
and ( n52511 , n52483 , n52509 );
or ( n52512 , n52500 , n52510 , n52511 );
and ( n52513 , n48108 , n47178 );
and ( n52514 , n47962 , n47176 );
nor ( n52515 , n52513 , n52514 );
xnor ( n52516 , n52515 , n47039 );
and ( n52517 , n48709 , n46712 );
and ( n52518 , n48632 , n46710 );
nor ( n52519 , n52517 , n52518 );
xnor ( n52520 , n52519 , n46587 );
or ( n52521 , n52516 , n52520 );
and ( n52522 , n51298 , n45777 );
and ( n52523 , n51077 , n45775 );
nor ( n52524 , n52522 , n52523 );
xnor ( n52525 , n52524 , n45734 );
and ( n52526 , n52332 , n20852 );
and ( n52527 , n52082 , n20850 );
nor ( n52528 , n52526 , n52527 );
xnor ( n52529 , n52528 , n20860 );
and ( n52530 , n52525 , n52529 );
and ( n52531 , n52521 , n52530 );
buf ( n52532 , n17543 );
buf ( n52533 , n52532 );
buf ( n52534 , n17545 );
buf ( n52535 , n52534 );
and ( n52536 , n52533 , n52535 );
not ( n52537 , n52536 );
and ( n52538 , n52005 , n52537 );
not ( n52539 , n52538 );
and ( n52540 , n20844 , n52269 );
and ( n52541 , n20855 , n52267 );
nor ( n52542 , n52540 , n52541 );
xnor ( n52543 , n52542 , n52008 );
and ( n52544 , n52539 , n52543 );
and ( n52545 , n45712 , n51750 );
and ( n52546 , n20864 , n51748 );
nor ( n52547 , n52545 , n52546 );
xnor ( n52548 , n52547 , n51520 );
and ( n52549 , n52543 , n52548 );
and ( n52550 , n52539 , n52548 );
or ( n52551 , n52544 , n52549 , n52550 );
and ( n52552 , n52530 , n52551 );
and ( n52553 , n52521 , n52551 );
or ( n52554 , n52531 , n52552 , n52553 );
and ( n52555 , n52512 , n52554 );
and ( n52556 , n45794 , n51221 );
and ( n52557 , n45763 , n51219 );
nor ( n52558 , n52556 , n52557 );
xnor ( n52559 , n52558 , n51000 );
and ( n52560 , n45907 , n50783 );
and ( n52561 , n45843 , n50781 );
nor ( n52562 , n52560 , n52561 );
xnor ( n52563 , n52562 , n50557 );
and ( n52564 , n52559 , n52563 );
and ( n52565 , n46041 , n50338 );
and ( n52566 , n45963 , n50336 );
nor ( n52567 , n52565 , n52566 );
xnor ( n52568 , n52567 , n50111 );
and ( n52569 , n52563 , n52568 );
and ( n52570 , n52559 , n52568 );
or ( n52571 , n52564 , n52569 , n52570 );
and ( n52572 , n46169 , n49896 );
and ( n52573 , n46100 , n49894 );
nor ( n52574 , n52572 , n52573 );
xnor ( n52575 , n52574 , n49711 );
and ( n52576 , n46345 , n49513 );
and ( n52577 , n46264 , n49511 );
nor ( n52578 , n52576 , n52577 );
xnor ( n52579 , n52578 , n49310 );
and ( n52580 , n52575 , n52579 );
and ( n52581 , n46530 , n49121 );
and ( n52582 , n46445 , n49119 );
nor ( n52583 , n52581 , n52582 );
xnor ( n52584 , n52583 , n48932 );
and ( n52585 , n52579 , n52584 );
and ( n52586 , n52575 , n52584 );
or ( n52587 , n52580 , n52585 , n52586 );
and ( n52588 , n52571 , n52587 );
and ( n52589 , n47778 , n47429 );
and ( n52590 , n47647 , n47427 );
nor ( n52591 , n52589 , n52590 );
xnor ( n52592 , n52591 , n47309 );
and ( n52593 , n49115 , n46496 );
and ( n52594 , n48988 , n46494 );
nor ( n52595 , n52593 , n52594 );
xnor ( n52596 , n52595 , n46402 );
and ( n52597 , n52592 , n52596 );
and ( n52598 , n49570 , n46306 );
and ( n52599 , n49374 , n46304 );
nor ( n52600 , n52598 , n52599 );
xnor ( n52601 , n52600 , n46228 );
and ( n52602 , n52596 , n52601 );
and ( n52603 , n52592 , n52601 );
or ( n52604 , n52597 , n52602 , n52603 );
and ( n52605 , n52587 , n52604 );
and ( n52606 , n52571 , n52604 );
or ( n52607 , n52588 , n52605 , n52606 );
and ( n52608 , n52554 , n52607 );
and ( n52609 , n52512 , n52607 );
or ( n52610 , n52555 , n52608 , n52609 );
buf ( n52611 , n20786 );
buf ( n52612 , n52611 );
and ( n52613 , n52612 , n20846 );
xor ( n52614 , n26756 , n45608 );
buf ( n52615 , n52614 );
buf ( n52616 , n52615 );
buf ( n52617 , n52616 );
and ( n52618 , n52613 , n52617 );
buf ( n52619 , n52618 );
xor ( n52620 , n52272 , n52276 );
xor ( n52621 , n52620 , n52281 );
and ( n52622 , n52619 , n52621 );
xor ( n52623 , n52292 , n52296 );
xor ( n52624 , n52623 , n52301 );
and ( n52625 , n52621 , n52624 );
and ( n52626 , n52619 , n52624 );
or ( n52627 , n52622 , n52625 , n52626 );
buf ( n52628 , n52191 );
xor ( n52629 , n52628 , n52192 );
and ( n52630 , n52627 , n52629 );
xor ( n52631 , n52217 , n52233 );
xor ( n52632 , n52631 , n52243 );
and ( n52633 , n52629 , n52632 );
and ( n52634 , n52627 , n52632 );
or ( n52635 , n52630 , n52633 , n52634 );
and ( n52636 , n52610 , n52635 );
xor ( n52637 , n52255 , n52264 );
xor ( n52638 , n52637 , n52284 );
xor ( n52639 , n52304 , n52320 );
xor ( n52640 , n52639 , n52336 );
and ( n52641 , n52638 , n52640 );
xor ( n52642 , n52344 , n52346 );
xor ( n52643 , n52642 , n52349 );
and ( n52644 , n52640 , n52643 );
and ( n52645 , n52638 , n52643 );
or ( n52646 , n52641 , n52644 , n52645 );
and ( n52647 , n52635 , n52646 );
and ( n52648 , n52610 , n52646 );
or ( n52649 , n52636 , n52647 , n52648 );
and ( n52650 , n52481 , n52649 );
and ( n52651 , n52425 , n52649 );
or ( n52652 , n52482 , n52650 , n52651 );
and ( n52653 , n52423 , n52652 );
xor ( n52654 , n52183 , n52188 );
xor ( n52655 , n52654 , n52194 );
xor ( n52656 , n52246 , n52287 );
xor ( n52657 , n52656 , n52339 );
and ( n52658 , n52655 , n52657 );
xor ( n52659 , n52352 , n52354 );
xor ( n52660 , n52659 , n52357 );
and ( n52661 , n52657 , n52660 );
and ( n52662 , n52655 , n52660 );
or ( n52663 , n52658 , n52661 , n52662 );
xor ( n52664 , n52178 , n52180 );
xor ( n52665 , n52664 , n52197 );
and ( n52666 , n52663 , n52665 );
xor ( n52667 , n52342 , n52360 );
xor ( n52668 , n52667 , n52371 );
and ( n52669 , n52665 , n52668 );
and ( n52670 , n52663 , n52668 );
or ( n52671 , n52666 , n52669 , n52670 );
and ( n52672 , n52652 , n52671 );
and ( n52673 , n52423 , n52671 );
or ( n52674 , n52653 , n52672 , n52673 );
and ( n52675 , n52421 , n52674 );
xor ( n52676 , n52377 , n52395 );
xor ( n52677 , n52676 , n52398 );
and ( n52678 , n52674 , n52677 );
and ( n52679 , n52421 , n52677 );
or ( n52680 , n52675 , n52678 , n52679 );
xor ( n52681 , n52174 , n52401 );
xor ( n52682 , n52681 , n52404 );
and ( n52683 , n52680 , n52682 );
xor ( n52684 , n52176 , n52200 );
xor ( n52685 , n52684 , n52374 );
xor ( n52686 , n52387 , n52389 );
xor ( n52687 , n52686 , n52392 );
and ( n52688 , n52685 , n52687 );
xor ( n52689 , n52379 , n52381 );
xor ( n52690 , n52689 , n52384 );
xor ( n52691 , n52363 , n52365 );
xor ( n52692 , n52691 , n52368 );
xor ( n52693 , n52308 , n52312 );
xor ( n52694 , n52693 , n52317 );
xor ( n52695 , n52325 , n52329 );
xor ( n52696 , n52695 , n52333 );
and ( n52697 , n52694 , n52696 );
xnor ( n52698 , n52453 , n52457 );
and ( n52699 , n52696 , n52698 );
and ( n52700 , n52694 , n52698 );
or ( n52701 , n52697 , n52699 , n52700 );
and ( n52702 , n47090 , n48394 );
and ( n52703 , n46969 , n48392 );
nor ( n52704 , n52702 , n52703 );
xnor ( n52705 , n52704 , n48220 );
and ( n52706 , n48272 , n47178 );
and ( n52707 , n48108 , n47176 );
nor ( n52708 , n52706 , n52707 );
xnor ( n52709 , n52708 , n47039 );
and ( n52710 , n52705 , n52709 );
and ( n52711 , n48988 , n46712 );
and ( n52712 , n48709 , n46710 );
nor ( n52713 , n52711 , n52712 );
xnor ( n52714 , n52713 , n46587 );
and ( n52715 , n52709 , n52714 );
and ( n52716 , n52705 , n52714 );
or ( n52717 , n52710 , n52715 , n52716 );
and ( n52718 , n50404 , n45990 );
and ( n52719 , n50195 , n45988 );
nor ( n52720 , n52718 , n52719 );
xnor ( n52721 , n52720 , n45939 );
or ( n52722 , n52717 , n52721 );
xor ( n52723 , n52441 , n52445 );
xor ( n52724 , n52723 , n52450 );
xor ( n52725 , n52487 , n52491 );
xor ( n52726 , n52725 , n52496 );
and ( n52727 , n52724 , n52726 );
xnor ( n52728 , n52504 , n52508 );
and ( n52729 , n52726 , n52728 );
and ( n52730 , n52724 , n52728 );
or ( n52731 , n52727 , n52729 , n52730 );
and ( n52732 , n52722 , n52731 );
xnor ( n52733 , n52516 , n52520 );
xor ( n52734 , n52525 , n52529 );
and ( n52735 , n52733 , n52734 );
and ( n52736 , n50625 , n45990 );
and ( n52737 , n50404 , n45988 );
nor ( n52738 , n52736 , n52737 );
xnor ( n52739 , n52738 , n45939 );
and ( n52740 , n51077 , n45886 );
and ( n52741 , n50726 , n45884 );
nor ( n52742 , n52740 , n52741 );
xnor ( n52743 , n52742 , n45824 );
and ( n52744 , n52739 , n52743 );
and ( n52745 , n52612 , n20852 );
and ( n52746 , n52332 , n20850 );
nor ( n52747 , n52745 , n52746 );
xnor ( n52748 , n52747 , n20860 );
and ( n52749 , n52743 , n52748 );
and ( n52750 , n52739 , n52748 );
or ( n52751 , n52744 , n52749 , n52750 );
and ( n52752 , n52734 , n52751 );
and ( n52753 , n52733 , n52751 );
or ( n52754 , n52735 , n52752 , n52753 );
and ( n52755 , n52731 , n52754 );
and ( n52756 , n52722 , n52754 );
or ( n52757 , n52732 , n52755 , n52756 );
and ( n52758 , n52701 , n52757 );
and ( n52759 , n49781 , n46306 );
and ( n52760 , n49570 , n46304 );
nor ( n52761 , n52759 , n52760 );
xnor ( n52762 , n52761 , n46228 );
and ( n52763 , n50195 , n46135 );
and ( n52764 , n49976 , n46133 );
nor ( n52765 , n52763 , n52764 );
xnor ( n52766 , n52765 , n46067 );
and ( n52767 , n52762 , n52766 );
and ( n52768 , n51510 , n45777 );
and ( n52769 , n51298 , n45775 );
nor ( n52770 , n52768 , n52769 );
xnor ( n52771 , n52770 , n45734 );
and ( n52772 , n52766 , n52771 );
and ( n52773 , n52762 , n52771 );
or ( n52774 , n52767 , n52772 , n52773 );
and ( n52775 , n47962 , n47429 );
and ( n52776 , n47778 , n47427 );
nor ( n52777 , n52775 , n52776 );
xnor ( n52778 , n52777 , n47309 );
and ( n52779 , n48632 , n46911 );
and ( n52780 , n48384 , n46909 );
nor ( n52781 , n52779 , n52780 );
xnor ( n52782 , n52781 , n46802 );
or ( n52783 , n52778 , n52782 );
and ( n52784 , n52774 , n52783 );
and ( n52785 , n47351 , n48042 );
and ( n52786 , n47216 , n48040 );
nor ( n52787 , n52785 , n52786 );
xnor ( n52788 , n52787 , n47921 );
buf ( n52789 , n20788 );
buf ( n52790 , n52789 );
and ( n52791 , n52790 , n20846 );
or ( n52792 , n52788 , n52791 );
and ( n52793 , n52783 , n52792 );
and ( n52794 , n52774 , n52792 );
or ( n52795 , n52784 , n52793 , n52794 );
xor ( n52796 , n52005 , n52533 );
xor ( n52797 , n52533 , n52535 );
not ( n52798 , n52797 );
and ( n52799 , n52796 , n52798 );
and ( n52800 , n20855 , n52799 );
not ( n52801 , n52800 );
xnor ( n52802 , n52801 , n52538 );
and ( n52803 , n20864 , n52269 );
and ( n52804 , n20844 , n52267 );
nor ( n52805 , n52803 , n52804 );
xnor ( n52806 , n52805 , n52008 );
and ( n52807 , n52802 , n52806 );
and ( n52808 , n45763 , n51750 );
and ( n52809 , n45712 , n51748 );
nor ( n52810 , n52808 , n52809 );
xnor ( n52811 , n52810 , n51520 );
and ( n52812 , n52806 , n52811 );
and ( n52813 , n52802 , n52811 );
or ( n52814 , n52807 , n52812 , n52813 );
and ( n52815 , n45843 , n51221 );
and ( n52816 , n45794 , n51219 );
nor ( n52817 , n52815 , n52816 );
xnor ( n52818 , n52817 , n51000 );
and ( n52819 , n45963 , n50783 );
and ( n52820 , n45907 , n50781 );
nor ( n52821 , n52819 , n52820 );
xnor ( n52822 , n52821 , n50557 );
and ( n52823 , n52818 , n52822 );
and ( n52824 , n46100 , n50338 );
and ( n52825 , n46041 , n50336 );
nor ( n52826 , n52824 , n52825 );
xnor ( n52827 , n52826 , n50111 );
and ( n52828 , n52822 , n52827 );
and ( n52829 , n52818 , n52827 );
or ( n52830 , n52823 , n52828 , n52829 );
and ( n52831 , n52814 , n52830 );
and ( n52832 , n46264 , n49896 );
and ( n52833 , n46169 , n49894 );
nor ( n52834 , n52832 , n52833 );
xnor ( n52835 , n52834 , n49711 );
and ( n52836 , n46445 , n49513 );
and ( n52837 , n46345 , n49511 );
nor ( n52838 , n52836 , n52837 );
xnor ( n52839 , n52838 , n49310 );
and ( n52840 , n52835 , n52839 );
and ( n52841 , n46577 , n49121 );
and ( n52842 , n46530 , n49119 );
nor ( n52843 , n52841 , n52842 );
xnor ( n52844 , n52843 , n48932 );
and ( n52845 , n52839 , n52844 );
and ( n52846 , n52835 , n52844 );
or ( n52847 , n52840 , n52845 , n52846 );
and ( n52848 , n52830 , n52847 );
and ( n52849 , n52814 , n52847 );
or ( n52850 , n52831 , n52848 , n52849 );
and ( n52851 , n52795 , n52850 );
and ( n52852 , n46843 , n48740 );
and ( n52853 , n46750 , n48738 );
nor ( n52854 , n52852 , n52853 );
xnor ( n52855 , n52854 , n48571 );
and ( n52856 , n47647 , n47734 );
and ( n52857 , n47474 , n47732 );
nor ( n52858 , n52856 , n52857 );
xnor ( n52859 , n52858 , n47606 );
and ( n52860 , n52855 , n52859 );
and ( n52861 , n49374 , n46496 );
and ( n52862 , n49115 , n46494 );
nor ( n52863 , n52861 , n52862 );
xnor ( n52864 , n52863 , n46402 );
and ( n52865 , n52859 , n52864 );
and ( n52866 , n52855 , n52864 );
or ( n52867 , n52860 , n52865 , n52866 );
and ( n52868 , n52082 , n45702 );
and ( n52869 , n51734 , n45700 );
nor ( n52870 , n52868 , n52869 );
xnor ( n52871 , n52870 , n20841 );
xor ( n52872 , n27474 , n45606 );
buf ( n52873 , n52872 );
buf ( n52874 , n52873 );
buf ( n52875 , n52874 );
and ( n52876 , n52871 , n52875 );
buf ( n52877 , n52876 );
and ( n52878 , n52867 , n52877 );
xor ( n52879 , n52539 , n52543 );
xor ( n52880 , n52879 , n52548 );
and ( n52881 , n52877 , n52880 );
and ( n52882 , n52867 , n52880 );
or ( n52883 , n52878 , n52881 , n52882 );
and ( n52884 , n52850 , n52883 );
and ( n52885 , n52795 , n52883 );
or ( n52886 , n52851 , n52884 , n52885 );
and ( n52887 , n52757 , n52886 );
and ( n52888 , n52701 , n52886 );
or ( n52889 , n52758 , n52887 , n52888 );
and ( n52890 , n52692 , n52889 );
xor ( n52891 , n52559 , n52563 );
xor ( n52892 , n52891 , n52568 );
xor ( n52893 , n52575 , n52579 );
xor ( n52894 , n52893 , n52584 );
and ( n52895 , n52892 , n52894 );
xor ( n52896 , n52592 , n52596 );
xor ( n52897 , n52896 , n52601 );
and ( n52898 , n52894 , n52897 );
and ( n52899 , n52892 , n52897 );
or ( n52900 , n52895 , n52898 , n52899 );
buf ( n52901 , n52462 );
xor ( n52902 , n52901 , n52464 );
and ( n52903 , n52900 , n52902 );
xor ( n52904 , n52469 , n52470 );
xor ( n52905 , n52904 , n52472 );
and ( n52906 , n52902 , n52905 );
and ( n52907 , n52900 , n52905 );
or ( n52908 , n52903 , n52906 , n52907 );
xor ( n52909 , n52483 , n52499 );
xor ( n52910 , n52909 , n52509 );
xor ( n52911 , n52521 , n52530 );
xor ( n52912 , n52911 , n52551 );
and ( n52913 , n52910 , n52912 );
xor ( n52914 , n52571 , n52587 );
xor ( n52915 , n52914 , n52604 );
and ( n52916 , n52912 , n52915 );
and ( n52917 , n52910 , n52915 );
or ( n52918 , n52913 , n52916 , n52917 );
and ( n52919 , n52908 , n52918 );
xor ( n52920 , n52429 , n52431 );
xor ( n52921 , n52920 , n52433 );
and ( n52922 , n52918 , n52921 );
and ( n52923 , n52908 , n52921 );
or ( n52924 , n52919 , n52922 , n52923 );
and ( n52925 , n52889 , n52924 );
and ( n52926 , n52692 , n52924 );
or ( n52927 , n52890 , n52925 , n52926 );
and ( n52928 , n52690 , n52927 );
xor ( n52929 , n52458 , n52466 );
xor ( n52930 , n52929 , n52475 );
xor ( n52931 , n52512 , n52554 );
xor ( n52932 , n52931 , n52607 );
and ( n52933 , n52930 , n52932 );
xor ( n52934 , n52627 , n52629 );
xor ( n52935 , n52934 , n52632 );
and ( n52936 , n52932 , n52935 );
and ( n52937 , n52930 , n52935 );
or ( n52938 , n52933 , n52936 , n52937 );
xor ( n52939 , n52427 , n52436 );
xor ( n52940 , n52939 , n52478 );
and ( n52941 , n52938 , n52940 );
xor ( n52942 , n52610 , n52635 );
xor ( n52943 , n52942 , n52646 );
and ( n52944 , n52940 , n52943 );
and ( n52945 , n52938 , n52943 );
or ( n52946 , n52941 , n52944 , n52945 );
and ( n52947 , n52927 , n52946 );
and ( n52948 , n52690 , n52946 );
or ( n52949 , n52928 , n52947 , n52948 );
and ( n52950 , n52687 , n52949 );
and ( n52951 , n52685 , n52949 );
or ( n52952 , n52688 , n52950 , n52951 );
xor ( n52953 , n52421 , n52674 );
xor ( n52954 , n52953 , n52677 );
and ( n52955 , n52952 , n52954 );
xor ( n52956 , n52423 , n52652 );
xor ( n52957 , n52956 , n52671 );
xor ( n52958 , n52425 , n52481 );
xor ( n52959 , n52958 , n52649 );
xor ( n52960 , n52663 , n52665 );
xor ( n52961 , n52960 , n52668 );
and ( n52962 , n52959 , n52961 );
xor ( n52963 , n52655 , n52657 );
xor ( n52964 , n52963 , n52660 );
xor ( n52965 , n52638 , n52640 );
xor ( n52966 , n52965 , n52643 );
xor ( n52967 , n52619 , n52621 );
xor ( n52968 , n52967 , n52624 );
xor ( n52969 , n52613 , n52617 );
buf ( n52970 , n52969 );
xnor ( n52971 , n52717 , n52721 );
and ( n52972 , n52970 , n52971 );
and ( n52973 , n49976 , n46306 );
and ( n52974 , n49781 , n46304 );
nor ( n52975 , n52973 , n52974 );
xnor ( n52976 , n52975 , n46228 );
and ( n52977 , n51298 , n45886 );
and ( n52978 , n51077 , n45884 );
nor ( n52979 , n52977 , n52978 );
xnor ( n52980 , n52979 , n45824 );
and ( n52981 , n52976 , n52980 );
and ( n52982 , n51734 , n45777 );
and ( n52983 , n51510 , n45775 );
nor ( n52984 , n52982 , n52983 );
xnor ( n52985 , n52984 , n45734 );
and ( n52986 , n52980 , n52985 );
and ( n52987 , n52976 , n52985 );
or ( n52988 , n52981 , n52986 , n52987 );
xor ( n52989 , n52762 , n52766 );
xor ( n52990 , n52989 , n52771 );
and ( n52991 , n52988 , n52990 );
and ( n52992 , n52971 , n52991 );
and ( n52993 , n52970 , n52991 );
or ( n52994 , n52972 , n52992 , n52993 );
and ( n52995 , n52968 , n52994 );
xor ( n52996 , n52705 , n52709 );
xor ( n52997 , n52996 , n52714 );
xor ( n52998 , n52739 , n52743 );
xor ( n52999 , n52998 , n52748 );
and ( n53000 , n52997 , n52999 );
xnor ( n53001 , n52778 , n52782 );
and ( n53002 , n52999 , n53001 );
and ( n53003 , n52997 , n53001 );
or ( n53004 , n53000 , n53002 , n53003 );
xnor ( n53005 , n52788 , n52791 );
and ( n53006 , n47216 , n48394 );
and ( n53007 , n47090 , n48392 );
nor ( n53008 , n53006 , n53007 );
xnor ( n53009 , n53008 , n48220 );
and ( n53010 , n48709 , n46911 );
and ( n53011 , n48632 , n46909 );
nor ( n53012 , n53010 , n53011 );
xnor ( n53013 , n53012 , n46802 );
and ( n53014 , n53009 , n53013 );
and ( n53015 , n49115 , n46712 );
and ( n53016 , n48988 , n46710 );
nor ( n53017 , n53015 , n53016 );
xnor ( n53018 , n53017 , n46587 );
and ( n53019 , n53013 , n53018 );
and ( n53020 , n53009 , n53018 );
or ( n53021 , n53014 , n53019 , n53020 );
and ( n53022 , n53005 , n53021 );
and ( n53023 , n52332 , n45702 );
and ( n53024 , n52082 , n45700 );
nor ( n53025 , n53023 , n53024 );
xnor ( n53026 , n53025 , n20841 );
and ( n53027 , n52790 , n20852 );
and ( n53028 , n52612 , n20850 );
nor ( n53029 , n53027 , n53028 );
xnor ( n53030 , n53029 , n20860 );
or ( n53031 , n53026 , n53030 );
and ( n53032 , n53021 , n53031 );
and ( n53033 , n53005 , n53031 );
or ( n53034 , n53022 , n53032 , n53033 );
and ( n53035 , n53004 , n53034 );
and ( n53036 , n48108 , n47429 );
and ( n53037 , n47962 , n47427 );
nor ( n53038 , n53036 , n53037 );
xnor ( n53039 , n53038 , n47309 );
buf ( n53040 , n20790 );
buf ( n53041 , n53040 );
and ( n53042 , n53041 , n20846 );
or ( n53043 , n53039 , n53042 );
and ( n53044 , n46969 , n48740 );
and ( n53045 , n46843 , n48738 );
nor ( n53046 , n53044 , n53045 );
xnor ( n53047 , n53046 , n48571 );
and ( n53048 , n47778 , n47734 );
and ( n53049 , n47647 , n47732 );
nor ( n53050 , n53048 , n53049 );
xnor ( n53051 , n53050 , n47606 );
or ( n53052 , n53047 , n53051 );
and ( n53053 , n53043 , n53052 );
buf ( n53054 , n17547 );
buf ( n53055 , n53054 );
buf ( n53056 , n17549 );
buf ( n53057 , n53056 );
and ( n53058 , n53055 , n53057 );
not ( n53059 , n53058 );
and ( n53060 , n52535 , n53059 );
not ( n53061 , n53060 );
and ( n53062 , n20844 , n52799 );
and ( n53063 , n20855 , n52797 );
nor ( n53064 , n53062 , n53063 );
xnor ( n53065 , n53064 , n52538 );
and ( n53066 , n53061 , n53065 );
and ( n53067 , n45712 , n52269 );
and ( n53068 , n20864 , n52267 );
nor ( n53069 , n53067 , n53068 );
xnor ( n53070 , n53069 , n52008 );
and ( n53071 , n53065 , n53070 );
and ( n53072 , n53061 , n53070 );
or ( n53073 , n53066 , n53071 , n53072 );
and ( n53074 , n53052 , n53073 );
and ( n53075 , n53043 , n53073 );
or ( n53076 , n53053 , n53074 , n53075 );
and ( n53077 , n53034 , n53076 );
and ( n53078 , n53004 , n53076 );
or ( n53079 , n53035 , n53077 , n53078 );
and ( n53080 , n52994 , n53079 );
and ( n53081 , n52968 , n53079 );
or ( n53082 , n52995 , n53080 , n53081 );
and ( n53083 , n52966 , n53082 );
and ( n53084 , n45794 , n51750 );
and ( n53085 , n45763 , n51748 );
nor ( n53086 , n53084 , n53085 );
xnor ( n53087 , n53086 , n51520 );
and ( n53088 , n45907 , n51221 );
and ( n53089 , n45843 , n51219 );
nor ( n53090 , n53088 , n53089 );
xnor ( n53091 , n53090 , n51000 );
and ( n53092 , n53087 , n53091 );
and ( n53093 , n46041 , n50783 );
and ( n53094 , n45963 , n50781 );
nor ( n53095 , n53093 , n53094 );
xnor ( n53096 , n53095 , n50557 );
and ( n53097 , n53091 , n53096 );
and ( n53098 , n53087 , n53096 );
or ( n53099 , n53092 , n53097 , n53098 );
and ( n53100 , n46169 , n50338 );
and ( n53101 , n46100 , n50336 );
nor ( n53102 , n53100 , n53101 );
xnor ( n53103 , n53102 , n50111 );
and ( n53104 , n46345 , n49896 );
and ( n53105 , n46264 , n49894 );
nor ( n53106 , n53104 , n53105 );
xnor ( n53107 , n53106 , n49711 );
and ( n53108 , n53103 , n53107 );
and ( n53109 , n46530 , n49513 );
and ( n53110 , n46445 , n49511 );
nor ( n53111 , n53109 , n53110 );
xnor ( n53112 , n53111 , n49310 );
and ( n53113 , n53107 , n53112 );
and ( n53114 , n53103 , n53112 );
or ( n53115 , n53108 , n53113 , n53114 );
and ( n53116 , n53099 , n53115 );
and ( n53117 , n46750 , n49121 );
and ( n53118 , n46577 , n49119 );
nor ( n53119 , n53117 , n53118 );
xnor ( n53120 , n53119 , n48932 );
and ( n53121 , n47474 , n48042 );
and ( n53122 , n47351 , n48040 );
nor ( n53123 , n53121 , n53122 );
xnor ( n53124 , n53123 , n47921 );
and ( n53125 , n53120 , n53124 );
and ( n53126 , n48384 , n47178 );
and ( n53127 , n48272 , n47176 );
nor ( n53128 , n53126 , n53127 );
xnor ( n53129 , n53128 , n47039 );
and ( n53130 , n53124 , n53129 );
and ( n53131 , n53120 , n53129 );
or ( n53132 , n53125 , n53130 , n53131 );
and ( n53133 , n53115 , n53132 );
and ( n53134 , n53099 , n53132 );
or ( n53135 , n53116 , n53133 , n53134 );
and ( n53136 , n49570 , n46496 );
and ( n53137 , n49374 , n46494 );
nor ( n53138 , n53136 , n53137 );
xnor ( n53139 , n53138 , n46402 );
and ( n53140 , n50404 , n46135 );
and ( n53141 , n50195 , n46133 );
nor ( n53142 , n53140 , n53141 );
xnor ( n53143 , n53142 , n46067 );
and ( n53144 , n53139 , n53143 );
xor ( n53145 , n28430 , n45604 );
buf ( n53146 , n53145 );
buf ( n53147 , n53146 );
buf ( n53148 , n53147 );
and ( n53149 , n53143 , n53148 );
and ( n53150 , n53139 , n53148 );
or ( n53151 , n53144 , n53149 , n53150 );
xor ( n53152 , n52802 , n52806 );
xor ( n53153 , n53152 , n52811 );
and ( n53154 , n53151 , n53153 );
xor ( n53155 , n52818 , n52822 );
xor ( n53156 , n53155 , n52827 );
and ( n53157 , n53153 , n53156 );
and ( n53158 , n53151 , n53156 );
or ( n53159 , n53154 , n53157 , n53158 );
and ( n53160 , n53135 , n53159 );
xor ( n53161 , n52835 , n52839 );
xor ( n53162 , n53161 , n52844 );
xor ( n53163 , n52855 , n52859 );
xor ( n53164 , n53163 , n52864 );
and ( n53165 , n53162 , n53164 );
xor ( n53166 , n52871 , n52875 );
buf ( n53167 , n53166 );
and ( n53168 , n53164 , n53167 );
and ( n53169 , n53162 , n53167 );
or ( n53170 , n53165 , n53168 , n53169 );
and ( n53171 , n53159 , n53170 );
and ( n53172 , n53135 , n53170 );
or ( n53173 , n53160 , n53171 , n53172 );
xor ( n53174 , n52724 , n52726 );
xor ( n53175 , n53174 , n52728 );
xor ( n53176 , n52733 , n52734 );
xor ( n53177 , n53176 , n52751 );
and ( n53178 , n53175 , n53177 );
xor ( n53179 , n52774 , n52783 );
xor ( n53180 , n53179 , n52792 );
and ( n53181 , n53177 , n53180 );
and ( n53182 , n53175 , n53180 );
or ( n53183 , n53178 , n53181 , n53182 );
and ( n53184 , n53173 , n53183 );
xor ( n53185 , n52814 , n52830 );
xor ( n53186 , n53185 , n52847 );
xor ( n53187 , n52867 , n52877 );
xor ( n53188 , n53187 , n52880 );
and ( n53189 , n53186 , n53188 );
xor ( n53190 , n52892 , n52894 );
xor ( n53191 , n53190 , n52897 );
and ( n53192 , n53188 , n53191 );
and ( n53193 , n53186 , n53191 );
or ( n53194 , n53189 , n53192 , n53193 );
and ( n53195 , n53183 , n53194 );
and ( n53196 , n53173 , n53194 );
or ( n53197 , n53184 , n53195 , n53196 );
and ( n53198 , n53082 , n53197 );
and ( n53199 , n52966 , n53197 );
or ( n53200 , n53083 , n53198 , n53199 );
and ( n53201 , n52964 , n53200 );
xor ( n53202 , n52694 , n52696 );
xor ( n53203 , n53202 , n52698 );
xor ( n53204 , n52722 , n52731 );
xor ( n53205 , n53204 , n52754 );
and ( n53206 , n53203 , n53205 );
xor ( n53207 , n52795 , n52850 );
xor ( n53208 , n53207 , n52883 );
and ( n53209 , n53205 , n53208 );
and ( n53210 , n53203 , n53208 );
or ( n53211 , n53206 , n53209 , n53210 );
xor ( n53212 , n52701 , n52757 );
xor ( n53213 , n53212 , n52886 );
and ( n53214 , n53211 , n53213 );
xor ( n53215 , n52908 , n52918 );
xor ( n53216 , n53215 , n52921 );
and ( n53217 , n53213 , n53216 );
and ( n53218 , n53211 , n53216 );
or ( n53219 , n53214 , n53217 , n53218 );
and ( n53220 , n53200 , n53219 );
and ( n53221 , n52964 , n53219 );
or ( n53222 , n53201 , n53220 , n53221 );
and ( n53223 , n52961 , n53222 );
and ( n53224 , n52959 , n53222 );
or ( n53225 , n52962 , n53223 , n53224 );
and ( n53226 , n52957 , n53225 );
xor ( n53227 , n52685 , n52687 );
xor ( n53228 , n53227 , n52949 );
and ( n53229 , n53225 , n53228 );
and ( n53230 , n52957 , n53228 );
or ( n53231 , n53226 , n53229 , n53230 );
and ( n53232 , n52954 , n53231 );
and ( n53233 , n52952 , n53231 );
or ( n53234 , n52955 , n53232 , n53233 );
and ( n53235 , n52682 , n53234 );
and ( n53236 , n52680 , n53234 );
or ( n53237 , n52683 , n53235 , n53236 );
and ( n53238 , n52419 , n53237 );
xor ( n53239 , n52419 , n53237 );
xor ( n53240 , n52680 , n52682 );
xor ( n53241 , n53240 , n53234 );
xor ( n53242 , n52952 , n52954 );
xor ( n53243 , n53242 , n53231 );
xor ( n53244 , n52690 , n52927 );
xor ( n53245 , n53244 , n52946 );
xor ( n53246 , n52692 , n52889 );
xor ( n53247 , n53246 , n52924 );
xor ( n53248 , n52938 , n52940 );
xor ( n53249 , n53248 , n52943 );
and ( n53250 , n53247 , n53249 );
xor ( n53251 , n52930 , n52932 );
xor ( n53252 , n53251 , n52935 );
xor ( n53253 , n52900 , n52902 );
xor ( n53254 , n53253 , n52905 );
xor ( n53255 , n52910 , n52912 );
xor ( n53256 , n53255 , n52915 );
and ( n53257 , n53254 , n53256 );
xor ( n53258 , n52988 , n52990 );
and ( n53259 , n48632 , n47178 );
and ( n53260 , n48384 , n47176 );
nor ( n53261 , n53259 , n53260 );
xnor ( n53262 , n53261 , n47039 );
and ( n53263 , n48988 , n46911 );
and ( n53264 , n48709 , n46909 );
nor ( n53265 , n53263 , n53264 );
xnor ( n53266 , n53265 , n46802 );
and ( n53267 , n53262 , n53266 );
and ( n53268 , n49374 , n46712 );
and ( n53269 , n49115 , n46710 );
nor ( n53270 , n53268 , n53269 );
xnor ( n53271 , n53270 , n46587 );
and ( n53272 , n53266 , n53271 );
and ( n53273 , n53262 , n53271 );
or ( n53274 , n53267 , n53272 , n53273 );
and ( n53275 , n50726 , n45990 );
and ( n53276 , n50625 , n45988 );
nor ( n53277 , n53275 , n53276 );
xnor ( n53278 , n53277 , n45939 );
and ( n53279 , n53274 , n53278 );
and ( n53280 , n53258 , n53279 );
xor ( n53281 , n52976 , n52980 );
xor ( n53282 , n53281 , n52985 );
xor ( n53283 , n53009 , n53013 );
xor ( n53284 , n53283 , n53018 );
and ( n53285 , n53282 , n53284 );
buf ( n53286 , n53285 );
and ( n53287 , n53279 , n53286 );
and ( n53288 , n53258 , n53286 );
or ( n53289 , n53280 , n53287 , n53288 );
xnor ( n53290 , n53026 , n53030 );
xnor ( n53291 , n53039 , n53042 );
and ( n53292 , n53290 , n53291 );
xnor ( n53293 , n53047 , n53051 );
and ( n53294 , n53291 , n53293 );
and ( n53295 , n53290 , n53293 );
or ( n53296 , n53292 , n53294 , n53295 );
and ( n53297 , n50195 , n46306 );
and ( n53298 , n49976 , n46304 );
nor ( n53299 , n53297 , n53298 );
xnor ( n53300 , n53299 , n46228 );
and ( n53301 , n50625 , n46135 );
and ( n53302 , n50404 , n46133 );
nor ( n53303 , n53301 , n53302 );
xnor ( n53304 , n53303 , n46067 );
and ( n53305 , n53300 , n53304 );
and ( n53306 , n52082 , n45777 );
and ( n53307 , n51734 , n45775 );
nor ( n53308 , n53306 , n53307 );
xnor ( n53309 , n53308 , n45734 );
and ( n53310 , n53304 , n53309 );
and ( n53311 , n53300 , n53309 );
or ( n53312 , n53305 , n53310 , n53311 );
and ( n53313 , n47090 , n48740 );
and ( n53314 , n46969 , n48738 );
nor ( n53315 , n53313 , n53314 );
xnor ( n53316 , n53315 , n48571 );
and ( n53317 , n47962 , n47734 );
and ( n53318 , n47778 , n47732 );
nor ( n53319 , n53317 , n53318 );
xnor ( n53320 , n53319 , n47606 );
or ( n53321 , n53316 , n53320 );
and ( n53322 , n53312 , n53321 );
and ( n53323 , n47351 , n48394 );
and ( n53324 , n47216 , n48392 );
nor ( n53325 , n53323 , n53324 );
xnor ( n53326 , n53325 , n48220 );
buf ( n53327 , n20792 );
buf ( n53328 , n53327 );
and ( n53329 , n53328 , n20846 );
or ( n53330 , n53326 , n53329 );
and ( n53331 , n53321 , n53330 );
and ( n53332 , n53312 , n53330 );
or ( n53333 , n53322 , n53331 , n53332 );
and ( n53334 , n53296 , n53333 );
and ( n53335 , n47647 , n48042 );
and ( n53336 , n47474 , n48040 );
nor ( n53337 , n53335 , n53336 );
xnor ( n53338 , n53337 , n47921 );
and ( n53339 , n48272 , n47429 );
and ( n53340 , n48108 , n47427 );
nor ( n53341 , n53339 , n53340 );
xnor ( n53342 , n53341 , n47309 );
or ( n53343 , n53338 , n53342 );
and ( n53344 , n51510 , n45886 );
and ( n53345 , n51298 , n45884 );
nor ( n53346 , n53344 , n53345 );
xnor ( n53347 , n53346 , n45824 );
and ( n53348 , n52612 , n45702 );
and ( n53349 , n52332 , n45700 );
nor ( n53350 , n53348 , n53349 );
xnor ( n53351 , n53350 , n20841 );
and ( n53352 , n53347 , n53351 );
and ( n53353 , n53343 , n53352 );
xor ( n53354 , n52535 , n53055 );
xor ( n53355 , n53055 , n53057 );
not ( n53356 , n53355 );
and ( n53357 , n53354 , n53356 );
and ( n53358 , n20855 , n53357 );
not ( n53359 , n53358 );
xnor ( n53360 , n53359 , n53060 );
and ( n53361 , n20864 , n52799 );
and ( n53362 , n20844 , n52797 );
nor ( n53363 , n53361 , n53362 );
xnor ( n53364 , n53363 , n52538 );
and ( n53365 , n53360 , n53364 );
and ( n53366 , n45763 , n52269 );
and ( n53367 , n45712 , n52267 );
nor ( n53368 , n53366 , n53367 );
xnor ( n53369 , n53368 , n52008 );
and ( n53370 , n53364 , n53369 );
and ( n53371 , n53360 , n53369 );
or ( n53372 , n53365 , n53370 , n53371 );
and ( n53373 , n53352 , n53372 );
and ( n53374 , n53343 , n53372 );
or ( n53375 , n53353 , n53373 , n53374 );
and ( n53376 , n53333 , n53375 );
and ( n53377 , n53296 , n53375 );
or ( n53378 , n53334 , n53376 , n53377 );
and ( n53379 , n53289 , n53378 );
and ( n53380 , n45843 , n51750 );
and ( n53381 , n45794 , n51748 );
nor ( n53382 , n53380 , n53381 );
xnor ( n53383 , n53382 , n51520 );
and ( n53384 , n45963 , n51221 );
and ( n53385 , n45907 , n51219 );
nor ( n53386 , n53384 , n53385 );
xnor ( n53387 , n53386 , n51000 );
and ( n53388 , n53383 , n53387 );
and ( n53389 , n46100 , n50783 );
and ( n53390 , n46041 , n50781 );
nor ( n53391 , n53389 , n53390 );
xnor ( n53392 , n53391 , n50557 );
and ( n53393 , n53387 , n53392 );
and ( n53394 , n53383 , n53392 );
or ( n53395 , n53388 , n53393 , n53394 );
and ( n53396 , n46264 , n50338 );
and ( n53397 , n46169 , n50336 );
nor ( n53398 , n53396 , n53397 );
xnor ( n53399 , n53398 , n50111 );
and ( n53400 , n46445 , n49896 );
and ( n53401 , n46345 , n49894 );
nor ( n53402 , n53400 , n53401 );
xnor ( n53403 , n53402 , n49711 );
and ( n53404 , n53399 , n53403 );
and ( n53405 , n46577 , n49513 );
and ( n53406 , n46530 , n49511 );
nor ( n53407 , n53405 , n53406 );
xnor ( n53408 , n53407 , n49310 );
and ( n53409 , n53403 , n53408 );
and ( n53410 , n53399 , n53408 );
or ( n53411 , n53404 , n53409 , n53410 );
and ( n53412 , n53395 , n53411 );
and ( n53413 , n46843 , n49121 );
and ( n53414 , n46750 , n49119 );
nor ( n53415 , n53413 , n53414 );
xnor ( n53416 , n53415 , n48932 );
and ( n53417 , n49781 , n46496 );
and ( n53418 , n49570 , n46494 );
nor ( n53419 , n53417 , n53418 );
xnor ( n53420 , n53419 , n46402 );
and ( n53421 , n53416 , n53420 );
xor ( n53422 , n28432 , n45603 );
buf ( n53423 , n53422 );
buf ( n53424 , n53423 );
buf ( n53425 , n53424 );
and ( n53426 , n53420 , n53425 );
and ( n53427 , n53416 , n53425 );
or ( n53428 , n53421 , n53426 , n53427 );
and ( n53429 , n53411 , n53428 );
and ( n53430 , n53395 , n53428 );
or ( n53431 , n53412 , n53429 , n53430 );
xor ( n53432 , n53061 , n53065 );
xor ( n53433 , n53432 , n53070 );
xor ( n53434 , n53087 , n53091 );
xor ( n53435 , n53434 , n53096 );
and ( n53436 , n53433 , n53435 );
xor ( n53437 , n53103 , n53107 );
xor ( n53438 , n53437 , n53112 );
and ( n53439 , n53435 , n53438 );
and ( n53440 , n53433 , n53438 );
or ( n53441 , n53436 , n53439 , n53440 );
and ( n53442 , n53431 , n53441 );
xor ( n53443 , n52997 , n52999 );
xor ( n53444 , n53443 , n53001 );
and ( n53445 , n53441 , n53444 );
and ( n53446 , n53431 , n53444 );
or ( n53447 , n53442 , n53445 , n53446 );
and ( n53448 , n53378 , n53447 );
and ( n53449 , n53289 , n53447 );
or ( n53450 , n53379 , n53448 , n53449 );
and ( n53451 , n53256 , n53450 );
and ( n53452 , n53254 , n53450 );
or ( n53453 , n53257 , n53451 , n53452 );
and ( n53454 , n53252 , n53453 );
xor ( n53455 , n53005 , n53021 );
xor ( n53456 , n53455 , n53031 );
xor ( n53457 , n53043 , n53052 );
xor ( n53458 , n53457 , n53073 );
and ( n53459 , n53456 , n53458 );
xor ( n53460 , n53099 , n53115 );
xor ( n53461 , n53460 , n53132 );
and ( n53462 , n53458 , n53461 );
and ( n53463 , n53456 , n53461 );
or ( n53464 , n53459 , n53462 , n53463 );
xor ( n53465 , n52970 , n52971 );
xor ( n53466 , n53465 , n52991 );
and ( n53467 , n53464 , n53466 );
xor ( n53468 , n53004 , n53034 );
xor ( n53469 , n53468 , n53076 );
and ( n53470 , n53466 , n53469 );
and ( n53471 , n53464 , n53469 );
or ( n53472 , n53467 , n53470 , n53471 );
xor ( n53473 , n53135 , n53159 );
xor ( n53474 , n53473 , n53170 );
xor ( n53475 , n53175 , n53177 );
xor ( n53476 , n53475 , n53180 );
and ( n53477 , n53474 , n53476 );
xor ( n53478 , n53186 , n53188 );
xor ( n53479 , n53478 , n53191 );
and ( n53480 , n53476 , n53479 );
and ( n53481 , n53474 , n53479 );
or ( n53482 , n53477 , n53480 , n53481 );
and ( n53483 , n53472 , n53482 );
xor ( n53484 , n52968 , n52994 );
xor ( n53485 , n53484 , n53079 );
and ( n53486 , n53482 , n53485 );
and ( n53487 , n53472 , n53485 );
or ( n53488 , n53483 , n53486 , n53487 );
and ( n53489 , n53453 , n53488 );
and ( n53490 , n53252 , n53488 );
or ( n53491 , n53454 , n53489 , n53490 );
and ( n53492 , n53249 , n53491 );
and ( n53493 , n53247 , n53491 );
or ( n53494 , n53250 , n53492 , n53493 );
and ( n53495 , n53245 , n53494 );
xor ( n53496 , n52959 , n52961 );
xor ( n53497 , n53496 , n53222 );
and ( n53498 , n53494 , n53497 );
and ( n53499 , n53245 , n53497 );
or ( n53500 , n53495 , n53498 , n53499 );
xor ( n53501 , n52957 , n53225 );
xor ( n53502 , n53501 , n53228 );
and ( n53503 , n53500 , n53502 );
xor ( n53504 , n52964 , n53200 );
xor ( n53505 , n53504 , n53219 );
xor ( n53506 , n52966 , n53082 );
xor ( n53507 , n53506 , n53197 );
xor ( n53508 , n53211 , n53213 );
xor ( n53509 , n53508 , n53216 );
and ( n53510 , n53507 , n53509 );
xor ( n53511 , n53173 , n53183 );
xor ( n53512 , n53511 , n53194 );
xor ( n53513 , n53203 , n53205 );
xor ( n53514 , n53513 , n53208 );
and ( n53515 , n53512 , n53514 );
xor ( n53516 , n53151 , n53153 );
xor ( n53517 , n53516 , n53156 );
xor ( n53518 , n53162 , n53164 );
xor ( n53519 , n53518 , n53167 );
and ( n53520 , n53517 , n53519 );
xor ( n53521 , n53120 , n53124 );
xor ( n53522 , n53521 , n53129 );
xor ( n53523 , n53139 , n53143 );
xor ( n53524 , n53523 , n53148 );
and ( n53525 , n53522 , n53524 );
xor ( n53526 , n53274 , n53278 );
and ( n53527 , n53524 , n53526 );
and ( n53528 , n53522 , n53526 );
or ( n53529 , n53525 , n53527 , n53528 );
and ( n53530 , n53519 , n53529 );
and ( n53531 , n53517 , n53529 );
or ( n53532 , n53520 , n53530 , n53531 );
and ( n53533 , n47216 , n48740 );
and ( n53534 , n47090 , n48738 );
nor ( n53535 , n53533 , n53534 );
xnor ( n53536 , n53535 , n48571 );
and ( n53537 , n48108 , n47734 );
and ( n53538 , n47962 , n47732 );
nor ( n53539 , n53537 , n53538 );
xnor ( n53540 , n53539 , n47606 );
and ( n53541 , n53536 , n53540 );
and ( n53542 , n49115 , n46911 );
and ( n53543 , n48988 , n46909 );
nor ( n53544 , n53542 , n53543 );
xnor ( n53545 , n53544 , n46802 );
and ( n53546 , n53540 , n53545 );
and ( n53547 , n53536 , n53545 );
or ( n53548 , n53541 , n53546 , n53547 );
and ( n53549 , n51077 , n45990 );
and ( n53550 , n50726 , n45988 );
nor ( n53551 , n53549 , n53550 );
xnor ( n53552 , n53551 , n45939 );
and ( n53553 , n53548 , n53552 );
and ( n53554 , n53041 , n20852 );
and ( n53555 , n52790 , n20850 );
nor ( n53556 , n53554 , n53555 );
xnor ( n53557 , n53556 , n20860 );
and ( n53558 , n53552 , n53557 );
and ( n53559 , n53548 , n53557 );
or ( n53560 , n53553 , n53558 , n53559 );
xor ( n53561 , n53262 , n53266 );
xor ( n53562 , n53561 , n53271 );
xnor ( n53563 , n53316 , n53320 );
and ( n53564 , n53562 , n53563 );
buf ( n53565 , n53564 );
and ( n53566 , n53560 , n53565 );
xnor ( n53567 , n53326 , n53329 );
xnor ( n53568 , n53338 , n53342 );
and ( n53569 , n53567 , n53568 );
xor ( n53570 , n53347 , n53351 );
and ( n53571 , n53568 , n53570 );
and ( n53572 , n53567 , n53570 );
or ( n53573 , n53569 , n53571 , n53572 );
and ( n53574 , n53565 , n53573 );
and ( n53575 , n53560 , n53573 );
or ( n53576 , n53566 , n53574 , n53575 );
and ( n53577 , n50404 , n46306 );
and ( n53578 , n50195 , n46304 );
nor ( n53579 , n53577 , n53578 );
xnor ( n53580 , n53579 , n46228 );
and ( n53581 , n52332 , n45777 );
and ( n53582 , n52082 , n45775 );
nor ( n53583 , n53581 , n53582 );
xnor ( n53584 , n53583 , n45734 );
and ( n53585 , n53580 , n53584 );
and ( n53586 , n52790 , n45702 );
and ( n53587 , n52612 , n45700 );
nor ( n53588 , n53586 , n53587 );
xnor ( n53589 , n53588 , n20841 );
and ( n53590 , n53584 , n53589 );
and ( n53591 , n53580 , n53589 );
or ( n53592 , n53585 , n53590 , n53591 );
and ( n53593 , n50726 , n46135 );
and ( n53594 , n50625 , n46133 );
nor ( n53595 , n53593 , n53594 );
xnor ( n53596 , n53595 , n46067 );
and ( n53597 , n51298 , n45990 );
and ( n53598 , n51077 , n45988 );
nor ( n53599 , n53597 , n53598 );
xnor ( n53600 , n53599 , n45939 );
or ( n53601 , n53596 , n53600 );
and ( n53602 , n53592 , n53601 );
and ( n53603 , n47778 , n48042 );
and ( n53604 , n47647 , n48040 );
nor ( n53605 , n53603 , n53604 );
xnor ( n53606 , n53605 , n47921 );
and ( n53607 , n48384 , n47429 );
and ( n53608 , n48272 , n47427 );
nor ( n53609 , n53607 , n53608 );
xnor ( n53610 , n53609 , n47309 );
or ( n53611 , n53606 , n53610 );
and ( n53612 , n53601 , n53611 );
and ( n53613 , n53592 , n53611 );
or ( n53614 , n53602 , n53612 , n53613 );
and ( n53615 , n48709 , n47178 );
and ( n53616 , n48632 , n47176 );
nor ( n53617 , n53615 , n53616 );
xnor ( n53618 , n53617 , n47039 );
and ( n53619 , n49570 , n46712 );
and ( n53620 , n49374 , n46710 );
nor ( n53621 , n53619 , n53620 );
xnor ( n53622 , n53621 , n46587 );
or ( n53623 , n53618 , n53622 );
and ( n53624 , n51734 , n45886 );
and ( n53625 , n51510 , n45884 );
nor ( n53626 , n53624 , n53625 );
xnor ( n53627 , n53626 , n45824 );
and ( n53628 , n53328 , n20852 );
and ( n53629 , n53041 , n20850 );
nor ( n53630 , n53628 , n53629 );
xnor ( n53631 , n53630 , n20860 );
or ( n53632 , n53627 , n53631 );
and ( n53633 , n53623 , n53632 );
and ( n53634 , n47474 , n48394 );
and ( n53635 , n47351 , n48392 );
nor ( n53636 , n53634 , n53635 );
xnor ( n53637 , n53636 , n48220 );
buf ( n53638 , n20794 );
buf ( n53639 , n53638 );
and ( n53640 , n53639 , n20846 );
and ( n53641 , n53637 , n53640 );
and ( n53642 , n53632 , n53641 );
and ( n53643 , n53623 , n53641 );
or ( n53644 , n53633 , n53642 , n53643 );
and ( n53645 , n53614 , n53644 );
buf ( n53646 , n17551 );
buf ( n53647 , n53646 );
buf ( n53648 , n17553 );
buf ( n53649 , n53648 );
and ( n53650 , n53647 , n53649 );
not ( n53651 , n53650 );
and ( n53652 , n53057 , n53651 );
not ( n53653 , n53652 );
and ( n53654 , n20844 , n53357 );
and ( n53655 , n20855 , n53355 );
nor ( n53656 , n53654 , n53655 );
xnor ( n53657 , n53656 , n53060 );
and ( n53658 , n53653 , n53657 );
and ( n53659 , n45712 , n52799 );
and ( n53660 , n20864 , n52797 );
nor ( n53661 , n53659 , n53660 );
xnor ( n53662 , n53661 , n52538 );
and ( n53663 , n53657 , n53662 );
and ( n53664 , n53653 , n53662 );
or ( n53665 , n53658 , n53663 , n53664 );
and ( n53666 , n45794 , n52269 );
and ( n53667 , n45763 , n52267 );
nor ( n53668 , n53666 , n53667 );
xnor ( n53669 , n53668 , n52008 );
and ( n53670 , n45907 , n51750 );
and ( n53671 , n45843 , n51748 );
nor ( n53672 , n53670 , n53671 );
xnor ( n53673 , n53672 , n51520 );
and ( n53674 , n53669 , n53673 );
and ( n53675 , n46041 , n51221 );
and ( n53676 , n45963 , n51219 );
nor ( n53677 , n53675 , n53676 );
xnor ( n53678 , n53677 , n51000 );
and ( n53679 , n53673 , n53678 );
and ( n53680 , n53669 , n53678 );
or ( n53681 , n53674 , n53679 , n53680 );
and ( n53682 , n53665 , n53681 );
and ( n53683 , n46169 , n50783 );
and ( n53684 , n46100 , n50781 );
nor ( n53685 , n53683 , n53684 );
xnor ( n53686 , n53685 , n50557 );
and ( n53687 , n46345 , n50338 );
and ( n53688 , n46264 , n50336 );
nor ( n53689 , n53687 , n53688 );
xnor ( n53690 , n53689 , n50111 );
and ( n53691 , n53686 , n53690 );
and ( n53692 , n46530 , n49896 );
and ( n53693 , n46445 , n49894 );
nor ( n53694 , n53692 , n53693 );
xnor ( n53695 , n53694 , n49711 );
and ( n53696 , n53690 , n53695 );
and ( n53697 , n53686 , n53695 );
or ( n53698 , n53691 , n53696 , n53697 );
and ( n53699 , n53681 , n53698 );
and ( n53700 , n53665 , n53698 );
or ( n53701 , n53682 , n53699 , n53700 );
and ( n53702 , n53644 , n53701 );
and ( n53703 , n53614 , n53701 );
or ( n53704 , n53645 , n53702 , n53703 );
and ( n53705 , n53576 , n53704 );
and ( n53706 , n46750 , n49513 );
and ( n53707 , n46577 , n49511 );
nor ( n53708 , n53706 , n53707 );
xnor ( n53709 , n53708 , n49310 );
and ( n53710 , n46969 , n49121 );
and ( n53711 , n46843 , n49119 );
nor ( n53712 , n53710 , n53711 );
xnor ( n53713 , n53712 , n48932 );
and ( n53714 , n53709 , n53713 );
and ( n53715 , n49976 , n46496 );
and ( n53716 , n49781 , n46494 );
nor ( n53717 , n53715 , n53716 );
xnor ( n53718 , n53717 , n46402 );
and ( n53719 , n53713 , n53718 );
and ( n53720 , n53709 , n53718 );
or ( n53721 , n53714 , n53719 , n53720 );
xor ( n53722 , n53360 , n53364 );
xor ( n53723 , n53722 , n53369 );
and ( n53724 , n53721 , n53723 );
xor ( n53725 , n53383 , n53387 );
xor ( n53726 , n53725 , n53392 );
and ( n53727 , n53723 , n53726 );
and ( n53728 , n53721 , n53726 );
or ( n53729 , n53724 , n53727 , n53728 );
buf ( n53730 , n53282 );
xor ( n53731 , n53730 , n53284 );
and ( n53732 , n53729 , n53731 );
xor ( n53733 , n53290 , n53291 );
xor ( n53734 , n53733 , n53293 );
and ( n53735 , n53731 , n53734 );
and ( n53736 , n53729 , n53734 );
or ( n53737 , n53732 , n53735 , n53736 );
and ( n53738 , n53704 , n53737 );
and ( n53739 , n53576 , n53737 );
or ( n53740 , n53705 , n53738 , n53739 );
and ( n53741 , n53532 , n53740 );
xor ( n53742 , n53312 , n53321 );
xor ( n53743 , n53742 , n53330 );
xor ( n53744 , n53343 , n53352 );
xor ( n53745 , n53744 , n53372 );
and ( n53746 , n53743 , n53745 );
xor ( n53747 , n53395 , n53411 );
xor ( n53748 , n53747 , n53428 );
and ( n53749 , n53745 , n53748 );
and ( n53750 , n53743 , n53748 );
or ( n53751 , n53746 , n53749 , n53750 );
xor ( n53752 , n53258 , n53279 );
xor ( n53753 , n53752 , n53286 );
and ( n53754 , n53751 , n53753 );
xor ( n53755 , n53296 , n53333 );
xor ( n53756 , n53755 , n53375 );
and ( n53757 , n53753 , n53756 );
and ( n53758 , n53751 , n53756 );
or ( n53759 , n53754 , n53757 , n53758 );
and ( n53760 , n53740 , n53759 );
and ( n53761 , n53532 , n53759 );
or ( n53762 , n53741 , n53760 , n53761 );
and ( n53763 , n53514 , n53762 );
and ( n53764 , n53512 , n53762 );
or ( n53765 , n53515 , n53763 , n53764 );
and ( n53766 , n53509 , n53765 );
and ( n53767 , n53507 , n53765 );
or ( n53768 , n53510 , n53766 , n53767 );
and ( n53769 , n53505 , n53768 );
xor ( n53770 , n53247 , n53249 );
xor ( n53771 , n53770 , n53491 );
and ( n53772 , n53768 , n53771 );
and ( n53773 , n53505 , n53771 );
or ( n53774 , n53769 , n53772 , n53773 );
xor ( n53775 , n53245 , n53494 );
xor ( n53776 , n53775 , n53497 );
and ( n53777 , n53774 , n53776 );
xor ( n53778 , n53289 , n53378 );
xor ( n53779 , n53778 , n53447 );
xor ( n53780 , n53464 , n53466 );
xor ( n53781 , n53780 , n53469 );
and ( n53782 , n53779 , n53781 );
xor ( n53783 , n53474 , n53476 );
xor ( n53784 , n53783 , n53479 );
and ( n53785 , n53781 , n53784 );
and ( n53786 , n53779 , n53784 );
or ( n53787 , n53782 , n53785 , n53786 );
xor ( n53788 , n53254 , n53256 );
xor ( n53789 , n53788 , n53450 );
and ( n53790 , n53787 , n53789 );
xor ( n53791 , n53472 , n53482 );
xor ( n53792 , n53791 , n53485 );
and ( n53793 , n53789 , n53792 );
and ( n53794 , n53787 , n53792 );
or ( n53795 , n53790 , n53793 , n53794 );
xor ( n53796 , n53252 , n53453 );
xor ( n53797 , n53796 , n53488 );
and ( n53798 , n53795 , n53797 );
xor ( n53799 , n53431 , n53441 );
xor ( n53800 , n53799 , n53444 );
xor ( n53801 , n53456 , n53458 );
xor ( n53802 , n53801 , n53461 );
and ( n53803 , n53800 , n53802 );
xor ( n53804 , n53433 , n53435 );
xor ( n53805 , n53804 , n53438 );
xor ( n53806 , n53300 , n53304 );
xor ( n53807 , n53806 , n53309 );
xor ( n53808 , n53548 , n53552 );
xor ( n53809 , n53808 , n53557 );
or ( n53810 , n53807 , n53809 );
and ( n53811 , n53805 , n53810 );
xor ( n53812 , n53399 , n53403 );
xor ( n53813 , n53812 , n53408 );
xor ( n53814 , n53416 , n53420 );
xor ( n53815 , n53814 , n53425 );
and ( n53816 , n53813 , n53815 );
and ( n53817 , n47962 , n48042 );
and ( n53818 , n47778 , n48040 );
nor ( n53819 , n53817 , n53818 );
xnor ( n53820 , n53819 , n47921 );
and ( n53821 , n48632 , n47429 );
and ( n53822 , n48384 , n47427 );
nor ( n53823 , n53821 , n53822 );
xnor ( n53824 , n53823 , n47309 );
and ( n53825 , n53820 , n53824 );
and ( n53826 , n49374 , n46911 );
and ( n53827 , n49115 , n46909 );
nor ( n53828 , n53826 , n53827 );
xnor ( n53829 , n53828 , n46802 );
and ( n53830 , n53824 , n53829 );
and ( n53831 , n53820 , n53829 );
or ( n53832 , n53825 , n53830 , n53831 );
xor ( n53833 , n53536 , n53540 );
xor ( n53834 , n53833 , n53545 );
or ( n53835 , n53832 , n53834 );
and ( n53836 , n53815 , n53835 );
and ( n53837 , n53813 , n53835 );
or ( n53838 , n53816 , n53836 , n53837 );
and ( n53839 , n53810 , n53838 );
and ( n53840 , n53805 , n53838 );
or ( n53841 , n53811 , n53839 , n53840 );
and ( n53842 , n53802 , n53841 );
and ( n53843 , n53800 , n53841 );
or ( n53844 , n53803 , n53842 , n53843 );
xor ( n53845 , n28433 , n45602 );
buf ( n53846 , n53845 );
buf ( n53847 , n53846 );
buf ( n53848 , n53847 );
xor ( n53849 , n53580 , n53584 );
xor ( n53850 , n53849 , n53589 );
and ( n53851 , n53848 , n53850 );
buf ( n53852 , n53851 );
xnor ( n53853 , n53596 , n53600 );
xnor ( n53854 , n53606 , n53610 );
and ( n53855 , n53853 , n53854 );
xnor ( n53856 , n53618 , n53622 );
and ( n53857 , n53854 , n53856 );
and ( n53858 , n53853 , n53856 );
or ( n53859 , n53855 , n53857 , n53858 );
and ( n53860 , n53852 , n53859 );
xnor ( n53861 , n53627 , n53631 );
xor ( n53862 , n53637 , n53640 );
and ( n53863 , n53861 , n53862 );
and ( n53864 , n50625 , n46306 );
and ( n53865 , n50404 , n46304 );
nor ( n53866 , n53864 , n53865 );
xnor ( n53867 , n53866 , n46228 );
and ( n53868 , n52082 , n45886 );
and ( n53869 , n51734 , n45884 );
nor ( n53870 , n53868 , n53869 );
xnor ( n53871 , n53870 , n45824 );
and ( n53872 , n53867 , n53871 );
and ( n53873 , n53041 , n45702 );
and ( n53874 , n52790 , n45700 );
nor ( n53875 , n53873 , n53874 );
xnor ( n53876 , n53875 , n20841 );
and ( n53877 , n53871 , n53876 );
and ( n53878 , n53867 , n53876 );
or ( n53879 , n53872 , n53877 , n53878 );
and ( n53880 , n53862 , n53879 );
and ( n53881 , n53861 , n53879 );
or ( n53882 , n53863 , n53880 , n53881 );
and ( n53883 , n53859 , n53882 );
and ( n53884 , n53852 , n53882 );
or ( n53885 , n53860 , n53883 , n53884 );
and ( n53886 , n46445 , n50338 );
and ( n53887 , n46345 , n50336 );
nor ( n53888 , n53886 , n53887 );
xnor ( n53889 , n53888 , n50111 );
and ( n53890 , n46577 , n49896 );
and ( n53891 , n46530 , n49894 );
nor ( n53892 , n53890 , n53891 );
xnor ( n53893 , n53892 , n49711 );
or ( n53894 , n53889 , n53893 );
and ( n53895 , n51077 , n46135 );
and ( n53896 , n50726 , n46133 );
nor ( n53897 , n53895 , n53896 );
xnor ( n53898 , n53897 , n46067 );
and ( n53899 , n52612 , n45777 );
and ( n53900 , n52332 , n45775 );
nor ( n53901 , n53899 , n53900 );
xnor ( n53902 , n53901 , n45734 );
or ( n53903 , n53898 , n53902 );
and ( n53904 , n53894 , n53903 );
and ( n53905 , n48988 , n47178 );
and ( n53906 , n48709 , n47176 );
nor ( n53907 , n53905 , n53906 );
xnor ( n53908 , n53907 , n47039 );
and ( n53909 , n49781 , n46712 );
and ( n53910 , n49570 , n46710 );
nor ( n53911 , n53909 , n53910 );
xnor ( n53912 , n53911 , n46587 );
or ( n53913 , n53908 , n53912 );
and ( n53914 , n53903 , n53913 );
and ( n53915 , n53894 , n53913 );
or ( n53916 , n53904 , n53914 , n53915 );
and ( n53917 , n47647 , n48394 );
and ( n53918 , n47474 , n48392 );
nor ( n53919 , n53917 , n53918 );
xnor ( n53920 , n53919 , n48220 );
buf ( n53921 , n20796 );
buf ( n53922 , n53921 );
and ( n53923 , n53922 , n20846 );
and ( n53924 , n53920 , n53923 );
xor ( n53925 , n53057 , n53647 );
xor ( n53926 , n53647 , n53649 );
not ( n53927 , n53926 );
and ( n53928 , n53925 , n53927 );
and ( n53929 , n20855 , n53928 );
not ( n53930 , n53929 );
xnor ( n53931 , n53930 , n53652 );
and ( n53932 , n20864 , n53357 );
and ( n53933 , n20844 , n53355 );
nor ( n53934 , n53932 , n53933 );
xnor ( n53935 , n53934 , n53060 );
and ( n53936 , n53931 , n53935 );
and ( n53937 , n45763 , n52799 );
and ( n53938 , n45712 , n52797 );
nor ( n53939 , n53937 , n53938 );
xnor ( n53940 , n53939 , n52538 );
and ( n53941 , n53935 , n53940 );
and ( n53942 , n53931 , n53940 );
or ( n53943 , n53936 , n53941 , n53942 );
and ( n53944 , n53924 , n53943 );
and ( n53945 , n45843 , n52269 );
and ( n53946 , n45794 , n52267 );
nor ( n53947 , n53945 , n53946 );
xnor ( n53948 , n53947 , n52008 );
and ( n53949 , n45963 , n51750 );
and ( n53950 , n45907 , n51748 );
nor ( n53951 , n53949 , n53950 );
xnor ( n53952 , n53951 , n51520 );
and ( n53953 , n53948 , n53952 );
and ( n53954 , n46100 , n51221 );
and ( n53955 , n46041 , n51219 );
nor ( n53956 , n53954 , n53955 );
xnor ( n53957 , n53956 , n51000 );
and ( n53958 , n53952 , n53957 );
and ( n53959 , n53948 , n53957 );
or ( n53960 , n53953 , n53958 , n53959 );
and ( n53961 , n53943 , n53960 );
and ( n53962 , n53924 , n53960 );
or ( n53963 , n53944 , n53961 , n53962 );
and ( n53964 , n53916 , n53963 );
and ( n53965 , n46264 , n50783 );
and ( n53966 , n46169 , n50781 );
nor ( n53967 , n53965 , n53966 );
xnor ( n53968 , n53967 , n50557 );
and ( n53969 , n46843 , n49513 );
and ( n53970 , n46750 , n49511 );
nor ( n53971 , n53969 , n53970 );
xnor ( n53972 , n53971 , n49310 );
and ( n53973 , n53968 , n53972 );
and ( n53974 , n47090 , n49121 );
and ( n53975 , n46969 , n49119 );
nor ( n53976 , n53974 , n53975 );
xnor ( n53977 , n53976 , n48932 );
and ( n53978 , n53972 , n53977 );
and ( n53979 , n53968 , n53977 );
or ( n53980 , n53973 , n53978 , n53979 );
and ( n53981 , n47351 , n48740 );
and ( n53982 , n47216 , n48738 );
nor ( n53983 , n53981 , n53982 );
xnor ( n53984 , n53983 , n48571 );
and ( n53985 , n48272 , n47734 );
and ( n53986 , n48108 , n47732 );
nor ( n53987 , n53985 , n53986 );
xnor ( n53988 , n53987 , n47606 );
and ( n53989 , n53984 , n53988 );
and ( n53990 , n50195 , n46496 );
and ( n53991 , n49976 , n46494 );
nor ( n53992 , n53990 , n53991 );
xnor ( n53993 , n53992 , n46402 );
and ( n53994 , n53988 , n53993 );
and ( n53995 , n53984 , n53993 );
or ( n53996 , n53989 , n53994 , n53995 );
and ( n53997 , n53980 , n53996 );
xor ( n53998 , n53653 , n53657 );
xor ( n53999 , n53998 , n53662 );
and ( n54000 , n53996 , n53999 );
and ( n54001 , n53980 , n53999 );
or ( n54002 , n53997 , n54000 , n54001 );
and ( n54003 , n53963 , n54002 );
and ( n54004 , n53916 , n54002 );
or ( n54005 , n53964 , n54003 , n54004 );
and ( n54006 , n53885 , n54005 );
xor ( n54007 , n53669 , n53673 );
xor ( n54008 , n54007 , n53678 );
xor ( n54009 , n53686 , n53690 );
xor ( n54010 , n54009 , n53695 );
and ( n54011 , n54008 , n54010 );
xor ( n54012 , n53709 , n53713 );
xor ( n54013 , n54012 , n53718 );
and ( n54014 , n54010 , n54013 );
and ( n54015 , n54008 , n54013 );
or ( n54016 , n54011 , n54014 , n54015 );
buf ( n54017 , n53562 );
xor ( n54018 , n54017 , n53563 );
and ( n54019 , n54016 , n54018 );
xor ( n54020 , n53567 , n53568 );
xor ( n54021 , n54020 , n53570 );
and ( n54022 , n54018 , n54021 );
and ( n54023 , n54016 , n54021 );
or ( n54024 , n54019 , n54022 , n54023 );
and ( n54025 , n54005 , n54024 );
and ( n54026 , n53885 , n54024 );
or ( n54027 , n54006 , n54025 , n54026 );
xor ( n54028 , n53592 , n53601 );
xor ( n54029 , n54028 , n53611 );
xor ( n54030 , n53623 , n53632 );
xor ( n54031 , n54030 , n53641 );
and ( n54032 , n54029 , n54031 );
xor ( n54033 , n53665 , n53681 );
xor ( n54034 , n54033 , n53698 );
and ( n54035 , n54031 , n54034 );
and ( n54036 , n54029 , n54034 );
or ( n54037 , n54032 , n54035 , n54036 );
xor ( n54038 , n53522 , n53524 );
xor ( n54039 , n54038 , n53526 );
and ( n54040 , n54037 , n54039 );
xor ( n54041 , n53560 , n53565 );
xor ( n54042 , n54041 , n53573 );
and ( n54043 , n54039 , n54042 );
and ( n54044 , n54037 , n54042 );
or ( n54045 , n54040 , n54043 , n54044 );
and ( n54046 , n54027 , n54045 );
xor ( n54047 , n53614 , n53644 );
xor ( n54048 , n54047 , n53701 );
xor ( n54049 , n53729 , n53731 );
xor ( n54050 , n54049 , n53734 );
and ( n54051 , n54048 , n54050 );
xor ( n54052 , n53743 , n53745 );
xor ( n54053 , n54052 , n53748 );
and ( n54054 , n54050 , n54053 );
and ( n54055 , n54048 , n54053 );
or ( n54056 , n54051 , n54054 , n54055 );
and ( n54057 , n54045 , n54056 );
and ( n54058 , n54027 , n54056 );
or ( n54059 , n54046 , n54057 , n54058 );
and ( n54060 , n53844 , n54059 );
xor ( n54061 , n53517 , n53519 );
xor ( n54062 , n54061 , n53529 );
xor ( n54063 , n53576 , n53704 );
xor ( n54064 , n54063 , n53737 );
and ( n54065 , n54062 , n54064 );
xor ( n54066 , n53751 , n53753 );
xor ( n54067 , n54066 , n53756 );
and ( n54068 , n54064 , n54067 );
and ( n54069 , n54062 , n54067 );
or ( n54070 , n54065 , n54068 , n54069 );
and ( n54071 , n54059 , n54070 );
and ( n54072 , n53844 , n54070 );
or ( n54073 , n54060 , n54071 , n54072 );
xor ( n54074 , n53512 , n53514 );
xor ( n54075 , n54074 , n53762 );
and ( n54076 , n54073 , n54075 );
xor ( n54077 , n53787 , n53789 );
xor ( n54078 , n54077 , n53792 );
and ( n54079 , n54075 , n54078 );
and ( n54080 , n54073 , n54078 );
or ( n54081 , n54076 , n54079 , n54080 );
and ( n54082 , n53797 , n54081 );
and ( n54083 , n53795 , n54081 );
or ( n54084 , n53798 , n54082 , n54083 );
xor ( n54085 , n53505 , n53768 );
xor ( n54086 , n54085 , n53771 );
and ( n54087 , n54084 , n54086 );
xor ( n54088 , n53507 , n53509 );
xor ( n54089 , n54088 , n53765 );
xor ( n54090 , n53795 , n53797 );
xor ( n54091 , n54090 , n54081 );
and ( n54092 , n54089 , n54091 );
xor ( n54093 , n53532 , n53740 );
xor ( n54094 , n54093 , n53759 );
xor ( n54095 , n53779 , n53781 );
xor ( n54096 , n54095 , n53784 );
and ( n54097 , n54094 , n54096 );
xor ( n54098 , n53721 , n53723 );
xor ( n54099 , n54098 , n53726 );
xnor ( n54100 , n53807 , n53809 );
and ( n54101 , n54099 , n54100 );
xnor ( n54102 , n53832 , n53834 );
and ( n54103 , n48108 , n48042 );
and ( n54104 , n47962 , n48040 );
nor ( n54105 , n54103 , n54104 );
xnor ( n54106 , n54105 , n47921 );
and ( n54107 , n48709 , n47429 );
and ( n54108 , n48632 , n47427 );
nor ( n54109 , n54107 , n54108 );
xnor ( n54110 , n54109 , n47309 );
and ( n54111 , n54106 , n54110 );
and ( n54112 , n49115 , n47178 );
and ( n54113 , n48988 , n47176 );
nor ( n54114 , n54112 , n54113 );
xnor ( n54115 , n54114 , n47039 );
and ( n54116 , n54110 , n54115 );
and ( n54117 , n54106 , n54115 );
or ( n54118 , n54111 , n54116 , n54117 );
and ( n54119 , n51510 , n45990 );
and ( n54120 , n51298 , n45988 );
nor ( n54121 , n54119 , n54120 );
xnor ( n54122 , n54121 , n45939 );
and ( n54123 , n54118 , n54122 );
and ( n54124 , n53639 , n20852 );
and ( n54125 , n53328 , n20850 );
nor ( n54126 , n54124 , n54125 );
xnor ( n54127 , n54126 , n20860 );
and ( n54128 , n54122 , n54127 );
and ( n54129 , n54118 , n54127 );
or ( n54130 , n54123 , n54128 , n54129 );
and ( n54131 , n54102 , n54130 );
and ( n54132 , n51298 , n46135 );
and ( n54133 , n51077 , n46133 );
nor ( n54134 , n54132 , n54133 );
xnor ( n54135 , n54134 , n46067 );
and ( n54136 , n52790 , n45777 );
and ( n54137 , n52612 , n45775 );
nor ( n54138 , n54136 , n54137 );
xnor ( n54139 , n54138 , n45734 );
and ( n54140 , n54135 , n54139 );
and ( n54141 , n53328 , n45702 );
and ( n54142 , n53041 , n45700 );
nor ( n54143 , n54141 , n54142 );
xnor ( n54144 , n54143 , n20841 );
and ( n54145 , n54139 , n54144 );
and ( n54146 , n54135 , n54144 );
or ( n54147 , n54140 , n54145 , n54146 );
xor ( n54148 , n53867 , n53871 );
xor ( n54149 , n54148 , n53876 );
or ( n54150 , n54147 , n54149 );
and ( n54151 , n54130 , n54150 );
and ( n54152 , n54102 , n54150 );
or ( n54153 , n54131 , n54151 , n54152 );
and ( n54154 , n54100 , n54153 );
and ( n54155 , n54099 , n54153 );
or ( n54156 , n54101 , n54154 , n54155 );
xor ( n54157 , n28436 , n45600 );
buf ( n54158 , n54157 );
buf ( n54159 , n54158 );
buf ( n54160 , n54159 );
xor ( n54161 , n53820 , n53824 );
xor ( n54162 , n54161 , n53829 );
and ( n54163 , n54160 , n54162 );
buf ( n54164 , n54163 );
xnor ( n54165 , n53889 , n53893 );
xnor ( n54166 , n53898 , n53902 );
and ( n54167 , n54165 , n54166 );
xnor ( n54168 , n53908 , n53912 );
and ( n54169 , n54166 , n54168 );
and ( n54170 , n54165 , n54168 );
or ( n54171 , n54167 , n54169 , n54170 );
and ( n54172 , n54164 , n54171 );
xor ( n54173 , n53920 , n53923 );
and ( n54174 , n47474 , n48740 );
and ( n54175 , n47351 , n48738 );
nor ( n54176 , n54174 , n54175 );
xnor ( n54177 , n54176 , n48571 );
and ( n54178 , n48384 , n47734 );
and ( n54179 , n48272 , n47732 );
nor ( n54180 , n54178 , n54179 );
xnor ( n54181 , n54180 , n47606 );
and ( n54182 , n54177 , n54181 );
and ( n54183 , n49976 , n46712 );
and ( n54184 , n49781 , n46710 );
nor ( n54185 , n54183 , n54184 );
xnor ( n54186 , n54185 , n46587 );
and ( n54187 , n54181 , n54186 );
and ( n54188 , n54177 , n54186 );
or ( n54189 , n54182 , n54187 , n54188 );
and ( n54190 , n54173 , n54189 );
and ( n54191 , n50726 , n46306 );
and ( n54192 , n50625 , n46304 );
nor ( n54193 , n54191 , n54192 );
xnor ( n54194 , n54193 , n46228 );
and ( n54195 , n52332 , n45886 );
and ( n54196 , n52082 , n45884 );
nor ( n54197 , n54195 , n54196 );
xnor ( n54198 , n54197 , n45824 );
and ( n54199 , n54194 , n54198 );
and ( n54200 , n53922 , n20852 );
and ( n54201 , n53639 , n20850 );
nor ( n54202 , n54200 , n54201 );
xnor ( n54203 , n54202 , n20860 );
and ( n54204 , n54198 , n54203 );
and ( n54205 , n54194 , n54203 );
or ( n54206 , n54199 , n54204 , n54205 );
and ( n54207 , n54189 , n54206 );
and ( n54208 , n54173 , n54206 );
or ( n54209 , n54190 , n54207 , n54208 );
and ( n54210 , n54171 , n54209 );
and ( n54211 , n54164 , n54209 );
or ( n54212 , n54172 , n54210 , n54211 );
and ( n54213 , n46530 , n50338 );
and ( n54214 , n46445 , n50336 );
nor ( n54215 , n54213 , n54214 );
xnor ( n54216 , n54215 , n50111 );
and ( n54217 , n46750 , n49896 );
and ( n54218 , n46577 , n49894 );
nor ( n54219 , n54217 , n54218 );
xnor ( n54220 , n54219 , n49711 );
or ( n54221 , n54216 , n54220 );
and ( n54222 , n49570 , n46911 );
and ( n54223 , n49374 , n46909 );
nor ( n54224 , n54222 , n54223 );
xnor ( n54225 , n54224 , n46802 );
buf ( n54226 , n20798 );
buf ( n54227 , n54226 );
and ( n54228 , n54227 , n20846 );
or ( n54229 , n54225 , n54228 );
and ( n54230 , n54221 , n54229 );
buf ( n54231 , n17555 );
buf ( n54232 , n54231 );
buf ( n54233 , n17557 );
buf ( n54234 , n54233 );
and ( n54235 , n54232 , n54234 );
not ( n54236 , n54235 );
and ( n54237 , n53649 , n54236 );
not ( n54238 , n54237 );
and ( n54239 , n20844 , n53928 );
and ( n54240 , n20855 , n53926 );
nor ( n54241 , n54239 , n54240 );
xnor ( n54242 , n54241 , n53652 );
and ( n54243 , n54238 , n54242 );
and ( n54244 , n45712 , n53357 );
and ( n54245 , n20864 , n53355 );
nor ( n54246 , n54244 , n54245 );
xnor ( n54247 , n54246 , n53060 );
and ( n54248 , n54242 , n54247 );
and ( n54249 , n54238 , n54247 );
or ( n54250 , n54243 , n54248 , n54249 );
and ( n54251 , n54229 , n54250 );
and ( n54252 , n54221 , n54250 );
or ( n54253 , n54230 , n54251 , n54252 );
and ( n54254 , n45794 , n52799 );
and ( n54255 , n45763 , n52797 );
nor ( n54256 , n54254 , n54255 );
xnor ( n54257 , n54256 , n52538 );
and ( n54258 , n45907 , n52269 );
and ( n54259 , n45843 , n52267 );
nor ( n54260 , n54258 , n54259 );
xnor ( n54261 , n54260 , n52008 );
and ( n54262 , n54257 , n54261 );
and ( n54263 , n46041 , n51750 );
and ( n54264 , n45963 , n51748 );
nor ( n54265 , n54263 , n54264 );
xnor ( n54266 , n54265 , n51520 );
and ( n54267 , n54261 , n54266 );
and ( n54268 , n54257 , n54266 );
or ( n54269 , n54262 , n54267 , n54268 );
and ( n54270 , n46169 , n51221 );
and ( n54271 , n46100 , n51219 );
nor ( n54272 , n54270 , n54271 );
xnor ( n54273 , n54272 , n51000 );
and ( n54274 , n46345 , n50783 );
and ( n54275 , n46264 , n50781 );
nor ( n54276 , n54274 , n54275 );
xnor ( n54277 , n54276 , n50557 );
and ( n54278 , n54273 , n54277 );
and ( n54279 , n46969 , n49513 );
and ( n54280 , n46843 , n49511 );
nor ( n54281 , n54279 , n54280 );
xnor ( n54282 , n54281 , n49310 );
and ( n54283 , n54277 , n54282 );
and ( n54284 , n54273 , n54282 );
or ( n54285 , n54278 , n54283 , n54284 );
and ( n54286 , n54269 , n54285 );
and ( n54287 , n47216 , n49121 );
and ( n54288 , n47090 , n49119 );
nor ( n54289 , n54287 , n54288 );
xnor ( n54290 , n54289 , n48932 );
and ( n54291 , n47778 , n48394 );
and ( n54292 , n47647 , n48392 );
nor ( n54293 , n54291 , n54292 );
xnor ( n54294 , n54293 , n48220 );
and ( n54295 , n54290 , n54294 );
and ( n54296 , n50404 , n46496 );
and ( n54297 , n50195 , n46494 );
nor ( n54298 , n54296 , n54297 );
xnor ( n54299 , n54298 , n46402 );
and ( n54300 , n54294 , n54299 );
and ( n54301 , n54290 , n54299 );
or ( n54302 , n54295 , n54300 , n54301 );
and ( n54303 , n54285 , n54302 );
and ( n54304 , n54269 , n54302 );
or ( n54305 , n54286 , n54303 , n54304 );
and ( n54306 , n54253 , n54305 );
and ( n54307 , n51734 , n45990 );
and ( n54308 , n51510 , n45988 );
nor ( n54309 , n54307 , n54308 );
xnor ( n54310 , n54309 , n45939 );
xor ( n54311 , n34201 , n45598 );
buf ( n54312 , n54311 );
buf ( n54313 , n54312 );
buf ( n54314 , n54313 );
and ( n54315 , n54310 , n54314 );
buf ( n54316 , n54315 );
xor ( n54317 , n53931 , n53935 );
xor ( n54318 , n54317 , n53940 );
and ( n54319 , n54316 , n54318 );
xor ( n54320 , n53948 , n53952 );
xor ( n54321 , n54320 , n53957 );
and ( n54322 , n54318 , n54321 );
and ( n54323 , n54316 , n54321 );
or ( n54324 , n54319 , n54322 , n54323 );
and ( n54325 , n54305 , n54324 );
and ( n54326 , n54253 , n54324 );
or ( n54327 , n54306 , n54325 , n54326 );
and ( n54328 , n54212 , n54327 );
buf ( n54329 , n53848 );
xor ( n54330 , n54329 , n53850 );
xor ( n54331 , n53853 , n53854 );
xor ( n54332 , n54331 , n53856 );
and ( n54333 , n54330 , n54332 );
xor ( n54334 , n53861 , n53862 );
xor ( n54335 , n54334 , n53879 );
and ( n54336 , n54332 , n54335 );
and ( n54337 , n54330 , n54335 );
or ( n54338 , n54333 , n54336 , n54337 );
and ( n54339 , n54327 , n54338 );
and ( n54340 , n54212 , n54338 );
or ( n54341 , n54328 , n54339 , n54340 );
and ( n54342 , n54156 , n54341 );
xor ( n54343 , n53894 , n53903 );
xor ( n54344 , n54343 , n53913 );
xor ( n54345 , n53924 , n53943 );
xor ( n54346 , n54345 , n53960 );
and ( n54347 , n54344 , n54346 );
xor ( n54348 , n53980 , n53996 );
xor ( n54349 , n54348 , n53999 );
and ( n54350 , n54346 , n54349 );
and ( n54351 , n54344 , n54349 );
or ( n54352 , n54347 , n54350 , n54351 );
xor ( n54353 , n53813 , n53815 );
xor ( n54354 , n54353 , n53835 );
and ( n54355 , n54352 , n54354 );
xor ( n54356 , n53852 , n53859 );
xor ( n54357 , n54356 , n53882 );
and ( n54358 , n54354 , n54357 );
and ( n54359 , n54352 , n54357 );
or ( n54360 , n54355 , n54358 , n54359 );
and ( n54361 , n54341 , n54360 );
and ( n54362 , n54156 , n54360 );
or ( n54363 , n54342 , n54361 , n54362 );
xor ( n54364 , n53916 , n53963 );
xor ( n54365 , n54364 , n54002 );
xor ( n54366 , n54016 , n54018 );
xor ( n54367 , n54366 , n54021 );
and ( n54368 , n54365 , n54367 );
xor ( n54369 , n54029 , n54031 );
xor ( n54370 , n54369 , n54034 );
and ( n54371 , n54367 , n54370 );
and ( n54372 , n54365 , n54370 );
or ( n54373 , n54368 , n54371 , n54372 );
xor ( n54374 , n53805 , n53810 );
xor ( n54375 , n54374 , n53838 );
and ( n54376 , n54373 , n54375 );
xor ( n54377 , n53885 , n54005 );
xor ( n54378 , n54377 , n54024 );
and ( n54379 , n54375 , n54378 );
and ( n54380 , n54373 , n54378 );
or ( n54381 , n54376 , n54379 , n54380 );
and ( n54382 , n54363 , n54381 );
xor ( n54383 , n53800 , n53802 );
xor ( n54384 , n54383 , n53841 );
and ( n54385 , n54381 , n54384 );
and ( n54386 , n54363 , n54384 );
or ( n54387 , n54382 , n54385 , n54386 );
and ( n54388 , n54096 , n54387 );
and ( n54389 , n54094 , n54387 );
or ( n54390 , n54097 , n54388 , n54389 );
xor ( n54391 , n54073 , n54075 );
xor ( n54392 , n54391 , n54078 );
and ( n54393 , n54390 , n54392 );
xor ( n54394 , n53844 , n54059 );
xor ( n54395 , n54394 , n54070 );
xor ( n54396 , n54027 , n54045 );
xor ( n54397 , n54396 , n54056 );
xor ( n54398 , n54062 , n54064 );
xor ( n54399 , n54398 , n54067 );
and ( n54400 , n54397 , n54399 );
xor ( n54401 , n54037 , n54039 );
xor ( n54402 , n54401 , n54042 );
xor ( n54403 , n54048 , n54050 );
xor ( n54404 , n54403 , n54053 );
and ( n54405 , n54402 , n54404 );
xor ( n54406 , n54008 , n54010 );
xor ( n54407 , n54406 , n54013 );
xor ( n54408 , n53968 , n53972 );
xor ( n54409 , n54408 , n53977 );
xor ( n54410 , n53984 , n53988 );
xor ( n54411 , n54410 , n53993 );
and ( n54412 , n54409 , n54411 );
xor ( n54413 , n54118 , n54122 );
xor ( n54414 , n54413 , n54127 );
and ( n54415 , n54411 , n54414 );
and ( n54416 , n54409 , n54414 );
or ( n54417 , n54412 , n54415 , n54416 );
and ( n54418 , n54407 , n54417 );
xnor ( n54419 , n54147 , n54149 );
xor ( n54420 , n54106 , n54110 );
xor ( n54421 , n54420 , n54115 );
xor ( n54422 , n54177 , n54181 );
xor ( n54423 , n54422 , n54186 );
or ( n54424 , n54421 , n54423 );
and ( n54425 , n54419 , n54424 );
and ( n54426 , n51077 , n46306 );
and ( n54427 , n50726 , n46304 );
nor ( n54428 , n54426 , n54427 );
xnor ( n54429 , n54428 , n46228 );
and ( n54430 , n52612 , n45886 );
and ( n54431 , n52332 , n45884 );
nor ( n54432 , n54430 , n54431 );
xnor ( n54433 , n54432 , n45824 );
and ( n54434 , n54429 , n54433 );
and ( n54435 , n53639 , n45702 );
and ( n54436 , n53328 , n45700 );
nor ( n54437 , n54435 , n54436 );
xnor ( n54438 , n54437 , n20841 );
and ( n54439 , n54433 , n54438 );
and ( n54440 , n54429 , n54438 );
or ( n54441 , n54434 , n54439 , n54440 );
xor ( n54442 , n54194 , n54198 );
xor ( n54443 , n54442 , n54203 );
or ( n54444 , n54441 , n54443 );
and ( n54445 , n54424 , n54444 );
and ( n54446 , n54419 , n54444 );
or ( n54447 , n54425 , n54445 , n54446 );
and ( n54448 , n54417 , n54447 );
and ( n54449 , n54407 , n54447 );
or ( n54450 , n54418 , n54448 , n54449 );
xor ( n54451 , n54135 , n54139 );
xor ( n54452 , n54451 , n54144 );
xnor ( n54453 , n54216 , n54220 );
and ( n54454 , n54452 , n54453 );
xnor ( n54455 , n54225 , n54228 );
and ( n54456 , n54453 , n54455 );
and ( n54457 , n54452 , n54455 );
or ( n54458 , n54454 , n54456 , n54457 );
and ( n54459 , n48272 , n48042 );
and ( n54460 , n48108 , n48040 );
nor ( n54461 , n54459 , n54460 );
xnor ( n54462 , n54461 , n47921 );
and ( n54463 , n49374 , n47178 );
and ( n54464 , n49115 , n47176 );
nor ( n54465 , n54463 , n54464 );
xnor ( n54466 , n54465 , n47039 );
and ( n54467 , n54462 , n54466 );
and ( n54468 , n49781 , n46911 );
and ( n54469 , n49570 , n46909 );
nor ( n54470 , n54468 , n54469 );
xnor ( n54471 , n54470 , n46802 );
and ( n54472 , n54466 , n54471 );
and ( n54473 , n54462 , n54471 );
or ( n54474 , n54467 , n54472 , n54473 );
and ( n54475 , n46264 , n51221 );
and ( n54476 , n46169 , n51219 );
nor ( n54477 , n54475 , n54476 );
xnor ( n54478 , n54477 , n51000 );
and ( n54479 , n46445 , n50783 );
and ( n54480 , n46345 , n50781 );
nor ( n54481 , n54479 , n54480 );
xnor ( n54482 , n54481 , n50557 );
or ( n54483 , n54478 , n54482 );
and ( n54484 , n54474 , n54483 );
and ( n54485 , n47962 , n48394 );
and ( n54486 , n47778 , n48392 );
nor ( n54487 , n54485 , n54486 );
xnor ( n54488 , n54487 , n48220 );
and ( n54489 , n50195 , n46712 );
and ( n54490 , n49976 , n46710 );
nor ( n54491 , n54489 , n54490 );
xnor ( n54492 , n54491 , n46587 );
or ( n54493 , n54488 , n54492 );
and ( n54494 , n54483 , n54493 );
and ( n54495 , n54474 , n54493 );
or ( n54496 , n54484 , n54494 , n54495 );
and ( n54497 , n54458 , n54496 );
and ( n54498 , n51510 , n46135 );
and ( n54499 , n51298 , n46133 );
nor ( n54500 , n54498 , n54499 );
xnor ( n54501 , n54500 , n46067 );
and ( n54502 , n52082 , n45990 );
and ( n54503 , n51734 , n45988 );
nor ( n54504 , n54502 , n54503 );
xnor ( n54505 , n54504 , n45939 );
or ( n54506 , n54501 , n54505 );
and ( n54507 , n47647 , n48740 );
and ( n54508 , n47474 , n48738 );
nor ( n54509 , n54507 , n54508 );
xnor ( n54510 , n54509 , n48571 );
and ( n54511 , n48632 , n47734 );
and ( n54512 , n48384 , n47732 );
nor ( n54513 , n54511 , n54512 );
xnor ( n54514 , n54513 , n47606 );
or ( n54515 , n54510 , n54514 );
and ( n54516 , n54506 , n54515 );
and ( n54517 , n53041 , n45777 );
and ( n54518 , n52790 , n45775 );
nor ( n54519 , n54517 , n54518 );
xnor ( n54520 , n54519 , n45734 );
and ( n54521 , n54227 , n20852 );
and ( n54522 , n53922 , n20850 );
nor ( n54523 , n54521 , n54522 );
xnor ( n54524 , n54523 , n20860 );
or ( n54525 , n54520 , n54524 );
and ( n54526 , n54515 , n54525 );
and ( n54527 , n54506 , n54525 );
or ( n54528 , n54516 , n54526 , n54527 );
and ( n54529 , n54496 , n54528 );
and ( n54530 , n54458 , n54528 );
or ( n54531 , n54497 , n54529 , n54530 );
xor ( n54532 , n53649 , n54232 );
xor ( n54533 , n54232 , n54234 );
not ( n54534 , n54533 );
and ( n54535 , n54532 , n54534 );
and ( n54536 , n20855 , n54535 );
not ( n54537 , n54536 );
xnor ( n54538 , n54537 , n54237 );
and ( n54539 , n20864 , n53928 );
and ( n54540 , n20844 , n53926 );
nor ( n54541 , n54539 , n54540 );
xnor ( n54542 , n54541 , n53652 );
and ( n54543 , n54538 , n54542 );
and ( n54544 , n45763 , n53357 );
and ( n54545 , n45712 , n53355 );
nor ( n54546 , n54544 , n54545 );
xnor ( n54547 , n54546 , n53060 );
and ( n54548 , n54542 , n54547 );
and ( n54549 , n54538 , n54547 );
or ( n54550 , n54543 , n54548 , n54549 );
and ( n54551 , n45843 , n52799 );
and ( n54552 , n45794 , n52797 );
nor ( n54553 , n54551 , n54552 );
xnor ( n54554 , n54553 , n52538 );
and ( n54555 , n45963 , n52269 );
and ( n54556 , n45907 , n52267 );
nor ( n54557 , n54555 , n54556 );
xnor ( n54558 , n54557 , n52008 );
and ( n54559 , n54554 , n54558 );
and ( n54560 , n46100 , n51750 );
and ( n54561 , n46041 , n51748 );
nor ( n54562 , n54560 , n54561 );
xnor ( n54563 , n54562 , n51520 );
and ( n54564 , n54558 , n54563 );
and ( n54565 , n54554 , n54563 );
or ( n54566 , n54559 , n54564 , n54565 );
and ( n54567 , n54550 , n54566 );
and ( n54568 , n46577 , n50338 );
and ( n54569 , n46530 , n50336 );
nor ( n54570 , n54568 , n54569 );
xnor ( n54571 , n54570 , n50111 );
and ( n54572 , n46843 , n49896 );
and ( n54573 , n46750 , n49894 );
nor ( n54574 , n54572 , n54573 );
xnor ( n54575 , n54574 , n49711 );
and ( n54576 , n54571 , n54575 );
and ( n54577 , n47090 , n49513 );
and ( n54578 , n46969 , n49511 );
nor ( n54579 , n54577 , n54578 );
xnor ( n54580 , n54579 , n49310 );
and ( n54581 , n54575 , n54580 );
and ( n54582 , n54571 , n54580 );
or ( n54583 , n54576 , n54581 , n54582 );
and ( n54584 , n54566 , n54583 );
and ( n54585 , n54550 , n54583 );
or ( n54586 , n54567 , n54584 , n54585 );
and ( n54587 , n47351 , n49121 );
and ( n54588 , n47216 , n49119 );
nor ( n54589 , n54587 , n54588 );
xnor ( n54590 , n54589 , n48932 );
and ( n54591 , n48988 , n47429 );
and ( n54592 , n48709 , n47427 );
nor ( n54593 , n54591 , n54592 );
xnor ( n54594 , n54593 , n47309 );
and ( n54595 , n54590 , n54594 );
and ( n54596 , n50625 , n46496 );
and ( n54597 , n50404 , n46494 );
nor ( n54598 , n54596 , n54597 );
xnor ( n54599 , n54598 , n46402 );
and ( n54600 , n54594 , n54599 );
and ( n54601 , n54590 , n54599 );
or ( n54602 , n54595 , n54600 , n54601 );
buf ( n54603 , n20800 );
buf ( n54604 , n54603 );
and ( n54605 , n54604 , n20846 );
xor ( n54606 , n34202 , n45597 );
buf ( n54607 , n54606 );
buf ( n54608 , n54607 );
buf ( n54609 , n54608 );
and ( n54610 , n54605 , n54609 );
buf ( n54611 , n54610 );
and ( n54612 , n54602 , n54611 );
xor ( n54613 , n54238 , n54242 );
xor ( n54614 , n54613 , n54247 );
and ( n54615 , n54611 , n54614 );
and ( n54616 , n54602 , n54614 );
or ( n54617 , n54612 , n54615 , n54616 );
and ( n54618 , n54586 , n54617 );
xor ( n54619 , n54257 , n54261 );
xor ( n54620 , n54619 , n54266 );
xor ( n54621 , n54273 , n54277 );
xor ( n54622 , n54621 , n54282 );
and ( n54623 , n54620 , n54622 );
xor ( n54624 , n54290 , n54294 );
xor ( n54625 , n54624 , n54299 );
and ( n54626 , n54622 , n54625 );
and ( n54627 , n54620 , n54625 );
or ( n54628 , n54623 , n54626 , n54627 );
and ( n54629 , n54617 , n54628 );
and ( n54630 , n54586 , n54628 );
or ( n54631 , n54618 , n54629 , n54630 );
and ( n54632 , n54531 , n54631 );
buf ( n54633 , n54160 );
xor ( n54634 , n54633 , n54162 );
xor ( n54635 , n54165 , n54166 );
xor ( n54636 , n54635 , n54168 );
and ( n54637 , n54634 , n54636 );
xor ( n54638 , n54173 , n54189 );
xor ( n54639 , n54638 , n54206 );
and ( n54640 , n54636 , n54639 );
and ( n54641 , n54634 , n54639 );
or ( n54642 , n54637 , n54640 , n54641 );
and ( n54643 , n54631 , n54642 );
and ( n54644 , n54531 , n54642 );
or ( n54645 , n54632 , n54643 , n54644 );
and ( n54646 , n54450 , n54645 );
xor ( n54647 , n54221 , n54229 );
xor ( n54648 , n54647 , n54250 );
xor ( n54649 , n54269 , n54285 );
xor ( n54650 , n54649 , n54302 );
and ( n54651 , n54648 , n54650 );
xor ( n54652 , n54316 , n54318 );
xor ( n54653 , n54652 , n54321 );
and ( n54654 , n54650 , n54653 );
and ( n54655 , n54648 , n54653 );
or ( n54656 , n54651 , n54654 , n54655 );
xor ( n54657 , n54102 , n54130 );
xor ( n54658 , n54657 , n54150 );
and ( n54659 , n54656 , n54658 );
xor ( n54660 , n54164 , n54171 );
xor ( n54661 , n54660 , n54209 );
and ( n54662 , n54658 , n54661 );
and ( n54663 , n54656 , n54661 );
or ( n54664 , n54659 , n54662 , n54663 );
and ( n54665 , n54645 , n54664 );
and ( n54666 , n54450 , n54664 );
or ( n54667 , n54646 , n54665 , n54666 );
and ( n54668 , n54404 , n54667 );
and ( n54669 , n54402 , n54667 );
or ( n54670 , n54405 , n54668 , n54669 );
and ( n54671 , n54399 , n54670 );
and ( n54672 , n54397 , n54670 );
or ( n54673 , n54400 , n54671 , n54672 );
and ( n54674 , n54395 , n54673 );
xor ( n54675 , n54094 , n54096 );
xor ( n54676 , n54675 , n54387 );
and ( n54677 , n54673 , n54676 );
and ( n54678 , n54395 , n54676 );
or ( n54679 , n54674 , n54677 , n54678 );
and ( n54680 , n54392 , n54679 );
and ( n54681 , n54390 , n54679 );
or ( n54682 , n54393 , n54680 , n54681 );
and ( n54683 , n54091 , n54682 );
and ( n54684 , n54089 , n54682 );
or ( n54685 , n54092 , n54683 , n54684 );
and ( n54686 , n54086 , n54685 );
and ( n54687 , n54084 , n54685 );
or ( n54688 , n54087 , n54686 , n54687 );
and ( n54689 , n53776 , n54688 );
and ( n54690 , n53774 , n54688 );
or ( n54691 , n53777 , n54689 , n54690 );
and ( n54692 , n53502 , n54691 );
and ( n54693 , n53500 , n54691 );
or ( n54694 , n53503 , n54692 , n54693 );
or ( n54695 , n53243 , n54694 );
and ( n54696 , n53241 , n54695 );
xor ( n54697 , n53241 , n54695 );
xnor ( n54698 , n53243 , n54694 );
xor ( n54699 , n53500 , n53502 );
xor ( n54700 , n54699 , n54691 );
xor ( n54701 , n53774 , n53776 );
xor ( n54702 , n54701 , n54688 );
not ( n54703 , n54702 );
xor ( n54704 , n54084 , n54086 );
xor ( n54705 , n54704 , n54685 );
xor ( n54706 , n54089 , n54091 );
xor ( n54707 , n54706 , n54682 );
xor ( n54708 , n54390 , n54392 );
xor ( n54709 , n54708 , n54679 );
xor ( n54710 , n54253 , n54305 );
xor ( n54711 , n54710 , n54324 );
xor ( n54712 , n54330 , n54332 );
xor ( n54713 , n54712 , n54335 );
and ( n54714 , n54711 , n54713 );
xor ( n54715 , n54344 , n54346 );
xor ( n54716 , n54715 , n54349 );
and ( n54717 , n54713 , n54716 );
and ( n54718 , n54711 , n54716 );
or ( n54719 , n54714 , n54717 , n54718 );
xor ( n54720 , n54099 , n54100 );
xor ( n54721 , n54720 , n54153 );
and ( n54722 , n54719 , n54721 );
xor ( n54723 , n54212 , n54327 );
xor ( n54724 , n54723 , n54338 );
and ( n54725 , n54721 , n54724 );
and ( n54726 , n54719 , n54724 );
or ( n54727 , n54722 , n54725 , n54726 );
xor ( n54728 , n54156 , n54341 );
xor ( n54729 , n54728 , n54360 );
and ( n54730 , n54727 , n54729 );
xor ( n54731 , n54373 , n54375 );
xor ( n54732 , n54731 , n54378 );
and ( n54733 , n54729 , n54732 );
and ( n54734 , n54727 , n54732 );
or ( n54735 , n54730 , n54733 , n54734 );
xor ( n54736 , n54363 , n54381 );
xor ( n54737 , n54736 , n54384 );
and ( n54738 , n54735 , n54737 );
xor ( n54739 , n54352 , n54354 );
xor ( n54740 , n54739 , n54357 );
xor ( n54741 , n54365 , n54367 );
xor ( n54742 , n54741 , n54370 );
and ( n54743 , n54740 , n54742 );
xor ( n54744 , n54310 , n54314 );
buf ( n54745 , n54744 );
xnor ( n54746 , n54421 , n54423 );
and ( n54747 , n54745 , n54746 );
xnor ( n54748 , n54441 , n54443 );
and ( n54749 , n54746 , n54748 );
and ( n54750 , n54745 , n54748 );
or ( n54751 , n54747 , n54749 , n54750 );
xnor ( n54752 , n54501 , n54505 );
xnor ( n54753 , n54510 , n54514 );
or ( n54754 , n54752 , n54753 );
and ( n54755 , n48709 , n47734 );
and ( n54756 , n48632 , n47732 );
nor ( n54757 , n54755 , n54756 );
xnor ( n54758 , n54757 , n47606 );
and ( n54759 , n49570 , n47178 );
and ( n54760 , n49374 , n47176 );
nor ( n54761 , n54759 , n54760 );
xnor ( n54762 , n54761 , n47039 );
and ( n54763 , n54758 , n54762 );
and ( n54764 , n49976 , n46911 );
and ( n54765 , n49781 , n46909 );
nor ( n54766 , n54764 , n54765 );
xnor ( n54767 , n54766 , n46802 );
and ( n54768 , n54762 , n54767 );
and ( n54769 , n54758 , n54767 );
or ( n54770 , n54763 , n54768 , n54769 );
xor ( n54771 , n54462 , n54466 );
xor ( n54772 , n54771 , n54471 );
or ( n54773 , n54770 , n54772 );
and ( n54774 , n54754 , n54773 );
xor ( n54775 , n54429 , n54433 );
xor ( n54776 , n54775 , n54438 );
xnor ( n54777 , n54478 , n54482 );
and ( n54778 , n54776 , n54777 );
xnor ( n54779 , n54488 , n54492 );
and ( n54780 , n54777 , n54779 );
and ( n54781 , n54776 , n54779 );
or ( n54782 , n54778 , n54780 , n54781 );
and ( n54783 , n54773 , n54782 );
and ( n54784 , n54754 , n54782 );
or ( n54785 , n54774 , n54783 , n54784 );
and ( n54786 , n54751 , n54785 );
xnor ( n54787 , n54520 , n54524 );
and ( n54788 , n51298 , n46306 );
and ( n54789 , n51077 , n46304 );
nor ( n54790 , n54788 , n54789 );
xnor ( n54791 , n54790 , n46228 );
and ( n54792 , n52332 , n45990 );
and ( n54793 , n52082 , n45988 );
nor ( n54794 , n54792 , n54793 );
xnor ( n54795 , n54794 , n45939 );
and ( n54796 , n54791 , n54795 );
and ( n54797 , n54604 , n20852 );
and ( n54798 , n54227 , n20850 );
nor ( n54799 , n54797 , n54798 );
xnor ( n54800 , n54799 , n20860 );
and ( n54801 , n54795 , n54800 );
and ( n54802 , n54791 , n54800 );
or ( n54803 , n54796 , n54801 , n54802 );
and ( n54804 , n54787 , n54803 );
and ( n54805 , n46750 , n50338 );
and ( n54806 , n46577 , n50336 );
nor ( n54807 , n54805 , n54806 );
xnor ( n54808 , n54807 , n50111 );
and ( n54809 , n46969 , n49896 );
and ( n54810 , n46843 , n49894 );
nor ( n54811 , n54809 , n54810 );
xnor ( n54812 , n54811 , n49711 );
or ( n54813 , n54808 , n54812 );
and ( n54814 , n54803 , n54813 );
and ( n54815 , n54787 , n54813 );
or ( n54816 , n54804 , n54814 , n54815 );
and ( n54817 , n51734 , n46135 );
and ( n54818 , n51510 , n46133 );
nor ( n54819 , n54817 , n54818 );
xnor ( n54820 , n54819 , n46067 );
and ( n54821 , n53922 , n45702 );
and ( n54822 , n53639 , n45700 );
nor ( n54823 , n54821 , n54822 );
xnor ( n54824 , n54823 , n20841 );
or ( n54825 , n54820 , n54824 );
and ( n54826 , n48108 , n48394 );
and ( n54827 , n47962 , n48392 );
nor ( n54828 , n54826 , n54827 );
xnor ( n54829 , n54828 , n48220 );
and ( n54830 , n50404 , n46712 );
and ( n54831 , n50195 , n46710 );
nor ( n54832 , n54830 , n54831 );
xnor ( n54833 , n54832 , n46587 );
or ( n54834 , n54829 , n54833 );
and ( n54835 , n54825 , n54834 );
and ( n54836 , n48384 , n48042 );
and ( n54837 , n48272 , n48040 );
nor ( n54838 , n54836 , n54837 );
xnor ( n54839 , n54838 , n47921 );
and ( n54840 , n49115 , n47429 );
and ( n54841 , n48988 , n47427 );
nor ( n54842 , n54840 , n54841 );
xnor ( n54843 , n54842 , n47309 );
or ( n54844 , n54839 , n54843 );
and ( n54845 , n54834 , n54844 );
and ( n54846 , n54825 , n54844 );
or ( n54847 , n54835 , n54845 , n54846 );
and ( n54848 , n54816 , n54847 );
and ( n54849 , n52790 , n45886 );
and ( n54850 , n52612 , n45884 );
nor ( n54851 , n54849 , n54850 );
xnor ( n54852 , n54851 , n45824 );
and ( n54853 , n53328 , n45777 );
and ( n54854 , n53041 , n45775 );
nor ( n54855 , n54853 , n54854 );
xnor ( n54856 , n54855 , n45734 );
and ( n54857 , n54852 , n54856 );
buf ( n54858 , n17559 );
buf ( n54859 , n54858 );
buf ( n54860 , n17561 );
buf ( n54861 , n54860 );
and ( n54862 , n54859 , n54861 );
not ( n54863 , n54862 );
and ( n54864 , n54234 , n54863 );
not ( n54865 , n54864 );
and ( n54866 , n20844 , n54535 );
and ( n54867 , n20855 , n54533 );
nor ( n54868 , n54866 , n54867 );
xnor ( n54869 , n54868 , n54237 );
and ( n54870 , n54865 , n54869 );
and ( n54871 , n45712 , n53928 );
and ( n54872 , n20864 , n53926 );
nor ( n54873 , n54871 , n54872 );
xnor ( n54874 , n54873 , n53652 );
and ( n54875 , n54869 , n54874 );
and ( n54876 , n54865 , n54874 );
or ( n54877 , n54870 , n54875 , n54876 );
and ( n54878 , n54857 , n54877 );
and ( n54879 , n45794 , n53357 );
and ( n54880 , n45763 , n53355 );
nor ( n54881 , n54879 , n54880 );
xnor ( n54882 , n54881 , n53060 );
and ( n54883 , n45907 , n52799 );
and ( n54884 , n45843 , n52797 );
nor ( n54885 , n54883 , n54884 );
xnor ( n54886 , n54885 , n52538 );
and ( n54887 , n54882 , n54886 );
and ( n54888 , n46041 , n52269 );
and ( n54889 , n45963 , n52267 );
nor ( n54890 , n54888 , n54889 );
xnor ( n54891 , n54890 , n52008 );
and ( n54892 , n54886 , n54891 );
and ( n54893 , n54882 , n54891 );
or ( n54894 , n54887 , n54892 , n54893 );
and ( n54895 , n54877 , n54894 );
and ( n54896 , n54857 , n54894 );
or ( n54897 , n54878 , n54895 , n54896 );
and ( n54898 , n54847 , n54897 );
and ( n54899 , n54816 , n54897 );
or ( n54900 , n54848 , n54898 , n54899 );
and ( n54901 , n54785 , n54900 );
and ( n54902 , n54751 , n54900 );
or ( n54903 , n54786 , n54901 , n54902 );
and ( n54904 , n46169 , n51750 );
and ( n54905 , n46100 , n51748 );
nor ( n54906 , n54904 , n54905 );
xnor ( n54907 , n54906 , n51520 );
and ( n54908 , n46345 , n51221 );
and ( n54909 , n46264 , n51219 );
nor ( n54910 , n54908 , n54909 );
xnor ( n54911 , n54910 , n51000 );
and ( n54912 , n54907 , n54911 );
and ( n54913 , n46530 , n50783 );
and ( n54914 , n46445 , n50781 );
nor ( n54915 , n54913 , n54914 );
xnor ( n54916 , n54915 , n50557 );
and ( n54917 , n54911 , n54916 );
and ( n54918 , n54907 , n54916 );
or ( n54919 , n54912 , n54917 , n54918 );
and ( n54920 , n47216 , n49513 );
and ( n54921 , n47090 , n49511 );
nor ( n54922 , n54920 , n54921 );
xnor ( n54923 , n54922 , n49310 );
and ( n54924 , n47474 , n49121 );
and ( n54925 , n47351 , n49119 );
nor ( n54926 , n54924 , n54925 );
xnor ( n54927 , n54926 , n48932 );
and ( n54928 , n54923 , n54927 );
and ( n54929 , n47778 , n48740 );
and ( n54930 , n47647 , n48738 );
nor ( n54931 , n54929 , n54930 );
xnor ( n54932 , n54931 , n48571 );
and ( n54933 , n54927 , n54932 );
and ( n54934 , n54923 , n54932 );
or ( n54935 , n54928 , n54933 , n54934 );
and ( n54936 , n54919 , n54935 );
and ( n54937 , n50726 , n46496 );
and ( n54938 , n50625 , n46494 );
nor ( n54939 , n54937 , n54938 );
xnor ( n54940 , n54939 , n46402 );
buf ( n54941 , n20802 );
buf ( n54942 , n54941 );
and ( n54943 , n54942 , n20846 );
and ( n54944 , n54940 , n54943 );
xor ( n54945 , n34203 , n45596 );
buf ( n54946 , n54945 );
buf ( n54947 , n54946 );
buf ( n54948 , n54947 );
and ( n54949 , n54943 , n54948 );
and ( n54950 , n54940 , n54948 );
or ( n54951 , n54944 , n54949 , n54950 );
and ( n54952 , n54935 , n54951 );
and ( n54953 , n54919 , n54951 );
or ( n54954 , n54936 , n54952 , n54953 );
xor ( n54955 , n54538 , n54542 );
xor ( n54956 , n54955 , n54547 );
xor ( n54957 , n54554 , n54558 );
xor ( n54958 , n54957 , n54563 );
and ( n54959 , n54956 , n54958 );
xor ( n54960 , n54571 , n54575 );
xor ( n54961 , n54960 , n54580 );
and ( n54962 , n54958 , n54961 );
and ( n54963 , n54956 , n54961 );
or ( n54964 , n54959 , n54962 , n54963 );
and ( n54965 , n54954 , n54964 );
xor ( n54966 , n54452 , n54453 );
xor ( n54967 , n54966 , n54455 );
and ( n54968 , n54964 , n54967 );
and ( n54969 , n54954 , n54967 );
or ( n54970 , n54965 , n54968 , n54969 );
xor ( n54971 , n54474 , n54483 );
xor ( n54972 , n54971 , n54493 );
xor ( n54973 , n54506 , n54515 );
xor ( n54974 , n54973 , n54525 );
and ( n54975 , n54972 , n54974 );
xor ( n54976 , n54550 , n54566 );
xor ( n54977 , n54976 , n54583 );
and ( n54978 , n54974 , n54977 );
and ( n54979 , n54972 , n54977 );
or ( n54980 , n54975 , n54978 , n54979 );
and ( n54981 , n54970 , n54980 );
xor ( n54982 , n54409 , n54411 );
xor ( n54983 , n54982 , n54414 );
and ( n54984 , n54980 , n54983 );
and ( n54985 , n54970 , n54983 );
or ( n54986 , n54981 , n54984 , n54985 );
and ( n54987 , n54903 , n54986 );
xor ( n54988 , n54419 , n54424 );
xor ( n54989 , n54988 , n54444 );
xor ( n54990 , n54458 , n54496 );
xor ( n54991 , n54990 , n54528 );
and ( n54992 , n54989 , n54991 );
xor ( n54993 , n54586 , n54617 );
xor ( n54994 , n54993 , n54628 );
and ( n54995 , n54991 , n54994 );
and ( n54996 , n54989 , n54994 );
or ( n54997 , n54992 , n54995 , n54996 );
and ( n54998 , n54986 , n54997 );
and ( n54999 , n54903 , n54997 );
or ( n55000 , n54987 , n54998 , n54999 );
and ( n55001 , n54742 , n55000 );
and ( n55002 , n54740 , n55000 );
or ( n55003 , n54743 , n55001 , n55002 );
xor ( n55004 , n54407 , n54417 );
xor ( n55005 , n55004 , n54447 );
xor ( n55006 , n54531 , n54631 );
xor ( n55007 , n55006 , n54642 );
and ( n55008 , n55005 , n55007 );
xor ( n55009 , n54656 , n54658 );
xor ( n55010 , n55009 , n54661 );
and ( n55011 , n55007 , n55010 );
and ( n55012 , n55005 , n55010 );
or ( n55013 , n55008 , n55011 , n55012 );
xor ( n55014 , n54450 , n54645 );
xor ( n55015 , n55014 , n54664 );
and ( n55016 , n55013 , n55015 );
xor ( n55017 , n54719 , n54721 );
xor ( n55018 , n55017 , n54724 );
and ( n55019 , n55015 , n55018 );
and ( n55020 , n55013 , n55018 );
or ( n55021 , n55016 , n55019 , n55020 );
and ( n55022 , n55003 , n55021 );
xor ( n55023 , n54402 , n54404 );
xor ( n55024 , n55023 , n54667 );
and ( n55025 , n55021 , n55024 );
and ( n55026 , n55003 , n55024 );
or ( n55027 , n55022 , n55025 , n55026 );
and ( n55028 , n54737 , n55027 );
and ( n55029 , n54735 , n55027 );
or ( n55030 , n54738 , n55028 , n55029 );
xor ( n55031 , n54395 , n54673 );
xor ( n55032 , n55031 , n54676 );
and ( n55033 , n55030 , n55032 );
xor ( n55034 , n54397 , n54399 );
xor ( n55035 , n55034 , n54670 );
xor ( n55036 , n54727 , n54729 );
xor ( n55037 , n55036 , n54732 );
xor ( n55038 , n54711 , n54713 );
xor ( n55039 , n55038 , n54716 );
xor ( n55040 , n54634 , n54636 );
xor ( n55041 , n55040 , n54639 );
xor ( n55042 , n54648 , n54650 );
xor ( n55043 , n55042 , n54653 );
and ( n55044 , n55041 , n55043 );
xor ( n55045 , n54602 , n54611 );
xor ( n55046 , n55045 , n54614 );
xor ( n55047 , n54620 , n54622 );
xor ( n55048 , n55047 , n54625 );
and ( n55049 , n55046 , n55048 );
xor ( n55050 , n54590 , n54594 );
xor ( n55051 , n55050 , n54599 );
xor ( n55052 , n54605 , n54609 );
buf ( n55053 , n55052 );
and ( n55054 , n55051 , n55053 );
xnor ( n55055 , n54752 , n54753 );
and ( n55056 , n55053 , n55055 );
and ( n55057 , n55051 , n55055 );
or ( n55058 , n55054 , n55056 , n55057 );
and ( n55059 , n55048 , n55058 );
and ( n55060 , n55046 , n55058 );
or ( n55061 , n55049 , n55059 , n55060 );
and ( n55062 , n55043 , n55061 );
and ( n55063 , n55041 , n55061 );
or ( n55064 , n55044 , n55062 , n55063 );
and ( n55065 , n55039 , n55064 );
xnor ( n55066 , n54770 , n54772 );
xor ( n55067 , n54758 , n54762 );
xor ( n55068 , n55067 , n54767 );
xor ( n55069 , n54791 , n54795 );
xor ( n55070 , n55069 , n54800 );
and ( n55071 , n55068 , n55070 );
buf ( n55072 , n55071 );
and ( n55073 , n55066 , n55072 );
xnor ( n55074 , n54808 , n54812 );
xnor ( n55075 , n54820 , n54824 );
and ( n55076 , n55074 , n55075 );
xnor ( n55077 , n54829 , n54833 );
and ( n55078 , n55075 , n55077 );
and ( n55079 , n55074 , n55077 );
or ( n55080 , n55076 , n55078 , n55079 );
and ( n55081 , n55072 , n55080 );
and ( n55082 , n55066 , n55080 );
or ( n55083 , n55073 , n55081 , n55082 );
xnor ( n55084 , n54839 , n54843 );
xor ( n55085 , n54852 , n54856 );
and ( n55086 , n55084 , n55085 );
and ( n55087 , n48272 , n48394 );
and ( n55088 , n48108 , n48392 );
nor ( n55089 , n55087 , n55088 );
xnor ( n55090 , n55089 , n48220 );
and ( n55091 , n48988 , n47734 );
and ( n55092 , n48709 , n47732 );
nor ( n55093 , n55091 , n55092 );
xnor ( n55094 , n55093 , n47606 );
and ( n55095 , n55090 , n55094 );
and ( n55096 , n49781 , n47178 );
and ( n55097 , n49570 , n47176 );
nor ( n55098 , n55096 , n55097 );
xnor ( n55099 , n55098 , n47039 );
and ( n55100 , n55094 , n55099 );
and ( n55101 , n55090 , n55099 );
or ( n55102 , n55095 , n55100 , n55101 );
and ( n55103 , n55085 , n55102 );
and ( n55104 , n55084 , n55102 );
or ( n55105 , n55086 , n55103 , n55104 );
and ( n55106 , n46264 , n51750 );
and ( n55107 , n46169 , n51748 );
nor ( n55108 , n55106 , n55107 );
xnor ( n55109 , n55108 , n51520 );
and ( n55110 , n46445 , n51221 );
and ( n55111 , n46345 , n51219 );
nor ( n55112 , n55110 , n55111 );
xnor ( n55113 , n55112 , n51000 );
or ( n55114 , n55109 , n55113 );
and ( n55115 , n53041 , n45886 );
and ( n55116 , n52790 , n45884 );
nor ( n55117 , n55115 , n55116 );
xnor ( n55118 , n55117 , n45824 );
and ( n55119 , n53639 , n45777 );
and ( n55120 , n53328 , n45775 );
nor ( n55121 , n55119 , n55120 );
xnor ( n55122 , n55121 , n45734 );
or ( n55123 , n55118 , n55122 );
and ( n55124 , n55114 , n55123 );
and ( n55125 , n51510 , n46306 );
and ( n55126 , n51298 , n46304 );
nor ( n55127 , n55125 , n55126 );
xnor ( n55128 , n55127 , n46228 );
and ( n55129 , n52612 , n45990 );
and ( n55130 , n52332 , n45988 );
nor ( n55131 , n55129 , n55130 );
xnor ( n55132 , n55131 , n45939 );
or ( n55133 , n55128 , n55132 );
and ( n55134 , n55123 , n55133 );
and ( n55135 , n55114 , n55133 );
or ( n55136 , n55124 , n55134 , n55135 );
and ( n55137 , n55105 , n55136 );
and ( n55138 , n54942 , n20852 );
and ( n55139 , n54604 , n20850 );
nor ( n55140 , n55138 , n55139 );
xnor ( n55141 , n55140 , n20860 );
buf ( n55142 , n20804 );
buf ( n55143 , n55142 );
and ( n55144 , n55143 , n20846 );
or ( n55145 , n55141 , n55144 );
and ( n55146 , n52082 , n46135 );
and ( n55147 , n51734 , n46133 );
nor ( n55148 , n55146 , n55147 );
xnor ( n55149 , n55148 , n46067 );
and ( n55150 , n54227 , n45702 );
and ( n55151 , n53922 , n45700 );
nor ( n55152 , n55150 , n55151 );
xnor ( n55153 , n55152 , n20841 );
or ( n55154 , n55149 , n55153 );
and ( n55155 , n55145 , n55154 );
xor ( n55156 , n54234 , n54859 );
xor ( n55157 , n54859 , n54861 );
not ( n55158 , n55157 );
and ( n55159 , n55156 , n55158 );
and ( n55160 , n20855 , n55159 );
not ( n55161 , n55160 );
xnor ( n55162 , n55161 , n54864 );
and ( n55163 , n20864 , n54535 );
and ( n55164 , n20844 , n54533 );
nor ( n55165 , n55163 , n55164 );
xnor ( n55166 , n55165 , n54237 );
and ( n55167 , n55162 , n55166 );
and ( n55168 , n45763 , n53928 );
and ( n55169 , n45712 , n53926 );
nor ( n55170 , n55168 , n55169 );
xnor ( n55171 , n55170 , n53652 );
and ( n55172 , n55166 , n55171 );
and ( n55173 , n55162 , n55171 );
or ( n55174 , n55167 , n55172 , n55173 );
and ( n55175 , n55154 , n55174 );
and ( n55176 , n55145 , n55174 );
or ( n55177 , n55155 , n55175 , n55176 );
and ( n55178 , n55136 , n55177 );
and ( n55179 , n55105 , n55177 );
or ( n55180 , n55137 , n55178 , n55179 );
and ( n55181 , n55083 , n55180 );
and ( n55182 , n45843 , n53357 );
and ( n55183 , n45794 , n53355 );
nor ( n55184 , n55182 , n55183 );
xnor ( n55185 , n55184 , n53060 );
and ( n55186 , n45963 , n52799 );
and ( n55187 , n45907 , n52797 );
nor ( n55188 , n55186 , n55187 );
xnor ( n55189 , n55188 , n52538 );
and ( n55190 , n55185 , n55189 );
and ( n55191 , n46100 , n52269 );
and ( n55192 , n46041 , n52267 );
nor ( n55193 , n55191 , n55192 );
xnor ( n55194 , n55193 , n52008 );
and ( n55195 , n55189 , n55194 );
and ( n55196 , n55185 , n55194 );
or ( n55197 , n55190 , n55195 , n55196 );
and ( n55198 , n46577 , n50783 );
and ( n55199 , n46530 , n50781 );
nor ( n55200 , n55198 , n55199 );
xnor ( n55201 , n55200 , n50557 );
and ( n55202 , n47090 , n49896 );
and ( n55203 , n46969 , n49894 );
nor ( n55204 , n55202 , n55203 );
xnor ( n55205 , n55204 , n49711 );
and ( n55206 , n55201 , n55205 );
and ( n55207 , n47351 , n49513 );
and ( n55208 , n47216 , n49511 );
nor ( n55209 , n55207 , n55208 );
xnor ( n55210 , n55209 , n49310 );
and ( n55211 , n55205 , n55210 );
and ( n55212 , n55201 , n55210 );
or ( n55213 , n55206 , n55211 , n55212 );
and ( n55214 , n55197 , n55213 );
and ( n55215 , n47647 , n49121 );
and ( n55216 , n47474 , n49119 );
nor ( n55217 , n55215 , n55216 );
xnor ( n55218 , n55217 , n48932 );
and ( n55219 , n47962 , n48740 );
and ( n55220 , n47778 , n48738 );
nor ( n55221 , n55219 , n55220 );
xnor ( n55222 , n55221 , n48571 );
and ( n55223 , n55218 , n55222 );
and ( n55224 , n48632 , n48042 );
and ( n55225 , n48384 , n48040 );
nor ( n55226 , n55224 , n55225 );
xnor ( n55227 , n55226 , n47921 );
and ( n55228 , n55222 , n55227 );
and ( n55229 , n55218 , n55227 );
or ( n55230 , n55223 , n55228 , n55229 );
and ( n55231 , n55213 , n55230 );
and ( n55232 , n55197 , n55230 );
or ( n55233 , n55214 , n55231 , n55232 );
and ( n55234 , n49374 , n47429 );
and ( n55235 , n49115 , n47427 );
nor ( n55236 , n55234 , n55235 );
xnor ( n55237 , n55236 , n47309 );
and ( n55238 , n50195 , n46911 );
and ( n55239 , n49976 , n46909 );
nor ( n55240 , n55238 , n55239 );
xnor ( n55241 , n55240 , n46802 );
and ( n55242 , n55237 , n55241 );
and ( n55243 , n50625 , n46712 );
and ( n55244 , n50404 , n46710 );
nor ( n55245 , n55243 , n55244 );
xnor ( n55246 , n55245 , n46587 );
and ( n55247 , n55241 , n55246 );
and ( n55248 , n55237 , n55246 );
or ( n55249 , n55242 , n55247 , n55248 );
and ( n55250 , n51077 , n46496 );
and ( n55251 , n50726 , n46494 );
nor ( n55252 , n55250 , n55251 );
xnor ( n55253 , n55252 , n46402 );
xor ( n55254 , n34206 , n45594 );
buf ( n55255 , n55254 );
buf ( n55256 , n55255 );
buf ( n55257 , n55256 );
and ( n55258 , n55253 , n55257 );
buf ( n55259 , n55258 );
and ( n55260 , n55249 , n55259 );
xor ( n55261 , n54865 , n54869 );
xor ( n55262 , n55261 , n54874 );
and ( n55263 , n55259 , n55262 );
and ( n55264 , n55249 , n55262 );
or ( n55265 , n55260 , n55263 , n55264 );
and ( n55266 , n55233 , n55265 );
xor ( n55267 , n54882 , n54886 );
xor ( n55268 , n55267 , n54891 );
xor ( n55269 , n54907 , n54911 );
xor ( n55270 , n55269 , n54916 );
and ( n55271 , n55268 , n55270 );
xor ( n55272 , n54923 , n54927 );
xor ( n55273 , n55272 , n54932 );
and ( n55274 , n55270 , n55273 );
and ( n55275 , n55268 , n55273 );
or ( n55276 , n55271 , n55274 , n55275 );
and ( n55277 , n55265 , n55276 );
and ( n55278 , n55233 , n55276 );
or ( n55279 , n55266 , n55277 , n55278 );
and ( n55280 , n55180 , n55279 );
and ( n55281 , n55083 , n55279 );
or ( n55282 , n55181 , n55280 , n55281 );
xor ( n55283 , n54776 , n54777 );
xor ( n55284 , n55283 , n54779 );
xor ( n55285 , n54787 , n54803 );
xor ( n55286 , n55285 , n54813 );
and ( n55287 , n55284 , n55286 );
xor ( n55288 , n54825 , n54834 );
xor ( n55289 , n55288 , n54844 );
and ( n55290 , n55286 , n55289 );
and ( n55291 , n55284 , n55289 );
or ( n55292 , n55287 , n55290 , n55291 );
xor ( n55293 , n54857 , n54877 );
xor ( n55294 , n55293 , n54894 );
xor ( n55295 , n54919 , n54935 );
xor ( n55296 , n55295 , n54951 );
and ( n55297 , n55294 , n55296 );
xor ( n55298 , n54956 , n54958 );
xor ( n55299 , n55298 , n54961 );
and ( n55300 , n55296 , n55299 );
and ( n55301 , n55294 , n55299 );
or ( n55302 , n55297 , n55300 , n55301 );
and ( n55303 , n55292 , n55302 );
xor ( n55304 , n54745 , n54746 );
xor ( n55305 , n55304 , n54748 );
and ( n55306 , n55302 , n55305 );
and ( n55307 , n55292 , n55305 );
or ( n55308 , n55303 , n55306 , n55307 );
and ( n55309 , n55282 , n55308 );
xor ( n55310 , n54754 , n54773 );
xor ( n55311 , n55310 , n54782 );
xor ( n55312 , n54816 , n54847 );
xor ( n55313 , n55312 , n54897 );
and ( n55314 , n55311 , n55313 );
xor ( n55315 , n54954 , n54964 );
xor ( n55316 , n55315 , n54967 );
and ( n55317 , n55313 , n55316 );
and ( n55318 , n55311 , n55316 );
or ( n55319 , n55314 , n55317 , n55318 );
and ( n55320 , n55308 , n55319 );
and ( n55321 , n55282 , n55319 );
or ( n55322 , n55309 , n55320 , n55321 );
and ( n55323 , n55064 , n55322 );
and ( n55324 , n55039 , n55322 );
or ( n55325 , n55065 , n55323 , n55324 );
xor ( n55326 , n54751 , n54785 );
xor ( n55327 , n55326 , n54900 );
xor ( n55328 , n54970 , n54980 );
xor ( n55329 , n55328 , n54983 );
and ( n55330 , n55327 , n55329 );
xor ( n55331 , n54989 , n54991 );
xor ( n55332 , n55331 , n54994 );
and ( n55333 , n55329 , n55332 );
and ( n55334 , n55327 , n55332 );
or ( n55335 , n55330 , n55333 , n55334 );
xor ( n55336 , n54903 , n54986 );
xor ( n55337 , n55336 , n54997 );
and ( n55338 , n55335 , n55337 );
xor ( n55339 , n55005 , n55007 );
xor ( n55340 , n55339 , n55010 );
and ( n55341 , n55337 , n55340 );
and ( n55342 , n55335 , n55340 );
or ( n55343 , n55338 , n55341 , n55342 );
and ( n55344 , n55325 , n55343 );
xor ( n55345 , n54740 , n54742 );
xor ( n55346 , n55345 , n55000 );
and ( n55347 , n55343 , n55346 );
and ( n55348 , n55325 , n55346 );
or ( n55349 , n55344 , n55347 , n55348 );
and ( n55350 , n55037 , n55349 );
xor ( n55351 , n55003 , n55021 );
xor ( n55352 , n55351 , n55024 );
and ( n55353 , n55349 , n55352 );
and ( n55354 , n55037 , n55352 );
or ( n55355 , n55350 , n55353 , n55354 );
and ( n55356 , n55035 , n55355 );
xor ( n55357 , n54735 , n54737 );
xor ( n55358 , n55357 , n55027 );
and ( n55359 , n55355 , n55358 );
and ( n55360 , n55035 , n55358 );
or ( n55361 , n55356 , n55359 , n55360 );
and ( n55362 , n55032 , n55361 );
and ( n55363 , n55030 , n55361 );
or ( n55364 , n55033 , n55362 , n55363 );
or ( n55365 , n54709 , n55364 );
or ( n55366 , n54707 , n55365 );
and ( n55367 , n54705 , n55366 );
xor ( n55368 , n54705 , n55366 );
xnor ( n55369 , n54707 , n55365 );
xnor ( n55370 , n54709 , n55364 );
xor ( n55371 , n55030 , n55032 );
xor ( n55372 , n55371 , n55361 );
xor ( n55373 , n55035 , n55355 );
xor ( n55374 , n55373 , n55358 );
xor ( n55375 , n55013 , n55015 );
xor ( n55376 , n55375 , n55018 );
xor ( n55377 , n54972 , n54974 );
xor ( n55378 , n55377 , n54977 );
xor ( n55379 , n54940 , n54943 );
xor ( n55380 , n55379 , n54948 );
and ( n55381 , n46345 , n51750 );
and ( n55382 , n46264 , n51748 );
nor ( n55383 , n55381 , n55382 );
xnor ( n55384 , n55383 , n51520 );
and ( n55385 , n46530 , n51221 );
and ( n55386 , n46445 , n51219 );
nor ( n55387 , n55385 , n55386 );
xnor ( n55388 , n55387 , n51000 );
and ( n55389 , n55384 , n55388 );
and ( n55390 , n46750 , n50783 );
and ( n55391 , n46577 , n50781 );
nor ( n55392 , n55390 , n55391 );
xnor ( n55393 , n55392 , n50557 );
and ( n55394 , n55388 , n55393 );
and ( n55395 , n55384 , n55393 );
or ( n55396 , n55389 , n55394 , n55395 );
and ( n55397 , n46843 , n50338 );
and ( n55398 , n46750 , n50336 );
nor ( n55399 , n55397 , n55398 );
xnor ( n55400 , n55399 , n50111 );
or ( n55401 , n55396 , n55400 );
and ( n55402 , n55380 , n55401 );
and ( n55403 , n51734 , n46306 );
and ( n55404 , n51510 , n46304 );
nor ( n55405 , n55403 , n55404 );
xnor ( n55406 , n55405 , n46228 );
and ( n55407 , n53328 , n45886 );
and ( n55408 , n53041 , n45884 );
nor ( n55409 , n55407 , n55408 );
xnor ( n55410 , n55409 , n45824 );
and ( n55411 , n55406 , n55410 );
and ( n55412 , n53922 , n45777 );
and ( n55413 , n53639 , n45775 );
nor ( n55414 , n55412 , n55413 );
xnor ( n55415 , n55414 , n45734 );
and ( n55416 , n55410 , n55415 );
and ( n55417 , n55406 , n55415 );
or ( n55418 , n55411 , n55416 , n55417 );
and ( n55419 , n52332 , n46135 );
and ( n55420 , n52082 , n46133 );
nor ( n55421 , n55419 , n55420 );
xnor ( n55422 , n55421 , n46067 );
and ( n55423 , n52790 , n45990 );
and ( n55424 , n52612 , n45988 );
nor ( n55425 , n55423 , n55424 );
xnor ( n55426 , n55425 , n45939 );
and ( n55427 , n55422 , n55426 );
and ( n55428 , n54604 , n45702 );
and ( n55429 , n54227 , n45700 );
nor ( n55430 , n55428 , n55429 );
xnor ( n55431 , n55430 , n20841 );
and ( n55432 , n55426 , n55431 );
and ( n55433 , n55422 , n55431 );
or ( n55434 , n55427 , n55432 , n55433 );
or ( n55435 , n55418 , n55434 );
and ( n55436 , n55401 , n55435 );
and ( n55437 , n55380 , n55435 );
or ( n55438 , n55402 , n55436 , n55437 );
and ( n55439 , n49976 , n47178 );
and ( n55440 , n49781 , n47176 );
nor ( n55441 , n55439 , n55440 );
xnor ( n55442 , n55441 , n47039 );
and ( n55443 , n50404 , n46911 );
and ( n55444 , n50195 , n46909 );
nor ( n55445 , n55443 , n55444 );
xnor ( n55446 , n55445 , n46802 );
and ( n55447 , n55442 , n55446 );
and ( n55448 , n50726 , n46712 );
and ( n55449 , n50625 , n46710 );
nor ( n55450 , n55448 , n55449 );
xnor ( n55451 , n55450 , n46587 );
and ( n55452 , n55446 , n55451 );
and ( n55453 , n55442 , n55451 );
or ( n55454 , n55447 , n55452 , n55453 );
and ( n55455 , n48709 , n48042 );
and ( n55456 , n48632 , n48040 );
nor ( n55457 , n55455 , n55456 );
xnor ( n55458 , n55457 , n47921 );
and ( n55459 , n49115 , n47734 );
and ( n55460 , n48988 , n47732 );
nor ( n55461 , n55459 , n55460 );
xnor ( n55462 , n55461 , n47606 );
and ( n55463 , n55458 , n55462 );
and ( n55464 , n49570 , n47429 );
and ( n55465 , n49374 , n47427 );
nor ( n55466 , n55464 , n55465 );
xnor ( n55467 , n55466 , n47309 );
and ( n55468 , n55462 , n55467 );
and ( n55469 , n55458 , n55467 );
or ( n55470 , n55463 , n55468 , n55469 );
and ( n55471 , n55454 , n55470 );
xor ( n55472 , n55090 , n55094 );
xor ( n55473 , n55472 , n55099 );
xnor ( n55474 , n55109 , n55113 );
and ( n55475 , n55473 , n55474 );
xnor ( n55476 , n55118 , n55122 );
and ( n55477 , n55474 , n55476 );
and ( n55478 , n55473 , n55476 );
or ( n55479 , n55475 , n55477 , n55478 );
and ( n55480 , n55471 , n55479 );
xnor ( n55481 , n55128 , n55132 );
xnor ( n55482 , n55141 , n55144 );
and ( n55483 , n55481 , n55482 );
xnor ( n55484 , n55149 , n55153 );
and ( n55485 , n55482 , n55484 );
and ( n55486 , n55481 , n55484 );
or ( n55487 , n55483 , n55485 , n55486 );
and ( n55488 , n55479 , n55487 );
and ( n55489 , n55471 , n55487 );
or ( n55490 , n55480 , n55488 , n55489 );
and ( n55491 , n55438 , n55490 );
and ( n55492 , n55143 , n20852 );
and ( n55493 , n54942 , n20850 );
nor ( n55494 , n55492 , n55493 );
xnor ( n55495 , n55494 , n20860 );
buf ( n55496 , n20806 );
buf ( n55497 , n55496 );
and ( n55498 , n55497 , n20846 );
or ( n55499 , n55495 , n55498 );
buf ( n55500 , n17563 );
buf ( n55501 , n55500 );
buf ( n55502 , n17565 );
buf ( n55503 , n55502 );
and ( n55504 , n55501 , n55503 );
not ( n55505 , n55504 );
and ( n55506 , n54861 , n55505 );
not ( n55507 , n55506 );
and ( n55508 , n20844 , n55159 );
and ( n55509 , n20855 , n55157 );
nor ( n55510 , n55508 , n55509 );
xnor ( n55511 , n55510 , n54864 );
and ( n55512 , n55507 , n55511 );
and ( n55513 , n45712 , n54535 );
and ( n55514 , n20864 , n54533 );
nor ( n55515 , n55513 , n55514 );
xnor ( n55516 , n55515 , n54237 );
and ( n55517 , n55511 , n55516 );
and ( n55518 , n55507 , n55516 );
or ( n55519 , n55512 , n55517 , n55518 );
and ( n55520 , n55499 , n55519 );
and ( n55521 , n45794 , n53928 );
and ( n55522 , n45763 , n53926 );
nor ( n55523 , n55521 , n55522 );
xnor ( n55524 , n55523 , n53652 );
and ( n55525 , n45907 , n53357 );
and ( n55526 , n45843 , n53355 );
nor ( n55527 , n55525 , n55526 );
xnor ( n55528 , n55527 , n53060 );
and ( n55529 , n55524 , n55528 );
and ( n55530 , n46041 , n52799 );
and ( n55531 , n45963 , n52797 );
nor ( n55532 , n55530 , n55531 );
xnor ( n55533 , n55532 , n52538 );
and ( n55534 , n55528 , n55533 );
and ( n55535 , n55524 , n55533 );
or ( n55536 , n55529 , n55534 , n55535 );
and ( n55537 , n55519 , n55536 );
and ( n55538 , n55499 , n55536 );
or ( n55539 , n55520 , n55537 , n55538 );
and ( n55540 , n46169 , n52269 );
and ( n55541 , n46100 , n52267 );
nor ( n55542 , n55540 , n55541 );
xnor ( n55543 , n55542 , n52008 );
and ( n55544 , n46969 , n50338 );
and ( n55545 , n46843 , n50336 );
nor ( n55546 , n55544 , n55545 );
xnor ( n55547 , n55546 , n50111 );
and ( n55548 , n55543 , n55547 );
and ( n55549 , n47216 , n49896 );
and ( n55550 , n47090 , n49894 );
nor ( n55551 , n55549 , n55550 );
xnor ( n55552 , n55551 , n49711 );
and ( n55553 , n55547 , n55552 );
and ( n55554 , n55543 , n55552 );
or ( n55555 , n55548 , n55553 , n55554 );
and ( n55556 , n47778 , n49121 );
and ( n55557 , n47647 , n49119 );
nor ( n55558 , n55556 , n55557 );
xnor ( n55559 , n55558 , n48932 );
and ( n55560 , n48108 , n48740 );
and ( n55561 , n47962 , n48738 );
nor ( n55562 , n55560 , n55561 );
xnor ( n55563 , n55562 , n48571 );
and ( n55564 , n55559 , n55563 );
and ( n55565 , n48384 , n48394 );
and ( n55566 , n48272 , n48392 );
nor ( n55567 , n55565 , n55566 );
xnor ( n55568 , n55567 , n48220 );
and ( n55569 , n55563 , n55568 );
and ( n55570 , n55559 , n55568 );
or ( n55571 , n55564 , n55569 , n55570 );
and ( n55572 , n55555 , n55571 );
and ( n55573 , n51298 , n46496 );
and ( n55574 , n51077 , n46494 );
nor ( n55575 , n55573 , n55574 );
xnor ( n55576 , n55575 , n46402 );
xor ( n55577 , n35242 , n45592 );
buf ( n55578 , n55577 );
buf ( n55579 , n55578 );
buf ( n55580 , n55579 );
and ( n55581 , n55576 , n55580 );
buf ( n55582 , n55581 );
and ( n55583 , n55571 , n55582 );
and ( n55584 , n55555 , n55582 );
or ( n55585 , n55572 , n55583 , n55584 );
and ( n55586 , n55539 , n55585 );
xor ( n55587 , n55162 , n55166 );
xor ( n55588 , n55587 , n55171 );
xor ( n55589 , n55185 , n55189 );
xor ( n55590 , n55589 , n55194 );
and ( n55591 , n55588 , n55590 );
xor ( n55592 , n55201 , n55205 );
xor ( n55593 , n55592 , n55210 );
and ( n55594 , n55590 , n55593 );
and ( n55595 , n55588 , n55593 );
or ( n55596 , n55591 , n55594 , n55595 );
and ( n55597 , n55585 , n55596 );
and ( n55598 , n55539 , n55596 );
or ( n55599 , n55586 , n55597 , n55598 );
and ( n55600 , n55490 , n55599 );
and ( n55601 , n55438 , n55599 );
or ( n55602 , n55491 , n55600 , n55601 );
and ( n55603 , n55378 , n55602 );
xor ( n55604 , n55218 , n55222 );
xor ( n55605 , n55604 , n55227 );
xor ( n55606 , n55237 , n55241 );
xor ( n55607 , n55606 , n55246 );
and ( n55608 , n55605 , n55607 );
xor ( n55609 , n55253 , n55257 );
buf ( n55610 , n55609 );
and ( n55611 , n55607 , n55610 );
and ( n55612 , n55605 , n55610 );
or ( n55613 , n55608 , n55611 , n55612 );
buf ( n55614 , n55068 );
xor ( n55615 , n55614 , n55070 );
and ( n55616 , n55613 , n55615 );
xor ( n55617 , n55074 , n55075 );
xor ( n55618 , n55617 , n55077 );
and ( n55619 , n55615 , n55618 );
and ( n55620 , n55613 , n55618 );
or ( n55621 , n55616 , n55619 , n55620 );
xor ( n55622 , n55084 , n55085 );
xor ( n55623 , n55622 , n55102 );
xor ( n55624 , n55114 , n55123 );
xor ( n55625 , n55624 , n55133 );
and ( n55626 , n55623 , n55625 );
xor ( n55627 , n55145 , n55154 );
xor ( n55628 , n55627 , n55174 );
and ( n55629 , n55625 , n55628 );
and ( n55630 , n55623 , n55628 );
or ( n55631 , n55626 , n55629 , n55630 );
and ( n55632 , n55621 , n55631 );
xor ( n55633 , n55197 , n55213 );
xor ( n55634 , n55633 , n55230 );
xor ( n55635 , n55249 , n55259 );
xor ( n55636 , n55635 , n55262 );
and ( n55637 , n55634 , n55636 );
xor ( n55638 , n55268 , n55270 );
xor ( n55639 , n55638 , n55273 );
and ( n55640 , n55636 , n55639 );
and ( n55641 , n55634 , n55639 );
or ( n55642 , n55637 , n55640 , n55641 );
and ( n55643 , n55631 , n55642 );
and ( n55644 , n55621 , n55642 );
or ( n55645 , n55632 , n55643 , n55644 );
and ( n55646 , n55602 , n55645 );
and ( n55647 , n55378 , n55645 );
or ( n55648 , n55603 , n55646 , n55647 );
xor ( n55649 , n55051 , n55053 );
xor ( n55650 , n55649 , n55055 );
xor ( n55651 , n55066 , n55072 );
xor ( n55652 , n55651 , n55080 );
and ( n55653 , n55650 , n55652 );
xor ( n55654 , n55105 , n55136 );
xor ( n55655 , n55654 , n55177 );
and ( n55656 , n55652 , n55655 );
and ( n55657 , n55650 , n55655 );
or ( n55658 , n55653 , n55656 , n55657 );
xor ( n55659 , n55233 , n55265 );
xor ( n55660 , n55659 , n55276 );
xor ( n55661 , n55284 , n55286 );
xor ( n55662 , n55661 , n55289 );
and ( n55663 , n55660 , n55662 );
xor ( n55664 , n55294 , n55296 );
xor ( n55665 , n55664 , n55299 );
and ( n55666 , n55662 , n55665 );
and ( n55667 , n55660 , n55665 );
or ( n55668 , n55663 , n55666 , n55667 );
and ( n55669 , n55658 , n55668 );
xor ( n55670 , n55046 , n55048 );
xor ( n55671 , n55670 , n55058 );
and ( n55672 , n55668 , n55671 );
and ( n55673 , n55658 , n55671 );
or ( n55674 , n55669 , n55672 , n55673 );
and ( n55675 , n55648 , n55674 );
xor ( n55676 , n55083 , n55180 );
xor ( n55677 , n55676 , n55279 );
xor ( n55678 , n55292 , n55302 );
xor ( n55679 , n55678 , n55305 );
and ( n55680 , n55677 , n55679 );
xor ( n55681 , n55311 , n55313 );
xor ( n55682 , n55681 , n55316 );
and ( n55683 , n55679 , n55682 );
and ( n55684 , n55677 , n55682 );
or ( n55685 , n55680 , n55683 , n55684 );
and ( n55686 , n55674 , n55685 );
and ( n55687 , n55648 , n55685 );
or ( n55688 , n55675 , n55686 , n55687 );
xor ( n55689 , n55041 , n55043 );
xor ( n55690 , n55689 , n55061 );
xor ( n55691 , n55282 , n55308 );
xor ( n55692 , n55691 , n55319 );
and ( n55693 , n55690 , n55692 );
xor ( n55694 , n55327 , n55329 );
xor ( n55695 , n55694 , n55332 );
and ( n55696 , n55692 , n55695 );
and ( n55697 , n55690 , n55695 );
or ( n55698 , n55693 , n55696 , n55697 );
and ( n55699 , n55688 , n55698 );
xor ( n55700 , n55039 , n55064 );
xor ( n55701 , n55700 , n55322 );
and ( n55702 , n55698 , n55701 );
and ( n55703 , n55688 , n55701 );
or ( n55704 , n55699 , n55702 , n55703 );
and ( n55705 , n55376 , n55704 );
xor ( n55706 , n55325 , n55343 );
xor ( n55707 , n55706 , n55346 );
and ( n55708 , n55704 , n55707 );
and ( n55709 , n55376 , n55707 );
or ( n55710 , n55705 , n55708 , n55709 );
xor ( n55711 , n55037 , n55349 );
xor ( n55712 , n55711 , n55352 );
and ( n55713 , n55710 , n55712 );
xor ( n55714 , n55335 , n55337 );
xor ( n55715 , n55714 , n55340 );
xnor ( n55716 , n55396 , n55400 );
xnor ( n55717 , n55418 , n55434 );
and ( n55718 , n55716 , n55717 );
xor ( n55719 , n55454 , n55470 );
and ( n55720 , n55717 , n55719 );
and ( n55721 , n55716 , n55719 );
or ( n55722 , n55718 , n55720 , n55721 );
and ( n55723 , n47474 , n49513 );
and ( n55724 , n47351 , n49511 );
nor ( n55725 , n55723 , n55724 );
xnor ( n55726 , n55725 , n49310 );
xor ( n55727 , n55384 , n55388 );
xor ( n55728 , n55727 , n55393 );
or ( n55729 , n55726 , n55728 );
and ( n55730 , n53041 , n45990 );
and ( n55731 , n52790 , n45988 );
nor ( n55732 , n55730 , n55731 );
xnor ( n55733 , n55732 , n45939 );
and ( n55734 , n54942 , n45702 );
and ( n55735 , n54604 , n45700 );
nor ( n55736 , n55734 , n55735 );
xnor ( n55737 , n55736 , n20841 );
and ( n55738 , n55733 , n55737 );
and ( n55739 , n55497 , n20852 );
and ( n55740 , n55143 , n20850 );
nor ( n55741 , n55739 , n55740 );
xnor ( n55742 , n55741 , n20860 );
and ( n55743 , n55737 , n55742 );
and ( n55744 , n55733 , n55742 );
or ( n55745 , n55738 , n55743 , n55744 );
and ( n55746 , n52612 , n46135 );
and ( n55747 , n52332 , n46133 );
nor ( n55748 , n55746 , n55747 );
xnor ( n55749 , n55748 , n46067 );
and ( n55750 , n54227 , n45777 );
and ( n55751 , n53922 , n45775 );
nor ( n55752 , n55750 , n55751 );
xnor ( n55753 , n55752 , n45734 );
and ( n55754 , n55749 , n55753 );
buf ( n55755 , n20808 );
buf ( n55756 , n55755 );
and ( n55757 , n55756 , n20846 );
and ( n55758 , n55753 , n55757 );
and ( n55759 , n55749 , n55757 );
or ( n55760 , n55754 , n55758 , n55759 );
or ( n55761 , n55745 , n55760 );
and ( n55762 , n55729 , n55761 );
xor ( n55763 , n55406 , n55410 );
xor ( n55764 , n55763 , n55415 );
xor ( n55765 , n55442 , n55446 );
xor ( n55766 , n55765 , n55451 );
and ( n55767 , n55764 , n55766 );
xor ( n55768 , n55458 , n55462 );
xor ( n55769 , n55768 , n55467 );
and ( n55770 , n55766 , n55769 );
and ( n55771 , n55764 , n55769 );
or ( n55772 , n55767 , n55770 , n55771 );
and ( n55773 , n55761 , n55772 );
and ( n55774 , n55729 , n55772 );
or ( n55775 , n55762 , n55773 , n55774 );
and ( n55776 , n55722 , n55775 );
xor ( n55777 , n55422 , n55426 );
xor ( n55778 , n55777 , n55431 );
xnor ( n55779 , n55495 , n55498 );
and ( n55780 , n55778 , n55779 );
and ( n55781 , n46264 , n52269 );
and ( n55782 , n46169 , n52267 );
nor ( n55783 , n55781 , n55782 );
xnor ( n55784 , n55783 , n52008 );
and ( n55785 , n46445 , n51750 );
and ( n55786 , n46345 , n51748 );
nor ( n55787 , n55785 , n55786 );
xnor ( n55788 , n55787 , n51520 );
and ( n55789 , n55784 , n55788 );
and ( n55790 , n46577 , n51221 );
and ( n55791 , n46530 , n51219 );
nor ( n55792 , n55790 , n55791 );
xnor ( n55793 , n55792 , n51000 );
and ( n55794 , n55788 , n55793 );
and ( n55795 , n55784 , n55793 );
or ( n55796 , n55789 , n55794 , n55795 );
and ( n55797 , n55779 , n55796 );
and ( n55798 , n55778 , n55796 );
or ( n55799 , n55780 , n55797 , n55798 );
and ( n55800 , n48988 , n48042 );
and ( n55801 , n48709 , n48040 );
nor ( n55802 , n55800 , n55801 );
xnor ( n55803 , n55802 , n47921 );
and ( n55804 , n49781 , n47429 );
and ( n55805 , n49570 , n47427 );
nor ( n55806 , n55804 , n55805 );
xnor ( n55807 , n55806 , n47309 );
and ( n55808 , n55803 , n55807 );
and ( n55809 , n50195 , n47178 );
and ( n55810 , n49976 , n47176 );
nor ( n55811 , n55809 , n55810 );
xnor ( n55812 , n55811 , n47039 );
and ( n55813 , n55807 , n55812 );
and ( n55814 , n55803 , n55812 );
or ( n55815 , n55808 , n55813 , n55814 );
and ( n55816 , n47090 , n50338 );
and ( n55817 , n46969 , n50336 );
nor ( n55818 , n55816 , n55817 );
xnor ( n55819 , n55818 , n50111 );
and ( n55820 , n47351 , n49896 );
and ( n55821 , n47216 , n49894 );
nor ( n55822 , n55820 , n55821 );
xnor ( n55823 , n55822 , n49711 );
or ( n55824 , n55819 , n55823 );
and ( n55825 , n55815 , n55824 );
and ( n55826 , n52082 , n46306 );
and ( n55827 , n51734 , n46304 );
nor ( n55828 , n55826 , n55827 );
xnor ( n55829 , n55828 , n46228 );
and ( n55830 , n53639 , n45886 );
and ( n55831 , n53328 , n45884 );
nor ( n55832 , n55830 , n55831 );
xnor ( n55833 , n55832 , n45824 );
or ( n55834 , n55829 , n55833 );
and ( n55835 , n55824 , n55834 );
and ( n55836 , n55815 , n55834 );
or ( n55837 , n55825 , n55835 , n55836 );
and ( n55838 , n55799 , n55837 );
and ( n55839 , n50625 , n46911 );
and ( n55840 , n50404 , n46909 );
nor ( n55841 , n55839 , n55840 );
xnor ( n55842 , n55841 , n46802 );
and ( n55843 , n51077 , n46712 );
and ( n55844 , n50726 , n46710 );
nor ( n55845 , n55843 , n55844 );
xnor ( n55846 , n55845 , n46587 );
and ( n55847 , n55842 , n55846 );
xor ( n55848 , n54861 , n55501 );
xor ( n55849 , n55501 , n55503 );
not ( n55850 , n55849 );
and ( n55851 , n55848 , n55850 );
and ( n55852 , n20855 , n55851 );
not ( n55853 , n55852 );
xnor ( n55854 , n55853 , n55506 );
and ( n55855 , n20864 , n55159 );
and ( n55856 , n20844 , n55157 );
nor ( n55857 , n55855 , n55856 );
xnor ( n55858 , n55857 , n54864 );
and ( n55859 , n55854 , n55858 );
and ( n55860 , n45763 , n54535 );
and ( n55861 , n45712 , n54533 );
nor ( n55862 , n55860 , n55861 );
xnor ( n55863 , n55862 , n54237 );
and ( n55864 , n55858 , n55863 );
and ( n55865 , n55854 , n55863 );
or ( n55866 , n55859 , n55864 , n55865 );
and ( n55867 , n55847 , n55866 );
and ( n55868 , n45843 , n53928 );
and ( n55869 , n45794 , n53926 );
nor ( n55870 , n55868 , n55869 );
xnor ( n55871 , n55870 , n53652 );
and ( n55872 , n45963 , n53357 );
and ( n55873 , n45907 , n53355 );
nor ( n55874 , n55872 , n55873 );
xnor ( n55875 , n55874 , n53060 );
and ( n55876 , n55871 , n55875 );
and ( n55877 , n46100 , n52799 );
and ( n55878 , n46041 , n52797 );
nor ( n55879 , n55877 , n55878 );
xnor ( n55880 , n55879 , n52538 );
and ( n55881 , n55875 , n55880 );
and ( n55882 , n55871 , n55880 );
or ( n55883 , n55876 , n55881 , n55882 );
and ( n55884 , n55866 , n55883 );
and ( n55885 , n55847 , n55883 );
or ( n55886 , n55867 , n55884 , n55885 );
and ( n55887 , n55837 , n55886 );
and ( n55888 , n55799 , n55886 );
or ( n55889 , n55838 , n55887 , n55888 );
and ( n55890 , n55775 , n55889 );
and ( n55891 , n55722 , n55889 );
or ( n55892 , n55776 , n55890 , n55891 );
and ( n55893 , n46843 , n50783 );
and ( n55894 , n46750 , n50781 );
nor ( n55895 , n55893 , n55894 );
xnor ( n55896 , n55895 , n50557 );
and ( n55897 , n47647 , n49513 );
and ( n55898 , n47474 , n49511 );
nor ( n55899 , n55897 , n55898 );
xnor ( n55900 , n55899 , n49310 );
and ( n55901 , n55896 , n55900 );
and ( n55902 , n47962 , n49121 );
and ( n55903 , n47778 , n49119 );
nor ( n55904 , n55902 , n55903 );
xnor ( n55905 , n55904 , n48932 );
and ( n55906 , n55900 , n55905 );
and ( n55907 , n55896 , n55905 );
or ( n55908 , n55901 , n55906 , n55907 );
and ( n55909 , n48272 , n48740 );
and ( n55910 , n48108 , n48738 );
nor ( n55911 , n55909 , n55910 );
xnor ( n55912 , n55911 , n48571 );
and ( n55913 , n48632 , n48394 );
and ( n55914 , n48384 , n48392 );
nor ( n55915 , n55913 , n55914 );
xnor ( n55916 , n55915 , n48220 );
and ( n55917 , n55912 , n55916 );
and ( n55918 , n49374 , n47734 );
and ( n55919 , n49115 , n47732 );
nor ( n55920 , n55918 , n55919 );
xnor ( n55921 , n55920 , n47606 );
and ( n55922 , n55916 , n55921 );
and ( n55923 , n55912 , n55921 );
or ( n55924 , n55917 , n55922 , n55923 );
and ( n55925 , n55908 , n55924 );
and ( n55926 , n51510 , n46496 );
and ( n55927 , n51298 , n46494 );
nor ( n55928 , n55926 , n55927 );
xnor ( n55929 , n55928 , n46402 );
xor ( n55930 , n35244 , n45591 );
buf ( n55931 , n55930 );
buf ( n55932 , n55931 );
buf ( n55933 , n55932 );
and ( n55934 , n55929 , n55933 );
buf ( n55935 , n55934 );
and ( n55936 , n55924 , n55935 );
and ( n55937 , n55908 , n55935 );
or ( n55938 , n55925 , n55936 , n55937 );
xor ( n55939 , n55507 , n55511 );
xor ( n55940 , n55939 , n55516 );
xor ( n55941 , n55524 , n55528 );
xor ( n55942 , n55941 , n55533 );
and ( n55943 , n55940 , n55942 );
xor ( n55944 , n55543 , n55547 );
xor ( n55945 , n55944 , n55552 );
and ( n55946 , n55942 , n55945 );
and ( n55947 , n55940 , n55945 );
or ( n55948 , n55943 , n55946 , n55947 );
and ( n55949 , n55938 , n55948 );
xor ( n55950 , n55473 , n55474 );
xor ( n55951 , n55950 , n55476 );
and ( n55952 , n55948 , n55951 );
and ( n55953 , n55938 , n55951 );
or ( n55954 , n55949 , n55952 , n55953 );
xor ( n55955 , n55481 , n55482 );
xor ( n55956 , n55955 , n55484 );
xor ( n55957 , n55499 , n55519 );
xor ( n55958 , n55957 , n55536 );
and ( n55959 , n55956 , n55958 );
xor ( n55960 , n55555 , n55571 );
xor ( n55961 , n55960 , n55582 );
and ( n55962 , n55958 , n55961 );
and ( n55963 , n55956 , n55961 );
or ( n55964 , n55959 , n55962 , n55963 );
and ( n55965 , n55954 , n55964 );
xor ( n55966 , n55380 , n55401 );
xor ( n55967 , n55966 , n55435 );
and ( n55968 , n55964 , n55967 );
and ( n55969 , n55954 , n55967 );
or ( n55970 , n55965 , n55968 , n55969 );
and ( n55971 , n55892 , n55970 );
xor ( n55972 , n55471 , n55479 );
xor ( n55973 , n55972 , n55487 );
xor ( n55974 , n55539 , n55585 );
xor ( n55975 , n55974 , n55596 );
and ( n55976 , n55973 , n55975 );
xor ( n55977 , n55613 , n55615 );
xor ( n55978 , n55977 , n55618 );
and ( n55979 , n55975 , n55978 );
and ( n55980 , n55973 , n55978 );
or ( n55981 , n55976 , n55979 , n55980 );
and ( n55982 , n55970 , n55981 );
and ( n55983 , n55892 , n55981 );
or ( n55984 , n55971 , n55982 , n55983 );
xor ( n55985 , n55438 , n55490 );
xor ( n55986 , n55985 , n55599 );
xor ( n55987 , n55621 , n55631 );
xor ( n55988 , n55987 , n55642 );
and ( n55989 , n55986 , n55988 );
xor ( n55990 , n55650 , n55652 );
xor ( n55991 , n55990 , n55655 );
and ( n55992 , n55988 , n55991 );
and ( n55993 , n55986 , n55991 );
or ( n55994 , n55989 , n55992 , n55993 );
and ( n55995 , n55984 , n55994 );
xor ( n55996 , n55378 , n55602 );
xor ( n55997 , n55996 , n55645 );
and ( n55998 , n55994 , n55997 );
and ( n55999 , n55984 , n55997 );
or ( n56000 , n55995 , n55998 , n55999 );
xor ( n56001 , n55648 , n55674 );
xor ( n56002 , n56001 , n55685 );
and ( n56003 , n56000 , n56002 );
xor ( n56004 , n55690 , n55692 );
xor ( n56005 , n56004 , n55695 );
and ( n56006 , n56002 , n56005 );
and ( n56007 , n56000 , n56005 );
or ( n56008 , n56003 , n56006 , n56007 );
and ( n56009 , n55715 , n56008 );
xor ( n56010 , n55688 , n55698 );
xor ( n56011 , n56010 , n55701 );
and ( n56012 , n56008 , n56011 );
and ( n56013 , n55715 , n56011 );
or ( n56014 , n56009 , n56012 , n56013 );
xor ( n56015 , n55376 , n55704 );
xor ( n56016 , n56015 , n55707 );
and ( n56017 , n56014 , n56016 );
xor ( n56018 , n55715 , n56008 );
xor ( n56019 , n56018 , n56011 );
xor ( n56020 , n55658 , n55668 );
xor ( n56021 , n56020 , n55671 );
xor ( n56022 , n55677 , n55679 );
xor ( n56023 , n56022 , n55682 );
and ( n56024 , n56021 , n56023 );
xor ( n56025 , n55660 , n55662 );
xor ( n56026 , n56025 , n55665 );
xor ( n56027 , n55623 , n55625 );
xor ( n56028 , n56027 , n55628 );
xor ( n56029 , n55634 , n55636 );
xor ( n56030 , n56029 , n55639 );
and ( n56031 , n56028 , n56030 );
xor ( n56032 , n55588 , n55590 );
xor ( n56033 , n56032 , n55593 );
xor ( n56034 , n55605 , n55607 );
xor ( n56035 , n56034 , n55610 );
and ( n56036 , n56033 , n56035 );
xor ( n56037 , n55559 , n55563 );
xor ( n56038 , n56037 , n55568 );
xor ( n56039 , n55576 , n55580 );
buf ( n56040 , n56039 );
and ( n56041 , n56038 , n56040 );
xnor ( n56042 , n55726 , n55728 );
and ( n56043 , n56040 , n56042 );
and ( n56044 , n56038 , n56042 );
or ( n56045 , n56041 , n56043 , n56044 );
and ( n56046 , n56035 , n56045 );
and ( n56047 , n56033 , n56045 );
or ( n56048 , n56036 , n56046 , n56047 );
and ( n56049 , n56030 , n56048 );
and ( n56050 , n56028 , n56048 );
or ( n56051 , n56031 , n56049 , n56050 );
and ( n56052 , n56026 , n56051 );
xnor ( n56053 , n55745 , n55760 );
and ( n56054 , n50404 , n47178 );
and ( n56055 , n50195 , n47176 );
nor ( n56056 , n56054 , n56055 );
xnor ( n56057 , n56056 , n47039 );
and ( n56058 , n50726 , n46911 );
and ( n56059 , n50625 , n46909 );
nor ( n56060 , n56058 , n56059 );
xnor ( n56061 , n56060 , n46802 );
and ( n56062 , n56057 , n56061 );
and ( n56063 , n51298 , n46712 );
and ( n56064 , n51077 , n46710 );
nor ( n56065 , n56063 , n56064 );
xnor ( n56066 , n56065 , n46587 );
and ( n56067 , n56061 , n56066 );
and ( n56068 , n56057 , n56066 );
or ( n56069 , n56062 , n56067 , n56068 );
and ( n56070 , n48709 , n48394 );
and ( n56071 , n48632 , n48392 );
nor ( n56072 , n56070 , n56071 );
xnor ( n56073 , n56072 , n48220 );
and ( n56074 , n49115 , n48042 );
and ( n56075 , n48988 , n48040 );
nor ( n56076 , n56074 , n56075 );
xnor ( n56077 , n56076 , n47921 );
and ( n56078 , n56073 , n56077 );
and ( n56079 , n49976 , n47429 );
and ( n56080 , n49781 , n47427 );
nor ( n56081 , n56079 , n56080 );
xnor ( n56082 , n56081 , n47309 );
and ( n56083 , n56077 , n56082 );
and ( n56084 , n56073 , n56082 );
or ( n56085 , n56078 , n56083 , n56084 );
or ( n56086 , n56069 , n56085 );
and ( n56087 , n56053 , n56086 );
xor ( n56088 , n55733 , n55737 );
xor ( n56089 , n56088 , n55742 );
xor ( n56090 , n55749 , n55753 );
xor ( n56091 , n56090 , n55757 );
or ( n56092 , n56089 , n56091 );
and ( n56093 , n56086 , n56092 );
and ( n56094 , n56053 , n56092 );
or ( n56095 , n56087 , n56093 , n56094 );
xor ( n56096 , n55784 , n55788 );
xor ( n56097 , n56096 , n55793 );
xor ( n56098 , n55803 , n55807 );
xor ( n56099 , n56098 , n55812 );
and ( n56100 , n56097 , n56099 );
xnor ( n56101 , n55819 , n55823 );
and ( n56102 , n56099 , n56101 );
and ( n56103 , n56097 , n56101 );
or ( n56104 , n56100 , n56102 , n56103 );
xnor ( n56105 , n55829 , n55833 );
xor ( n56106 , n55842 , n55846 );
and ( n56107 , n56105 , n56106 );
and ( n56108 , n52790 , n46135 );
and ( n56109 , n52612 , n46133 );
nor ( n56110 , n56108 , n56109 );
xnor ( n56111 , n56110 , n46067 );
and ( n56112 , n53328 , n45990 );
and ( n56113 , n53041 , n45988 );
nor ( n56114 , n56112 , n56113 );
xnor ( n56115 , n56114 , n45939 );
and ( n56116 , n56111 , n56115 );
and ( n56117 , n53922 , n45886 );
and ( n56118 , n53639 , n45884 );
nor ( n56119 , n56117 , n56118 );
xnor ( n56120 , n56119 , n45824 );
and ( n56121 , n56115 , n56120 );
and ( n56122 , n56111 , n56120 );
or ( n56123 , n56116 , n56121 , n56122 );
and ( n56124 , n56106 , n56123 );
and ( n56125 , n56105 , n56123 );
or ( n56126 , n56107 , n56124 , n56125 );
and ( n56127 , n56104 , n56126 );
and ( n56128 , n47216 , n50338 );
and ( n56129 , n47090 , n50336 );
nor ( n56130 , n56128 , n56129 );
xnor ( n56131 , n56130 , n50111 );
and ( n56132 , n47474 , n49896 );
and ( n56133 , n47351 , n49894 );
nor ( n56134 , n56132 , n56133 );
xnor ( n56135 , n56134 , n49711 );
or ( n56136 , n56131 , n56135 );
and ( n56137 , n46345 , n52269 );
and ( n56138 , n46264 , n52267 );
nor ( n56139 , n56137 , n56138 );
xnor ( n56140 , n56139 , n52008 );
and ( n56141 , n46530 , n51750 );
and ( n56142 , n46445 , n51748 );
nor ( n56143 , n56141 , n56142 );
xnor ( n56144 , n56143 , n51520 );
or ( n56145 , n56140 , n56144 );
and ( n56146 , n56136 , n56145 );
and ( n56147 , n48384 , n48740 );
and ( n56148 , n48272 , n48738 );
nor ( n56149 , n56147 , n56148 );
xnor ( n56150 , n56149 , n48571 );
and ( n56151 , n49570 , n47734 );
and ( n56152 , n49374 , n47732 );
nor ( n56153 , n56151 , n56152 );
xnor ( n56154 , n56153 , n47606 );
or ( n56155 , n56150 , n56154 );
and ( n56156 , n56145 , n56155 );
and ( n56157 , n56136 , n56155 );
or ( n56158 , n56146 , n56156 , n56157 );
and ( n56159 , n56126 , n56158 );
and ( n56160 , n56104 , n56158 );
or ( n56161 , n56127 , n56159 , n56160 );
and ( n56162 , n56095 , n56161 );
and ( n56163 , n52332 , n46306 );
and ( n56164 , n52082 , n46304 );
nor ( n56165 , n56163 , n56164 );
xnor ( n56166 , n56165 , n46228 );
and ( n56167 , n54604 , n45777 );
and ( n56168 , n54227 , n45775 );
nor ( n56169 , n56167 , n56168 );
xnor ( n56170 , n56169 , n45734 );
or ( n56171 , n56166 , n56170 );
buf ( n56172 , n17567 );
buf ( n56173 , n56172 );
buf ( n56174 , n17570 );
buf ( n56175 , n56174 );
and ( n56176 , n56173 , n56175 );
not ( n56177 , n56176 );
and ( n56178 , n55503 , n56177 );
not ( n56179 , n56178 );
and ( n56180 , n20844 , n55851 );
and ( n56181 , n20855 , n55849 );
nor ( n56182 , n56180 , n56181 );
xnor ( n56183 , n56182 , n55506 );
and ( n56184 , n56179 , n56183 );
and ( n56185 , n45712 , n55159 );
and ( n56186 , n20864 , n55157 );
nor ( n56187 , n56185 , n56186 );
xnor ( n56188 , n56187 , n54864 );
and ( n56189 , n56183 , n56188 );
and ( n56190 , n56179 , n56188 );
or ( n56191 , n56184 , n56189 , n56190 );
and ( n56192 , n56171 , n56191 );
and ( n56193 , n45794 , n54535 );
and ( n56194 , n45763 , n54533 );
nor ( n56195 , n56193 , n56194 );
xnor ( n56196 , n56195 , n54237 );
and ( n56197 , n45907 , n53928 );
and ( n56198 , n45843 , n53926 );
nor ( n56199 , n56197 , n56198 );
xnor ( n56200 , n56199 , n53652 );
and ( n56201 , n56196 , n56200 );
and ( n56202 , n46041 , n53357 );
and ( n56203 , n45963 , n53355 );
nor ( n56204 , n56202 , n56203 );
xnor ( n56205 , n56204 , n53060 );
and ( n56206 , n56200 , n56205 );
and ( n56207 , n56196 , n56205 );
or ( n56208 , n56201 , n56206 , n56207 );
and ( n56209 , n56191 , n56208 );
and ( n56210 , n56171 , n56208 );
or ( n56211 , n56192 , n56209 , n56210 );
and ( n56212 , n46169 , n52799 );
and ( n56213 , n46100 , n52797 );
nor ( n56214 , n56212 , n56213 );
xnor ( n56215 , n56214 , n52538 );
and ( n56216 , n46750 , n51221 );
and ( n56217 , n46577 , n51219 );
nor ( n56218 , n56216 , n56217 );
xnor ( n56219 , n56218 , n51000 );
and ( n56220 , n56215 , n56219 );
and ( n56221 , n46969 , n50783 );
and ( n56222 , n46843 , n50781 );
nor ( n56223 , n56221 , n56222 );
xnor ( n56224 , n56223 , n50557 );
and ( n56225 , n56219 , n56224 );
and ( n56226 , n56215 , n56224 );
or ( n56227 , n56220 , n56225 , n56226 );
and ( n56228 , n47778 , n49513 );
and ( n56229 , n47647 , n49511 );
nor ( n56230 , n56228 , n56229 );
xnor ( n56231 , n56230 , n49310 );
and ( n56232 , n48108 , n49121 );
and ( n56233 , n47962 , n49119 );
nor ( n56234 , n56232 , n56233 );
xnor ( n56235 , n56234 , n48932 );
and ( n56236 , n56231 , n56235 );
and ( n56237 , n51734 , n46496 );
and ( n56238 , n51510 , n46494 );
nor ( n56239 , n56237 , n56238 );
xnor ( n56240 , n56239 , n46402 );
and ( n56241 , n56235 , n56240 );
and ( n56242 , n56231 , n56240 );
or ( n56243 , n56236 , n56241 , n56242 );
and ( n56244 , n56227 , n56243 );
and ( n56245 , n55143 , n45702 );
and ( n56246 , n54942 , n45700 );
nor ( n56247 , n56245 , n56246 );
xnor ( n56248 , n56247 , n20841 );
and ( n56249 , n55756 , n20852 );
and ( n56250 , n55497 , n20850 );
nor ( n56251 , n56249 , n56250 );
xnor ( n56252 , n56251 , n20860 );
and ( n56253 , n56248 , n56252 );
buf ( n56254 , n20810 );
buf ( n56255 , n56254 );
and ( n56256 , n56255 , n20846 );
and ( n56257 , n56252 , n56256 );
and ( n56258 , n56248 , n56256 );
or ( n56259 , n56253 , n56257 , n56258 );
and ( n56260 , n56243 , n56259 );
and ( n56261 , n56227 , n56259 );
or ( n56262 , n56244 , n56260 , n56261 );
and ( n56263 , n56211 , n56262 );
xor ( n56264 , n55854 , n55858 );
xor ( n56265 , n56264 , n55863 );
xor ( n56266 , n55871 , n55875 );
xor ( n56267 , n56266 , n55880 );
and ( n56268 , n56265 , n56267 );
xor ( n56269 , n55896 , n55900 );
xor ( n56270 , n56269 , n55905 );
and ( n56271 , n56267 , n56270 );
and ( n56272 , n56265 , n56270 );
or ( n56273 , n56268 , n56271 , n56272 );
and ( n56274 , n56262 , n56273 );
and ( n56275 , n56211 , n56273 );
or ( n56276 , n56263 , n56274 , n56275 );
and ( n56277 , n56161 , n56276 );
and ( n56278 , n56095 , n56276 );
or ( n56279 , n56162 , n56277 , n56278 );
xor ( n56280 , n55764 , n55766 );
xor ( n56281 , n56280 , n55769 );
xor ( n56282 , n55778 , n55779 );
xor ( n56283 , n56282 , n55796 );
and ( n56284 , n56281 , n56283 );
xor ( n56285 , n55815 , n55824 );
xor ( n56286 , n56285 , n55834 );
and ( n56287 , n56283 , n56286 );
and ( n56288 , n56281 , n56286 );
or ( n56289 , n56284 , n56287 , n56288 );
xor ( n56290 , n55847 , n55866 );
xor ( n56291 , n56290 , n55883 );
xor ( n56292 , n55908 , n55924 );
xor ( n56293 , n56292 , n55935 );
and ( n56294 , n56291 , n56293 );
xor ( n56295 , n55940 , n55942 );
xor ( n56296 , n56295 , n55945 );
and ( n56297 , n56293 , n56296 );
and ( n56298 , n56291 , n56296 );
or ( n56299 , n56294 , n56297 , n56298 );
and ( n56300 , n56289 , n56299 );
xor ( n56301 , n55716 , n55717 );
xor ( n56302 , n56301 , n55719 );
and ( n56303 , n56299 , n56302 );
and ( n56304 , n56289 , n56302 );
or ( n56305 , n56300 , n56303 , n56304 );
and ( n56306 , n56279 , n56305 );
xor ( n56307 , n55729 , n55761 );
xor ( n56308 , n56307 , n55772 );
xor ( n56309 , n55799 , n55837 );
xor ( n56310 , n56309 , n55886 );
and ( n56311 , n56308 , n56310 );
xor ( n56312 , n55938 , n55948 );
xor ( n56313 , n56312 , n55951 );
and ( n56314 , n56310 , n56313 );
and ( n56315 , n56308 , n56313 );
or ( n56316 , n56311 , n56314 , n56315 );
and ( n56317 , n56305 , n56316 );
and ( n56318 , n56279 , n56316 );
or ( n56319 , n56306 , n56317 , n56318 );
and ( n56320 , n56051 , n56319 );
and ( n56321 , n56026 , n56319 );
or ( n56322 , n56052 , n56320 , n56321 );
and ( n56323 , n56023 , n56322 );
and ( n56324 , n56021 , n56322 );
or ( n56325 , n56024 , n56323 , n56324 );
xor ( n56326 , n56000 , n56002 );
xor ( n56327 , n56326 , n56005 );
and ( n56328 , n56325 , n56327 );
xor ( n56329 , n55722 , n55775 );
xor ( n56330 , n56329 , n55889 );
xor ( n56331 , n55954 , n55964 );
xor ( n56332 , n56331 , n55967 );
and ( n56333 , n56330 , n56332 );
xor ( n56334 , n55973 , n55975 );
xor ( n56335 , n56334 , n55978 );
and ( n56336 , n56332 , n56335 );
and ( n56337 , n56330 , n56335 );
or ( n56338 , n56333 , n56336 , n56337 );
xor ( n56339 , n55892 , n55970 );
xor ( n56340 , n56339 , n55981 );
and ( n56341 , n56338 , n56340 );
xor ( n56342 , n55986 , n55988 );
xor ( n56343 , n56342 , n55991 );
and ( n56344 , n56340 , n56343 );
and ( n56345 , n56338 , n56343 );
or ( n56346 , n56341 , n56344 , n56345 );
xor ( n56347 , n55984 , n55994 );
xor ( n56348 , n56347 , n55997 );
and ( n56349 , n56346 , n56348 );
xor ( n56350 , n55956 , n55958 );
xor ( n56351 , n56350 , n55961 );
xor ( n56352 , n55912 , n55916 );
xor ( n56353 , n56352 , n55921 );
xor ( n56354 , n55929 , n55933 );
buf ( n56355 , n56354 );
and ( n56356 , n56353 , n56355 );
xnor ( n56357 , n56069 , n56085 );
and ( n56358 , n56355 , n56357 );
and ( n56359 , n56353 , n56357 );
or ( n56360 , n56356 , n56358 , n56359 );
xnor ( n56361 , n56089 , n56091 );
and ( n56362 , n53639 , n45990 );
and ( n56363 , n53328 , n45988 );
nor ( n56364 , n56362 , n56363 );
xnor ( n56365 , n56364 , n45939 );
and ( n56366 , n54227 , n45886 );
and ( n56367 , n53922 , n45884 );
nor ( n56368 , n56366 , n56367 );
xnor ( n56369 , n56368 , n45824 );
and ( n56370 , n56365 , n56369 );
and ( n56371 , n54942 , n45777 );
and ( n56372 , n54604 , n45775 );
nor ( n56373 , n56371 , n56372 );
xnor ( n56374 , n56373 , n45734 );
and ( n56375 , n56369 , n56374 );
and ( n56376 , n56365 , n56374 );
or ( n56377 , n56370 , n56375 , n56376 );
and ( n56378 , n53041 , n46135 );
and ( n56379 , n52790 , n46133 );
nor ( n56380 , n56378 , n56379 );
xnor ( n56381 , n56380 , n46067 );
and ( n56382 , n55497 , n45702 );
and ( n56383 , n55143 , n45700 );
nor ( n56384 , n56382 , n56383 );
xnor ( n56385 , n56384 , n20841 );
and ( n56386 , n56381 , n56385 );
buf ( n56387 , n20812 );
buf ( n56388 , n56387 );
and ( n56389 , n56388 , n20846 );
and ( n56390 , n56385 , n56389 );
and ( n56391 , n56381 , n56389 );
or ( n56392 , n56386 , n56390 , n56391 );
or ( n56393 , n56377 , n56392 );
and ( n56394 , n56361 , n56393 );
xor ( n56395 , n35246 , n45590 );
buf ( n56396 , n56395 );
buf ( n56397 , n56396 );
buf ( n56398 , n56397 );
xor ( n56399 , n56057 , n56061 );
xor ( n56400 , n56399 , n56066 );
and ( n56401 , n56398 , n56400 );
buf ( n56402 , n56401 );
and ( n56403 , n56393 , n56402 );
and ( n56404 , n56361 , n56402 );
or ( n56405 , n56394 , n56403 , n56404 );
and ( n56406 , n56360 , n56405 );
xor ( n56407 , n56073 , n56077 );
xor ( n56408 , n56407 , n56082 );
xor ( n56409 , n56111 , n56115 );
xor ( n56410 , n56409 , n56120 );
and ( n56411 , n56408 , n56410 );
xnor ( n56412 , n56131 , n56135 );
and ( n56413 , n56410 , n56412 );
and ( n56414 , n56408 , n56412 );
or ( n56415 , n56411 , n56413 , n56414 );
xnor ( n56416 , n56140 , n56144 );
xnor ( n56417 , n56150 , n56154 );
and ( n56418 , n56416 , n56417 );
xnor ( n56419 , n56166 , n56170 );
and ( n56420 , n56417 , n56419 );
and ( n56421 , n56416 , n56419 );
or ( n56422 , n56418 , n56420 , n56421 );
and ( n56423 , n56415 , n56422 );
and ( n56424 , n48988 , n48394 );
and ( n56425 , n48709 , n48392 );
nor ( n56426 , n56424 , n56425 );
xnor ( n56427 , n56426 , n48220 );
and ( n56428 , n49374 , n48042 );
and ( n56429 , n49115 , n48040 );
nor ( n56430 , n56428 , n56429 );
xnor ( n56431 , n56430 , n47921 );
and ( n56432 , n56427 , n56431 );
and ( n56433 , n50195 , n47429 );
and ( n56434 , n49976 , n47427 );
nor ( n56435 , n56433 , n56434 );
xnor ( n56436 , n56435 , n47309 );
and ( n56437 , n56431 , n56436 );
and ( n56438 , n56427 , n56436 );
or ( n56439 , n56432 , n56437 , n56438 );
and ( n56440 , n46843 , n51221 );
and ( n56441 , n46750 , n51219 );
nor ( n56442 , n56440 , n56441 );
xnor ( n56443 , n56442 , n51000 );
and ( n56444 , n47090 , n50783 );
and ( n56445 , n46969 , n50781 );
nor ( n56446 , n56444 , n56445 );
xnor ( n56447 , n56446 , n50557 );
or ( n56448 , n56443 , n56447 );
and ( n56449 , n56439 , n56448 );
and ( n56450 , n46577 , n51750 );
and ( n56451 , n46530 , n51748 );
nor ( n56452 , n56450 , n56451 );
xnor ( n56453 , n56452 , n51520 );
and ( n56454 , n47351 , n50338 );
and ( n56455 , n47216 , n50336 );
nor ( n56456 , n56454 , n56455 );
xnor ( n56457 , n56456 , n50111 );
or ( n56458 , n56453 , n56457 );
and ( n56459 , n56448 , n56458 );
and ( n56460 , n56439 , n56458 );
or ( n56461 , n56449 , n56459 , n56460 );
and ( n56462 , n56422 , n56461 );
and ( n56463 , n56415 , n56461 );
or ( n56464 , n56423 , n56462 , n56463 );
and ( n56465 , n56405 , n56464 );
and ( n56466 , n56360 , n56464 );
or ( n56467 , n56406 , n56465 , n56466 );
and ( n56468 , n56351 , n56467 );
and ( n56469 , n48632 , n48740 );
and ( n56470 , n48384 , n48738 );
nor ( n56471 , n56469 , n56470 );
xnor ( n56472 , n56471 , n48571 );
and ( n56473 , n51510 , n46712 );
and ( n56474 , n51298 , n46710 );
nor ( n56475 , n56473 , n56474 );
xnor ( n56476 , n56475 , n46587 );
or ( n56477 , n56472 , n56476 );
and ( n56478 , n50625 , n47178 );
and ( n56479 , n50404 , n47176 );
nor ( n56480 , n56478 , n56479 );
xnor ( n56481 , n56480 , n47039 );
and ( n56482 , n51077 , n46911 );
and ( n56483 , n50726 , n46909 );
nor ( n56484 , n56482 , n56483 );
xnor ( n56485 , n56484 , n46802 );
or ( n56486 , n56481 , n56485 );
and ( n56487 , n56477 , n56486 );
and ( n56488 , n52612 , n46306 );
and ( n56489 , n52332 , n46304 );
nor ( n56490 , n56488 , n56489 );
xnor ( n56491 , n56490 , n46228 );
and ( n56492 , n56255 , n20852 );
and ( n56493 , n55756 , n20850 );
nor ( n56494 , n56492 , n56493 );
xnor ( n56495 , n56494 , n20860 );
or ( n56496 , n56491 , n56495 );
and ( n56497 , n56486 , n56496 );
and ( n56498 , n56477 , n56496 );
or ( n56499 , n56487 , n56497 , n56498 );
xor ( n56500 , n55503 , n56173 );
xor ( n56501 , n56173 , n56175 );
not ( n56502 , n56501 );
and ( n56503 , n56500 , n56502 );
and ( n56504 , n20855 , n56503 );
not ( n56505 , n56504 );
xnor ( n56506 , n56505 , n56178 );
and ( n56507 , n20864 , n55851 );
and ( n56508 , n20844 , n55849 );
nor ( n56509 , n56507 , n56508 );
xnor ( n56510 , n56509 , n55506 );
and ( n56511 , n56506 , n56510 );
and ( n56512 , n45763 , n55159 );
and ( n56513 , n45712 , n55157 );
nor ( n56514 , n56512 , n56513 );
xnor ( n56515 , n56514 , n54864 );
and ( n56516 , n56510 , n56515 );
and ( n56517 , n56506 , n56515 );
or ( n56518 , n56511 , n56516 , n56517 );
and ( n56519 , n45843 , n54535 );
and ( n56520 , n45794 , n54533 );
nor ( n56521 , n56519 , n56520 );
xnor ( n56522 , n56521 , n54237 );
and ( n56523 , n45963 , n53928 );
and ( n56524 , n45907 , n53926 );
nor ( n56525 , n56523 , n56524 );
xnor ( n56526 , n56525 , n53652 );
and ( n56527 , n56522 , n56526 );
and ( n56528 , n46100 , n53357 );
and ( n56529 , n46041 , n53355 );
nor ( n56530 , n56528 , n56529 );
xnor ( n56531 , n56530 , n53060 );
and ( n56532 , n56526 , n56531 );
and ( n56533 , n56522 , n56531 );
or ( n56534 , n56527 , n56532 , n56533 );
and ( n56535 , n56518 , n56534 );
and ( n56536 , n46264 , n52799 );
and ( n56537 , n46169 , n52797 );
nor ( n56538 , n56536 , n56537 );
xnor ( n56539 , n56538 , n52538 );
and ( n56540 , n46445 , n52269 );
and ( n56541 , n46345 , n52267 );
nor ( n56542 , n56540 , n56541 );
xnor ( n56543 , n56542 , n52008 );
and ( n56544 , n56539 , n56543 );
and ( n56545 , n47647 , n49896 );
and ( n56546 , n47474 , n49894 );
nor ( n56547 , n56545 , n56546 );
xnor ( n56548 , n56547 , n49711 );
and ( n56549 , n56543 , n56548 );
and ( n56550 , n56539 , n56548 );
or ( n56551 , n56544 , n56549 , n56550 );
and ( n56552 , n56534 , n56551 );
and ( n56553 , n56518 , n56551 );
or ( n56554 , n56535 , n56552 , n56553 );
and ( n56555 , n56499 , n56554 );
and ( n56556 , n47962 , n49513 );
and ( n56557 , n47778 , n49511 );
nor ( n56558 , n56556 , n56557 );
xnor ( n56559 , n56558 , n49310 );
and ( n56560 , n48272 , n49121 );
and ( n56561 , n48108 , n49119 );
nor ( n56562 , n56560 , n56561 );
xnor ( n56563 , n56562 , n48932 );
and ( n56564 , n56559 , n56563 );
and ( n56565 , n49781 , n47734 );
and ( n56566 , n49570 , n47732 );
nor ( n56567 , n56565 , n56566 );
xnor ( n56568 , n56567 , n47606 );
and ( n56569 , n56563 , n56568 );
and ( n56570 , n56559 , n56568 );
or ( n56571 , n56564 , n56569 , n56570 );
and ( n56572 , n52082 , n46496 );
and ( n56573 , n51734 , n46494 );
nor ( n56574 , n56572 , n56573 );
xnor ( n56575 , n56574 , n46402 );
xor ( n56576 , n35248 , n45589 );
buf ( n56577 , n56576 );
buf ( n56578 , n56577 );
buf ( n56579 , n56578 );
and ( n56580 , n56575 , n56579 );
buf ( n56581 , n56580 );
and ( n56582 , n56571 , n56581 );
xor ( n56583 , n56179 , n56183 );
xor ( n56584 , n56583 , n56188 );
and ( n56585 , n56581 , n56584 );
and ( n56586 , n56571 , n56584 );
or ( n56587 , n56582 , n56585 , n56586 );
and ( n56588 , n56554 , n56587 );
and ( n56589 , n56499 , n56587 );
or ( n56590 , n56555 , n56588 , n56589 );
xor ( n56591 , n56196 , n56200 );
xor ( n56592 , n56591 , n56205 );
xor ( n56593 , n56215 , n56219 );
xor ( n56594 , n56593 , n56224 );
and ( n56595 , n56592 , n56594 );
xor ( n56596 , n56231 , n56235 );
xor ( n56597 , n56596 , n56240 );
and ( n56598 , n56594 , n56597 );
and ( n56599 , n56592 , n56597 );
or ( n56600 , n56595 , n56598 , n56599 );
xor ( n56601 , n56097 , n56099 );
xor ( n56602 , n56601 , n56101 );
and ( n56603 , n56600 , n56602 );
xor ( n56604 , n56105 , n56106 );
xor ( n56605 , n56604 , n56123 );
and ( n56606 , n56602 , n56605 );
and ( n56607 , n56600 , n56605 );
or ( n56608 , n56603 , n56606 , n56607 );
and ( n56609 , n56590 , n56608 );
xor ( n56610 , n56136 , n56145 );
xor ( n56611 , n56610 , n56155 );
xor ( n56612 , n56171 , n56191 );
xor ( n56613 , n56612 , n56208 );
and ( n56614 , n56611 , n56613 );
xor ( n56615 , n56227 , n56243 );
xor ( n56616 , n56615 , n56259 );
and ( n56617 , n56613 , n56616 );
and ( n56618 , n56611 , n56616 );
or ( n56619 , n56614 , n56617 , n56618 );
and ( n56620 , n56608 , n56619 );
and ( n56621 , n56590 , n56619 );
or ( n56622 , n56609 , n56620 , n56621 );
and ( n56623 , n56467 , n56622 );
and ( n56624 , n56351 , n56622 );
or ( n56625 , n56468 , n56623 , n56624 );
xor ( n56626 , n56038 , n56040 );
xor ( n56627 , n56626 , n56042 );
xor ( n56628 , n56053 , n56086 );
xor ( n56629 , n56628 , n56092 );
and ( n56630 , n56627 , n56629 );
xor ( n56631 , n56104 , n56126 );
xor ( n56632 , n56631 , n56158 );
and ( n56633 , n56629 , n56632 );
and ( n56634 , n56627 , n56632 );
or ( n56635 , n56630 , n56633 , n56634 );
xor ( n56636 , n56211 , n56262 );
xor ( n56637 , n56636 , n56273 );
xor ( n56638 , n56281 , n56283 );
xor ( n56639 , n56638 , n56286 );
and ( n56640 , n56637 , n56639 );
xor ( n56641 , n56291 , n56293 );
xor ( n56642 , n56641 , n56296 );
and ( n56643 , n56639 , n56642 );
and ( n56644 , n56637 , n56642 );
or ( n56645 , n56640 , n56643 , n56644 );
and ( n56646 , n56635 , n56645 );
xor ( n56647 , n56033 , n56035 );
xor ( n56648 , n56647 , n56045 );
and ( n56649 , n56645 , n56648 );
and ( n56650 , n56635 , n56648 );
or ( n56651 , n56646 , n56649 , n56650 );
and ( n56652 , n56625 , n56651 );
xor ( n56653 , n56095 , n56161 );
xor ( n56654 , n56653 , n56276 );
xor ( n56655 , n56289 , n56299 );
xor ( n56656 , n56655 , n56302 );
and ( n56657 , n56654 , n56656 );
xor ( n56658 , n56308 , n56310 );
xor ( n56659 , n56658 , n56313 );
and ( n56660 , n56656 , n56659 );
and ( n56661 , n56654 , n56659 );
or ( n56662 , n56657 , n56660 , n56661 );
and ( n56663 , n56651 , n56662 );
and ( n56664 , n56625 , n56662 );
or ( n56665 , n56652 , n56663 , n56664 );
xor ( n56666 , n56028 , n56030 );
xor ( n56667 , n56666 , n56048 );
xor ( n56668 , n56279 , n56305 );
xor ( n56669 , n56668 , n56316 );
and ( n56670 , n56667 , n56669 );
xor ( n56671 , n56330 , n56332 );
xor ( n56672 , n56671 , n56335 );
and ( n56673 , n56669 , n56672 );
and ( n56674 , n56667 , n56672 );
or ( n56675 , n56670 , n56673 , n56674 );
and ( n56676 , n56665 , n56675 );
xor ( n56677 , n56026 , n56051 );
xor ( n56678 , n56677 , n56319 );
and ( n56679 , n56675 , n56678 );
and ( n56680 , n56665 , n56678 );
or ( n56681 , n56676 , n56679 , n56680 );
and ( n56682 , n56348 , n56681 );
and ( n56683 , n56346 , n56681 );
or ( n56684 , n56349 , n56682 , n56683 );
and ( n56685 , n56327 , n56684 );
and ( n56686 , n56325 , n56684 );
or ( n56687 , n56328 , n56685 , n56686 );
or ( n56688 , n56019 , n56687 );
and ( n56689 , n56016 , n56688 );
and ( n56690 , n56014 , n56688 );
or ( n56691 , n56017 , n56689 , n56690 );
and ( n56692 , n55712 , n56691 );
and ( n56693 , n55710 , n56691 );
or ( n56694 , n55713 , n56692 , n56693 );
or ( n56695 , n55374 , n56694 );
and ( n56696 , n55372 , n56695 );
xor ( n56697 , n55372 , n56695 );
xnor ( n56698 , n55374 , n56694 );
xor ( n56699 , n55710 , n55712 );
xor ( n56700 , n56699 , n56691 );
not ( n56701 , n56700 );
xor ( n56702 , n56014 , n56016 );
xor ( n56703 , n56702 , n56688 );
xnor ( n56704 , n56019 , n56687 );
xor ( n56705 , n56021 , n56023 );
xor ( n56706 , n56705 , n56322 );
xor ( n56707 , n56338 , n56340 );
xor ( n56708 , n56707 , n56343 );
xor ( n56709 , n56265 , n56267 );
xor ( n56710 , n56709 , n56270 );
xor ( n56711 , n56248 , n56252 );
xor ( n56712 , n56711 , n56256 );
xnor ( n56713 , n56377 , n56392 );
and ( n56714 , n56712 , n56713 );
xor ( n56715 , n56365 , n56369 );
xor ( n56716 , n56715 , n56374 );
xor ( n56717 , n56381 , n56385 );
xor ( n56718 , n56717 , n56389 );
or ( n56719 , n56716 , n56718 );
and ( n56720 , n56713 , n56719 );
and ( n56721 , n56712 , n56719 );
or ( n56722 , n56714 , n56720 , n56721 );
and ( n56723 , n56710 , n56722 );
xor ( n56724 , n56427 , n56431 );
xor ( n56725 , n56724 , n56436 );
xnor ( n56726 , n56443 , n56447 );
and ( n56727 , n56725 , n56726 );
xnor ( n56728 , n56453 , n56457 );
and ( n56729 , n56726 , n56728 );
and ( n56730 , n56725 , n56728 );
or ( n56731 , n56727 , n56729 , n56730 );
xnor ( n56732 , n56472 , n56476 );
xnor ( n56733 , n56481 , n56485 );
and ( n56734 , n56732 , n56733 );
xnor ( n56735 , n56491 , n56495 );
and ( n56736 , n56733 , n56735 );
and ( n56737 , n56732 , n56735 );
or ( n56738 , n56734 , n56736 , n56737 );
and ( n56739 , n56731 , n56738 );
and ( n56740 , n49570 , n48042 );
and ( n56741 , n49374 , n48040 );
nor ( n56742 , n56740 , n56741 );
xnor ( n56743 , n56742 , n47921 );
and ( n56744 , n50726 , n47178 );
and ( n56745 , n50625 , n47176 );
nor ( n56746 , n56744 , n56745 );
xnor ( n56747 , n56746 , n47039 );
and ( n56748 , n56743 , n56747 );
and ( n56749 , n51734 , n46712 );
and ( n56750 , n51510 , n46710 );
nor ( n56751 , n56749 , n56750 );
xnor ( n56752 , n56751 , n46587 );
and ( n56753 , n56747 , n56752 );
and ( n56754 , n56743 , n56752 );
or ( n56755 , n56748 , n56753 , n56754 );
and ( n56756 , n48709 , n48740 );
and ( n56757 , n48632 , n48738 );
nor ( n56758 , n56756 , n56757 );
xnor ( n56759 , n56758 , n48571 );
and ( n56760 , n49976 , n47734 );
and ( n56761 , n49781 , n47732 );
nor ( n56762 , n56760 , n56761 );
xnor ( n56763 , n56762 , n47606 );
and ( n56764 , n56759 , n56763 );
and ( n56765 , n50404 , n47429 );
and ( n56766 , n50195 , n47427 );
nor ( n56767 , n56765 , n56766 );
xnor ( n56768 , n56767 , n47309 );
and ( n56769 , n56763 , n56768 );
and ( n56770 , n56759 , n56768 );
or ( n56771 , n56764 , n56769 , n56770 );
and ( n56772 , n56755 , n56771 );
and ( n56773 , n47474 , n50338 );
and ( n56774 , n47351 , n50336 );
nor ( n56775 , n56773 , n56774 );
xnor ( n56776 , n56775 , n50111 );
and ( n56777 , n47778 , n49896 );
and ( n56778 , n47647 , n49894 );
nor ( n56779 , n56777 , n56778 );
xnor ( n56780 , n56779 , n49711 );
or ( n56781 , n56776 , n56780 );
and ( n56782 , n56771 , n56781 );
and ( n56783 , n56755 , n56781 );
or ( n56784 , n56772 , n56782 , n56783 );
and ( n56785 , n56738 , n56784 );
and ( n56786 , n56731 , n56784 );
or ( n56787 , n56739 , n56785 , n56786 );
and ( n56788 , n56722 , n56787 );
and ( n56789 , n56710 , n56787 );
or ( n56790 , n56723 , n56788 , n56789 );
and ( n56791 , n49115 , n48394 );
and ( n56792 , n48988 , n48392 );
nor ( n56793 , n56791 , n56792 );
xnor ( n56794 , n56793 , n48220 );
and ( n56795 , n51298 , n46911 );
and ( n56796 , n51077 , n46909 );
nor ( n56797 , n56795 , n56796 );
xnor ( n56798 , n56797 , n46802 );
or ( n56799 , n56794 , n56798 );
and ( n56800 , n53328 , n46135 );
and ( n56801 , n53041 , n46133 );
nor ( n56802 , n56800 , n56801 );
xnor ( n56803 , n56802 , n46067 );
and ( n56804 , n55756 , n45702 );
and ( n56805 , n55497 , n45700 );
nor ( n56806 , n56804 , n56805 );
xnor ( n56807 , n56806 , n20841 );
or ( n56808 , n56803 , n56807 );
and ( n56809 , n56799 , n56808 );
and ( n56810 , n53922 , n45990 );
and ( n56811 , n53639 , n45988 );
nor ( n56812 , n56810 , n56811 );
xnor ( n56813 , n56812 , n45939 );
and ( n56814 , n56388 , n20852 );
and ( n56815 , n56255 , n20850 );
nor ( n56816 , n56814 , n56815 );
xnor ( n56817 , n56816 , n20860 );
or ( n56818 , n56813 , n56817 );
and ( n56819 , n56808 , n56818 );
and ( n56820 , n56799 , n56818 );
or ( n56821 , n56809 , n56819 , n56820 );
not ( n56822 , n56175 );
and ( n56823 , n20844 , n56503 );
and ( n56824 , n20855 , n56501 );
nor ( n56825 , n56823 , n56824 );
xnor ( n56826 , n56825 , n56178 );
and ( n56827 , n56822 , n56826 );
and ( n56828 , n45712 , n55851 );
and ( n56829 , n20864 , n55849 );
nor ( n56830 , n56828 , n56829 );
xnor ( n56831 , n56830 , n55506 );
and ( n56832 , n56826 , n56831 );
and ( n56833 , n56822 , n56831 );
or ( n56834 , n56827 , n56832 , n56833 );
and ( n56835 , n45794 , n55159 );
and ( n56836 , n45763 , n55157 );
nor ( n56837 , n56835 , n56836 );
xnor ( n56838 , n56837 , n54864 );
and ( n56839 , n45907 , n54535 );
and ( n56840 , n45843 , n54533 );
nor ( n56841 , n56839 , n56840 );
xnor ( n56842 , n56841 , n54237 );
and ( n56843 , n56838 , n56842 );
and ( n56844 , n46041 , n53928 );
and ( n56845 , n45963 , n53926 );
nor ( n56846 , n56844 , n56845 );
xnor ( n56847 , n56846 , n53652 );
and ( n56848 , n56842 , n56847 );
and ( n56849 , n56838 , n56847 );
or ( n56850 , n56843 , n56848 , n56849 );
and ( n56851 , n56834 , n56850 );
and ( n56852 , n46169 , n53357 );
and ( n56853 , n46100 , n53355 );
nor ( n56854 , n56852 , n56853 );
xnor ( n56855 , n56854 , n53060 );
and ( n56856 , n46345 , n52799 );
and ( n56857 , n46264 , n52797 );
nor ( n56858 , n56856 , n56857 );
xnor ( n56859 , n56858 , n52538 );
and ( n56860 , n56855 , n56859 );
and ( n56861 , n46530 , n52269 );
and ( n56862 , n46445 , n52267 );
nor ( n56863 , n56861 , n56862 );
xnor ( n56864 , n56863 , n52008 );
and ( n56865 , n56859 , n56864 );
and ( n56866 , n56855 , n56864 );
or ( n56867 , n56860 , n56865 , n56866 );
and ( n56868 , n56850 , n56867 );
and ( n56869 , n56834 , n56867 );
or ( n56870 , n56851 , n56868 , n56869 );
and ( n56871 , n56821 , n56870 );
and ( n56872 , n46750 , n51750 );
and ( n56873 , n46577 , n51748 );
nor ( n56874 , n56872 , n56873 );
xnor ( n56875 , n56874 , n51520 );
and ( n56876 , n46969 , n51221 );
and ( n56877 , n46843 , n51219 );
nor ( n56878 , n56876 , n56877 );
xnor ( n56879 , n56878 , n51000 );
and ( n56880 , n56875 , n56879 );
and ( n56881 , n47216 , n50783 );
and ( n56882 , n47090 , n50781 );
nor ( n56883 , n56881 , n56882 );
xnor ( n56884 , n56883 , n50557 );
and ( n56885 , n56879 , n56884 );
and ( n56886 , n56875 , n56884 );
or ( n56887 , n56880 , n56885 , n56886 );
and ( n56888 , n48108 , n49513 );
and ( n56889 , n47962 , n49511 );
nor ( n56890 , n56888 , n56889 );
xnor ( n56891 , n56890 , n49310 );
and ( n56892 , n48384 , n49121 );
and ( n56893 , n48272 , n49119 );
nor ( n56894 , n56892 , n56893 );
xnor ( n56895 , n56894 , n48932 );
and ( n56896 , n56891 , n56895 );
and ( n56897 , n52332 , n46496 );
and ( n56898 , n52082 , n46494 );
nor ( n56899 , n56897 , n56898 );
xnor ( n56900 , n56899 , n46402 );
and ( n56901 , n56895 , n56900 );
and ( n56902 , n56891 , n56900 );
or ( n56903 , n56896 , n56901 , n56902 );
and ( n56904 , n56887 , n56903 );
and ( n56905 , n52790 , n46306 );
and ( n56906 , n52612 , n46304 );
nor ( n56907 , n56905 , n56906 );
xnor ( n56908 , n56907 , n46228 );
and ( n56909 , n54604 , n45886 );
and ( n56910 , n54227 , n45884 );
nor ( n56911 , n56909 , n56910 );
xnor ( n56912 , n56911 , n45824 );
and ( n56913 , n56908 , n56912 );
buf ( n56914 , n20814 );
buf ( n56915 , n56914 );
and ( n56916 , n56915 , n20846 );
and ( n56917 , n56912 , n56916 );
and ( n56918 , n56908 , n56916 );
or ( n56919 , n56913 , n56917 , n56918 );
and ( n56920 , n56903 , n56919 );
and ( n56921 , n56887 , n56919 );
or ( n56922 , n56904 , n56920 , n56921 );
and ( n56923 , n56870 , n56922 );
and ( n56924 , n56821 , n56922 );
or ( n56925 , n56871 , n56923 , n56924 );
xor ( n56926 , n56506 , n56510 );
xor ( n56927 , n56926 , n56515 );
xor ( n56928 , n56522 , n56526 );
xor ( n56929 , n56928 , n56531 );
and ( n56930 , n56927 , n56929 );
xor ( n56931 , n56539 , n56543 );
xor ( n56932 , n56931 , n56548 );
and ( n56933 , n56929 , n56932 );
and ( n56934 , n56927 , n56932 );
or ( n56935 , n56930 , n56933 , n56934 );
buf ( n56936 , n56398 );
xor ( n56937 , n56936 , n56400 );
and ( n56938 , n56935 , n56937 );
xor ( n56939 , n56408 , n56410 );
xor ( n56940 , n56939 , n56412 );
and ( n56941 , n56937 , n56940 );
and ( n56942 , n56935 , n56940 );
or ( n56943 , n56938 , n56941 , n56942 );
and ( n56944 , n56925 , n56943 );
xor ( n56945 , n56416 , n56417 );
xor ( n56946 , n56945 , n56419 );
xor ( n56947 , n56439 , n56448 );
xor ( n56948 , n56947 , n56458 );
and ( n56949 , n56946 , n56948 );
xor ( n56950 , n56477 , n56486 );
xor ( n56951 , n56950 , n56496 );
and ( n56952 , n56948 , n56951 );
and ( n56953 , n56946 , n56951 );
or ( n56954 , n56949 , n56952 , n56953 );
and ( n56955 , n56943 , n56954 );
and ( n56956 , n56925 , n56954 );
or ( n56957 , n56944 , n56955 , n56956 );
and ( n56958 , n56790 , n56957 );
xor ( n56959 , n56518 , n56534 );
xor ( n56960 , n56959 , n56551 );
xor ( n56961 , n56571 , n56581 );
xor ( n56962 , n56961 , n56584 );
and ( n56963 , n56960 , n56962 );
xor ( n56964 , n56592 , n56594 );
xor ( n56965 , n56964 , n56597 );
and ( n56966 , n56962 , n56965 );
and ( n56967 , n56960 , n56965 );
or ( n56968 , n56963 , n56966 , n56967 );
xor ( n56969 , n56353 , n56355 );
xor ( n56970 , n56969 , n56357 );
and ( n56971 , n56968 , n56970 );
xor ( n56972 , n56361 , n56393 );
xor ( n56973 , n56972 , n56402 );
and ( n56974 , n56970 , n56973 );
and ( n56975 , n56968 , n56973 );
or ( n56976 , n56971 , n56974 , n56975 );
and ( n56977 , n56957 , n56976 );
and ( n56978 , n56790 , n56976 );
or ( n56979 , n56958 , n56977 , n56978 );
xor ( n56980 , n56415 , n56422 );
xor ( n56981 , n56980 , n56461 );
xor ( n56982 , n56499 , n56554 );
xor ( n56983 , n56982 , n56587 );
and ( n56984 , n56981 , n56983 );
xor ( n56985 , n56600 , n56602 );
xor ( n56986 , n56985 , n56605 );
and ( n56987 , n56983 , n56986 );
and ( n56988 , n56981 , n56986 );
or ( n56989 , n56984 , n56987 , n56988 );
xor ( n56990 , n56360 , n56405 );
xor ( n56991 , n56990 , n56464 );
and ( n56992 , n56989 , n56991 );
xor ( n56993 , n56590 , n56608 );
xor ( n56994 , n56993 , n56619 );
and ( n56995 , n56991 , n56994 );
and ( n56996 , n56989 , n56994 );
or ( n56997 , n56992 , n56995 , n56996 );
and ( n56998 , n56979 , n56997 );
xor ( n56999 , n56351 , n56467 );
xor ( n57000 , n56999 , n56622 );
and ( n57001 , n56997 , n57000 );
and ( n57002 , n56979 , n57000 );
or ( n57003 , n56998 , n57001 , n57002 );
xor ( n57004 , n56625 , n56651 );
xor ( n57005 , n57004 , n56662 );
and ( n57006 , n57003 , n57005 );
xor ( n57007 , n56667 , n56669 );
xor ( n57008 , n57007 , n56672 );
and ( n57009 , n57005 , n57008 );
and ( n57010 , n57003 , n57008 );
or ( n57011 , n57006 , n57009 , n57010 );
and ( n57012 , n56708 , n57011 );
xor ( n57013 , n56665 , n56675 );
xor ( n57014 , n57013 , n56678 );
and ( n57015 , n57011 , n57014 );
and ( n57016 , n56708 , n57014 );
or ( n57017 , n57012 , n57015 , n57016 );
and ( n57018 , n56706 , n57017 );
xor ( n57019 , n56346 , n56348 );
xor ( n57020 , n57019 , n56681 );
and ( n57021 , n57017 , n57020 );
and ( n57022 , n56706 , n57020 );
or ( n57023 , n57018 , n57021 , n57022 );
xor ( n57024 , n56325 , n56327 );
xor ( n57025 , n57024 , n56684 );
and ( n57026 , n57023 , n57025 );
xor ( n57027 , n57023 , n57025 );
xor ( n57028 , n56706 , n57017 );
xor ( n57029 , n57028 , n57020 );
xor ( n57030 , n56708 , n57011 );
xor ( n57031 , n57030 , n57014 );
xor ( n57032 , n56635 , n56645 );
xor ( n57033 , n57032 , n56648 );
xor ( n57034 , n56654 , n56656 );
xor ( n57035 , n57034 , n56659 );
and ( n57036 , n57033 , n57035 );
xor ( n57037 , n56627 , n56629 );
xor ( n57038 , n57037 , n56632 );
xor ( n57039 , n56637 , n56639 );
xor ( n57040 , n57039 , n56642 );
and ( n57041 , n57038 , n57040 );
xor ( n57042 , n56611 , n56613 );
xor ( n57043 , n57042 , n56616 );
xor ( n57044 , n56559 , n56563 );
xor ( n57045 , n57044 , n56568 );
xor ( n57046 , n56575 , n56579 );
buf ( n57047 , n57046 );
and ( n57048 , n57045 , n57047 );
xnor ( n57049 , n56716 , n56718 );
and ( n57050 , n57047 , n57049 );
and ( n57051 , n57045 , n57049 );
or ( n57052 , n57048 , n57050 , n57051 );
and ( n57053 , n48988 , n48740 );
and ( n57054 , n48709 , n48738 );
nor ( n57055 , n57053 , n57054 );
xnor ( n57056 , n57055 , n48571 );
and ( n57057 , n50195 , n47734 );
and ( n57058 , n49976 , n47732 );
nor ( n57059 , n57057 , n57058 );
xnor ( n57060 , n57059 , n47606 );
and ( n57061 , n57056 , n57060 );
buf ( n57062 , n20816 );
buf ( n57063 , n57062 );
and ( n57064 , n57063 , n20846 );
and ( n57065 , n57060 , n57064 );
and ( n57066 , n57056 , n57064 );
or ( n57067 , n57061 , n57065 , n57066 );
and ( n57068 , n55143 , n45777 );
and ( n57069 , n54942 , n45775 );
nor ( n57070 , n57068 , n57069 );
xnor ( n57071 , n57070 , n45734 );
and ( n57072 , n57067 , n57071 );
xor ( n57073 , n56759 , n56763 );
xor ( n57074 , n57073 , n56768 );
and ( n57075 , n57071 , n57074 );
and ( n57076 , n57067 , n57074 );
or ( n57077 , n57072 , n57075 , n57076 );
xor ( n57078 , n35500 , n45587 );
buf ( n57079 , n57078 );
buf ( n57080 , n57079 );
buf ( n57081 , n57080 );
xor ( n57082 , n56743 , n56747 );
xor ( n57083 , n57082 , n56752 );
and ( n57084 , n57081 , n57083 );
buf ( n57085 , n57084 );
and ( n57086 , n57077 , n57085 );
xnor ( n57087 , n56776 , n56780 );
xnor ( n57088 , n56794 , n56798 );
and ( n57089 , n57087 , n57088 );
xnor ( n57090 , n56803 , n56807 );
and ( n57091 , n57088 , n57090 );
and ( n57092 , n57087 , n57090 );
or ( n57093 , n57089 , n57091 , n57092 );
and ( n57094 , n57085 , n57093 );
and ( n57095 , n57077 , n57093 );
or ( n57096 , n57086 , n57094 , n57095 );
and ( n57097 , n57052 , n57096 );
xnor ( n57098 , n56813 , n56817 );
and ( n57099 , n46577 , n52269 );
and ( n57100 , n46530 , n52267 );
nor ( n57101 , n57099 , n57100 );
xnor ( n57102 , n57101 , n52008 );
and ( n57103 , n46843 , n51750 );
and ( n57104 , n46750 , n51748 );
nor ( n57105 , n57103 , n57104 );
xnor ( n57106 , n57105 , n51520 );
and ( n57107 , n57102 , n57106 );
and ( n57108 , n47351 , n50783 );
and ( n57109 , n47216 , n50781 );
nor ( n57110 , n57108 , n57109 );
xnor ( n57111 , n57110 , n50557 );
and ( n57112 , n57106 , n57111 );
and ( n57113 , n57102 , n57111 );
or ( n57114 , n57107 , n57112 , n57113 );
and ( n57115 , n57098 , n57114 );
and ( n57116 , n49374 , n48394 );
and ( n57117 , n49115 , n48392 );
nor ( n57118 , n57116 , n57117 );
xnor ( n57119 , n57118 , n48220 );
and ( n57120 , n50625 , n47429 );
and ( n57121 , n50404 , n47427 );
nor ( n57122 , n57120 , n57121 );
xnor ( n57123 , n57122 , n47309 );
and ( n57124 , n57119 , n57123 );
and ( n57125 , n52082 , n46712 );
and ( n57126 , n51734 , n46710 );
nor ( n57127 , n57125 , n57126 );
xnor ( n57128 , n57127 , n46587 );
and ( n57129 , n57123 , n57128 );
and ( n57130 , n57119 , n57128 );
or ( n57131 , n57124 , n57129 , n57130 );
and ( n57132 , n57114 , n57131 );
and ( n57133 , n57098 , n57131 );
or ( n57134 , n57115 , n57132 , n57133 );
and ( n57135 , n54227 , n45990 );
and ( n57136 , n53922 , n45988 );
nor ( n57137 , n57135 , n57136 );
xnor ( n57138 , n57137 , n45939 );
and ( n57139 , n55497 , n45777 );
and ( n57140 , n55143 , n45775 );
nor ( n57141 , n57139 , n57140 );
xnor ( n57142 , n57141 , n45734 );
and ( n57143 , n57138 , n57142 );
and ( n57144 , n56255 , n45702 );
and ( n57145 , n55756 , n45700 );
nor ( n57146 , n57144 , n57145 );
xnor ( n57147 , n57146 , n20841 );
and ( n57148 , n57142 , n57147 );
and ( n57149 , n57138 , n57147 );
or ( n57150 , n57143 , n57148 , n57149 );
and ( n57151 , n47647 , n50338 );
and ( n57152 , n47474 , n50336 );
nor ( n57153 , n57151 , n57152 );
xnor ( n57154 , n57153 , n50111 );
and ( n57155 , n47962 , n49896 );
and ( n57156 , n47778 , n49894 );
nor ( n57157 , n57155 , n57156 );
xnor ( n57158 , n57157 , n49711 );
or ( n57159 , n57154 , n57158 );
and ( n57160 , n57150 , n57159 );
and ( n57161 , n49781 , n48042 );
and ( n57162 , n49570 , n48040 );
nor ( n57163 , n57161 , n57162 );
xnor ( n57164 , n57163 , n47921 );
and ( n57165 , n51510 , n46911 );
and ( n57166 , n51298 , n46909 );
nor ( n57167 , n57165 , n57166 );
xnor ( n57168 , n57167 , n46802 );
or ( n57169 , n57164 , n57168 );
and ( n57170 , n57159 , n57169 );
and ( n57171 , n57150 , n57169 );
or ( n57172 , n57160 , n57170 , n57171 );
and ( n57173 , n57134 , n57172 );
and ( n57174 , n53041 , n46306 );
and ( n57175 , n52790 , n46304 );
nor ( n57176 , n57174 , n57175 );
xnor ( n57177 , n57176 , n46228 );
and ( n57178 , n53639 , n46135 );
and ( n57179 , n53328 , n46133 );
nor ( n57180 , n57178 , n57179 );
xnor ( n57181 , n57180 , n46067 );
or ( n57182 , n57177 , n57181 );
buf ( n57183 , n17572 );
buf ( n57184 , n57183 );
xor ( n57185 , n56175 , n57184 );
not ( n57186 , n57184 );
and ( n57187 , n57185 , n57186 );
and ( n57188 , n20855 , n57187 );
not ( n57189 , n57188 );
xnor ( n57190 , n57189 , n56175 );
and ( n57191 , n20864 , n56503 );
and ( n57192 , n20844 , n56501 );
nor ( n57193 , n57191 , n57192 );
xnor ( n57194 , n57193 , n56178 );
and ( n57195 , n57190 , n57194 );
and ( n57196 , n45763 , n55851 );
and ( n57197 , n45712 , n55849 );
nor ( n57198 , n57196 , n57197 );
xnor ( n57199 , n57198 , n55506 );
and ( n57200 , n57194 , n57199 );
and ( n57201 , n57190 , n57199 );
or ( n57202 , n57195 , n57200 , n57201 );
and ( n57203 , n57182 , n57202 );
and ( n57204 , n45843 , n55159 );
and ( n57205 , n45794 , n55157 );
nor ( n57206 , n57204 , n57205 );
xnor ( n57207 , n57206 , n54864 );
and ( n57208 , n45963 , n54535 );
and ( n57209 , n45907 , n54533 );
nor ( n57210 , n57208 , n57209 );
xnor ( n57211 , n57210 , n54237 );
and ( n57212 , n57207 , n57211 );
and ( n57213 , n46100 , n53928 );
and ( n57214 , n46041 , n53926 );
nor ( n57215 , n57213 , n57214 );
xnor ( n57216 , n57215 , n53652 );
and ( n57217 , n57211 , n57216 );
and ( n57218 , n57207 , n57216 );
or ( n57219 , n57212 , n57217 , n57218 );
and ( n57220 , n57202 , n57219 );
and ( n57221 , n57182 , n57219 );
or ( n57222 , n57203 , n57220 , n57221 );
and ( n57223 , n57172 , n57222 );
and ( n57224 , n57134 , n57222 );
or ( n57225 , n57173 , n57223 , n57224 );
and ( n57226 , n57096 , n57225 );
and ( n57227 , n57052 , n57225 );
or ( n57228 , n57097 , n57226 , n57227 );
and ( n57229 , n57043 , n57228 );
and ( n57230 , n46264 , n53357 );
and ( n57231 , n46169 , n53355 );
nor ( n57232 , n57230 , n57231 );
xnor ( n57233 , n57232 , n53060 );
and ( n57234 , n46445 , n52799 );
and ( n57235 , n46345 , n52797 );
nor ( n57236 , n57234 , n57235 );
xnor ( n57237 , n57236 , n52538 );
and ( n57238 , n57233 , n57237 );
and ( n57239 , n47090 , n51221 );
and ( n57240 , n46969 , n51219 );
nor ( n57241 , n57239 , n57240 );
xnor ( n57242 , n57241 , n51000 );
and ( n57243 , n57237 , n57242 );
and ( n57244 , n57233 , n57242 );
or ( n57245 , n57238 , n57243 , n57244 );
and ( n57246 , n48272 , n49513 );
and ( n57247 , n48108 , n49511 );
nor ( n57248 , n57246 , n57247 );
xnor ( n57249 , n57248 , n49310 );
and ( n57250 , n48632 , n49121 );
and ( n57251 , n48384 , n49119 );
nor ( n57252 , n57250 , n57251 );
xnor ( n57253 , n57252 , n48932 );
and ( n57254 , n57249 , n57253 );
and ( n57255 , n51077 , n47178 );
and ( n57256 , n50726 , n47176 );
nor ( n57257 , n57255 , n57256 );
xnor ( n57258 , n57257 , n47039 );
and ( n57259 , n57253 , n57258 );
and ( n57260 , n57249 , n57258 );
or ( n57261 , n57254 , n57259 , n57260 );
and ( n57262 , n57245 , n57261 );
and ( n57263 , n52612 , n46496 );
and ( n57264 , n52332 , n46494 );
nor ( n57265 , n57263 , n57264 );
xnor ( n57266 , n57265 , n46402 );
and ( n57267 , n56915 , n20852 );
and ( n57268 , n56388 , n20850 );
nor ( n57269 , n57267 , n57268 );
xnor ( n57270 , n57269 , n20860 );
and ( n57271 , n57266 , n57270 );
xor ( n57272 , n39385 , n45585 );
buf ( n57273 , n57272 );
buf ( n57274 , n57273 );
buf ( n57275 , n57274 );
and ( n57276 , n57270 , n57275 );
and ( n57277 , n57266 , n57275 );
or ( n57278 , n57271 , n57276 , n57277 );
and ( n57279 , n57261 , n57278 );
and ( n57280 , n57245 , n57278 );
or ( n57281 , n57262 , n57279 , n57280 );
xor ( n57282 , n56822 , n56826 );
xor ( n57283 , n57282 , n56831 );
xor ( n57284 , n56838 , n56842 );
xor ( n57285 , n57284 , n56847 );
and ( n57286 , n57283 , n57285 );
xor ( n57287 , n56855 , n56859 );
xor ( n57288 , n57287 , n56864 );
and ( n57289 , n57285 , n57288 );
and ( n57290 , n57283 , n57288 );
or ( n57291 , n57286 , n57289 , n57290 );
and ( n57292 , n57281 , n57291 );
xor ( n57293 , n56875 , n56879 );
xor ( n57294 , n57293 , n56884 );
xor ( n57295 , n56891 , n56895 );
xor ( n57296 , n57295 , n56900 );
and ( n57297 , n57294 , n57296 );
xor ( n57298 , n56908 , n56912 );
xor ( n57299 , n57298 , n56916 );
and ( n57300 , n57296 , n57299 );
and ( n57301 , n57294 , n57299 );
or ( n57302 , n57297 , n57300 , n57301 );
and ( n57303 , n57291 , n57302 );
and ( n57304 , n57281 , n57302 );
or ( n57305 , n57292 , n57303 , n57304 );
xor ( n57306 , n56725 , n56726 );
xor ( n57307 , n57306 , n56728 );
xor ( n57308 , n56732 , n56733 );
xor ( n57309 , n57308 , n56735 );
and ( n57310 , n57307 , n57309 );
xor ( n57311 , n56755 , n56771 );
xor ( n57312 , n57311 , n56781 );
and ( n57313 , n57309 , n57312 );
and ( n57314 , n57307 , n57312 );
or ( n57315 , n57310 , n57313 , n57314 );
and ( n57316 , n57305 , n57315 );
xor ( n57317 , n56799 , n56808 );
xor ( n57318 , n57317 , n56818 );
xor ( n57319 , n56834 , n56850 );
xor ( n57320 , n57319 , n56867 );
and ( n57321 , n57318 , n57320 );
xor ( n57322 , n56887 , n56903 );
xor ( n57323 , n57322 , n56919 );
and ( n57324 , n57320 , n57323 );
and ( n57325 , n57318 , n57323 );
or ( n57326 , n57321 , n57324 , n57325 );
and ( n57327 , n57315 , n57326 );
and ( n57328 , n57305 , n57326 );
or ( n57329 , n57316 , n57327 , n57328 );
and ( n57330 , n57228 , n57329 );
and ( n57331 , n57043 , n57329 );
or ( n57332 , n57229 , n57330 , n57331 );
and ( n57333 , n57040 , n57332 );
and ( n57334 , n57038 , n57332 );
or ( n57335 , n57041 , n57333 , n57334 );
and ( n57336 , n57035 , n57335 );
and ( n57337 , n57033 , n57335 );
or ( n57338 , n57036 , n57336 , n57337 );
xor ( n57339 , n57003 , n57005 );
xor ( n57340 , n57339 , n57008 );
and ( n57341 , n57338 , n57340 );
xor ( n57342 , n56712 , n56713 );
xor ( n57343 , n57342 , n56719 );
xor ( n57344 , n56731 , n56738 );
xor ( n57345 , n57344 , n56784 );
and ( n57346 , n57343 , n57345 );
xor ( n57347 , n56821 , n56870 );
xor ( n57348 , n57347 , n56922 );
and ( n57349 , n57345 , n57348 );
and ( n57350 , n57343 , n57348 );
or ( n57351 , n57346 , n57349 , n57350 );
xor ( n57352 , n56935 , n56937 );
xor ( n57353 , n57352 , n56940 );
xor ( n57354 , n56946 , n56948 );
xor ( n57355 , n57354 , n56951 );
and ( n57356 , n57353 , n57355 );
xor ( n57357 , n56960 , n56962 );
xor ( n57358 , n57357 , n56965 );
and ( n57359 , n57355 , n57358 );
and ( n57360 , n57353 , n57358 );
or ( n57361 , n57356 , n57359 , n57360 );
and ( n57362 , n57351 , n57361 );
xor ( n57363 , n56710 , n56722 );
xor ( n57364 , n57363 , n56787 );
and ( n57365 , n57361 , n57364 );
and ( n57366 , n57351 , n57364 );
or ( n57367 , n57362 , n57365 , n57366 );
xor ( n57368 , n56925 , n56943 );
xor ( n57369 , n57368 , n56954 );
xor ( n57370 , n56968 , n56970 );
xor ( n57371 , n57370 , n56973 );
and ( n57372 , n57369 , n57371 );
xor ( n57373 , n56981 , n56983 );
xor ( n57374 , n57373 , n56986 );
and ( n57375 , n57371 , n57374 );
and ( n57376 , n57369 , n57374 );
or ( n57377 , n57372 , n57375 , n57376 );
and ( n57378 , n57367 , n57377 );
xor ( n57379 , n56790 , n56957 );
xor ( n57380 , n57379 , n56976 );
and ( n57381 , n57377 , n57380 );
and ( n57382 , n57367 , n57380 );
or ( n57383 , n57378 , n57381 , n57382 );
xor ( n57384 , n56979 , n56997 );
xor ( n57385 , n57384 , n57000 );
and ( n57386 , n57383 , n57385 );
xor ( n57387 , n56989 , n56991 );
xor ( n57388 , n57387 , n56994 );
xor ( n57389 , n56927 , n56929 );
xor ( n57390 , n57389 , n56932 );
xor ( n57391 , n57067 , n57071 );
xor ( n57392 , n57391 , n57074 );
and ( n57393 , n54942 , n45886 );
and ( n57394 , n54604 , n45884 );
nor ( n57395 , n57393 , n57394 );
xnor ( n57396 , n57395 , n45824 );
xor ( n57397 , n57056 , n57060 );
xor ( n57398 , n57397 , n57064 );
or ( n57399 , n57396 , n57398 );
and ( n57400 , n57392 , n57399 );
xor ( n57401 , n57102 , n57106 );
xor ( n57402 , n57401 , n57111 );
xor ( n57403 , n57119 , n57123 );
xor ( n57404 , n57403 , n57128 );
and ( n57405 , n57402 , n57404 );
buf ( n57406 , n57405 );
and ( n57407 , n57399 , n57406 );
and ( n57408 , n57392 , n57406 );
or ( n57409 , n57400 , n57407 , n57408 );
and ( n57410 , n57390 , n57409 );
xor ( n57411 , n57138 , n57142 );
xor ( n57412 , n57411 , n57147 );
xnor ( n57413 , n57154 , n57158 );
and ( n57414 , n57412 , n57413 );
xnor ( n57415 , n57164 , n57168 );
and ( n57416 , n57413 , n57415 );
and ( n57417 , n57412 , n57415 );
or ( n57418 , n57414 , n57416 , n57417 );
xnor ( n57419 , n57177 , n57181 );
and ( n57420 , n53328 , n46306 );
and ( n57421 , n53041 , n46304 );
nor ( n57422 , n57420 , n57421 );
xnor ( n57423 , n57422 , n46228 );
and ( n57424 , n54604 , n45990 );
and ( n57425 , n54227 , n45988 );
nor ( n57426 , n57424 , n57425 );
xnor ( n57427 , n57426 , n45939 );
and ( n57428 , n57423 , n57427 );
and ( n57429 , n56388 , n45702 );
and ( n57430 , n56255 , n45700 );
nor ( n57431 , n57429 , n57430 );
xnor ( n57432 , n57431 , n20841 );
and ( n57433 , n57427 , n57432 );
and ( n57434 , n57423 , n57432 );
or ( n57435 , n57428 , n57433 , n57434 );
and ( n57436 , n57419 , n57435 );
and ( n57437 , n49976 , n48042 );
and ( n57438 , n49781 , n48040 );
nor ( n57439 , n57437 , n57438 );
xnor ( n57440 , n57439 , n47921 );
and ( n57441 , n52332 , n46712 );
and ( n57442 , n52082 , n46710 );
nor ( n57443 , n57441 , n57442 );
xnor ( n57444 , n57443 , n46587 );
and ( n57445 , n57440 , n57444 );
and ( n57446 , n57063 , n20850 );
not ( n57447 , n57446 );
and ( n57448 , n57447 , n20860 );
and ( n57449 , n57444 , n57448 );
and ( n57450 , n57440 , n57448 );
or ( n57451 , n57445 , n57449 , n57450 );
and ( n57452 , n57435 , n57451 );
and ( n57453 , n57419 , n57451 );
or ( n57454 , n57436 , n57452 , n57453 );
and ( n57455 , n57418 , n57454 );
and ( n57456 , n46969 , n51750 );
and ( n57457 , n46843 , n51748 );
nor ( n57458 , n57456 , n57457 );
xnor ( n57459 , n57458 , n51520 );
and ( n57460 , n47216 , n51221 );
and ( n57461 , n47090 , n51219 );
nor ( n57462 , n57460 , n57461 );
xnor ( n57463 , n57462 , n51000 );
or ( n57464 , n57459 , n57463 );
and ( n57465 , n49115 , n48740 );
and ( n57466 , n48988 , n48738 );
nor ( n57467 , n57465 , n57466 );
xnor ( n57468 , n57467 , n48571 );
and ( n57469 , n50404 , n47734 );
and ( n57470 , n50195 , n47732 );
nor ( n57471 , n57469 , n57470 );
xnor ( n57472 , n57471 , n47606 );
or ( n57473 , n57468 , n57472 );
and ( n57474 , n57464 , n57473 );
and ( n57475 , n55756 , n45777 );
and ( n57476 , n55497 , n45775 );
nor ( n57477 , n57475 , n57476 );
xnor ( n57478 , n57477 , n45734 );
and ( n57479 , n57063 , n20852 );
and ( n57480 , n56915 , n20850 );
nor ( n57481 , n57479 , n57480 );
xnor ( n57482 , n57481 , n20860 );
or ( n57483 , n57478 , n57482 );
and ( n57484 , n57473 , n57483 );
and ( n57485 , n57464 , n57483 );
or ( n57486 , n57474 , n57484 , n57485 );
and ( n57487 , n57454 , n57486 );
and ( n57488 , n57418 , n57486 );
or ( n57489 , n57455 , n57487 , n57488 );
and ( n57490 , n57409 , n57489 );
and ( n57491 , n57390 , n57489 );
or ( n57492 , n57410 , n57490 , n57491 );
and ( n57493 , n53922 , n46135 );
and ( n57494 , n53639 , n46133 );
nor ( n57495 , n57493 , n57494 );
xnor ( n57496 , n57495 , n46067 );
and ( n57497 , n55143 , n45886 );
and ( n57498 , n54942 , n45884 );
nor ( n57499 , n57497 , n57498 );
xnor ( n57500 , n57499 , n45824 );
or ( n57501 , n57496 , n57500 );
and ( n57502 , n46750 , n52269 );
and ( n57503 , n46577 , n52267 );
nor ( n57504 , n57502 , n57503 );
xnor ( n57505 , n57504 , n52008 );
and ( n57506 , n47474 , n50783 );
and ( n57507 , n47351 , n50781 );
nor ( n57508 , n57506 , n57507 );
xnor ( n57509 , n57508 , n50557 );
and ( n57510 , n57505 , n57509 );
and ( n57511 , n57501 , n57510 );
and ( n57512 , n49570 , n48394 );
and ( n57513 , n49374 , n48392 );
nor ( n57514 , n57512 , n57513 );
xnor ( n57515 , n57514 , n48220 );
and ( n57516 , n51298 , n47178 );
and ( n57517 , n51077 , n47176 );
nor ( n57518 , n57516 , n57517 );
xnor ( n57519 , n57518 , n47039 );
and ( n57520 , n57515 , n57519 );
and ( n57521 , n57510 , n57520 );
and ( n57522 , n57501 , n57520 );
or ( n57523 , n57511 , n57521 , n57522 );
and ( n57524 , n20844 , n57187 );
and ( n57525 , n20855 , n57184 );
nor ( n57526 , n57524 , n57525 );
xnor ( n57527 , n57526 , n56175 );
and ( n57528 , n45712 , n56503 );
and ( n57529 , n20864 , n56501 );
nor ( n57530 , n57528 , n57529 );
xnor ( n57531 , n57530 , n56178 );
and ( n57532 , n57527 , n57531 );
and ( n57533 , n45794 , n55851 );
and ( n57534 , n45763 , n55849 );
nor ( n57535 , n57533 , n57534 );
xnor ( n57536 , n57535 , n55506 );
and ( n57537 , n57531 , n57536 );
and ( n57538 , n57527 , n57536 );
or ( n57539 , n57532 , n57537 , n57538 );
and ( n57540 , n45907 , n55159 );
and ( n57541 , n45843 , n55157 );
nor ( n57542 , n57540 , n57541 );
xnor ( n57543 , n57542 , n54864 );
and ( n57544 , n46041 , n54535 );
and ( n57545 , n45963 , n54533 );
nor ( n57546 , n57544 , n57545 );
xnor ( n57547 , n57546 , n54237 );
and ( n57548 , n57543 , n57547 );
and ( n57549 , n46169 , n53928 );
and ( n57550 , n46100 , n53926 );
nor ( n57551 , n57549 , n57550 );
xnor ( n57552 , n57551 , n53652 );
and ( n57553 , n57547 , n57552 );
and ( n57554 , n57543 , n57552 );
or ( n57555 , n57548 , n57553 , n57554 );
and ( n57556 , n57539 , n57555 );
and ( n57557 , n46345 , n53357 );
and ( n57558 , n46264 , n53355 );
nor ( n57559 , n57557 , n57558 );
xnor ( n57560 , n57559 , n53060 );
and ( n57561 , n46530 , n52799 );
and ( n57562 , n46445 , n52797 );
nor ( n57563 , n57561 , n57562 );
xnor ( n57564 , n57563 , n52538 );
and ( n57565 , n57560 , n57564 );
and ( n57566 , n47778 , n50338 );
and ( n57567 , n47647 , n50336 );
nor ( n57568 , n57566 , n57567 );
xnor ( n57569 , n57568 , n50111 );
and ( n57570 , n57564 , n57569 );
and ( n57571 , n57560 , n57569 );
or ( n57572 , n57565 , n57570 , n57571 );
and ( n57573 , n57555 , n57572 );
and ( n57574 , n57539 , n57572 );
or ( n57575 , n57556 , n57573 , n57574 );
and ( n57576 , n57523 , n57575 );
and ( n57577 , n48384 , n49513 );
and ( n57578 , n48272 , n49511 );
nor ( n57579 , n57577 , n57578 );
xnor ( n57580 , n57579 , n49310 );
and ( n57581 , n48709 , n49121 );
and ( n57582 , n48632 , n49119 );
nor ( n57583 , n57581 , n57582 );
xnor ( n57584 , n57583 , n48932 );
and ( n57585 , n57580 , n57584 );
and ( n57586 , n50726 , n47429 );
and ( n57587 , n50625 , n47427 );
nor ( n57588 , n57586 , n57587 );
xnor ( n57589 , n57588 , n47309 );
and ( n57590 , n57584 , n57589 );
and ( n57591 , n57580 , n57589 );
or ( n57592 , n57585 , n57590 , n57591 );
and ( n57593 , n51734 , n46911 );
and ( n57594 , n51510 , n46909 );
nor ( n57595 , n57593 , n57594 );
xnor ( n57596 , n57595 , n46802 );
and ( n57597 , n52790 , n46496 );
and ( n57598 , n52612 , n46494 );
nor ( n57599 , n57597 , n57598 );
xnor ( n57600 , n57599 , n46402 );
and ( n57601 , n57596 , n57600 );
xor ( n57602 , n39387 , n45584 );
buf ( n57603 , n57602 );
buf ( n57604 , n57603 );
buf ( n57605 , n57604 );
and ( n57606 , n57600 , n57605 );
and ( n57607 , n57596 , n57605 );
or ( n57608 , n57601 , n57606 , n57607 );
and ( n57609 , n57592 , n57608 );
xor ( n57610 , n57190 , n57194 );
xor ( n57611 , n57610 , n57199 );
and ( n57612 , n57608 , n57611 );
and ( n57613 , n57592 , n57611 );
or ( n57614 , n57609 , n57612 , n57613 );
and ( n57615 , n57575 , n57614 );
and ( n57616 , n57523 , n57614 );
or ( n57617 , n57576 , n57615 , n57616 );
xor ( n57618 , n57207 , n57211 );
xor ( n57619 , n57618 , n57216 );
xor ( n57620 , n57233 , n57237 );
xor ( n57621 , n57620 , n57242 );
and ( n57622 , n57619 , n57621 );
xor ( n57623 , n57249 , n57253 );
xor ( n57624 , n57623 , n57258 );
and ( n57625 , n57621 , n57624 );
and ( n57626 , n57619 , n57624 );
or ( n57627 , n57622 , n57625 , n57626 );
buf ( n57628 , n57081 );
xor ( n57629 , n57628 , n57083 );
and ( n57630 , n57627 , n57629 );
xor ( n57631 , n57087 , n57088 );
xor ( n57632 , n57631 , n57090 );
and ( n57633 , n57629 , n57632 );
and ( n57634 , n57627 , n57632 );
or ( n57635 , n57630 , n57633 , n57634 );
and ( n57636 , n57617 , n57635 );
xor ( n57637 , n57098 , n57114 );
xor ( n57638 , n57637 , n57131 );
xor ( n57639 , n57150 , n57159 );
xor ( n57640 , n57639 , n57169 );
and ( n57641 , n57638 , n57640 );
xor ( n57642 , n57182 , n57202 );
xor ( n57643 , n57642 , n57219 );
and ( n57644 , n57640 , n57643 );
and ( n57645 , n57638 , n57643 );
or ( n57646 , n57641 , n57644 , n57645 );
and ( n57647 , n57635 , n57646 );
and ( n57648 , n57617 , n57646 );
or ( n57649 , n57636 , n57647 , n57648 );
and ( n57650 , n57492 , n57649 );
xor ( n57651 , n57245 , n57261 );
xor ( n57652 , n57651 , n57278 );
xor ( n57653 , n57283 , n57285 );
xor ( n57654 , n57653 , n57288 );
and ( n57655 , n57652 , n57654 );
xor ( n57656 , n57294 , n57296 );
xor ( n57657 , n57656 , n57299 );
and ( n57658 , n57654 , n57657 );
and ( n57659 , n57652 , n57657 );
or ( n57660 , n57655 , n57658 , n57659 );
xor ( n57661 , n57045 , n57047 );
xor ( n57662 , n57661 , n57049 );
and ( n57663 , n57660 , n57662 );
xor ( n57664 , n57077 , n57085 );
xor ( n57665 , n57664 , n57093 );
and ( n57666 , n57662 , n57665 );
and ( n57667 , n57660 , n57665 );
or ( n57668 , n57663 , n57666 , n57667 );
and ( n57669 , n57649 , n57668 );
and ( n57670 , n57492 , n57668 );
or ( n57671 , n57650 , n57669 , n57670 );
xor ( n57672 , n57134 , n57172 );
xor ( n57673 , n57672 , n57222 );
xor ( n57674 , n57281 , n57291 );
xor ( n57675 , n57674 , n57302 );
and ( n57676 , n57673 , n57675 );
xor ( n57677 , n57307 , n57309 );
xor ( n57678 , n57677 , n57312 );
and ( n57679 , n57675 , n57678 );
and ( n57680 , n57673 , n57678 );
or ( n57681 , n57676 , n57679 , n57680 );
xor ( n57682 , n57052 , n57096 );
xor ( n57683 , n57682 , n57225 );
and ( n57684 , n57681 , n57683 );
xor ( n57685 , n57305 , n57315 );
xor ( n57686 , n57685 , n57326 );
and ( n57687 , n57683 , n57686 );
and ( n57688 , n57681 , n57686 );
or ( n57689 , n57684 , n57687 , n57688 );
and ( n57690 , n57671 , n57689 );
xor ( n57691 , n57043 , n57228 );
xor ( n57692 , n57691 , n57329 );
and ( n57693 , n57689 , n57692 );
and ( n57694 , n57671 , n57692 );
or ( n57695 , n57690 , n57693 , n57694 );
and ( n57696 , n57388 , n57695 );
xor ( n57697 , n57038 , n57040 );
xor ( n57698 , n57697 , n57332 );
and ( n57699 , n57695 , n57698 );
and ( n57700 , n57388 , n57698 );
or ( n57701 , n57696 , n57699 , n57700 );
and ( n57702 , n57385 , n57701 );
and ( n57703 , n57383 , n57701 );
or ( n57704 , n57386 , n57702 , n57703 );
and ( n57705 , n57340 , n57704 );
and ( n57706 , n57338 , n57704 );
or ( n57707 , n57341 , n57705 , n57706 );
and ( n57708 , n57031 , n57707 );
xor ( n57709 , n57033 , n57035 );
xor ( n57710 , n57709 , n57335 );
xor ( n57711 , n57367 , n57377 );
xor ( n57712 , n57711 , n57380 );
xor ( n57713 , n57351 , n57361 );
xor ( n57714 , n57713 , n57364 );
xor ( n57715 , n57369 , n57371 );
xor ( n57716 , n57715 , n57374 );
and ( n57717 , n57714 , n57716 );
xor ( n57718 , n57343 , n57345 );
xor ( n57719 , n57718 , n57348 );
xor ( n57720 , n57353 , n57355 );
xor ( n57721 , n57720 , n57358 );
and ( n57722 , n57719 , n57721 );
xor ( n57723 , n57318 , n57320 );
xor ( n57724 , n57723 , n57323 );
xor ( n57725 , n57266 , n57270 );
xor ( n57726 , n57725 , n57275 );
xnor ( n57727 , n57396 , n57398 );
and ( n57728 , n57726 , n57727 );
and ( n57729 , n47090 , n51750 );
and ( n57730 , n46969 , n51748 );
nor ( n57731 , n57729 , n57730 );
xnor ( n57732 , n57731 , n51520 );
and ( n57733 , n47351 , n51221 );
and ( n57734 , n47216 , n51219 );
nor ( n57735 , n57733 , n57734 );
xnor ( n57736 , n57735 , n51000 );
and ( n57737 , n57732 , n57736 );
and ( n57738 , n47647 , n50783 );
and ( n57739 , n47474 , n50781 );
nor ( n57740 , n57738 , n57739 );
xnor ( n57741 , n57740 , n50557 );
and ( n57742 , n57736 , n57741 );
and ( n57743 , n57732 , n57741 );
or ( n57744 , n57737 , n57742 , n57743 );
and ( n57745 , n48108 , n49896 );
and ( n57746 , n47962 , n49894 );
nor ( n57747 , n57745 , n57746 );
xnor ( n57748 , n57747 , n49711 );
or ( n57749 , n57744 , n57748 );
and ( n57750 , n57727 , n57749 );
and ( n57751 , n57726 , n57749 );
or ( n57752 , n57728 , n57750 , n57751 );
xor ( n57753 , n57423 , n57427 );
xor ( n57754 , n57753 , n57432 );
xor ( n57755 , n57440 , n57444 );
xor ( n57756 , n57755 , n57448 );
and ( n57757 , n57754 , n57756 );
buf ( n57758 , n57757 );
xnor ( n57759 , n57459 , n57463 );
xnor ( n57760 , n57468 , n57472 );
and ( n57761 , n57759 , n57760 );
xnor ( n57762 , n57478 , n57482 );
and ( n57763 , n57760 , n57762 );
and ( n57764 , n57759 , n57762 );
or ( n57765 , n57761 , n57763 , n57764 );
and ( n57766 , n57758 , n57765 );
xnor ( n57767 , n57496 , n57500 );
xor ( n57768 , n57505 , n57509 );
and ( n57769 , n57767 , n57768 );
xor ( n57770 , n57515 , n57519 );
and ( n57771 , n57768 , n57770 );
and ( n57772 , n57767 , n57770 );
or ( n57773 , n57769 , n57771 , n57772 );
and ( n57774 , n57765 , n57773 );
and ( n57775 , n57758 , n57773 );
or ( n57776 , n57766 , n57774 , n57775 );
and ( n57777 , n57752 , n57776 );
and ( n57778 , n50195 , n48042 );
and ( n57779 , n49976 , n48040 );
nor ( n57780 , n57778 , n57779 );
xnor ( n57781 , n57780 , n47921 );
and ( n57782 , n51510 , n47178 );
and ( n57783 , n51298 , n47176 );
nor ( n57784 , n57782 , n57783 );
xnor ( n57785 , n57784 , n47039 );
and ( n57786 , n57781 , n57785 );
and ( n57787 , n52082 , n46911 );
and ( n57788 , n51734 , n46909 );
nor ( n57789 , n57787 , n57788 );
xnor ( n57790 , n57789 , n46802 );
and ( n57791 , n57785 , n57790 );
and ( n57792 , n57781 , n57790 );
or ( n57793 , n57786 , n57791 , n57792 );
and ( n57794 , n54942 , n45990 );
and ( n57795 , n54604 , n45988 );
nor ( n57796 , n57794 , n57795 );
xnor ( n57797 , n57796 , n45939 );
and ( n57798 , n55497 , n45886 );
and ( n57799 , n55143 , n45884 );
nor ( n57800 , n57798 , n57799 );
xnor ( n57801 , n57800 , n45824 );
and ( n57802 , n57797 , n57801 );
and ( n57803 , n56915 , n45702 );
and ( n57804 , n56388 , n45700 );
nor ( n57805 , n57803 , n57804 );
xnor ( n57806 , n57805 , n20841 );
and ( n57807 , n57801 , n57806 );
and ( n57808 , n57797 , n57806 );
or ( n57809 , n57802 , n57807 , n57808 );
and ( n57810 , n57793 , n57809 );
and ( n57811 , n46264 , n53928 );
and ( n57812 , n46169 , n53926 );
nor ( n57813 , n57811 , n57812 );
xnor ( n57814 , n57813 , n53652 );
and ( n57815 , n48272 , n49896 );
and ( n57816 , n48108 , n49894 );
nor ( n57817 , n57815 , n57816 );
xnor ( n57818 , n57817 , n49711 );
or ( n57819 , n57814 , n57818 );
and ( n57820 , n57809 , n57819 );
and ( n57821 , n57793 , n57819 );
or ( n57822 , n57810 , n57820 , n57821 );
and ( n57823 , n49374 , n48740 );
and ( n57824 , n49115 , n48738 );
nor ( n57825 , n57823 , n57824 );
xnor ( n57826 , n57825 , n48571 );
and ( n57827 , n51077 , n47429 );
and ( n57828 , n50726 , n47427 );
nor ( n57829 , n57827 , n57828 );
xnor ( n57830 , n57829 , n47309 );
or ( n57831 , n57826 , n57830 );
and ( n57832 , n49781 , n48394 );
and ( n57833 , n49570 , n48392 );
nor ( n57834 , n57832 , n57833 );
xnor ( n57835 , n57834 , n48220 );
and ( n57836 , n52612 , n46712 );
and ( n57837 , n52332 , n46710 );
nor ( n57838 , n57836 , n57837 );
xnor ( n57839 , n57838 , n46587 );
or ( n57840 , n57835 , n57839 );
and ( n57841 , n57831 , n57840 );
and ( n57842 , n53639 , n46306 );
and ( n57843 , n53328 , n46304 );
nor ( n57844 , n57842 , n57843 );
xnor ( n57845 , n57844 , n46228 );
and ( n57846 , n54227 , n46135 );
and ( n57847 , n53922 , n46133 );
nor ( n57848 , n57846 , n57847 );
xnor ( n57849 , n57848 , n46067 );
or ( n57850 , n57845 , n57849 );
and ( n57851 , n57840 , n57850 );
and ( n57852 , n57831 , n57850 );
or ( n57853 , n57841 , n57851 , n57852 );
and ( n57854 , n57822 , n57853 );
and ( n57855 , n20864 , n57187 );
and ( n57856 , n20844 , n57184 );
nor ( n57857 , n57855 , n57856 );
xnor ( n57858 , n57857 , n56175 );
and ( n57859 , n45763 , n56503 );
and ( n57860 , n45712 , n56501 );
nor ( n57861 , n57859 , n57860 );
xnor ( n57862 , n57861 , n56178 );
and ( n57863 , n57858 , n57862 );
and ( n57864 , n45843 , n55851 );
and ( n57865 , n45794 , n55849 );
nor ( n57866 , n57864 , n57865 );
xnor ( n57867 , n57866 , n55506 );
and ( n57868 , n57862 , n57867 );
and ( n57869 , n57858 , n57867 );
or ( n57870 , n57863 , n57868 , n57869 );
and ( n57871 , n45963 , n55159 );
and ( n57872 , n45907 , n55157 );
nor ( n57873 , n57871 , n57872 );
xnor ( n57874 , n57873 , n54864 );
and ( n57875 , n46100 , n54535 );
and ( n57876 , n46041 , n54533 );
nor ( n57877 , n57875 , n57876 );
xnor ( n57878 , n57877 , n54237 );
and ( n57879 , n57874 , n57878 );
and ( n57880 , n46445 , n53357 );
and ( n57881 , n46345 , n53355 );
nor ( n57882 , n57880 , n57881 );
xnor ( n57883 , n57882 , n53060 );
and ( n57884 , n57878 , n57883 );
and ( n57885 , n57874 , n57883 );
or ( n57886 , n57879 , n57884 , n57885 );
and ( n57887 , n57870 , n57886 );
and ( n57888 , n46577 , n52799 );
and ( n57889 , n46530 , n52797 );
nor ( n57890 , n57888 , n57889 );
xnor ( n57891 , n57890 , n52538 );
and ( n57892 , n46843 , n52269 );
and ( n57893 , n46750 , n52267 );
nor ( n57894 , n57892 , n57893 );
xnor ( n57895 , n57894 , n52008 );
and ( n57896 , n57891 , n57895 );
and ( n57897 , n47962 , n50338 );
and ( n57898 , n47778 , n50336 );
nor ( n57899 , n57897 , n57898 );
xnor ( n57900 , n57899 , n50111 );
and ( n57901 , n57895 , n57900 );
and ( n57902 , n57891 , n57900 );
or ( n57903 , n57896 , n57901 , n57902 );
and ( n57904 , n57886 , n57903 );
and ( n57905 , n57870 , n57903 );
or ( n57906 , n57887 , n57904 , n57905 );
and ( n57907 , n57853 , n57906 );
and ( n57908 , n57822 , n57906 );
or ( n57909 , n57854 , n57907 , n57908 );
and ( n57910 , n57776 , n57909 );
and ( n57911 , n57752 , n57909 );
or ( n57912 , n57777 , n57910 , n57911 );
and ( n57913 , n57724 , n57912 );
and ( n57914 , n48632 , n49513 );
and ( n57915 , n48384 , n49511 );
nor ( n57916 , n57914 , n57915 );
xnor ( n57917 , n57916 , n49310 );
and ( n57918 , n48988 , n49121 );
and ( n57919 , n48709 , n49119 );
nor ( n57920 , n57918 , n57919 );
xnor ( n57921 , n57920 , n48932 );
and ( n57922 , n57917 , n57921 );
and ( n57923 , n50625 , n47734 );
and ( n57924 , n50404 , n47732 );
nor ( n57925 , n57923 , n57924 );
xnor ( n57926 , n57925 , n47606 );
and ( n57927 , n57921 , n57926 );
and ( n57928 , n57917 , n57926 );
or ( n57929 , n57922 , n57927 , n57928 );
and ( n57930 , n53041 , n46496 );
and ( n57931 , n52790 , n46494 );
nor ( n57932 , n57930 , n57931 );
xnor ( n57933 , n57932 , n46402 );
and ( n57934 , n56255 , n45777 );
and ( n57935 , n55756 , n45775 );
nor ( n57936 , n57934 , n57935 );
xnor ( n57937 , n57936 , n45734 );
and ( n57938 , n57933 , n57937 );
and ( n57939 , n57937 , n57446 );
and ( n57940 , n57933 , n57446 );
or ( n57941 , n57938 , n57939 , n57940 );
and ( n57942 , n57929 , n57941 );
xor ( n57943 , n39390 , n45582 );
buf ( n57944 , n57943 );
buf ( n57945 , n57944 );
buf ( n57946 , n57945 );
buf ( n57947 , n20184 );
buf ( n57948 , n57947 );
buf ( n57949 , n57948 );
not ( n57950 , n57949 );
and ( n57951 , n57946 , n57950 );
buf ( n57952 , n57951 );
and ( n57953 , n57941 , n57952 );
and ( n57954 , n57929 , n57952 );
or ( n57955 , n57942 , n57953 , n57954 );
xor ( n57956 , n57527 , n57531 );
xor ( n57957 , n57956 , n57536 );
xor ( n57958 , n57543 , n57547 );
xor ( n57959 , n57958 , n57552 );
and ( n57960 , n57957 , n57959 );
xor ( n57961 , n57560 , n57564 );
xor ( n57962 , n57961 , n57569 );
and ( n57963 , n57959 , n57962 );
and ( n57964 , n57957 , n57962 );
or ( n57965 , n57960 , n57963 , n57964 );
and ( n57966 , n57955 , n57965 );
buf ( n57967 , n57402 );
xor ( n57968 , n57967 , n57404 );
and ( n57969 , n57965 , n57968 );
and ( n57970 , n57955 , n57968 );
or ( n57971 , n57966 , n57969 , n57970 );
xor ( n57972 , n57412 , n57413 );
xor ( n57973 , n57972 , n57415 );
xor ( n57974 , n57419 , n57435 );
xor ( n57975 , n57974 , n57451 );
and ( n57976 , n57973 , n57975 );
xor ( n57977 , n57464 , n57473 );
xor ( n57978 , n57977 , n57483 );
and ( n57979 , n57975 , n57978 );
and ( n57980 , n57973 , n57978 );
or ( n57981 , n57976 , n57979 , n57980 );
and ( n57982 , n57971 , n57981 );
xor ( n57983 , n57501 , n57510 );
xor ( n57984 , n57983 , n57520 );
xor ( n57985 , n57539 , n57555 );
xor ( n57986 , n57985 , n57572 );
and ( n57987 , n57984 , n57986 );
xor ( n57988 , n57592 , n57608 );
xor ( n57989 , n57988 , n57611 );
and ( n57990 , n57986 , n57989 );
and ( n57991 , n57984 , n57989 );
or ( n57992 , n57987 , n57990 , n57991 );
and ( n57993 , n57981 , n57992 );
and ( n57994 , n57971 , n57992 );
or ( n57995 , n57982 , n57993 , n57994 );
and ( n57996 , n57912 , n57995 );
and ( n57997 , n57724 , n57995 );
or ( n57998 , n57913 , n57996 , n57997 );
and ( n57999 , n57721 , n57998 );
and ( n58000 , n57719 , n57998 );
or ( n58001 , n57722 , n57999 , n58000 );
and ( n58002 , n57716 , n58001 );
and ( n58003 , n57714 , n58001 );
or ( n58004 , n57717 , n58002 , n58003 );
and ( n58005 , n57712 , n58004 );
xor ( n58006 , n57388 , n57695 );
xor ( n58007 , n58006 , n57698 );
and ( n58008 , n58004 , n58007 );
and ( n58009 , n57712 , n58007 );
or ( n58010 , n58005 , n58008 , n58009 );
and ( n58011 , n57710 , n58010 );
xor ( n58012 , n57383 , n57385 );
xor ( n58013 , n58012 , n57701 );
and ( n58014 , n58010 , n58013 );
and ( n58015 , n57710 , n58013 );
or ( n58016 , n58011 , n58014 , n58015 );
xor ( n58017 , n57338 , n57340 );
xor ( n58018 , n58017 , n57704 );
or ( n58019 , n58016 , n58018 );
and ( n58020 , n57707 , n58019 );
and ( n58021 , n57031 , n58019 );
or ( n58022 , n57708 , n58020 , n58021 );
and ( n58023 , n57029 , n58022 );
xor ( n58024 , n57029 , n58022 );
xor ( n58025 , n57031 , n57707 );
xor ( n58026 , n58025 , n58019 );
not ( n58027 , n58026 );
xnor ( n58028 , n58016 , n58018 );
xor ( n58029 , n57710 , n58010 );
xor ( n58030 , n58029 , n58013 );
xor ( n58031 , n57392 , n57399 );
xor ( n58032 , n58031 , n57406 );
xor ( n58033 , n57418 , n57454 );
xor ( n58034 , n58033 , n57486 );
and ( n58035 , n58032 , n58034 );
xor ( n58036 , n57523 , n57575 );
xor ( n58037 , n58036 , n57614 );
and ( n58038 , n58034 , n58037 );
and ( n58039 , n58032 , n58037 );
or ( n58040 , n58035 , n58038 , n58039 );
xor ( n58041 , n57627 , n57629 );
xor ( n58042 , n58041 , n57632 );
xor ( n58043 , n57638 , n57640 );
xor ( n58044 , n58043 , n57643 );
and ( n58045 , n58042 , n58044 );
xor ( n58046 , n57652 , n57654 );
xor ( n58047 , n58046 , n57657 );
and ( n58048 , n58044 , n58047 );
and ( n58049 , n58042 , n58047 );
or ( n58050 , n58045 , n58048 , n58049 );
and ( n58051 , n58040 , n58050 );
xor ( n58052 , n57390 , n57409 );
xor ( n58053 , n58052 , n57489 );
and ( n58054 , n58050 , n58053 );
and ( n58055 , n58040 , n58053 );
or ( n58056 , n58051 , n58054 , n58055 );
xor ( n58057 , n57617 , n57635 );
xor ( n58058 , n58057 , n57646 );
xor ( n58059 , n57660 , n57662 );
xor ( n58060 , n58059 , n57665 );
and ( n58061 , n58058 , n58060 );
xor ( n58062 , n57673 , n57675 );
xor ( n58063 , n58062 , n57678 );
and ( n58064 , n58060 , n58063 );
and ( n58065 , n58058 , n58063 );
or ( n58066 , n58061 , n58064 , n58065 );
and ( n58067 , n58056 , n58066 );
xor ( n58068 , n57492 , n57649 );
xor ( n58069 , n58068 , n57668 );
and ( n58070 , n58066 , n58069 );
and ( n58071 , n58056 , n58069 );
or ( n58072 , n58067 , n58070 , n58071 );
xor ( n58073 , n57671 , n57689 );
xor ( n58074 , n58073 , n57692 );
and ( n58075 , n58072 , n58074 );
xor ( n58076 , n57681 , n57683 );
xor ( n58077 , n58076 , n57686 );
xor ( n58078 , n57619 , n57621 );
xor ( n58079 , n58078 , n57624 );
xor ( n58080 , n57580 , n57584 );
xor ( n58081 , n58080 , n57589 );
xor ( n58082 , n57596 , n57600 );
xor ( n58083 , n58082 , n57605 );
and ( n58084 , n58081 , n58083 );
xnor ( n58085 , n57744 , n57748 );
and ( n58086 , n58083 , n58085 );
and ( n58087 , n58081 , n58085 );
or ( n58088 , n58084 , n58086 , n58087 );
and ( n58089 , n58079 , n58088 );
and ( n58090 , n49976 , n48394 );
and ( n58091 , n49781 , n48392 );
nor ( n58092 , n58090 , n58091 );
xnor ( n58093 , n58092 , n48220 );
and ( n58094 , n50404 , n48042 );
and ( n58095 , n50195 , n48040 );
nor ( n58096 , n58094 , n58095 );
xnor ( n58097 , n58096 , n47921 );
and ( n58098 , n58093 , n58097 );
and ( n58099 , n52790 , n46712 );
and ( n58100 , n52612 , n46710 );
nor ( n58101 , n58099 , n58100 );
xnor ( n58102 , n58101 , n46587 );
and ( n58103 , n58097 , n58102 );
and ( n58104 , n58093 , n58102 );
or ( n58105 , n58098 , n58103 , n58104 );
xor ( n58106 , n57781 , n57785 );
xor ( n58107 , n58106 , n57790 );
or ( n58108 , n58105 , n58107 );
xor ( n58109 , n57732 , n57736 );
xor ( n58110 , n58109 , n57741 );
xor ( n58111 , n57797 , n57801 );
xor ( n58112 , n58111 , n57806 );
and ( n58113 , n58110 , n58112 );
xnor ( n58114 , n57814 , n57818 );
and ( n58115 , n58112 , n58114 );
and ( n58116 , n58110 , n58114 );
or ( n58117 , n58113 , n58115 , n58116 );
and ( n58118 , n58108 , n58117 );
xnor ( n58119 , n57826 , n57830 );
xnor ( n58120 , n57835 , n57839 );
and ( n58121 , n58119 , n58120 );
xnor ( n58122 , n57845 , n57849 );
and ( n58123 , n58120 , n58122 );
and ( n58124 , n58119 , n58122 );
or ( n58125 , n58121 , n58123 , n58124 );
and ( n58126 , n58117 , n58125 );
and ( n58127 , n58108 , n58125 );
or ( n58128 , n58118 , n58126 , n58127 );
and ( n58129 , n58088 , n58128 );
and ( n58130 , n58079 , n58128 );
or ( n58131 , n58089 , n58129 , n58130 );
and ( n58132 , n55756 , n45886 );
and ( n58133 , n55497 , n45884 );
nor ( n58134 , n58132 , n58133 );
xnor ( n58135 , n58134 , n45824 );
and ( n58136 , n56388 , n45777 );
and ( n58137 , n56255 , n45775 );
nor ( n58138 , n58136 , n58137 );
xnor ( n58139 , n58138 , n45734 );
or ( n58140 , n58135 , n58139 );
and ( n58141 , n52332 , n46911 );
and ( n58142 , n52082 , n46909 );
nor ( n58143 , n58141 , n58142 );
xnor ( n58144 , n58143 , n46802 );
and ( n58145 , n57063 , n45700 );
not ( n58146 , n58145 );
and ( n58147 , n58146 , n20841 );
or ( n58148 , n58144 , n58147 );
and ( n58149 , n58140 , n58148 );
and ( n58150 , n46969 , n52269 );
and ( n58151 , n46843 , n52267 );
nor ( n58152 , n58150 , n58151 );
xnor ( n58153 , n58152 , n52008 );
and ( n58154 , n47778 , n50783 );
and ( n58155 , n47647 , n50781 );
nor ( n58156 , n58154 , n58155 );
xnor ( n58157 , n58156 , n50557 );
or ( n58158 , n58153 , n58157 );
and ( n58159 , n58148 , n58158 );
and ( n58160 , n58140 , n58158 );
or ( n58161 , n58149 , n58159 , n58160 );
and ( n58162 , n54604 , n46135 );
and ( n58163 , n54227 , n46133 );
nor ( n58164 , n58162 , n58163 );
xnor ( n58165 , n58164 , n46067 );
and ( n58166 , n57063 , n45702 );
and ( n58167 , n56915 , n45700 );
nor ( n58168 , n58166 , n58167 );
xnor ( n58169 , n58168 , n20841 );
or ( n58170 , n58165 , n58169 );
and ( n58171 , n49570 , n48740 );
and ( n58172 , n49374 , n48738 );
nor ( n58173 , n58171 , n58172 );
xnor ( n58174 , n58173 , n48571 );
and ( n58175 , n50726 , n47734 );
and ( n58176 , n50625 , n47732 );
nor ( n58177 , n58175 , n58176 );
xnor ( n58178 , n58177 , n47606 );
and ( n58179 , n58174 , n58178 );
and ( n58180 , n58170 , n58179 );
and ( n58181 , n51298 , n47429 );
and ( n58182 , n51077 , n47427 );
nor ( n58183 , n58181 , n58182 );
xnor ( n58184 , n58183 , n47309 );
and ( n58185 , n51734 , n47178 );
and ( n58186 , n51510 , n47176 );
nor ( n58187 , n58185 , n58186 );
xnor ( n58188 , n58187 , n47039 );
and ( n58189 , n58184 , n58188 );
and ( n58190 , n58179 , n58189 );
and ( n58191 , n58170 , n58189 );
or ( n58192 , n58180 , n58190 , n58191 );
and ( n58193 , n58161 , n58192 );
and ( n58194 , n45712 , n57187 );
and ( n58195 , n20864 , n57184 );
nor ( n58196 , n58194 , n58195 );
xnor ( n58197 , n58196 , n56175 );
and ( n58198 , n45794 , n56503 );
and ( n58199 , n45763 , n56501 );
nor ( n58200 , n58198 , n58199 );
xnor ( n58201 , n58200 , n56178 );
and ( n58202 , n58197 , n58201 );
and ( n58203 , n45907 , n55851 );
and ( n58204 , n45843 , n55849 );
nor ( n58205 , n58203 , n58204 );
xnor ( n58206 , n58205 , n55506 );
and ( n58207 , n58201 , n58206 );
and ( n58208 , n58197 , n58206 );
or ( n58209 , n58202 , n58207 , n58208 );
and ( n58210 , n46041 , n55159 );
and ( n58211 , n45963 , n55157 );
nor ( n58212 , n58210 , n58211 );
xnor ( n58213 , n58212 , n54864 );
and ( n58214 , n46169 , n54535 );
and ( n58215 , n46100 , n54533 );
nor ( n58216 , n58214 , n58215 );
xnor ( n58217 , n58216 , n54237 );
and ( n58218 , n58213 , n58217 );
and ( n58219 , n46530 , n53357 );
and ( n58220 , n46445 , n53355 );
nor ( n58221 , n58219 , n58220 );
xnor ( n58222 , n58221 , n53060 );
and ( n58223 , n58217 , n58222 );
and ( n58224 , n58213 , n58222 );
or ( n58225 , n58218 , n58223 , n58224 );
and ( n58226 , n58209 , n58225 );
and ( n58227 , n46750 , n52799 );
and ( n58228 , n46577 , n52797 );
nor ( n58229 , n58227 , n58228 );
xnor ( n58230 , n58229 , n52538 );
and ( n58231 , n47216 , n51750 );
and ( n58232 , n47090 , n51748 );
nor ( n58233 , n58231 , n58232 );
xnor ( n58234 , n58233 , n51520 );
and ( n58235 , n58230 , n58234 );
and ( n58236 , n47474 , n51221 );
and ( n58237 , n47351 , n51219 );
nor ( n58238 , n58236 , n58237 );
xnor ( n58239 , n58238 , n51000 );
and ( n58240 , n58234 , n58239 );
and ( n58241 , n58230 , n58239 );
or ( n58242 , n58235 , n58240 , n58241 );
and ( n58243 , n58225 , n58242 );
and ( n58244 , n58209 , n58242 );
or ( n58245 , n58226 , n58243 , n58244 );
and ( n58246 , n58192 , n58245 );
and ( n58247 , n58161 , n58245 );
or ( n58248 , n58193 , n58246 , n58247 );
and ( n58249 , n48108 , n50338 );
and ( n58250 , n47962 , n50336 );
nor ( n58251 , n58249 , n58250 );
xnor ( n58252 , n58251 , n50111 );
and ( n58253 , n48384 , n49896 );
and ( n58254 , n48272 , n49894 );
nor ( n58255 , n58253 , n58254 );
xnor ( n58256 , n58255 , n49711 );
and ( n58257 , n58252 , n58256 );
and ( n58258 , n48709 , n49513 );
and ( n58259 , n48632 , n49511 );
nor ( n58260 , n58258 , n58259 );
xnor ( n58261 , n58260 , n49310 );
and ( n58262 , n58256 , n58261 );
and ( n58263 , n58252 , n58261 );
or ( n58264 , n58257 , n58262 , n58263 );
and ( n58265 , n49115 , n49121 );
and ( n58266 , n48988 , n49119 );
nor ( n58267 , n58265 , n58266 );
xnor ( n58268 , n58267 , n48932 );
and ( n58269 , n53328 , n46496 );
and ( n58270 , n53041 , n46494 );
nor ( n58271 , n58269 , n58270 );
xnor ( n58272 , n58271 , n46402 );
and ( n58273 , n58268 , n58272 );
and ( n58274 , n53922 , n46306 );
and ( n58275 , n53639 , n46304 );
nor ( n58276 , n58274 , n58275 );
xnor ( n58277 , n58276 , n46228 );
and ( n58278 , n58272 , n58277 );
and ( n58279 , n58268 , n58277 );
or ( n58280 , n58273 , n58278 , n58279 );
and ( n58281 , n58264 , n58280 );
and ( n58282 , n55143 , n45990 );
and ( n58283 , n54942 , n45988 );
nor ( n58284 , n58282 , n58283 );
xnor ( n58285 , n58284 , n45939 );
xor ( n58286 , n39391 , n45581 );
buf ( n58287 , n58286 );
buf ( n58288 , n58287 );
buf ( n58289 , n58288 );
and ( n58290 , n58285 , n58289 );
buf ( n58291 , n20187 );
buf ( n58292 , n58291 );
buf ( n58293 , n20184 );
buf ( n58294 , n58293 );
and ( n58295 , n58292 , n58294 );
not ( n58296 , n58295 );
and ( n58297 , n58289 , n58296 );
and ( n58298 , n58285 , n58296 );
or ( n58299 , n58290 , n58297 , n58298 );
and ( n58300 , n58280 , n58299 );
and ( n58301 , n58264 , n58299 );
or ( n58302 , n58281 , n58300 , n58301 );
xor ( n58303 , n57858 , n57862 );
xor ( n58304 , n58303 , n57867 );
xor ( n58305 , n57874 , n57878 );
xor ( n58306 , n58305 , n57883 );
and ( n58307 , n58304 , n58306 );
xor ( n58308 , n57891 , n57895 );
xor ( n58309 , n58308 , n57900 );
and ( n58310 , n58306 , n58309 );
and ( n58311 , n58304 , n58309 );
or ( n58312 , n58307 , n58310 , n58311 );
and ( n58313 , n58302 , n58312 );
xor ( n58314 , n57917 , n57921 );
xor ( n58315 , n58314 , n57926 );
xor ( n58316 , n57933 , n57937 );
xor ( n58317 , n58316 , n57446 );
and ( n58318 , n58315 , n58317 );
xor ( n58319 , n57946 , n57950 );
buf ( n58320 , n58319 );
and ( n58321 , n58317 , n58320 );
and ( n58322 , n58315 , n58320 );
or ( n58323 , n58318 , n58321 , n58322 );
and ( n58324 , n58312 , n58323 );
and ( n58325 , n58302 , n58323 );
or ( n58326 , n58313 , n58324 , n58325 );
and ( n58327 , n58248 , n58326 );
buf ( n58328 , n57754 );
xor ( n58329 , n58328 , n57756 );
xor ( n58330 , n57759 , n57760 );
xor ( n58331 , n58330 , n57762 );
and ( n58332 , n58329 , n58331 );
xor ( n58333 , n57767 , n57768 );
xor ( n58334 , n58333 , n57770 );
and ( n58335 , n58331 , n58334 );
and ( n58336 , n58329 , n58334 );
or ( n58337 , n58332 , n58335 , n58336 );
and ( n58338 , n58326 , n58337 );
and ( n58339 , n58248 , n58337 );
or ( n58340 , n58327 , n58338 , n58339 );
and ( n58341 , n58131 , n58340 );
xor ( n58342 , n57793 , n57809 );
xor ( n58343 , n58342 , n57819 );
xor ( n58344 , n57831 , n57840 );
xor ( n58345 , n58344 , n57850 );
and ( n58346 , n58343 , n58345 );
xor ( n58347 , n57870 , n57886 );
xor ( n58348 , n58347 , n57903 );
and ( n58349 , n58345 , n58348 );
and ( n58350 , n58343 , n58348 );
or ( n58351 , n58346 , n58349 , n58350 );
xor ( n58352 , n57726 , n57727 );
xor ( n58353 , n58352 , n57749 );
and ( n58354 , n58351 , n58353 );
xor ( n58355 , n57758 , n57765 );
xor ( n58356 , n58355 , n57773 );
and ( n58357 , n58353 , n58356 );
and ( n58358 , n58351 , n58356 );
or ( n58359 , n58354 , n58357 , n58358 );
and ( n58360 , n58340 , n58359 );
and ( n58361 , n58131 , n58359 );
or ( n58362 , n58341 , n58360 , n58361 );
xor ( n58363 , n57822 , n57853 );
xor ( n58364 , n58363 , n57906 );
xor ( n58365 , n57955 , n57965 );
xor ( n58366 , n58365 , n57968 );
and ( n58367 , n58364 , n58366 );
xor ( n58368 , n57973 , n57975 );
xor ( n58369 , n58368 , n57978 );
and ( n58370 , n58366 , n58369 );
and ( n58371 , n58364 , n58369 );
or ( n58372 , n58367 , n58370 , n58371 );
xor ( n58373 , n57752 , n57776 );
xor ( n58374 , n58373 , n57909 );
and ( n58375 , n58372 , n58374 );
xor ( n58376 , n57971 , n57981 );
xor ( n58377 , n58376 , n57992 );
and ( n58378 , n58374 , n58377 );
and ( n58379 , n58372 , n58377 );
or ( n58380 , n58375 , n58378 , n58379 );
and ( n58381 , n58362 , n58380 );
xor ( n58382 , n57724 , n57912 );
xor ( n58383 , n58382 , n57995 );
and ( n58384 , n58380 , n58383 );
and ( n58385 , n58362 , n58383 );
or ( n58386 , n58381 , n58384 , n58385 );
and ( n58387 , n58077 , n58386 );
xor ( n58388 , n57719 , n57721 );
xor ( n58389 , n58388 , n57998 );
and ( n58390 , n58386 , n58389 );
and ( n58391 , n58077 , n58389 );
or ( n58392 , n58387 , n58390 , n58391 );
and ( n58393 , n58074 , n58392 );
and ( n58394 , n58072 , n58392 );
or ( n58395 , n58075 , n58393 , n58394 );
xor ( n58396 , n57712 , n58004 );
xor ( n58397 , n58396 , n58007 );
and ( n58398 , n58395 , n58397 );
xor ( n58399 , n57714 , n57716 );
xor ( n58400 , n58399 , n58001 );
xor ( n58401 , n58056 , n58066 );
xor ( n58402 , n58401 , n58069 );
xor ( n58403 , n58040 , n58050 );
xor ( n58404 , n58403 , n58053 );
xor ( n58405 , n58058 , n58060 );
xor ( n58406 , n58405 , n58063 );
and ( n58407 , n58404 , n58406 );
xor ( n58408 , n58032 , n58034 );
xor ( n58409 , n58408 , n58037 );
xor ( n58410 , n58042 , n58044 );
xor ( n58411 , n58410 , n58047 );
and ( n58412 , n58409 , n58411 );
xor ( n58413 , n57984 , n57986 );
xor ( n58414 , n58413 , n57989 );
xor ( n58415 , n57929 , n57941 );
xor ( n58416 , n58415 , n57952 );
xor ( n58417 , n57957 , n57959 );
xor ( n58418 , n58417 , n57962 );
and ( n58419 , n58416 , n58418 );
xnor ( n58420 , n58105 , n58107 );
and ( n58421 , n47351 , n51750 );
and ( n58422 , n47216 , n51748 );
nor ( n58423 , n58421 , n58422 );
xnor ( n58424 , n58423 , n51520 );
and ( n58425 , n47647 , n51221 );
and ( n58426 , n47474 , n51219 );
nor ( n58427 , n58425 , n58426 );
xnor ( n58428 , n58427 , n51000 );
and ( n58429 , n58424 , n58428 );
and ( n58430 , n47962 , n50783 );
and ( n58431 , n47778 , n50781 );
nor ( n58432 , n58430 , n58431 );
xnor ( n58433 , n58432 , n50557 );
and ( n58434 , n58428 , n58433 );
and ( n58435 , n58424 , n58433 );
or ( n58436 , n58429 , n58434 , n58435 );
and ( n58437 , n46345 , n53928 );
and ( n58438 , n46264 , n53926 );
nor ( n58439 , n58437 , n58438 );
xnor ( n58440 , n58439 , n53652 );
or ( n58441 , n58436 , n58440 );
and ( n58442 , n58420 , n58441 );
buf ( n58443 , n20187 );
buf ( n58444 , n58443 );
and ( n58445 , n57948 , n58444 );
not ( n58446 , n58445 );
xor ( n58447 , n58093 , n58097 );
xor ( n58448 , n58447 , n58102 );
and ( n58449 , n58446 , n58448 );
buf ( n58450 , n58449 );
and ( n58451 , n58441 , n58450 );
and ( n58452 , n58420 , n58450 );
or ( n58453 , n58442 , n58451 , n58452 );
and ( n58454 , n58418 , n58453 );
and ( n58455 , n58416 , n58453 );
or ( n58456 , n58419 , n58454 , n58455 );
and ( n58457 , n58414 , n58456 );
xnor ( n58458 , n58135 , n58139 );
xnor ( n58459 , n58144 , n58147 );
and ( n58460 , n58458 , n58459 );
xnor ( n58461 , n58153 , n58157 );
and ( n58462 , n58459 , n58461 );
and ( n58463 , n58458 , n58461 );
or ( n58464 , n58460 , n58462 , n58463 );
xnor ( n58465 , n58165 , n58169 );
xor ( n58466 , n58174 , n58178 );
and ( n58467 , n58465 , n58466 );
xor ( n58468 , n58184 , n58188 );
and ( n58469 , n58466 , n58468 );
and ( n58470 , n58465 , n58468 );
or ( n58471 , n58467 , n58469 , n58470 );
and ( n58472 , n58464 , n58471 );
and ( n58473 , n51510 , n47429 );
and ( n58474 , n51298 , n47427 );
nor ( n58475 , n58473 , n58474 );
xnor ( n58476 , n58475 , n47309 );
and ( n58477 , n52082 , n47178 );
and ( n58478 , n51734 , n47176 );
nor ( n58479 , n58477 , n58478 );
xnor ( n58480 , n58479 , n47039 );
and ( n58481 , n58476 , n58480 );
and ( n58482 , n58480 , n58145 );
and ( n58483 , n58476 , n58145 );
or ( n58484 , n58481 , n58482 , n58483 );
and ( n58485 , n54227 , n46306 );
and ( n58486 , n53922 , n46304 );
nor ( n58487 , n58485 , n58486 );
xnor ( n58488 , n58487 , n46228 );
and ( n58489 , n55497 , n45990 );
and ( n58490 , n55143 , n45988 );
nor ( n58491 , n58489 , n58490 );
xnor ( n58492 , n58491 , n45939 );
or ( n58493 , n58488 , n58492 );
and ( n58494 , n58484 , n58493 );
and ( n58495 , n46843 , n52799 );
and ( n58496 , n46750 , n52797 );
nor ( n58497 , n58495 , n58496 );
xnor ( n58498 , n58497 , n52538 );
and ( n58499 , n47090 , n52269 );
and ( n58500 , n46969 , n52267 );
nor ( n58501 , n58499 , n58500 );
xnor ( n58502 , n58501 , n52008 );
or ( n58503 , n58498 , n58502 );
and ( n58504 , n58493 , n58503 );
and ( n58505 , n58484 , n58503 );
or ( n58506 , n58494 , n58504 , n58505 );
and ( n58507 , n58471 , n58506 );
and ( n58508 , n58464 , n58506 );
or ( n58509 , n58472 , n58507 , n58508 );
and ( n58510 , n49781 , n48740 );
and ( n58511 , n49570 , n48738 );
nor ( n58512 , n58510 , n58511 );
xnor ( n58513 , n58512 , n48571 );
and ( n58514 , n51077 , n47734 );
and ( n58515 , n50726 , n47732 );
nor ( n58516 , n58514 , n58515 );
xnor ( n58517 , n58516 , n47606 );
or ( n58518 , n58513 , n58517 );
and ( n58519 , n46264 , n54535 );
and ( n58520 , n46169 , n54533 );
nor ( n58521 , n58519 , n58520 );
xnor ( n58522 , n58521 , n54237 );
and ( n58523 , n48272 , n50338 );
and ( n58524 , n48108 , n50336 );
nor ( n58525 , n58523 , n58524 );
xnor ( n58526 , n58525 , n50111 );
or ( n58527 , n58522 , n58526 );
and ( n58528 , n58518 , n58527 );
and ( n58529 , n50195 , n48394 );
and ( n58530 , n49976 , n48392 );
nor ( n58531 , n58529 , n58530 );
xnor ( n58532 , n58531 , n48220 );
and ( n58533 , n53041 , n46712 );
and ( n58534 , n52790 , n46710 );
nor ( n58535 , n58533 , n58534 );
xnor ( n58536 , n58535 , n46587 );
or ( n58537 , n58532 , n58536 );
and ( n58538 , n58527 , n58537 );
and ( n58539 , n58518 , n58537 );
or ( n58540 , n58528 , n58538 , n58539 );
buf ( n58541 , n20190 );
buf ( n58542 , n58541 );
and ( n58543 , n57948 , n58542 );
not ( n58544 , n58543 );
buf ( n58545 , n58292 );
not ( n58546 , n58545 );
or ( n58547 , n58544 , n58546 );
and ( n58548 , n45763 , n57187 );
and ( n58549 , n45712 , n57184 );
nor ( n58550 , n58548 , n58549 );
xnor ( n58551 , n58550 , n56175 );
and ( n58552 , n45843 , n56503 );
and ( n58553 , n45794 , n56501 );
nor ( n58554 , n58552 , n58553 );
xnor ( n58555 , n58554 , n56178 );
and ( n58556 , n58551 , n58555 );
and ( n58557 , n45963 , n55851 );
and ( n58558 , n45907 , n55849 );
nor ( n58559 , n58557 , n58558 );
xnor ( n58560 , n58559 , n55506 );
and ( n58561 , n58555 , n58560 );
and ( n58562 , n58551 , n58560 );
or ( n58563 , n58556 , n58561 , n58562 );
and ( n58564 , n58547 , n58563 );
and ( n58565 , n46100 , n55159 );
and ( n58566 , n46041 , n55157 );
nor ( n58567 , n58565 , n58566 );
xnor ( n58568 , n58567 , n54864 );
and ( n58569 , n46445 , n53928 );
and ( n58570 , n46345 , n53926 );
nor ( n58571 , n58569 , n58570 );
xnor ( n58572 , n58571 , n53652 );
and ( n58573 , n58568 , n58572 );
and ( n58574 , n46577 , n53357 );
and ( n58575 , n46530 , n53355 );
nor ( n58576 , n58574 , n58575 );
xnor ( n58577 , n58576 , n53060 );
and ( n58578 , n58572 , n58577 );
and ( n58579 , n58568 , n58577 );
or ( n58580 , n58573 , n58578 , n58579 );
and ( n58581 , n58563 , n58580 );
and ( n58582 , n58547 , n58580 );
or ( n58583 , n58564 , n58581 , n58582 );
and ( n58584 , n58540 , n58583 );
and ( n58585 , n49374 , n49121 );
and ( n58586 , n49115 , n49119 );
nor ( n58587 , n58585 , n58586 );
xnor ( n58588 , n58587 , n48932 );
and ( n58589 , n50625 , n48042 );
and ( n58590 , n50404 , n48040 );
nor ( n58591 , n58589 , n58590 );
xnor ( n58592 , n58591 , n47921 );
and ( n58593 , n58588 , n58592 );
and ( n58594 , n52612 , n46911 );
and ( n58595 , n52332 , n46909 );
nor ( n58596 , n58594 , n58595 );
xnor ( n58597 , n58596 , n46802 );
and ( n58598 , n58592 , n58597 );
and ( n58599 , n58588 , n58597 );
or ( n58600 , n58593 , n58598 , n58599 );
and ( n58601 , n53639 , n46496 );
and ( n58602 , n53328 , n46494 );
nor ( n58603 , n58601 , n58602 );
xnor ( n58604 , n58603 , n46402 );
and ( n58605 , n54942 , n46135 );
and ( n58606 , n54604 , n46133 );
nor ( n58607 , n58605 , n58606 );
xnor ( n58608 , n58607 , n46067 );
and ( n58609 , n58604 , n58608 );
and ( n58610 , n56255 , n45886 );
and ( n58611 , n55756 , n45884 );
nor ( n58612 , n58610 , n58611 );
xnor ( n58613 , n58612 , n45824 );
and ( n58614 , n58608 , n58613 );
and ( n58615 , n58604 , n58613 );
or ( n58616 , n58609 , n58614 , n58615 );
and ( n58617 , n58600 , n58616 );
and ( n58618 , n56915 , n45777 );
and ( n58619 , n56388 , n45775 );
nor ( n58620 , n58618 , n58619 );
xnor ( n58621 , n58620 , n45734 );
xor ( n58622 , n39394 , n45579 );
buf ( n58623 , n58622 );
buf ( n58624 , n58623 );
buf ( n58625 , n58624 );
and ( n58626 , n58621 , n58625 );
buf ( n58627 , n20190 );
buf ( n58628 , n58627 );
and ( n58629 , n58628 , n58294 );
not ( n58630 , n58629 );
and ( n58631 , n58625 , n58630 );
and ( n58632 , n58621 , n58630 );
or ( n58633 , n58626 , n58631 , n58632 );
and ( n58634 , n58616 , n58633 );
and ( n58635 , n58600 , n58633 );
or ( n58636 , n58617 , n58634 , n58635 );
and ( n58637 , n58583 , n58636 );
and ( n58638 , n58540 , n58636 );
or ( n58639 , n58584 , n58637 , n58638 );
and ( n58640 , n58509 , n58639 );
xor ( n58641 , n58197 , n58201 );
xor ( n58642 , n58641 , n58206 );
xor ( n58643 , n58213 , n58217 );
xor ( n58644 , n58643 , n58222 );
and ( n58645 , n58642 , n58644 );
xor ( n58646 , n58230 , n58234 );
xor ( n58647 , n58646 , n58239 );
and ( n58648 , n58644 , n58647 );
and ( n58649 , n58642 , n58647 );
or ( n58650 , n58645 , n58648 , n58649 );
xor ( n58651 , n58252 , n58256 );
xor ( n58652 , n58651 , n58261 );
xor ( n58653 , n58268 , n58272 );
xor ( n58654 , n58653 , n58277 );
and ( n58655 , n58652 , n58654 );
xor ( n58656 , n58285 , n58289 );
xor ( n58657 , n58656 , n58296 );
and ( n58658 , n58654 , n58657 );
and ( n58659 , n58652 , n58657 );
or ( n58660 , n58655 , n58658 , n58659 );
and ( n58661 , n58650 , n58660 );
xor ( n58662 , n58110 , n58112 );
xor ( n58663 , n58662 , n58114 );
and ( n58664 , n58660 , n58663 );
and ( n58665 , n58650 , n58663 );
or ( n58666 , n58661 , n58664 , n58665 );
and ( n58667 , n58639 , n58666 );
and ( n58668 , n58509 , n58666 );
or ( n58669 , n58640 , n58667 , n58668 );
and ( n58670 , n58456 , n58669 );
and ( n58671 , n58414 , n58669 );
or ( n58672 , n58457 , n58670 , n58671 );
and ( n58673 , n58411 , n58672 );
and ( n58674 , n58409 , n58672 );
or ( n58675 , n58412 , n58673 , n58674 );
and ( n58676 , n58406 , n58675 );
and ( n58677 , n58404 , n58675 );
or ( n58678 , n58407 , n58676 , n58677 );
and ( n58679 , n58402 , n58678 );
xor ( n58680 , n58077 , n58386 );
xor ( n58681 , n58680 , n58389 );
and ( n58682 , n58678 , n58681 );
and ( n58683 , n58402 , n58681 );
or ( n58684 , n58679 , n58682 , n58683 );
and ( n58685 , n58400 , n58684 );
xor ( n58686 , n58072 , n58074 );
xor ( n58687 , n58686 , n58392 );
and ( n58688 , n58684 , n58687 );
and ( n58689 , n58400 , n58687 );
or ( n58690 , n58685 , n58688 , n58689 );
and ( n58691 , n58397 , n58690 );
and ( n58692 , n58395 , n58690 );
or ( n58693 , n58398 , n58691 , n58692 );
and ( n58694 , n58030 , n58693 );
xor ( n58695 , n58030 , n58693 );
xor ( n58696 , n58395 , n58397 );
xor ( n58697 , n58696 , n58690 );
not ( n58698 , n58697 );
xor ( n58699 , n58400 , n58684 );
xor ( n58700 , n58699 , n58687 );
xor ( n58701 , n58119 , n58120 );
xor ( n58702 , n58701 , n58122 );
xor ( n58703 , n58140 , n58148 );
xor ( n58704 , n58703 , n58158 );
and ( n58705 , n58702 , n58704 );
xor ( n58706 , n58170 , n58179 );
xor ( n58707 , n58706 , n58189 );
and ( n58708 , n58704 , n58707 );
and ( n58709 , n58702 , n58707 );
or ( n58710 , n58705 , n58708 , n58709 );
xor ( n58711 , n58209 , n58225 );
xor ( n58712 , n58711 , n58242 );
xor ( n58713 , n58264 , n58280 );
xor ( n58714 , n58713 , n58299 );
and ( n58715 , n58712 , n58714 );
xor ( n58716 , n58304 , n58306 );
xor ( n58717 , n58716 , n58309 );
and ( n58718 , n58714 , n58717 );
and ( n58719 , n58712 , n58717 );
or ( n58720 , n58715 , n58718 , n58719 );
and ( n58721 , n58710 , n58720 );
xor ( n58722 , n58081 , n58083 );
xor ( n58723 , n58722 , n58085 );
and ( n58724 , n58720 , n58723 );
and ( n58725 , n58710 , n58723 );
or ( n58726 , n58721 , n58724 , n58725 );
xor ( n58727 , n58108 , n58117 );
xor ( n58728 , n58727 , n58125 );
xor ( n58729 , n58161 , n58192 );
xor ( n58730 , n58729 , n58245 );
and ( n58731 , n58728 , n58730 );
xor ( n58732 , n58302 , n58312 );
xor ( n58733 , n58732 , n58323 );
and ( n58734 , n58730 , n58733 );
and ( n58735 , n58728 , n58733 );
or ( n58736 , n58731 , n58734 , n58735 );
and ( n58737 , n58726 , n58736 );
xor ( n58738 , n58079 , n58088 );
xor ( n58739 , n58738 , n58128 );
and ( n58740 , n58736 , n58739 );
and ( n58741 , n58726 , n58739 );
or ( n58742 , n58737 , n58740 , n58741 );
xor ( n58743 , n58248 , n58326 );
xor ( n58744 , n58743 , n58337 );
xor ( n58745 , n58351 , n58353 );
xor ( n58746 , n58745 , n58356 );
and ( n58747 , n58744 , n58746 );
xor ( n58748 , n58364 , n58366 );
xor ( n58749 , n58748 , n58369 );
and ( n58750 , n58746 , n58749 );
and ( n58751 , n58744 , n58749 );
or ( n58752 , n58747 , n58750 , n58751 );
and ( n58753 , n58742 , n58752 );
xor ( n58754 , n58131 , n58340 );
xor ( n58755 , n58754 , n58359 );
and ( n58756 , n58752 , n58755 );
and ( n58757 , n58742 , n58755 );
or ( n58758 , n58753 , n58756 , n58757 );
xor ( n58759 , n58362 , n58380 );
xor ( n58760 , n58759 , n58383 );
and ( n58761 , n58758 , n58760 );
xor ( n58762 , n58372 , n58374 );
xor ( n58763 , n58762 , n58377 );
xor ( n58764 , n58329 , n58331 );
xor ( n58765 , n58764 , n58334 );
xor ( n58766 , n58343 , n58345 );
xor ( n58767 , n58766 , n58348 );
and ( n58768 , n58765 , n58767 );
xor ( n58769 , n58315 , n58317 );
xor ( n58770 , n58769 , n58320 );
xnor ( n58771 , n58436 , n58440 );
and ( n58772 , n46345 , n54535 );
and ( n58773 , n46264 , n54533 );
nor ( n58774 , n58772 , n58773 );
xnor ( n58775 , n58774 , n54237 );
and ( n58776 , n46530 , n53928 );
and ( n58777 , n46445 , n53926 );
nor ( n58778 , n58776 , n58777 );
xnor ( n58779 , n58778 , n53652 );
and ( n58780 , n58775 , n58779 );
and ( n58781 , n46750 , n53357 );
and ( n58782 , n46577 , n53355 );
nor ( n58783 , n58781 , n58782 );
xnor ( n58784 , n58783 , n53060 );
and ( n58785 , n58779 , n58784 );
and ( n58786 , n58775 , n58784 );
or ( n58787 , n58780 , n58785 , n58786 );
xor ( n58788 , n58424 , n58428 );
xor ( n58789 , n58788 , n58433 );
or ( n58790 , n58787 , n58789 );
and ( n58791 , n58771 , n58790 );
and ( n58792 , n46969 , n52799 );
and ( n58793 , n46843 , n52797 );
nor ( n58794 , n58792 , n58793 );
xnor ( n58795 , n58794 , n52538 );
and ( n58796 , n47216 , n52269 );
and ( n58797 , n47090 , n52267 );
nor ( n58798 , n58796 , n58797 );
xnor ( n58799 , n58798 , n52008 );
and ( n58800 , n58795 , n58799 );
and ( n58801 , n47778 , n51221 );
and ( n58802 , n47647 , n51219 );
nor ( n58803 , n58801 , n58802 );
xnor ( n58804 , n58803 , n51000 );
and ( n58805 , n58799 , n58804 );
and ( n58806 , n58795 , n58804 );
or ( n58807 , n58800 , n58805 , n58806 );
and ( n58808 , n48632 , n49896 );
and ( n58809 , n48384 , n49894 );
nor ( n58810 , n58808 , n58809 );
xnor ( n58811 , n58810 , n49711 );
and ( n58812 , n58807 , n58811 );
and ( n58813 , n58790 , n58812 );
and ( n58814 , n58771 , n58812 );
or ( n58815 , n58791 , n58813 , n58814 );
and ( n58816 , n58770 , n58815 );
xor ( n58817 , n58476 , n58480 );
xor ( n58818 , n58817 , n58145 );
xnor ( n58819 , n58488 , n58492 );
and ( n58820 , n58818 , n58819 );
buf ( n58821 , n58820 );
xnor ( n58822 , n58498 , n58502 );
xnor ( n58823 , n58513 , n58517 );
and ( n58824 , n58822 , n58823 );
xnor ( n58825 , n58522 , n58526 );
and ( n58826 , n58823 , n58825 );
and ( n58827 , n58822 , n58825 );
or ( n58828 , n58824 , n58826 , n58827 );
and ( n58829 , n58821 , n58828 );
xnor ( n58830 , n58532 , n58536 );
xnor ( n58831 , n58544 , n58546 );
and ( n58832 , n58830 , n58831 );
and ( n58833 , n50726 , n48042 );
and ( n58834 , n50625 , n48040 );
nor ( n58835 , n58833 , n58834 );
xnor ( n58836 , n58835 , n47921 );
and ( n58837 , n51734 , n47429 );
and ( n58838 , n51510 , n47427 );
nor ( n58839 , n58837 , n58838 );
xnor ( n58840 , n58839 , n47309 );
and ( n58841 , n58836 , n58840 );
and ( n58842 , n52790 , n46911 );
and ( n58843 , n52612 , n46909 );
nor ( n58844 , n58842 , n58843 );
xnor ( n58845 , n58844 , n46802 );
and ( n58846 , n58840 , n58845 );
and ( n58847 , n58836 , n58845 );
or ( n58848 , n58841 , n58846 , n58847 );
and ( n58849 , n58831 , n58848 );
and ( n58850 , n58830 , n58848 );
or ( n58851 , n58832 , n58849 , n58850 );
and ( n58852 , n58828 , n58851 );
and ( n58853 , n58821 , n58851 );
or ( n58854 , n58829 , n58852 , n58853 );
and ( n58855 , n58815 , n58854 );
and ( n58856 , n58770 , n58854 );
or ( n58857 , n58816 , n58855 , n58856 );
and ( n58858 , n58767 , n58857 );
and ( n58859 , n58765 , n58857 );
or ( n58860 , n58768 , n58858 , n58859 );
and ( n58861 , n53328 , n46712 );
and ( n58862 , n53041 , n46710 );
nor ( n58863 , n58861 , n58862 );
xnor ( n58864 , n58863 , n46587 );
and ( n58865 , n57063 , n45775 );
not ( n58866 , n58865 );
and ( n58867 , n58866 , n45734 );
or ( n58868 , n58864 , n58867 );
and ( n58869 , n55143 , n46135 );
and ( n58870 , n54942 , n46133 );
nor ( n58871 , n58869 , n58870 );
xnor ( n58872 , n58871 , n46067 );
and ( n58873 , n57063 , n45777 );
and ( n58874 , n56915 , n45775 );
nor ( n58875 , n58873 , n58874 );
xnor ( n58876 , n58875 , n45734 );
or ( n58877 , n58872 , n58876 );
and ( n58878 , n58868 , n58877 );
and ( n58879 , n54604 , n46306 );
and ( n58880 , n54227 , n46304 );
nor ( n58881 , n58879 , n58880 );
xnor ( n58882 , n58881 , n46228 );
and ( n58883 , n55756 , n45990 );
and ( n58884 , n55497 , n45988 );
nor ( n58885 , n58883 , n58884 );
xnor ( n58886 , n58885 , n45939 );
or ( n58887 , n58882 , n58886 );
and ( n58888 , n58877 , n58887 );
and ( n58889 , n58868 , n58887 );
or ( n58890 , n58878 , n58888 , n58889 );
and ( n58891 , n49976 , n48740 );
and ( n58892 , n49781 , n48738 );
nor ( n58893 , n58891 , n58892 );
xnor ( n58894 , n58893 , n48571 );
and ( n58895 , n51298 , n47734 );
and ( n58896 , n51077 , n47732 );
nor ( n58897 , n58895 , n58896 );
xnor ( n58898 , n58897 , n47606 );
or ( n58899 , n58894 , n58898 );
and ( n58900 , n47474 , n51750 );
and ( n58901 , n47351 , n51748 );
nor ( n58902 , n58900 , n58901 );
xnor ( n58903 , n58902 , n51520 );
and ( n58904 , n48108 , n50783 );
and ( n58905 , n47962 , n50781 );
nor ( n58906 , n58904 , n58905 );
xnor ( n58907 , n58906 , n50557 );
and ( n58908 , n58903 , n58907 );
and ( n58909 , n58899 , n58908 );
buf ( n58910 , n20193 );
buf ( n58911 , n58910 );
and ( n58912 , n57948 , n58911 );
not ( n58913 , n58912 );
buf ( n58914 , n20193 );
buf ( n58915 , n58914 );
and ( n58916 , n58915 , n58294 );
not ( n58917 , n58916 );
and ( n58918 , n58913 , n58917 );
and ( n58919 , n58908 , n58918 );
and ( n58920 , n58899 , n58918 );
or ( n58921 , n58909 , n58919 , n58920 );
and ( n58922 , n58890 , n58921 );
and ( n58923 , n45794 , n57187 );
and ( n58924 , n45763 , n57184 );
nor ( n58925 , n58923 , n58924 );
xnor ( n58926 , n58925 , n56175 );
and ( n58927 , n45907 , n56503 );
and ( n58928 , n45843 , n56501 );
nor ( n58929 , n58927 , n58928 );
xnor ( n58930 , n58929 , n56178 );
and ( n58931 , n58926 , n58930 );
and ( n58932 , n46041 , n55851 );
and ( n58933 , n45963 , n55849 );
nor ( n58934 , n58932 , n58933 );
xnor ( n58935 , n58934 , n55506 );
and ( n58936 , n58930 , n58935 );
and ( n58937 , n58926 , n58935 );
or ( n58938 , n58931 , n58936 , n58937 );
and ( n58939 , n46169 , n55159 );
and ( n58940 , n46100 , n55157 );
nor ( n58941 , n58939 , n58940 );
xnor ( n58942 , n58941 , n54864 );
and ( n58943 , n48709 , n49896 );
and ( n58944 , n48632 , n49894 );
nor ( n58945 , n58943 , n58944 );
xnor ( n58946 , n58945 , n49711 );
and ( n58947 , n58942 , n58946 );
and ( n58948 , n49115 , n49513 );
and ( n58949 , n48988 , n49511 );
nor ( n58950 , n58948 , n58949 );
xnor ( n58951 , n58950 , n49310 );
and ( n58952 , n58946 , n58951 );
and ( n58953 , n58942 , n58951 );
or ( n58954 , n58947 , n58952 , n58953 );
and ( n58955 , n58938 , n58954 );
and ( n58956 , n49570 , n49121 );
and ( n58957 , n49374 , n49119 );
nor ( n58958 , n58956 , n58957 );
xnor ( n58959 , n58958 , n48932 );
and ( n58960 , n50404 , n48394 );
and ( n58961 , n50195 , n48392 );
nor ( n58962 , n58960 , n58961 );
xnor ( n58963 , n58962 , n48220 );
and ( n58964 , n58959 , n58963 );
and ( n58965 , n52332 , n47178 );
and ( n58966 , n52082 , n47176 );
nor ( n58967 , n58965 , n58966 );
xnor ( n58968 , n58967 , n47039 );
and ( n58969 , n58963 , n58968 );
and ( n58970 , n58959 , n58968 );
or ( n58971 , n58964 , n58969 , n58970 );
and ( n58972 , n58954 , n58971 );
and ( n58973 , n58938 , n58971 );
or ( n58974 , n58955 , n58972 , n58973 );
and ( n58975 , n58921 , n58974 );
and ( n58976 , n58890 , n58974 );
or ( n58977 , n58922 , n58975 , n58976 );
and ( n58978 , n53922 , n46496 );
and ( n58979 , n53639 , n46494 );
nor ( n58980 , n58978 , n58979 );
xnor ( n58981 , n58980 , n46402 );
and ( n58982 , n56388 , n45886 );
and ( n58983 , n56255 , n45884 );
nor ( n58984 , n58982 , n58983 );
xnor ( n58985 , n58984 , n45824 );
and ( n58986 , n58981 , n58985 );
xor ( n58987 , n39397 , n45577 );
buf ( n58988 , n58987 );
buf ( n58989 , n58988 );
buf ( n58990 , n58989 );
and ( n58991 , n58985 , n58990 );
and ( n58992 , n58981 , n58990 );
or ( n58993 , n58986 , n58991 , n58992 );
and ( n58994 , n58628 , n58444 );
not ( n58995 , n58994 );
and ( n58996 , n58292 , n58542 );
not ( n58997 , n58996 );
and ( n58998 , n58995 , n58997 );
buf ( n58999 , n58998 );
and ( n59000 , n58993 , n58999 );
xor ( n59001 , n58551 , n58555 );
xor ( n59002 , n59001 , n58560 );
and ( n59003 , n58999 , n59002 );
and ( n59004 , n58993 , n59002 );
or ( n59005 , n59000 , n59003 , n59004 );
xor ( n59006 , n58568 , n58572 );
xor ( n59007 , n59006 , n58577 );
xor ( n59008 , n58588 , n58592 );
xor ( n59009 , n59008 , n58597 );
and ( n59010 , n59007 , n59009 );
xor ( n59011 , n58604 , n58608 );
xor ( n59012 , n59011 , n58613 );
and ( n59013 , n59009 , n59012 );
and ( n59014 , n59007 , n59012 );
or ( n59015 , n59010 , n59013 , n59014 );
and ( n59016 , n59005 , n59015 );
buf ( n59017 , n58446 );
xor ( n59018 , n59017 , n58448 );
and ( n59019 , n59015 , n59018 );
and ( n59020 , n59005 , n59018 );
or ( n59021 , n59016 , n59019 , n59020 );
and ( n59022 , n58977 , n59021 );
xor ( n59023 , n58458 , n58459 );
xor ( n59024 , n59023 , n58461 );
xor ( n59025 , n58465 , n58466 );
xor ( n59026 , n59025 , n58468 );
and ( n59027 , n59024 , n59026 );
xor ( n59028 , n58484 , n58493 );
xor ( n59029 , n59028 , n58503 );
and ( n59030 , n59026 , n59029 );
and ( n59031 , n59024 , n59029 );
or ( n59032 , n59027 , n59030 , n59031 );
and ( n59033 , n59021 , n59032 );
and ( n59034 , n58977 , n59032 );
or ( n59035 , n59022 , n59033 , n59034 );
xor ( n59036 , n58518 , n58527 );
xor ( n59037 , n59036 , n58537 );
xor ( n59038 , n58547 , n58563 );
xor ( n59039 , n59038 , n58580 );
and ( n59040 , n59037 , n59039 );
xor ( n59041 , n58600 , n58616 );
xor ( n59042 , n59041 , n58633 );
and ( n59043 , n59039 , n59042 );
and ( n59044 , n59037 , n59042 );
or ( n59045 , n59040 , n59043 , n59044 );
xor ( n59046 , n58420 , n58441 );
xor ( n59047 , n59046 , n58450 );
and ( n59048 , n59045 , n59047 );
xor ( n59049 , n58464 , n58471 );
xor ( n59050 , n59049 , n58506 );
and ( n59051 , n59047 , n59050 );
and ( n59052 , n59045 , n59050 );
or ( n59053 , n59048 , n59051 , n59052 );
and ( n59054 , n59035 , n59053 );
xor ( n59055 , n58540 , n58583 );
xor ( n59056 , n59055 , n58636 );
xor ( n59057 , n58650 , n58660 );
xor ( n59058 , n59057 , n58663 );
and ( n59059 , n59056 , n59058 );
xor ( n59060 , n58702 , n58704 );
xor ( n59061 , n59060 , n58707 );
and ( n59062 , n59058 , n59061 );
and ( n59063 , n59056 , n59061 );
or ( n59064 , n59059 , n59062 , n59063 );
and ( n59065 , n59053 , n59064 );
and ( n59066 , n59035 , n59064 );
or ( n59067 , n59054 , n59065 , n59066 );
and ( n59068 , n58860 , n59067 );
xor ( n59069 , n58416 , n58418 );
xor ( n59070 , n59069 , n58453 );
xor ( n59071 , n58509 , n58639 );
xor ( n59072 , n59071 , n58666 );
and ( n59073 , n59070 , n59072 );
xor ( n59074 , n58710 , n58720 );
xor ( n59075 , n59074 , n58723 );
and ( n59076 , n59072 , n59075 );
and ( n59077 , n59070 , n59075 );
or ( n59078 , n59073 , n59076 , n59077 );
and ( n59079 , n59067 , n59078 );
and ( n59080 , n58860 , n59078 );
or ( n59081 , n59068 , n59079 , n59080 );
and ( n59082 , n58763 , n59081 );
xor ( n59083 , n58414 , n58456 );
xor ( n59084 , n59083 , n58669 );
xor ( n59085 , n58726 , n58736 );
xor ( n59086 , n59085 , n58739 );
and ( n59087 , n59084 , n59086 );
xor ( n59088 , n58744 , n58746 );
xor ( n59089 , n59088 , n58749 );
and ( n59090 , n59086 , n59089 );
and ( n59091 , n59084 , n59089 );
or ( n59092 , n59087 , n59090 , n59091 );
and ( n59093 , n59081 , n59092 );
and ( n59094 , n58763 , n59092 );
or ( n59095 , n59082 , n59093 , n59094 );
and ( n59096 , n58760 , n59095 );
and ( n59097 , n58758 , n59095 );
or ( n59098 , n58761 , n59096 , n59097 );
xor ( n59099 , n58402 , n58678 );
xor ( n59100 , n59099 , n58681 );
and ( n59101 , n59098 , n59100 );
xor ( n59102 , n58404 , n58406 );
xor ( n59103 , n59102 , n58675 );
xor ( n59104 , n58409 , n58411 );
xor ( n59105 , n59104 , n58672 );
xor ( n59106 , n58742 , n58752 );
xor ( n59107 , n59106 , n58755 );
and ( n59108 , n59105 , n59107 );
xor ( n59109 , n58728 , n58730 );
xor ( n59110 , n59109 , n58733 );
xor ( n59111 , n58712 , n58714 );
xor ( n59112 , n59111 , n58717 );
xor ( n59113 , n58642 , n58644 );
xor ( n59114 , n59113 , n58647 );
xor ( n59115 , n58652 , n58654 );
xor ( n59116 , n59115 , n58657 );
and ( n59117 , n59114 , n59116 );
and ( n59118 , n48988 , n49513 );
and ( n59119 , n48709 , n49511 );
nor ( n59120 , n59118 , n59119 );
xnor ( n59121 , n59120 , n49310 );
not ( n59122 , n59121 );
xnor ( n59123 , n58787 , n58789 );
and ( n59124 , n59122 , n59123 );
and ( n59125 , n59116 , n59124 );
and ( n59126 , n59114 , n59124 );
or ( n59127 , n59117 , n59125 , n59126 );
and ( n59128 , n59112 , n59127 );
buf ( n59129 , n59121 );
xor ( n59130 , n58621 , n58625 );
xor ( n59131 , n59130 , n58630 );
xor ( n59132 , n58807 , n58811 );
and ( n59133 , n59131 , n59132 );
and ( n59134 , n47090 , n52799 );
and ( n59135 , n46969 , n52797 );
nor ( n59136 , n59134 , n59135 );
xnor ( n59137 , n59136 , n52538 );
and ( n59138 , n47351 , n52269 );
and ( n59139 , n47216 , n52267 );
nor ( n59140 , n59138 , n59139 );
xnor ( n59141 , n59140 , n52008 );
and ( n59142 , n59137 , n59141 );
and ( n59143 , n47962 , n51221 );
and ( n59144 , n47778 , n51219 );
nor ( n59145 , n59143 , n59144 );
xnor ( n59146 , n59145 , n51000 );
and ( n59147 , n59141 , n59146 );
and ( n59148 , n59137 , n59146 );
or ( n59149 , n59142 , n59147 , n59148 );
and ( n59150 , n48384 , n50338 );
and ( n59151 , n48272 , n50336 );
nor ( n59152 , n59150 , n59151 );
xnor ( n59153 , n59152 , n50111 );
or ( n59154 , n59149 , n59153 );
and ( n59155 , n59132 , n59154 );
and ( n59156 , n59131 , n59154 );
or ( n59157 , n59133 , n59155 , n59156 );
and ( n59158 , n59129 , n59157 );
xor ( n59159 , n58795 , n58799 );
xor ( n59160 , n59159 , n58804 );
xor ( n59161 , n58775 , n58779 );
xor ( n59162 , n59161 , n58784 );
and ( n59163 , n59160 , n59162 );
xor ( n59164 , n58836 , n58840 );
xor ( n59165 , n59164 , n58845 );
and ( n59166 , n59162 , n59165 );
and ( n59167 , n59160 , n59165 );
or ( n59168 , n59163 , n59166 , n59167 );
xnor ( n59169 , n58864 , n58867 );
xnor ( n59170 , n58872 , n58876 );
and ( n59171 , n59169 , n59170 );
xnor ( n59172 , n58882 , n58886 );
and ( n59173 , n59170 , n59172 );
and ( n59174 , n59169 , n59172 );
or ( n59175 , n59171 , n59173 , n59174 );
and ( n59176 , n59168 , n59175 );
xnor ( n59177 , n58894 , n58898 );
xor ( n59178 , n58903 , n58907 );
and ( n59179 , n59177 , n59178 );
xor ( n59180 , n58913 , n58917 );
and ( n59181 , n59178 , n59180 );
and ( n59182 , n59177 , n59180 );
or ( n59183 , n59179 , n59181 , n59182 );
and ( n59184 , n59175 , n59183 );
and ( n59185 , n59168 , n59183 );
or ( n59186 , n59176 , n59184 , n59185 );
and ( n59187 , n59157 , n59186 );
and ( n59188 , n59129 , n59186 );
or ( n59189 , n59158 , n59187 , n59188 );
and ( n59190 , n59127 , n59189 );
and ( n59191 , n59112 , n59189 );
or ( n59192 , n59128 , n59190 , n59191 );
and ( n59193 , n59110 , n59192 );
and ( n59194 , n52612 , n47178 );
and ( n59195 , n52332 , n47176 );
nor ( n59196 , n59194 , n59195 );
xnor ( n59197 , n59196 , n47039 );
and ( n59198 , n53041 , n46911 );
and ( n59199 , n52790 , n46909 );
nor ( n59200 , n59198 , n59199 );
xnor ( n59201 , n59200 , n46802 );
and ( n59202 , n59197 , n59201 );
and ( n59203 , n59201 , n58865 );
and ( n59204 , n59197 , n58865 );
or ( n59205 , n59202 , n59203 , n59204 );
buf ( n59206 , n20196 );
buf ( n59207 , n59206 );
and ( n59208 , n57948 , n59207 );
not ( n59209 , n59208 );
and ( n59210 , n58292 , n58911 );
and ( n59211 , n59209 , n59210 );
buf ( n59212 , n58628 );
not ( n59213 , n59212 );
and ( n59214 , n59210 , n59213 );
and ( n59215 , n59209 , n59213 );
or ( n59216 , n59211 , n59214 , n59215 );
and ( n59217 , n59205 , n59216 );
not ( n59218 , n59210 );
buf ( n59219 , n59218 );
and ( n59220 , n59216 , n59219 );
and ( n59221 , n59205 , n59219 );
or ( n59222 , n59217 , n59220 , n59221 );
and ( n59223 , n52082 , n47429 );
and ( n59224 , n51734 , n47427 );
nor ( n59225 , n59223 , n59224 );
xnor ( n59226 , n59225 , n47309 );
and ( n59227 , n53639 , n46712 );
and ( n59228 , n53328 , n46710 );
nor ( n59229 , n59227 , n59228 );
xnor ( n59230 , n59229 , n46587 );
or ( n59231 , n59226 , n59230 );
and ( n59232 , n46445 , n54535 );
and ( n59233 , n46345 , n54533 );
nor ( n59234 , n59232 , n59233 );
xnor ( n59235 , n59234 , n54237 );
and ( n59236 , n46577 , n53928 );
and ( n59237 , n46530 , n53926 );
nor ( n59238 , n59236 , n59237 );
xnor ( n59239 , n59238 , n53652 );
or ( n59240 , n59235 , n59239 );
and ( n59241 , n59231 , n59240 );
and ( n59242 , n46843 , n53357 );
and ( n59243 , n46750 , n53355 );
nor ( n59244 , n59242 , n59243 );
xnor ( n59245 , n59244 , n53060 );
and ( n59246 , n48272 , n50783 );
and ( n59247 , n48108 , n50781 );
nor ( n59248 , n59246 , n59247 );
xnor ( n59249 , n59248 , n50557 );
or ( n59250 , n59245 , n59249 );
and ( n59251 , n59240 , n59250 );
and ( n59252 , n59231 , n59250 );
or ( n59253 , n59241 , n59251 , n59252 );
and ( n59254 , n59222 , n59253 );
and ( n59255 , n54942 , n46306 );
and ( n59256 , n54604 , n46304 );
nor ( n59257 , n59255 , n59256 );
xnor ( n59258 , n59257 , n46228 );
and ( n59259 , n56255 , n45990 );
and ( n59260 , n55756 , n45988 );
nor ( n59261 , n59259 , n59260 );
xnor ( n59262 , n59261 , n45939 );
and ( n59263 , n59258 , n59262 );
and ( n59264 , n45843 , n57187 );
and ( n59265 , n45794 , n57184 );
nor ( n59266 , n59264 , n59265 );
xnor ( n59267 , n59266 , n56175 );
and ( n59268 , n45963 , n56503 );
and ( n59269 , n45907 , n56501 );
nor ( n59270 , n59268 , n59269 );
xnor ( n59271 , n59270 , n56178 );
and ( n59272 , n59267 , n59271 );
and ( n59273 , n46100 , n55851 );
and ( n59274 , n46041 , n55849 );
nor ( n59275 , n59273 , n59274 );
xnor ( n59276 , n59275 , n55506 );
and ( n59277 , n59271 , n59276 );
and ( n59278 , n59267 , n59276 );
or ( n59279 , n59272 , n59277 , n59278 );
and ( n59280 , n59263 , n59279 );
and ( n59281 , n46264 , n55159 );
and ( n59282 , n46169 , n55157 );
nor ( n59283 , n59281 , n59282 );
xnor ( n59284 , n59283 , n54864 );
and ( n59285 , n47647 , n51750 );
and ( n59286 , n47474 , n51748 );
nor ( n59287 , n59285 , n59286 );
xnor ( n59288 , n59287 , n51520 );
and ( n59289 , n59284 , n59288 );
and ( n59290 , n48632 , n50338 );
and ( n59291 , n48384 , n50336 );
nor ( n59292 , n59290 , n59291 );
xnor ( n59293 , n59292 , n50111 );
and ( n59294 , n59288 , n59293 );
and ( n59295 , n59284 , n59293 );
or ( n59296 , n59289 , n59294 , n59295 );
and ( n59297 , n59279 , n59296 );
and ( n59298 , n59263 , n59296 );
or ( n59299 , n59280 , n59297 , n59298 );
and ( n59300 , n59253 , n59299 );
and ( n59301 , n59222 , n59299 );
or ( n59302 , n59254 , n59300 , n59301 );
and ( n59303 , n48988 , n49896 );
and ( n59304 , n48709 , n49894 );
nor ( n59305 , n59303 , n59304 );
xnor ( n59306 , n59305 , n49711 );
and ( n59307 , n49374 , n49513 );
and ( n59308 , n49115 , n49511 );
nor ( n59309 , n59307 , n59308 );
xnor ( n59310 , n59309 , n49310 );
and ( n59311 , n59306 , n59310 );
and ( n59312 , n49781 , n49121 );
and ( n59313 , n49570 , n49119 );
nor ( n59314 , n59312 , n59313 );
xnor ( n59315 , n59314 , n48932 );
and ( n59316 , n59310 , n59315 );
and ( n59317 , n59306 , n59315 );
or ( n59318 , n59311 , n59316 , n59317 );
and ( n59319 , n50195 , n48740 );
and ( n59320 , n49976 , n48738 );
nor ( n59321 , n59319 , n59320 );
xnor ( n59322 , n59321 , n48571 );
and ( n59323 , n50625 , n48394 );
and ( n59324 , n50404 , n48392 );
nor ( n59325 , n59323 , n59324 );
xnor ( n59326 , n59325 , n48220 );
and ( n59327 , n59322 , n59326 );
and ( n59328 , n51077 , n48042 );
and ( n59329 , n50726 , n48040 );
nor ( n59330 , n59328 , n59329 );
xnor ( n59331 , n59330 , n47921 );
and ( n59332 , n59326 , n59331 );
and ( n59333 , n59322 , n59331 );
or ( n59334 , n59327 , n59332 , n59333 );
and ( n59335 , n59318 , n59334 );
and ( n59336 , n51510 , n47734 );
and ( n59337 , n51298 , n47732 );
nor ( n59338 , n59336 , n59337 );
xnor ( n59339 , n59338 , n47606 );
and ( n59340 , n54227 , n46496 );
and ( n59341 , n53922 , n46494 );
nor ( n59342 , n59340 , n59341 );
xnor ( n59343 , n59342 , n46402 );
and ( n59344 , n59339 , n59343 );
and ( n59345 , n55497 , n46135 );
and ( n59346 , n55143 , n46133 );
nor ( n59347 , n59345 , n59346 );
xnor ( n59348 , n59347 , n46067 );
and ( n59349 , n59343 , n59348 );
and ( n59350 , n59339 , n59348 );
or ( n59351 , n59344 , n59349 , n59350 );
and ( n59352 , n59334 , n59351 );
and ( n59353 , n59318 , n59351 );
or ( n59354 , n59335 , n59352 , n59353 );
and ( n59355 , n56915 , n45886 );
and ( n59356 , n56388 , n45884 );
nor ( n59357 , n59355 , n59356 );
xnor ( n59358 , n59357 , n45824 );
xor ( n59359 , n39400 , n45575 );
buf ( n59360 , n59359 );
buf ( n59361 , n59360 );
buf ( n59362 , n59361 );
and ( n59363 , n59358 , n59362 );
buf ( n59364 , n20196 );
buf ( n59365 , n59364 );
and ( n59366 , n59365 , n58294 );
not ( n59367 , n59366 );
and ( n59368 , n59362 , n59367 );
and ( n59369 , n59358 , n59367 );
or ( n59370 , n59363 , n59368 , n59369 );
xor ( n59371 , n58926 , n58930 );
xor ( n59372 , n59371 , n58935 );
and ( n59373 , n59370 , n59372 );
xor ( n59374 , n58942 , n58946 );
xor ( n59375 , n59374 , n58951 );
and ( n59376 , n59372 , n59375 );
and ( n59377 , n59370 , n59375 );
or ( n59378 , n59373 , n59376 , n59377 );
and ( n59379 , n59354 , n59378 );
xor ( n59380 , n58959 , n58963 );
xor ( n59381 , n59380 , n58968 );
xor ( n59382 , n58981 , n58985 );
xor ( n59383 , n59382 , n58990 );
and ( n59384 , n59381 , n59383 );
xor ( n59385 , n58995 , n58997 );
buf ( n59386 , n59385 );
and ( n59387 , n59383 , n59386 );
and ( n59388 , n59381 , n59386 );
or ( n59389 , n59384 , n59387 , n59388 );
and ( n59390 , n59378 , n59389 );
and ( n59391 , n59354 , n59389 );
or ( n59392 , n59379 , n59390 , n59391 );
and ( n59393 , n59302 , n59392 );
buf ( n59394 , n58818 );
xor ( n59395 , n59394 , n58819 );
xor ( n59396 , n58822 , n58823 );
xor ( n59397 , n59396 , n58825 );
and ( n59398 , n59395 , n59397 );
xor ( n59399 , n58830 , n58831 );
xor ( n59400 , n59399 , n58848 );
and ( n59401 , n59397 , n59400 );
and ( n59402 , n59395 , n59400 );
or ( n59403 , n59398 , n59401 , n59402 );
and ( n59404 , n59392 , n59403 );
and ( n59405 , n59302 , n59403 );
or ( n59406 , n59393 , n59404 , n59405 );
xor ( n59407 , n58868 , n58877 );
xor ( n59408 , n59407 , n58887 );
xor ( n59409 , n58899 , n58908 );
xor ( n59410 , n59409 , n58918 );
and ( n59411 , n59408 , n59410 );
xor ( n59412 , n58938 , n58954 );
xor ( n59413 , n59412 , n58971 );
and ( n59414 , n59410 , n59413 );
and ( n59415 , n59408 , n59413 );
or ( n59416 , n59411 , n59414 , n59415 );
xor ( n59417 , n58771 , n58790 );
xor ( n59418 , n59417 , n58812 );
and ( n59419 , n59416 , n59418 );
xor ( n59420 , n58821 , n58828 );
xor ( n59421 , n59420 , n58851 );
and ( n59422 , n59418 , n59421 );
and ( n59423 , n59416 , n59421 );
or ( n59424 , n59419 , n59422 , n59423 );
and ( n59425 , n59406 , n59424 );
xor ( n59426 , n58890 , n58921 );
xor ( n59427 , n59426 , n58974 );
xor ( n59428 , n59005 , n59015 );
xor ( n59429 , n59428 , n59018 );
and ( n59430 , n59427 , n59429 );
xor ( n59431 , n59024 , n59026 );
xor ( n59432 , n59431 , n59029 );
and ( n59433 , n59429 , n59432 );
and ( n59434 , n59427 , n59432 );
or ( n59435 , n59430 , n59433 , n59434 );
and ( n59436 , n59424 , n59435 );
and ( n59437 , n59406 , n59435 );
or ( n59438 , n59425 , n59436 , n59437 );
and ( n59439 , n59192 , n59438 );
and ( n59440 , n59110 , n59438 );
or ( n59441 , n59193 , n59439 , n59440 );
xor ( n59442 , n58770 , n58815 );
xor ( n59443 , n59442 , n58854 );
xor ( n59444 , n58977 , n59021 );
xor ( n59445 , n59444 , n59032 );
and ( n59446 , n59443 , n59445 );
xor ( n59447 , n59045 , n59047 );
xor ( n59448 , n59447 , n59050 );
and ( n59449 , n59445 , n59448 );
and ( n59450 , n59443 , n59448 );
or ( n59451 , n59446 , n59449 , n59450 );
xor ( n59452 , n58765 , n58767 );
xor ( n59453 , n59452 , n58857 );
and ( n59454 , n59451 , n59453 );
xor ( n59455 , n59035 , n59053 );
xor ( n59456 , n59455 , n59064 );
and ( n59457 , n59453 , n59456 );
and ( n59458 , n59451 , n59456 );
or ( n59459 , n59454 , n59457 , n59458 );
and ( n59460 , n59441 , n59459 );
xor ( n59461 , n58860 , n59067 );
xor ( n59462 , n59461 , n59078 );
and ( n59463 , n59459 , n59462 );
and ( n59464 , n59441 , n59462 );
or ( n59465 , n59460 , n59463 , n59464 );
and ( n59466 , n59107 , n59465 );
and ( n59467 , n59105 , n59465 );
or ( n59468 , n59108 , n59466 , n59467 );
and ( n59469 , n59103 , n59468 );
xor ( n59470 , n58758 , n58760 );
xor ( n59471 , n59470 , n59095 );
and ( n59472 , n59468 , n59471 );
and ( n59473 , n59103 , n59471 );
or ( n59474 , n59469 , n59472 , n59473 );
and ( n59475 , n59100 , n59474 );
and ( n59476 , n59098 , n59474 );
or ( n59477 , n59101 , n59475 , n59476 );
and ( n59478 , n58700 , n59477 );
xor ( n59479 , n58700 , n59477 );
xor ( n59480 , n59098 , n59100 );
xor ( n59481 , n59480 , n59474 );
xor ( n59482 , n58763 , n59081 );
xor ( n59483 , n59482 , n59092 );
xor ( n59484 , n59084 , n59086 );
xor ( n59485 , n59484 , n59089 );
xor ( n59486 , n59070 , n59072 );
xor ( n59487 , n59486 , n59075 );
xor ( n59488 , n59056 , n59058 );
xor ( n59489 , n59488 , n59061 );
xor ( n59490 , n59037 , n59039 );
xor ( n59491 , n59490 , n59042 );
xor ( n59492 , n58993 , n58999 );
xor ( n59493 , n59492 , n59002 );
xor ( n59494 , n59007 , n59009 );
xor ( n59495 , n59494 , n59012 );
and ( n59496 , n59493 , n59495 );
xor ( n59497 , n59122 , n59123 );
and ( n59498 , n59495 , n59497 );
and ( n59499 , n59493 , n59497 );
or ( n59500 , n59496 , n59498 , n59499 );
and ( n59501 , n59491 , n59500 );
xnor ( n59502 , n59149 , n59153 );
and ( n59503 , n58915 , n58444 );
not ( n59504 , n59503 );
xor ( n59505 , n59137 , n59141 );
xor ( n59506 , n59505 , n59146 );
and ( n59507 , n59504 , n59506 );
buf ( n59508 , n59507 );
and ( n59509 , n59502 , n59508 );
xor ( n59510 , n59197 , n59201 );
xor ( n59511 , n59510 , n58865 );
xor ( n59512 , n59209 , n59210 );
xor ( n59513 , n59512 , n59213 );
and ( n59514 , n59511 , n59513 );
xnor ( n59515 , n59226 , n59230 );
and ( n59516 , n59513 , n59515 );
and ( n59517 , n59511 , n59515 );
or ( n59518 , n59514 , n59516 , n59517 );
and ( n59519 , n59508 , n59518 );
and ( n59520 , n59502 , n59518 );
or ( n59521 , n59509 , n59519 , n59520 );
xnor ( n59522 , n59235 , n59239 );
xnor ( n59523 , n59245 , n59249 );
and ( n59524 , n59522 , n59523 );
xor ( n59525 , n59258 , n59262 );
and ( n59526 , n59523 , n59525 );
and ( n59527 , n59522 , n59525 );
or ( n59528 , n59524 , n59526 , n59527 );
and ( n59529 , n47474 , n52269 );
and ( n59530 , n47351 , n52267 );
nor ( n59531 , n59529 , n59530 );
xnor ( n59532 , n59531 , n52008 );
and ( n59533 , n47778 , n51750 );
and ( n59534 , n47647 , n51748 );
nor ( n59535 , n59533 , n59534 );
xnor ( n59536 , n59535 , n51520 );
and ( n59537 , n59532 , n59536 );
and ( n59538 , n48384 , n50783 );
and ( n59539 , n48272 , n50781 );
nor ( n59540 , n59538 , n59539 );
xnor ( n59541 , n59540 , n50557 );
and ( n59542 , n59536 , n59541 );
and ( n59543 , n59532 , n59541 );
or ( n59544 , n59537 , n59542 , n59543 );
and ( n59545 , n50726 , n48394 );
and ( n59546 , n50625 , n48392 );
nor ( n59547 , n59545 , n59546 );
xnor ( n59548 , n59547 , n48220 );
and ( n59549 , n53328 , n46911 );
and ( n59550 , n53041 , n46909 );
nor ( n59551 , n59549 , n59550 );
xnor ( n59552 , n59551 , n46802 );
and ( n59553 , n59548 , n59552 );
and ( n59554 , n53922 , n46712 );
and ( n59555 , n53639 , n46710 );
nor ( n59556 , n59554 , n59555 );
xnor ( n59557 , n59556 , n46587 );
and ( n59558 , n59552 , n59557 );
and ( n59559 , n59548 , n59557 );
or ( n59560 , n59553 , n59558 , n59559 );
and ( n59561 , n59544 , n59560 );
and ( n59562 , n48709 , n50338 );
and ( n59563 , n48632 , n50336 );
nor ( n59564 , n59562 , n59563 );
xnor ( n59565 , n59564 , n50111 );
and ( n59566 , n49115 , n49896 );
and ( n59567 , n48988 , n49894 );
nor ( n59568 , n59566 , n59567 );
xnor ( n59569 , n59568 , n49711 );
or ( n59570 , n59565 , n59569 );
and ( n59571 , n59560 , n59570 );
and ( n59572 , n59544 , n59570 );
or ( n59573 , n59561 , n59571 , n59572 );
and ( n59574 , n59528 , n59573 );
and ( n59575 , n46530 , n54535 );
and ( n59576 , n46445 , n54533 );
nor ( n59577 , n59575 , n59576 );
xnor ( n59578 , n59577 , n54237 );
and ( n59579 , n46750 , n53928 );
and ( n59580 , n46577 , n53926 );
nor ( n59581 , n59579 , n59580 );
xnor ( n59582 , n59581 , n53652 );
or ( n59583 , n59578 , n59582 );
and ( n59584 , n55143 , n46306 );
and ( n59585 , n54942 , n46304 );
nor ( n59586 , n59584 , n59585 );
xnor ( n59587 , n59586 , n46228 );
and ( n59588 , n56388 , n45990 );
and ( n59589 , n56255 , n45988 );
nor ( n59590 , n59588 , n59589 );
xnor ( n59591 , n59590 , n45939 );
or ( n59592 , n59587 , n59591 );
and ( n59593 , n59583 , n59592 );
and ( n59594 , n51298 , n48042 );
and ( n59595 , n51077 , n48040 );
nor ( n59596 , n59594 , n59595 );
xnor ( n59597 , n59596 , n47921 );
and ( n59598 , n52790 , n47178 );
and ( n59599 , n52612 , n47176 );
nor ( n59600 , n59598 , n59599 );
xnor ( n59601 , n59600 , n47039 );
and ( n59602 , n59597 , n59601 );
and ( n59603 , n59592 , n59602 );
and ( n59604 , n59583 , n59602 );
or ( n59605 , n59593 , n59603 , n59604 );
and ( n59606 , n59573 , n59605 );
and ( n59607 , n59528 , n59605 );
or ( n59608 , n59574 , n59606 , n59607 );
and ( n59609 , n59521 , n59608 );
buf ( n59610 , n20199 );
buf ( n59611 , n59610 );
and ( n59612 , n57948 , n59611 );
not ( n59613 , n59612 );
buf ( n59614 , n20199 );
buf ( n59615 , n59614 );
and ( n59616 , n59615 , n58294 );
not ( n59617 , n59616 );
and ( n59618 , n59613 , n59617 );
and ( n59619 , n58292 , n59207 );
not ( n59620 , n59619 );
and ( n59621 , n59365 , n58444 );
not ( n59622 , n59621 );
and ( n59623 , n59620 , n59622 );
and ( n59624 , n59618 , n59623 );
and ( n59625 , n58628 , n58911 );
not ( n59626 , n59625 );
and ( n59627 , n58915 , n58542 );
not ( n59628 , n59627 );
and ( n59629 , n59626 , n59628 );
and ( n59630 , n59623 , n59629 );
and ( n59631 , n59618 , n59629 );
or ( n59632 , n59624 , n59630 , n59631 );
and ( n59633 , n45907 , n57187 );
and ( n59634 , n45843 , n57184 );
nor ( n59635 , n59633 , n59634 );
xnor ( n59636 , n59635 , n56175 );
and ( n59637 , n46041 , n56503 );
and ( n59638 , n45963 , n56501 );
nor ( n59639 , n59637 , n59638 );
xnor ( n59640 , n59639 , n56178 );
and ( n59641 , n59636 , n59640 );
and ( n59642 , n46169 , n55851 );
and ( n59643 , n46100 , n55849 );
nor ( n59644 , n59642 , n59643 );
xnor ( n59645 , n59644 , n55506 );
and ( n59646 , n59640 , n59645 );
and ( n59647 , n59636 , n59645 );
or ( n59648 , n59641 , n59646 , n59647 );
and ( n59649 , n46345 , n55159 );
and ( n59650 , n46264 , n55157 );
nor ( n59651 , n59649 , n59650 );
xnor ( n59652 , n59651 , n54864 );
and ( n59653 , n46969 , n53357 );
and ( n59654 , n46843 , n53355 );
nor ( n59655 , n59653 , n59654 );
xnor ( n59656 , n59655 , n53060 );
and ( n59657 , n59652 , n59656 );
and ( n59658 , n47216 , n52799 );
and ( n59659 , n47090 , n52797 );
nor ( n59660 , n59658 , n59659 );
xnor ( n59661 , n59660 , n52538 );
and ( n59662 , n59656 , n59661 );
and ( n59663 , n59652 , n59661 );
or ( n59664 , n59657 , n59662 , n59663 );
and ( n59665 , n59648 , n59664 );
and ( n59666 , n48108 , n51221 );
and ( n59667 , n47962 , n51219 );
nor ( n59668 , n59666 , n59667 );
xnor ( n59669 , n59668 , n51000 );
and ( n59670 , n49570 , n49513 );
and ( n59671 , n49374 , n49511 );
nor ( n59672 , n59670 , n59671 );
xnor ( n59673 , n59672 , n49310 );
and ( n59674 , n59669 , n59673 );
and ( n59675 , n49976 , n49121 );
and ( n59676 , n49781 , n49119 );
nor ( n59677 , n59675 , n59676 );
xnor ( n59678 , n59677 , n48932 );
and ( n59679 , n59673 , n59678 );
and ( n59680 , n59669 , n59678 );
or ( n59681 , n59674 , n59679 , n59680 );
and ( n59682 , n59664 , n59681 );
and ( n59683 , n59648 , n59681 );
or ( n59684 , n59665 , n59682 , n59683 );
and ( n59685 , n59632 , n59684 );
and ( n59686 , n50404 , n48740 );
and ( n59687 , n50195 , n48738 );
nor ( n59688 , n59686 , n59687 );
xnor ( n59689 , n59688 , n48571 );
and ( n59690 , n51734 , n47734 );
and ( n59691 , n51510 , n47732 );
nor ( n59692 , n59690 , n59691 );
xnor ( n59693 , n59692 , n47606 );
and ( n59694 , n59689 , n59693 );
and ( n59695 , n52332 , n47429 );
and ( n59696 , n52082 , n47427 );
nor ( n59697 , n59695 , n59696 );
xnor ( n59698 , n59697 , n47309 );
and ( n59699 , n59693 , n59698 );
and ( n59700 , n59689 , n59698 );
or ( n59701 , n59694 , n59699 , n59700 );
and ( n59702 , n54604 , n46496 );
and ( n59703 , n54227 , n46494 );
nor ( n59704 , n59702 , n59703 );
xnor ( n59705 , n59704 , n46402 );
and ( n59706 , n55756 , n46135 );
and ( n59707 , n55497 , n46133 );
nor ( n59708 , n59706 , n59707 );
xnor ( n59709 , n59708 , n46067 );
and ( n59710 , n59705 , n59709 );
and ( n59711 , n57063 , n45886 );
and ( n59712 , n56915 , n45884 );
nor ( n59713 , n59711 , n59712 );
xnor ( n59714 , n59713 , n45824 );
and ( n59715 , n59709 , n59714 );
and ( n59716 , n59705 , n59714 );
or ( n59717 , n59710 , n59715 , n59716 );
and ( n59718 , n59701 , n59717 );
and ( n59719 , n57063 , n45884 );
not ( n59720 , n59719 );
and ( n59721 , n59720 , n45824 );
xor ( n59722 , n39401 , n45574 );
buf ( n59723 , n59722 );
buf ( n59724 , n59723 );
buf ( n59725 , n59724 );
and ( n59726 , n59721 , n59725 );
buf ( n59727 , n59726 );
and ( n59728 , n59717 , n59727 );
and ( n59729 , n59701 , n59727 );
or ( n59730 , n59718 , n59728 , n59729 );
and ( n59731 , n59684 , n59730 );
and ( n59732 , n59632 , n59730 );
or ( n59733 , n59685 , n59731 , n59732 );
and ( n59734 , n59608 , n59733 );
and ( n59735 , n59521 , n59733 );
or ( n59736 , n59609 , n59734 , n59735 );
and ( n59737 , n59500 , n59736 );
and ( n59738 , n59491 , n59736 );
or ( n59739 , n59501 , n59737 , n59738 );
and ( n59740 , n59489 , n59739 );
xor ( n59741 , n59267 , n59271 );
xor ( n59742 , n59741 , n59276 );
xor ( n59743 , n59284 , n59288 );
xor ( n59744 , n59743 , n59293 );
and ( n59745 , n59742 , n59744 );
xor ( n59746 , n59306 , n59310 );
xor ( n59747 , n59746 , n59315 );
and ( n59748 , n59744 , n59747 );
and ( n59749 , n59742 , n59747 );
or ( n59750 , n59745 , n59748 , n59749 );
xor ( n59751 , n59322 , n59326 );
xor ( n59752 , n59751 , n59331 );
xor ( n59753 , n59339 , n59343 );
xor ( n59754 , n59753 , n59348 );
and ( n59755 , n59752 , n59754 );
xor ( n59756 , n59358 , n59362 );
xor ( n59757 , n59756 , n59367 );
and ( n59758 , n59754 , n59757 );
and ( n59759 , n59752 , n59757 );
or ( n59760 , n59755 , n59758 , n59759 );
and ( n59761 , n59750 , n59760 );
xor ( n59762 , n59160 , n59162 );
xor ( n59763 , n59762 , n59165 );
and ( n59764 , n59760 , n59763 );
and ( n59765 , n59750 , n59763 );
or ( n59766 , n59761 , n59764 , n59765 );
xor ( n59767 , n59169 , n59170 );
xor ( n59768 , n59767 , n59172 );
xor ( n59769 , n59177 , n59178 );
xor ( n59770 , n59769 , n59180 );
and ( n59771 , n59768 , n59770 );
xor ( n59772 , n59205 , n59216 );
xor ( n59773 , n59772 , n59219 );
and ( n59774 , n59770 , n59773 );
and ( n59775 , n59768 , n59773 );
or ( n59776 , n59771 , n59774 , n59775 );
and ( n59777 , n59766 , n59776 );
xor ( n59778 , n59231 , n59240 );
xor ( n59779 , n59778 , n59250 );
xor ( n59780 , n59263 , n59279 );
xor ( n59781 , n59780 , n59296 );
and ( n59782 , n59779 , n59781 );
xor ( n59783 , n59318 , n59334 );
xor ( n59784 , n59783 , n59351 );
and ( n59785 , n59781 , n59784 );
and ( n59786 , n59779 , n59784 );
or ( n59787 , n59782 , n59785 , n59786 );
and ( n59788 , n59776 , n59787 );
and ( n59789 , n59766 , n59787 );
or ( n59790 , n59777 , n59788 , n59789 );
xor ( n59791 , n59131 , n59132 );
xor ( n59792 , n59791 , n59154 );
xor ( n59793 , n59168 , n59175 );
xor ( n59794 , n59793 , n59183 );
and ( n59795 , n59792 , n59794 );
xor ( n59796 , n59222 , n59253 );
xor ( n59797 , n59796 , n59299 );
and ( n59798 , n59794 , n59797 );
and ( n59799 , n59792 , n59797 );
or ( n59800 , n59795 , n59798 , n59799 );
and ( n59801 , n59790 , n59800 );
xor ( n59802 , n59354 , n59378 );
xor ( n59803 , n59802 , n59389 );
xor ( n59804 , n59395 , n59397 );
xor ( n59805 , n59804 , n59400 );
and ( n59806 , n59803 , n59805 );
xor ( n59807 , n59408 , n59410 );
xor ( n59808 , n59807 , n59413 );
and ( n59809 , n59805 , n59808 );
and ( n59810 , n59803 , n59808 );
or ( n59811 , n59806 , n59809 , n59810 );
and ( n59812 , n59800 , n59811 );
and ( n59813 , n59790 , n59811 );
or ( n59814 , n59801 , n59812 , n59813 );
and ( n59815 , n59739 , n59814 );
and ( n59816 , n59489 , n59814 );
or ( n59817 , n59740 , n59815 , n59816 );
and ( n59818 , n59487 , n59817 );
xor ( n59819 , n59114 , n59116 );
xor ( n59820 , n59819 , n59124 );
xor ( n59821 , n59129 , n59157 );
xor ( n59822 , n59821 , n59186 );
and ( n59823 , n59820 , n59822 );
xor ( n59824 , n59302 , n59392 );
xor ( n59825 , n59824 , n59403 );
and ( n59826 , n59822 , n59825 );
and ( n59827 , n59820 , n59825 );
or ( n59828 , n59823 , n59826 , n59827 );
xor ( n59829 , n59112 , n59127 );
xor ( n59830 , n59829 , n59189 );
and ( n59831 , n59828 , n59830 );
xor ( n59832 , n59406 , n59424 );
xor ( n59833 , n59832 , n59435 );
and ( n59834 , n59830 , n59833 );
and ( n59835 , n59828 , n59833 );
or ( n59836 , n59831 , n59834 , n59835 );
and ( n59837 , n59817 , n59836 );
and ( n59838 , n59487 , n59836 );
or ( n59839 , n59818 , n59837 , n59838 );
and ( n59840 , n59485 , n59839 );
xor ( n59841 , n59441 , n59459 );
xor ( n59842 , n59841 , n59462 );
and ( n59843 , n59839 , n59842 );
and ( n59844 , n59485 , n59842 );
or ( n59845 , n59840 , n59843 , n59844 );
and ( n59846 , n59483 , n59845 );
xor ( n59847 , n59105 , n59107 );
xor ( n59848 , n59847 , n59465 );
and ( n59849 , n59845 , n59848 );
and ( n59850 , n59483 , n59848 );
or ( n59851 , n59846 , n59849 , n59850 );
xor ( n59852 , n59103 , n59468 );
xor ( n59853 , n59852 , n59471 );
and ( n59854 , n59851 , n59853 );
xor ( n59855 , n59483 , n59845 );
xor ( n59856 , n59855 , n59848 );
xor ( n59857 , n59110 , n59192 );
xor ( n59858 , n59857 , n59438 );
xor ( n59859 , n59451 , n59453 );
xor ( n59860 , n59859 , n59456 );
and ( n59861 , n59858 , n59860 );
xor ( n59862 , n59443 , n59445 );
xor ( n59863 , n59862 , n59448 );
xor ( n59864 , n59416 , n59418 );
xor ( n59865 , n59864 , n59421 );
xor ( n59866 , n59427 , n59429 );
xor ( n59867 , n59866 , n59432 );
and ( n59868 , n59865 , n59867 );
xor ( n59869 , n59370 , n59372 );
xor ( n59870 , n59869 , n59375 );
xor ( n59871 , n59381 , n59383 );
xor ( n59872 , n59871 , n59386 );
and ( n59873 , n59870 , n59872 );
and ( n59874 , n46843 , n53928 );
and ( n59875 , n46750 , n53926 );
nor ( n59876 , n59874 , n59875 );
xnor ( n59877 , n59876 , n53652 );
and ( n59878 , n47090 , n53357 );
and ( n59879 , n46969 , n53355 );
nor ( n59880 , n59878 , n59879 );
xnor ( n59881 , n59880 , n53060 );
and ( n59882 , n59877 , n59881 );
and ( n59883 , n47962 , n51750 );
and ( n59884 , n47778 , n51748 );
nor ( n59885 , n59883 , n59884 );
xnor ( n59886 , n59885 , n51520 );
and ( n59887 , n59881 , n59886 );
and ( n59888 , n59877 , n59886 );
or ( n59889 , n59882 , n59887 , n59888 );
and ( n59890 , n46445 , n55159 );
and ( n59891 , n46345 , n55157 );
nor ( n59892 , n59890 , n59891 );
xnor ( n59893 , n59892 , n54864 );
and ( n59894 , n47351 , n52799 );
and ( n59895 , n47216 , n52797 );
nor ( n59896 , n59894 , n59895 );
xnor ( n59897 , n59896 , n52538 );
and ( n59898 , n59893 , n59897 );
and ( n59899 , n47647 , n52269 );
and ( n59900 , n47474 , n52267 );
nor ( n59901 , n59899 , n59900 );
xnor ( n59902 , n59901 , n52008 );
and ( n59903 , n59897 , n59902 );
and ( n59904 , n59893 , n59902 );
or ( n59905 , n59898 , n59903 , n59904 );
or ( n59906 , n59889 , n59905 );
buf ( n59907 , n20202 );
buf ( n59908 , n59907 );
and ( n59909 , n59908 , n58294 );
not ( n59910 , n59909 );
and ( n59911 , n59615 , n58444 );
not ( n59912 , n59911 );
and ( n59913 , n59910 , n59912 );
and ( n59914 , n59365 , n58542 );
not ( n59915 , n59914 );
and ( n59916 , n59912 , n59915 );
and ( n59917 , n59910 , n59915 );
or ( n59918 , n59913 , n59916 , n59917 );
buf ( n59919 , n20202 );
buf ( n59920 , n59919 );
and ( n59921 , n57948 , n59920 );
not ( n59922 , n59921 );
and ( n59923 , n58292 , n59611 );
not ( n59924 , n59923 );
and ( n59925 , n59922 , n59924 );
and ( n59926 , n58628 , n59207 );
not ( n59927 , n59926 );
and ( n59928 , n59924 , n59927 );
and ( n59929 , n59922 , n59927 );
or ( n59930 , n59925 , n59928 , n59929 );
and ( n59931 , n59918 , n59930 );
and ( n59932 , n59906 , n59931 );
xor ( n59933 , n59532 , n59536 );
xor ( n59934 , n59933 , n59541 );
xor ( n59935 , n59548 , n59552 );
xor ( n59936 , n59935 , n59557 );
and ( n59937 , n59934 , n59936 );
xnor ( n59938 , n59565 , n59569 );
and ( n59939 , n59936 , n59938 );
and ( n59940 , n59934 , n59938 );
or ( n59941 , n59937 , n59939 , n59940 );
and ( n59942 , n59931 , n59941 );
and ( n59943 , n59906 , n59941 );
or ( n59944 , n59932 , n59942 , n59943 );
and ( n59945 , n59872 , n59944 );
and ( n59946 , n59870 , n59944 );
or ( n59947 , n59873 , n59945 , n59946 );
xnor ( n59948 , n59578 , n59582 );
xnor ( n59949 , n59587 , n59591 );
and ( n59950 , n59948 , n59949 );
xor ( n59951 , n59597 , n59601 );
and ( n59952 , n59949 , n59951 );
and ( n59953 , n59948 , n59951 );
or ( n59954 , n59950 , n59952 , n59953 );
xor ( n59955 , n59613 , n59617 );
xor ( n59956 , n59620 , n59622 );
and ( n59957 , n59955 , n59956 );
xor ( n59958 , n59626 , n59628 );
and ( n59959 , n59956 , n59958 );
and ( n59960 , n59955 , n59958 );
or ( n59961 , n59957 , n59959 , n59960 );
and ( n59962 , n59954 , n59961 );
and ( n59963 , n51077 , n48394 );
and ( n59964 , n50726 , n48392 );
nor ( n59965 , n59963 , n59964 );
xnor ( n59966 , n59965 , n48220 );
and ( n59967 , n53041 , n47178 );
and ( n59968 , n52790 , n47176 );
nor ( n59969 , n59967 , n59968 );
xnor ( n59970 , n59969 , n47039 );
and ( n59971 , n59966 , n59970 );
and ( n59972 , n54227 , n46712 );
and ( n59973 , n53922 , n46710 );
nor ( n59974 , n59972 , n59973 );
xnor ( n59975 , n59974 , n46587 );
and ( n59976 , n59970 , n59975 );
and ( n59977 , n59966 , n59975 );
or ( n59978 , n59971 , n59976 , n59977 );
and ( n59979 , n46264 , n55851 );
and ( n59980 , n46169 , n55849 );
nor ( n59981 , n59979 , n59980 );
xnor ( n59982 , n59981 , n55506 );
and ( n59983 , n48988 , n50338 );
and ( n59984 , n48709 , n50336 );
nor ( n59985 , n59983 , n59984 );
xnor ( n59986 , n59985 , n50111 );
and ( n59987 , n59982 , n59986 );
and ( n59988 , n49374 , n49896 );
and ( n59989 , n49115 , n49894 );
nor ( n59990 , n59988 , n59989 );
xnor ( n59991 , n59990 , n49711 );
and ( n59992 , n59986 , n59991 );
and ( n59993 , n59982 , n59991 );
or ( n59994 , n59987 , n59992 , n59993 );
and ( n59995 , n59978 , n59994 );
and ( n59996 , n50625 , n48740 );
and ( n59997 , n50404 , n48738 );
nor ( n59998 , n59996 , n59997 );
xnor ( n59999 , n59998 , n48571 );
and ( n60000 , n52082 , n47734 );
and ( n60001 , n51734 , n47732 );
nor ( n60002 , n60000 , n60001 );
xnor ( n60003 , n60002 , n47606 );
or ( n60004 , n59999 , n60003 );
and ( n60005 , n59994 , n60004 );
and ( n60006 , n59978 , n60004 );
or ( n60007 , n59995 , n60005 , n60006 );
and ( n60008 , n59961 , n60007 );
and ( n60009 , n59954 , n60007 );
or ( n60010 , n59962 , n60008 , n60009 );
and ( n60011 , n48272 , n51221 );
and ( n60012 , n48108 , n51219 );
nor ( n60013 , n60011 , n60012 );
xnor ( n60014 , n60013 , n51000 );
and ( n60015 , n48632 , n50783 );
and ( n60016 , n48384 , n50781 );
nor ( n60017 , n60015 , n60016 );
xnor ( n60018 , n60017 , n50557 );
or ( n60019 , n60014 , n60018 );
and ( n60020 , n56255 , n46135 );
and ( n60021 , n55756 , n46133 );
nor ( n60022 , n60020 , n60021 );
xnor ( n60023 , n60022 , n46067 );
and ( n60024 , n56915 , n45990 );
and ( n60025 , n56388 , n45988 );
nor ( n60026 , n60024 , n60025 );
xnor ( n60027 , n60026 , n45939 );
or ( n60028 , n60023 , n60027 );
and ( n60029 , n60019 , n60028 );
and ( n60030 , n53639 , n46911 );
and ( n60031 , n53328 , n46909 );
nor ( n60032 , n60030 , n60031 );
xnor ( n60033 , n60032 , n46802 );
and ( n60034 , n60033 , n59719 );
and ( n60035 , n60028 , n60034 );
and ( n60036 , n60019 , n60034 );
or ( n60037 , n60029 , n60035 , n60036 );
and ( n60038 , n45963 , n57187 );
and ( n60039 , n45907 , n57184 );
nor ( n60040 , n60038 , n60039 );
xnor ( n60041 , n60040 , n56175 );
and ( n60042 , n46100 , n56503 );
and ( n60043 , n46041 , n56501 );
nor ( n60044 , n60042 , n60043 );
xnor ( n60045 , n60044 , n56178 );
and ( n60046 , n60041 , n60045 );
and ( n60047 , n46577 , n54535 );
and ( n60048 , n46530 , n54533 );
nor ( n60049 , n60047 , n60048 );
xnor ( n60050 , n60049 , n54237 );
and ( n60051 , n60045 , n60050 );
and ( n60052 , n60041 , n60050 );
or ( n60053 , n60046 , n60051 , n60052 );
and ( n60054 , n49781 , n49513 );
and ( n60055 , n49570 , n49511 );
nor ( n60056 , n60054 , n60055 );
xnor ( n60057 , n60056 , n49310 );
and ( n60058 , n50195 , n49121 );
and ( n60059 , n49976 , n49119 );
nor ( n60060 , n60058 , n60059 );
xnor ( n60061 , n60060 , n48932 );
and ( n60062 , n60057 , n60061 );
and ( n60063 , n51510 , n48042 );
and ( n60064 , n51298 , n48040 );
nor ( n60065 , n60063 , n60064 );
xnor ( n60066 , n60065 , n47921 );
and ( n60067 , n60061 , n60066 );
and ( n60068 , n60057 , n60066 );
or ( n60069 , n60062 , n60067 , n60068 );
and ( n60070 , n60053 , n60069 );
and ( n60071 , n52612 , n47429 );
and ( n60072 , n52332 , n47427 );
nor ( n60073 , n60071 , n60072 );
xnor ( n60074 , n60073 , n47309 );
and ( n60075 , n54942 , n46496 );
and ( n60076 , n54604 , n46494 );
nor ( n60077 , n60075 , n60076 );
xnor ( n60078 , n60077 , n46402 );
and ( n60079 , n60074 , n60078 );
and ( n60080 , n55497 , n46306 );
and ( n60081 , n55143 , n46304 );
nor ( n60082 , n60080 , n60081 );
xnor ( n60083 , n60082 , n46228 );
and ( n60084 , n60078 , n60083 );
and ( n60085 , n60074 , n60083 );
or ( n60086 , n60079 , n60084 , n60085 );
and ( n60087 , n60069 , n60086 );
and ( n60088 , n60053 , n60086 );
or ( n60089 , n60070 , n60087 , n60088 );
and ( n60090 , n60037 , n60089 );
xor ( n60091 , n39404 , n45572 );
buf ( n60092 , n60091 );
buf ( n60093 , n60092 );
buf ( n60094 , n60093 );
buf ( n60095 , n58915 );
not ( n60096 , n60095 );
and ( n60097 , n60094 , n60096 );
buf ( n60098 , n60097 );
xor ( n60099 , n59636 , n59640 );
xor ( n60100 , n60099 , n59645 );
and ( n60101 , n60098 , n60100 );
xor ( n60102 , n59652 , n59656 );
xor ( n60103 , n60102 , n59661 );
and ( n60104 , n60100 , n60103 );
and ( n60105 , n60098 , n60103 );
or ( n60106 , n60101 , n60104 , n60105 );
and ( n60107 , n60089 , n60106 );
and ( n60108 , n60037 , n60106 );
or ( n60109 , n60090 , n60107 , n60108 );
and ( n60110 , n60010 , n60109 );
xor ( n60111 , n59669 , n59673 );
xor ( n60112 , n60111 , n59678 );
xor ( n60113 , n59689 , n59693 );
xor ( n60114 , n60113 , n59698 );
and ( n60115 , n60112 , n60114 );
xor ( n60116 , n59705 , n59709 );
xor ( n60117 , n60116 , n59714 );
and ( n60118 , n60114 , n60117 );
and ( n60119 , n60112 , n60117 );
or ( n60120 , n60115 , n60118 , n60119 );
buf ( n60121 , n59504 );
xor ( n60122 , n60121 , n59506 );
and ( n60123 , n60120 , n60122 );
xor ( n60124 , n59511 , n59513 );
xor ( n60125 , n60124 , n59515 );
and ( n60126 , n60122 , n60125 );
and ( n60127 , n60120 , n60125 );
or ( n60128 , n60123 , n60126 , n60127 );
and ( n60129 , n60109 , n60128 );
and ( n60130 , n60010 , n60128 );
or ( n60131 , n60110 , n60129 , n60130 );
and ( n60132 , n59947 , n60131 );
xor ( n60133 , n59522 , n59523 );
xor ( n60134 , n60133 , n59525 );
xor ( n60135 , n59544 , n59560 );
xor ( n60136 , n60135 , n59570 );
and ( n60137 , n60134 , n60136 );
xor ( n60138 , n59583 , n59592 );
xor ( n60139 , n60138 , n59602 );
and ( n60140 , n60136 , n60139 );
and ( n60141 , n60134 , n60139 );
or ( n60142 , n60137 , n60140 , n60141 );
xor ( n60143 , n59618 , n59623 );
xor ( n60144 , n60143 , n59629 );
xor ( n60145 , n59648 , n59664 );
xor ( n60146 , n60145 , n59681 );
and ( n60147 , n60144 , n60146 );
xor ( n60148 , n59701 , n59717 );
xor ( n60149 , n60148 , n59727 );
and ( n60150 , n60146 , n60149 );
and ( n60151 , n60144 , n60149 );
or ( n60152 , n60147 , n60150 , n60151 );
and ( n60153 , n60142 , n60152 );
xor ( n60154 , n59502 , n59508 );
xor ( n60155 , n60154 , n59518 );
and ( n60156 , n60152 , n60155 );
and ( n60157 , n60142 , n60155 );
or ( n60158 , n60153 , n60156 , n60157 );
and ( n60159 , n60131 , n60158 );
and ( n60160 , n59947 , n60158 );
or ( n60161 , n60132 , n60159 , n60160 );
and ( n60162 , n59867 , n60161 );
and ( n60163 , n59865 , n60161 );
or ( n60164 , n59868 , n60162 , n60163 );
and ( n60165 , n59863 , n60164 );
xor ( n60166 , n59528 , n59573 );
xor ( n60167 , n60166 , n59605 );
xor ( n60168 , n59632 , n59684 );
xor ( n60169 , n60168 , n59730 );
and ( n60170 , n60167 , n60169 );
xor ( n60171 , n59750 , n59760 );
xor ( n60172 , n60171 , n59763 );
and ( n60173 , n60169 , n60172 );
and ( n60174 , n60167 , n60172 );
or ( n60175 , n60170 , n60173 , n60174 );
xor ( n60176 , n59493 , n59495 );
xor ( n60177 , n60176 , n59497 );
and ( n60178 , n60175 , n60177 );
xor ( n60179 , n59521 , n59608 );
xor ( n60180 , n60179 , n59733 );
and ( n60181 , n60177 , n60180 );
and ( n60182 , n60175 , n60180 );
or ( n60183 , n60178 , n60181 , n60182 );
xor ( n60184 , n59766 , n59776 );
xor ( n60185 , n60184 , n59787 );
xor ( n60186 , n59792 , n59794 );
xor ( n60187 , n60186 , n59797 );
and ( n60188 , n60185 , n60187 );
xor ( n60189 , n59803 , n59805 );
xor ( n60190 , n60189 , n59808 );
and ( n60191 , n60187 , n60190 );
and ( n60192 , n60185 , n60190 );
or ( n60193 , n60188 , n60191 , n60192 );
and ( n60194 , n60183 , n60193 );
xor ( n60195 , n59491 , n59500 );
xor ( n60196 , n60195 , n59736 );
and ( n60197 , n60193 , n60196 );
and ( n60198 , n60183 , n60196 );
or ( n60199 , n60194 , n60197 , n60198 );
and ( n60200 , n60164 , n60199 );
and ( n60201 , n59863 , n60199 );
or ( n60202 , n60165 , n60200 , n60201 );
and ( n60203 , n59860 , n60202 );
and ( n60204 , n59858 , n60202 );
or ( n60205 , n59861 , n60203 , n60204 );
xor ( n60206 , n59485 , n59839 );
xor ( n60207 , n60206 , n59842 );
and ( n60208 , n60205 , n60207 );
xor ( n60209 , n59487 , n59817 );
xor ( n60210 , n60209 , n59836 );
xor ( n60211 , n59489 , n59739 );
xor ( n60212 , n60211 , n59814 );
xor ( n60213 , n59828 , n59830 );
xor ( n60214 , n60213 , n59833 );
and ( n60215 , n60212 , n60214 );
xor ( n60216 , n59790 , n59800 );
xor ( n60217 , n60216 , n59811 );
xor ( n60218 , n59820 , n59822 );
xor ( n60219 , n60218 , n59825 );
and ( n60220 , n60217 , n60219 );
xor ( n60221 , n59768 , n59770 );
xor ( n60222 , n60221 , n59773 );
xor ( n60223 , n59779 , n59781 );
xor ( n60224 , n60223 , n59784 );
and ( n60225 , n60222 , n60224 );
xor ( n60226 , n59742 , n59744 );
xor ( n60227 , n60226 , n59747 );
xor ( n60228 , n59752 , n59754 );
xor ( n60229 , n60228 , n59757 );
and ( n60230 , n60227 , n60229 );
xor ( n60231 , n59721 , n59725 );
buf ( n60232 , n60231 );
xnor ( n60233 , n59889 , n59905 );
and ( n60234 , n60232 , n60233 );
xor ( n60235 , n59918 , n59930 );
and ( n60236 , n60233 , n60235 );
and ( n60237 , n60232 , n60235 );
or ( n60238 , n60234 , n60236 , n60237 );
and ( n60239 , n60229 , n60238 );
and ( n60240 , n60227 , n60238 );
or ( n60241 , n60230 , n60239 , n60240 );
and ( n60242 , n60224 , n60241 );
and ( n60243 , n60222 , n60241 );
or ( n60244 , n60225 , n60242 , n60243 );
and ( n60245 , n59908 , n58444 );
not ( n60246 , n60245 );
and ( n60247 , n59615 , n58542 );
not ( n60248 , n60247 );
and ( n60249 , n60246 , n60248 );
and ( n60250 , n58292 , n59920 );
not ( n60251 , n60250 );
and ( n60252 , n58628 , n59611 );
not ( n60253 , n60252 );
and ( n60254 , n60251 , n60253 );
and ( n60255 , n60249 , n60254 );
xor ( n60256 , n59910 , n59912 );
xor ( n60257 , n60256 , n59915 );
xor ( n60258 , n59922 , n59924 );
xor ( n60259 , n60258 , n59927 );
and ( n60260 , n60257 , n60259 );
and ( n60261 , n60255 , n60260 );
xor ( n60262 , n59966 , n59970 );
xor ( n60263 , n60262 , n59975 );
xor ( n60264 , n59877 , n59881 );
xor ( n60265 , n60264 , n59886 );
and ( n60266 , n60263 , n60265 );
xor ( n60267 , n59893 , n59897 );
xor ( n60268 , n60267 , n59902 );
and ( n60269 , n60265 , n60268 );
and ( n60270 , n60263 , n60268 );
or ( n60271 , n60266 , n60269 , n60270 );
and ( n60272 , n60260 , n60271 );
and ( n60273 , n60255 , n60271 );
or ( n60274 , n60261 , n60272 , n60273 );
xor ( n60275 , n59982 , n59986 );
xor ( n60276 , n60275 , n59991 );
xnor ( n60277 , n59999 , n60003 );
and ( n60278 , n60276 , n60277 );
xnor ( n60279 , n60014 , n60018 );
and ( n60280 , n60277 , n60279 );
and ( n60281 , n60276 , n60279 );
or ( n60282 , n60278 , n60280 , n60281 );
xnor ( n60283 , n60023 , n60027 );
xor ( n60284 , n60033 , n59719 );
and ( n60285 , n60283 , n60284 );
and ( n60286 , n46969 , n53928 );
and ( n60287 , n46843 , n53926 );
nor ( n60288 , n60286 , n60287 );
xnor ( n60289 , n60288 , n53652 );
and ( n60290 , n47216 , n53357 );
and ( n60291 , n47090 , n53355 );
nor ( n60292 , n60290 , n60291 );
xnor ( n60293 , n60292 , n53060 );
and ( n60294 , n60289 , n60293 );
and ( n60295 , n48709 , n50783 );
and ( n60296 , n48632 , n50781 );
nor ( n60297 , n60295 , n60296 );
xnor ( n60298 , n60297 , n50557 );
and ( n60299 , n60293 , n60298 );
and ( n60300 , n60289 , n60298 );
or ( n60301 , n60294 , n60299 , n60300 );
and ( n60302 , n60284 , n60301 );
and ( n60303 , n60283 , n60301 );
or ( n60304 , n60285 , n60302 , n60303 );
and ( n60305 , n60282 , n60304 );
and ( n60306 , n46750 , n54535 );
and ( n60307 , n46577 , n54533 );
nor ( n60308 , n60306 , n60307 );
xnor ( n60309 , n60308 , n54237 );
and ( n60310 , n47778 , n52269 );
and ( n60311 , n47647 , n52267 );
nor ( n60312 , n60310 , n60311 );
xnor ( n60313 , n60312 , n52008 );
and ( n60314 , n60309 , n60313 );
and ( n60315 , n48384 , n51221 );
and ( n60316 , n48272 , n51219 );
nor ( n60317 , n60315 , n60316 );
xnor ( n60318 , n60317 , n51000 );
and ( n60319 , n60313 , n60318 );
and ( n60320 , n60309 , n60318 );
or ( n60321 , n60314 , n60319 , n60320 );
and ( n60322 , n52790 , n47429 );
and ( n60323 , n52612 , n47427 );
nor ( n60324 , n60322 , n60323 );
xnor ( n60325 , n60324 , n47309 );
and ( n60326 , n53328 , n47178 );
and ( n60327 , n53041 , n47176 );
nor ( n60328 , n60326 , n60327 );
xnor ( n60329 , n60328 , n47039 );
and ( n60330 , n60325 , n60329 );
and ( n60331 , n54604 , n46712 );
and ( n60332 , n54227 , n46710 );
nor ( n60333 , n60331 , n60332 );
xnor ( n60334 , n60333 , n46587 );
and ( n60335 , n60329 , n60334 );
and ( n60336 , n60325 , n60334 );
or ( n60337 , n60330 , n60335 , n60336 );
and ( n60338 , n60321 , n60337 );
and ( n60339 , n55756 , n46306 );
and ( n60340 , n55497 , n46304 );
nor ( n60341 , n60339 , n60340 );
xnor ( n60342 , n60341 , n46228 );
and ( n60343 , n56388 , n46135 );
and ( n60344 , n56255 , n46133 );
nor ( n60345 , n60343 , n60344 );
xnor ( n60346 , n60345 , n46067 );
and ( n60347 , n60342 , n60346 );
and ( n60348 , n57063 , n45990 );
and ( n60349 , n56915 , n45988 );
nor ( n60350 , n60348 , n60349 );
xnor ( n60351 , n60350 , n45939 );
and ( n60352 , n60346 , n60351 );
and ( n60353 , n60342 , n60351 );
or ( n60354 , n60347 , n60352 , n60353 );
and ( n60355 , n60337 , n60354 );
and ( n60356 , n60321 , n60354 );
or ( n60357 , n60338 , n60355 , n60356 );
and ( n60358 , n60304 , n60357 );
and ( n60359 , n60282 , n60357 );
or ( n60360 , n60305 , n60358 , n60359 );
and ( n60361 , n60274 , n60360 );
and ( n60362 , n51298 , n48394 );
and ( n60363 , n51077 , n48392 );
nor ( n60364 , n60362 , n60363 );
xnor ( n60365 , n60364 , n48220 );
and ( n60366 , n51734 , n48042 );
and ( n60367 , n51510 , n48040 );
nor ( n60368 , n60366 , n60367 );
xnor ( n60369 , n60368 , n47921 );
and ( n60370 , n60365 , n60369 );
buf ( n60371 , n20205 );
buf ( n60372 , n60371 );
and ( n60373 , n57948 , n60372 );
not ( n60374 , n60373 );
buf ( n60375 , n20205 );
buf ( n60376 , n60375 );
and ( n60377 , n60376 , n58294 );
not ( n60378 , n60377 );
and ( n60379 , n60374 , n60378 );
and ( n60380 , n60370 , n60379 );
and ( n60381 , n58915 , n59207 );
not ( n60382 , n60381 );
and ( n60383 , n59365 , n58911 );
not ( n60384 , n60383 );
and ( n60385 , n60382 , n60384 );
and ( n60386 , n60379 , n60385 );
and ( n60387 , n60370 , n60385 );
or ( n60388 , n60380 , n60386 , n60387 );
and ( n60389 , n46041 , n57187 );
and ( n60390 , n45963 , n57184 );
nor ( n60391 , n60389 , n60390 );
xnor ( n60392 , n60391 , n56175 );
and ( n60393 , n46169 , n56503 );
and ( n60394 , n46100 , n56501 );
nor ( n60395 , n60393 , n60394 );
xnor ( n60396 , n60395 , n56178 );
and ( n60397 , n60392 , n60396 );
and ( n60398 , n46345 , n55851 );
and ( n60399 , n46264 , n55849 );
nor ( n60400 , n60398 , n60399 );
xnor ( n60401 , n60400 , n55506 );
and ( n60402 , n60396 , n60401 );
and ( n60403 , n60392 , n60401 );
or ( n60404 , n60397 , n60402 , n60403 );
and ( n60405 , n46530 , n55159 );
and ( n60406 , n46445 , n55157 );
nor ( n60407 , n60405 , n60406 );
xnor ( n60408 , n60407 , n54864 );
and ( n60409 , n47474 , n52799 );
and ( n60410 , n47351 , n52797 );
nor ( n60411 , n60409 , n60410 );
xnor ( n60412 , n60411 , n52538 );
and ( n60413 , n60408 , n60412 );
and ( n60414 , n48108 , n51750 );
and ( n60415 , n47962 , n51748 );
nor ( n60416 , n60414 , n60415 );
xnor ( n60417 , n60416 , n51520 );
and ( n60418 , n60412 , n60417 );
and ( n60419 , n60408 , n60417 );
or ( n60420 , n60413 , n60418 , n60419 );
and ( n60421 , n60404 , n60420 );
and ( n60422 , n49115 , n50338 );
and ( n60423 , n48988 , n50336 );
nor ( n60424 , n60422 , n60423 );
xnor ( n60425 , n60424 , n50111 );
and ( n60426 , n49570 , n49896 );
and ( n60427 , n49374 , n49894 );
nor ( n60428 , n60426 , n60427 );
xnor ( n60429 , n60428 , n49711 );
and ( n60430 , n60425 , n60429 );
and ( n60431 , n49976 , n49513 );
and ( n60432 , n49781 , n49511 );
nor ( n60433 , n60431 , n60432 );
xnor ( n60434 , n60433 , n49310 );
and ( n60435 , n60429 , n60434 );
and ( n60436 , n60425 , n60434 );
or ( n60437 , n60430 , n60435 , n60436 );
and ( n60438 , n60420 , n60437 );
and ( n60439 , n60404 , n60437 );
or ( n60440 , n60421 , n60438 , n60439 );
and ( n60441 , n60388 , n60440 );
and ( n60442 , n50404 , n49121 );
and ( n60443 , n50195 , n49119 );
nor ( n60444 , n60442 , n60443 );
xnor ( n60445 , n60444 , n48932 );
and ( n60446 , n50726 , n48740 );
and ( n60447 , n50625 , n48738 );
nor ( n60448 , n60446 , n60447 );
xnor ( n60449 , n60448 , n48571 );
and ( n60450 , n60445 , n60449 );
and ( n60451 , n52332 , n47734 );
and ( n60452 , n52082 , n47732 );
nor ( n60453 , n60451 , n60452 );
xnor ( n60454 , n60453 , n47606 );
and ( n60455 , n60449 , n60454 );
and ( n60456 , n60445 , n60454 );
or ( n60457 , n60450 , n60455 , n60456 );
and ( n60458 , n53922 , n46911 );
and ( n60459 , n53639 , n46909 );
nor ( n60460 , n60458 , n60459 );
xnor ( n60461 , n60460 , n46802 );
and ( n60462 , n55143 , n46496 );
and ( n60463 , n54942 , n46494 );
nor ( n60464 , n60462 , n60463 );
xnor ( n60465 , n60464 , n46402 );
and ( n60466 , n60461 , n60465 );
and ( n60467 , n57063 , n45988 );
not ( n60468 , n60467 );
and ( n60469 , n60468 , n45939 );
and ( n60470 , n60465 , n60469 );
and ( n60471 , n60461 , n60469 );
or ( n60472 , n60466 , n60470 , n60471 );
and ( n60473 , n60457 , n60472 );
xor ( n60474 , n60041 , n60045 );
xor ( n60475 , n60474 , n60050 );
and ( n60476 , n60472 , n60475 );
and ( n60477 , n60457 , n60475 );
or ( n60478 , n60473 , n60476 , n60477 );
and ( n60479 , n60440 , n60478 );
and ( n60480 , n60388 , n60478 );
or ( n60481 , n60441 , n60479 , n60480 );
and ( n60482 , n60360 , n60481 );
and ( n60483 , n60274 , n60481 );
or ( n60484 , n60361 , n60482 , n60483 );
xor ( n60485 , n60057 , n60061 );
xor ( n60486 , n60485 , n60066 );
xor ( n60487 , n60074 , n60078 );
xor ( n60488 , n60487 , n60083 );
and ( n60489 , n60486 , n60488 );
xor ( n60490 , n60094 , n60096 );
buf ( n60491 , n60490 );
and ( n60492 , n60488 , n60491 );
and ( n60493 , n60486 , n60491 );
or ( n60494 , n60489 , n60492 , n60493 );
xor ( n60495 , n59934 , n59936 );
xor ( n60496 , n60495 , n59938 );
and ( n60497 , n60494 , n60496 );
xor ( n60498 , n59948 , n59949 );
xor ( n60499 , n60498 , n59951 );
and ( n60500 , n60496 , n60499 );
and ( n60501 , n60494 , n60499 );
or ( n60502 , n60497 , n60500 , n60501 );
xor ( n60503 , n59955 , n59956 );
xor ( n60504 , n60503 , n59958 );
xor ( n60505 , n59978 , n59994 );
xor ( n60506 , n60505 , n60004 );
and ( n60507 , n60504 , n60506 );
xor ( n60508 , n60019 , n60028 );
xor ( n60509 , n60508 , n60034 );
and ( n60510 , n60506 , n60509 );
and ( n60511 , n60504 , n60509 );
or ( n60512 , n60507 , n60510 , n60511 );
and ( n60513 , n60502 , n60512 );
xor ( n60514 , n60053 , n60069 );
xor ( n60515 , n60514 , n60086 );
xor ( n60516 , n60098 , n60100 );
xor ( n60517 , n60516 , n60103 );
and ( n60518 , n60515 , n60517 );
xor ( n60519 , n60112 , n60114 );
xor ( n60520 , n60519 , n60117 );
and ( n60521 , n60517 , n60520 );
and ( n60522 , n60515 , n60520 );
or ( n60523 , n60518 , n60521 , n60522 );
and ( n60524 , n60512 , n60523 );
and ( n60525 , n60502 , n60523 );
or ( n60526 , n60513 , n60524 , n60525 );
and ( n60527 , n60484 , n60526 );
xor ( n60528 , n59906 , n59931 );
xor ( n60529 , n60528 , n59941 );
xor ( n60530 , n59954 , n59961 );
xor ( n60531 , n60530 , n60007 );
and ( n60532 , n60529 , n60531 );
xor ( n60533 , n60037 , n60089 );
xor ( n60534 , n60533 , n60106 );
and ( n60535 , n60531 , n60534 );
and ( n60536 , n60529 , n60534 );
or ( n60537 , n60532 , n60535 , n60536 );
and ( n60538 , n60526 , n60537 );
and ( n60539 , n60484 , n60537 );
or ( n60540 , n60527 , n60538 , n60539 );
and ( n60541 , n60244 , n60540 );
xor ( n60542 , n60120 , n60122 );
xor ( n60543 , n60542 , n60125 );
xor ( n60544 , n60134 , n60136 );
xor ( n60545 , n60544 , n60139 );
and ( n60546 , n60543 , n60545 );
xor ( n60547 , n60144 , n60146 );
xor ( n60548 , n60547 , n60149 );
and ( n60549 , n60545 , n60548 );
and ( n60550 , n60543 , n60548 );
or ( n60551 , n60546 , n60549 , n60550 );
xor ( n60552 , n59870 , n59872 );
xor ( n60553 , n60552 , n59944 );
and ( n60554 , n60551 , n60553 );
xor ( n60555 , n60010 , n60109 );
xor ( n60556 , n60555 , n60128 );
and ( n60557 , n60553 , n60556 );
and ( n60558 , n60551 , n60556 );
or ( n60559 , n60554 , n60557 , n60558 );
and ( n60560 , n60540 , n60559 );
and ( n60561 , n60244 , n60559 );
or ( n60562 , n60541 , n60560 , n60561 );
and ( n60563 , n60219 , n60562 );
and ( n60564 , n60217 , n60562 );
or ( n60565 , n60220 , n60563 , n60564 );
and ( n60566 , n60214 , n60565 );
and ( n60567 , n60212 , n60565 );
or ( n60568 , n60215 , n60566 , n60567 );
and ( n60569 , n60210 , n60568 );
xor ( n60570 , n59858 , n59860 );
xor ( n60571 , n60570 , n60202 );
and ( n60572 , n60568 , n60571 );
and ( n60573 , n60210 , n60571 );
or ( n60574 , n60569 , n60572 , n60573 );
and ( n60575 , n60207 , n60574 );
and ( n60576 , n60205 , n60574 );
or ( n60577 , n60208 , n60575 , n60576 );
and ( n60578 , n59856 , n60577 );
xor ( n60579 , n60205 , n60207 );
xor ( n60580 , n60579 , n60574 );
xor ( n60581 , n59947 , n60131 );
xor ( n60582 , n60581 , n60158 );
xor ( n60583 , n60175 , n60177 );
xor ( n60584 , n60583 , n60180 );
and ( n60585 , n60582 , n60584 );
xor ( n60586 , n60185 , n60187 );
xor ( n60587 , n60586 , n60190 );
and ( n60588 , n60584 , n60587 );
and ( n60589 , n60582 , n60587 );
or ( n60590 , n60585 , n60588 , n60589 );
xor ( n60591 , n59865 , n59867 );
xor ( n60592 , n60591 , n60161 );
and ( n60593 , n60590 , n60592 );
xor ( n60594 , n60183 , n60193 );
xor ( n60595 , n60594 , n60196 );
and ( n60596 , n60592 , n60595 );
and ( n60597 , n60590 , n60595 );
or ( n60598 , n60593 , n60596 , n60597 );
xor ( n60599 , n59863 , n60164 );
xor ( n60600 , n60599 , n60199 );
and ( n60601 , n60598 , n60600 );
xor ( n60602 , n60142 , n60152 );
xor ( n60603 , n60602 , n60155 );
xor ( n60604 , n60167 , n60169 );
xor ( n60605 , n60604 , n60172 );
and ( n60606 , n60603 , n60605 );
xor ( n60607 , n60249 , n60254 );
xor ( n60608 , n60257 , n60259 );
and ( n60609 , n60607 , n60608 );
xor ( n60610 , n60246 , n60248 );
xor ( n60611 , n60251 , n60253 );
and ( n60612 , n60610 , n60611 );
and ( n60613 , n60608 , n60612 );
and ( n60614 , n60607 , n60612 );
or ( n60615 , n60609 , n60613 , n60614 );
xor ( n60616 , n39406 , n45571 );
buf ( n60617 , n60616 );
buf ( n60618 , n60617 );
buf ( n60619 , n60618 );
xor ( n60620 , n60289 , n60293 );
xor ( n60621 , n60620 , n60298 );
and ( n60622 , n60619 , n60621 );
buf ( n60623 , n60622 );
xor ( n60624 , n60309 , n60313 );
xor ( n60625 , n60624 , n60318 );
xor ( n60626 , n60325 , n60329 );
xor ( n60627 , n60626 , n60334 );
and ( n60628 , n60625 , n60627 );
xor ( n60629 , n60342 , n60346 );
xor ( n60630 , n60629 , n60351 );
and ( n60631 , n60627 , n60630 );
and ( n60632 , n60625 , n60630 );
or ( n60633 , n60628 , n60631 , n60632 );
and ( n60634 , n60623 , n60633 );
xor ( n60635 , n60365 , n60369 );
xor ( n60636 , n60374 , n60378 );
and ( n60637 , n60635 , n60636 );
xor ( n60638 , n60382 , n60384 );
and ( n60639 , n60636 , n60638 );
and ( n60640 , n60635 , n60638 );
or ( n60641 , n60637 , n60639 , n60640 );
and ( n60642 , n60633 , n60641 );
and ( n60643 , n60623 , n60641 );
or ( n60644 , n60634 , n60642 , n60643 );
and ( n60645 , n60615 , n60644 );
and ( n60646 , n47351 , n53357 );
and ( n60647 , n47216 , n53355 );
nor ( n60648 , n60646 , n60647 );
xnor ( n60649 , n60648 , n53060 );
and ( n60650 , n47962 , n52269 );
and ( n60651 , n47778 , n52267 );
nor ( n60652 , n60650 , n60651 );
xnor ( n60653 , n60652 , n52008 );
and ( n60654 , n60649 , n60653 );
and ( n60655 , n48272 , n51750 );
and ( n60656 , n48108 , n51748 );
nor ( n60657 , n60655 , n60656 );
xnor ( n60658 , n60657 , n51520 );
and ( n60659 , n60653 , n60658 );
and ( n60660 , n60649 , n60658 );
or ( n60661 , n60654 , n60659 , n60660 );
and ( n60662 , n46843 , n54535 );
and ( n60663 , n46750 , n54533 );
nor ( n60664 , n60662 , n60663 );
xnor ( n60665 , n60664 , n54237 );
and ( n60666 , n48632 , n51221 );
and ( n60667 , n48384 , n51219 );
nor ( n60668 , n60666 , n60667 );
xnor ( n60669 , n60668 , n51000 );
and ( n60670 , n60665 , n60669 );
and ( n60671 , n48988 , n50783 );
and ( n60672 , n48709 , n50781 );
nor ( n60673 , n60671 , n60672 );
xnor ( n60674 , n60673 , n50557 );
and ( n60675 , n60669 , n60674 );
and ( n60676 , n60665 , n60674 );
or ( n60677 , n60670 , n60675 , n60676 );
and ( n60678 , n60661 , n60677 );
and ( n60679 , n46264 , n56503 );
and ( n60680 , n46169 , n56501 );
nor ( n60681 , n60679 , n60680 );
xnor ( n60682 , n60681 , n56178 );
and ( n60683 , n46445 , n55851 );
and ( n60684 , n46345 , n55849 );
nor ( n60685 , n60683 , n60684 );
xnor ( n60686 , n60685 , n55506 );
and ( n60687 , n60682 , n60686 );
and ( n60688 , n47090 , n53928 );
and ( n60689 , n46969 , n53926 );
nor ( n60690 , n60688 , n60689 );
xnor ( n60691 , n60690 , n53652 );
and ( n60692 , n60686 , n60691 );
and ( n60693 , n60682 , n60691 );
or ( n60694 , n60687 , n60692 , n60693 );
and ( n60695 , n60677 , n60694 );
and ( n60696 , n60661 , n60694 );
or ( n60697 , n60678 , n60695 , n60696 );
and ( n60698 , n54227 , n46911 );
and ( n60699 , n53922 , n46909 );
nor ( n60700 , n60698 , n60699 );
xnor ( n60701 , n60700 , n46802 );
and ( n60702 , n54942 , n46712 );
and ( n60703 , n54604 , n46710 );
nor ( n60704 , n60702 , n60703 );
xnor ( n60705 , n60704 , n46587 );
and ( n60706 , n60701 , n60705 );
and ( n60707 , n60705 , n60467 );
and ( n60708 , n60701 , n60467 );
or ( n60709 , n60706 , n60707 , n60708 );
buf ( n60710 , n20208 );
buf ( n60711 , n60710 );
and ( n60712 , n57948 , n60711 );
not ( n60713 , n60712 );
and ( n60714 , n58628 , n59920 );
not ( n60715 , n60714 );
and ( n60716 , n60713 , n60715 );
and ( n60717 , n58915 , n59611 );
not ( n60718 , n60717 );
and ( n60719 , n60715 , n60718 );
and ( n60720 , n60713 , n60718 );
or ( n60721 , n60716 , n60719 , n60720 );
and ( n60722 , n60709 , n60721 );
and ( n60723 , n58292 , n60372 );
not ( n60724 , n60723 );
and ( n60725 , n59908 , n58542 );
not ( n60726 , n60725 );
and ( n60727 , n60724 , n60726 );
and ( n60728 , n59615 , n58911 );
not ( n60729 , n60728 );
and ( n60730 , n60726 , n60729 );
and ( n60731 , n60724 , n60729 );
or ( n60732 , n60727 , n60730 , n60731 );
and ( n60733 , n60721 , n60732 );
and ( n60734 , n60709 , n60732 );
or ( n60735 , n60722 , n60733 , n60734 );
and ( n60736 , n60697 , n60735 );
and ( n60737 , n46100 , n57187 );
and ( n60738 , n46041 , n57184 );
nor ( n60739 , n60737 , n60738 );
xnor ( n60740 , n60739 , n56175 );
and ( n60741 , n46577 , n55159 );
and ( n60742 , n46530 , n55157 );
nor ( n60743 , n60741 , n60742 );
xnor ( n60744 , n60743 , n54864 );
and ( n60745 , n60740 , n60744 );
and ( n60746 , n47647 , n52799 );
and ( n60747 , n47474 , n52797 );
nor ( n60748 , n60746 , n60747 );
xnor ( n60749 , n60748 , n52538 );
and ( n60750 , n60744 , n60749 );
and ( n60751 , n60740 , n60749 );
or ( n60752 , n60745 , n60750 , n60751 );
and ( n60753 , n50625 , n49121 );
and ( n60754 , n50404 , n49119 );
nor ( n60755 , n60753 , n60754 );
xnor ( n60756 , n60755 , n48932 );
and ( n60757 , n51077 , n48740 );
and ( n60758 , n50726 , n48738 );
nor ( n60759 , n60757 , n60758 );
xnor ( n60760 , n60759 , n48571 );
and ( n60761 , n60756 , n60760 );
and ( n60762 , n51510 , n48394 );
and ( n60763 , n51298 , n48392 );
nor ( n60764 , n60762 , n60763 );
xnor ( n60765 , n60764 , n48220 );
and ( n60766 , n60760 , n60765 );
and ( n60767 , n60756 , n60765 );
or ( n60768 , n60761 , n60766 , n60767 );
and ( n60769 , n60752 , n60768 );
and ( n60770 , n52082 , n48042 );
and ( n60771 , n51734 , n48040 );
nor ( n60772 , n60770 , n60771 );
xnor ( n60773 , n60772 , n47921 );
and ( n60774 , n52612 , n47734 );
and ( n60775 , n52332 , n47732 );
nor ( n60776 , n60774 , n60775 );
xnor ( n60777 , n60776 , n47606 );
and ( n60778 , n60773 , n60777 );
and ( n60779 , n53041 , n47429 );
and ( n60780 , n52790 , n47427 );
nor ( n60781 , n60779 , n60780 );
xnor ( n60782 , n60781 , n47309 );
and ( n60783 , n60777 , n60782 );
and ( n60784 , n60773 , n60782 );
or ( n60785 , n60778 , n60783 , n60784 );
and ( n60786 , n60768 , n60785 );
and ( n60787 , n60752 , n60785 );
or ( n60788 , n60769 , n60786 , n60787 );
and ( n60789 , n60735 , n60788 );
and ( n60790 , n60697 , n60788 );
or ( n60791 , n60736 , n60789 , n60790 );
and ( n60792 , n60644 , n60791 );
and ( n60793 , n60615 , n60791 );
or ( n60794 , n60645 , n60792 , n60793 );
and ( n60795 , n53639 , n47178 );
and ( n60796 , n53328 , n47176 );
nor ( n60797 , n60795 , n60796 );
xnor ( n60798 , n60797 , n47039 );
and ( n60799 , n55497 , n46496 );
and ( n60800 , n55143 , n46494 );
nor ( n60801 , n60799 , n60800 );
xnor ( n60802 , n60801 , n46402 );
and ( n60803 , n60798 , n60802 );
and ( n60804 , n56255 , n46306 );
and ( n60805 , n55756 , n46304 );
nor ( n60806 , n60804 , n60805 );
xnor ( n60807 , n60806 , n46228 );
and ( n60808 , n60802 , n60807 );
and ( n60809 , n60798 , n60807 );
or ( n60810 , n60803 , n60808 , n60809 );
and ( n60811 , n56915 , n46135 );
and ( n60812 , n56388 , n46133 );
nor ( n60813 , n60811 , n60812 );
xnor ( n60814 , n60813 , n46067 );
xor ( n60815 , n39408 , n45570 );
buf ( n60816 , n60815 );
buf ( n60817 , n60816 );
buf ( n60818 , n60817 );
and ( n60819 , n60814 , n60818 );
buf ( n60820 , n20208 );
buf ( n60821 , n60820 );
and ( n60822 , n60821 , n58294 );
not ( n60823 , n60822 );
and ( n60824 , n60818 , n60823 );
and ( n60825 , n60814 , n60823 );
or ( n60826 , n60819 , n60824 , n60825 );
and ( n60827 , n60810 , n60826 );
xor ( n60828 , n60392 , n60396 );
xor ( n60829 , n60828 , n60401 );
and ( n60830 , n60826 , n60829 );
and ( n60831 , n60810 , n60829 );
or ( n60832 , n60827 , n60830 , n60831 );
xor ( n60833 , n60408 , n60412 );
xor ( n60834 , n60833 , n60417 );
xor ( n60835 , n60425 , n60429 );
xor ( n60836 , n60835 , n60434 );
and ( n60837 , n60834 , n60836 );
xor ( n60838 , n60445 , n60449 );
xor ( n60839 , n60838 , n60454 );
and ( n60840 , n60836 , n60839 );
and ( n60841 , n60834 , n60839 );
or ( n60842 , n60837 , n60840 , n60841 );
and ( n60843 , n60832 , n60842 );
xor ( n60844 , n60263 , n60265 );
xor ( n60845 , n60844 , n60268 );
and ( n60846 , n60842 , n60845 );
and ( n60847 , n60832 , n60845 );
or ( n60848 , n60843 , n60846 , n60847 );
xor ( n60849 , n60276 , n60277 );
xor ( n60850 , n60849 , n60279 );
xor ( n60851 , n60283 , n60284 );
xor ( n60852 , n60851 , n60301 );
and ( n60853 , n60850 , n60852 );
xor ( n60854 , n60321 , n60337 );
xor ( n60855 , n60854 , n60354 );
and ( n60856 , n60852 , n60855 );
and ( n60857 , n60850 , n60855 );
or ( n60858 , n60853 , n60856 , n60857 );
and ( n60859 , n60848 , n60858 );
xor ( n60860 , n60370 , n60379 );
xor ( n60861 , n60860 , n60385 );
xor ( n60862 , n60404 , n60420 );
xor ( n60863 , n60862 , n60437 );
and ( n60864 , n60861 , n60863 );
xor ( n60865 , n60457 , n60472 );
xor ( n60866 , n60865 , n60475 );
and ( n60867 , n60863 , n60866 );
and ( n60868 , n60861 , n60866 );
or ( n60869 , n60864 , n60867 , n60868 );
and ( n60870 , n60858 , n60869 );
and ( n60871 , n60848 , n60869 );
or ( n60872 , n60859 , n60870 , n60871 );
and ( n60873 , n60794 , n60872 );
xor ( n60874 , n60232 , n60233 );
xor ( n60875 , n60874 , n60235 );
xor ( n60876 , n60255 , n60260 );
xor ( n60877 , n60876 , n60271 );
and ( n60878 , n60875 , n60877 );
xor ( n60879 , n60282 , n60304 );
xor ( n60880 , n60879 , n60357 );
and ( n60881 , n60877 , n60880 );
and ( n60882 , n60875 , n60880 );
or ( n60883 , n60878 , n60881 , n60882 );
and ( n60884 , n60872 , n60883 );
and ( n60885 , n60794 , n60883 );
or ( n60886 , n60873 , n60884 , n60885 );
and ( n60887 , n60605 , n60886 );
and ( n60888 , n60603 , n60886 );
or ( n60889 , n60606 , n60887 , n60888 );
xor ( n60890 , n60388 , n60440 );
xor ( n60891 , n60890 , n60478 );
xor ( n60892 , n60494 , n60496 );
xor ( n60893 , n60892 , n60499 );
and ( n60894 , n60891 , n60893 );
xor ( n60895 , n60504 , n60506 );
xor ( n60896 , n60895 , n60509 );
and ( n60897 , n60893 , n60896 );
and ( n60898 , n60891 , n60896 );
or ( n60899 , n60894 , n60897 , n60898 );
xor ( n60900 , n60227 , n60229 );
xor ( n60901 , n60900 , n60238 );
and ( n60902 , n60899 , n60901 );
xor ( n60903 , n60274 , n60360 );
xor ( n60904 , n60903 , n60481 );
and ( n60905 , n60901 , n60904 );
and ( n60906 , n60899 , n60904 );
or ( n60907 , n60902 , n60905 , n60906 );
xor ( n60908 , n60502 , n60512 );
xor ( n60909 , n60908 , n60523 );
xor ( n60910 , n60529 , n60531 );
xor ( n60911 , n60910 , n60534 );
and ( n60912 , n60909 , n60911 );
xor ( n60913 , n60543 , n60545 );
xor ( n60914 , n60913 , n60548 );
and ( n60915 , n60911 , n60914 );
and ( n60916 , n60909 , n60914 );
or ( n60917 , n60912 , n60915 , n60916 );
and ( n60918 , n60907 , n60917 );
xor ( n60919 , n60222 , n60224 );
xor ( n60920 , n60919 , n60241 );
and ( n60921 , n60917 , n60920 );
and ( n60922 , n60907 , n60920 );
or ( n60923 , n60918 , n60921 , n60922 );
and ( n60924 , n60889 , n60923 );
xor ( n60925 , n60244 , n60540 );
xor ( n60926 , n60925 , n60559 );
and ( n60927 , n60923 , n60926 );
and ( n60928 , n60889 , n60926 );
or ( n60929 , n60924 , n60927 , n60928 );
xor ( n60930 , n60217 , n60219 );
xor ( n60931 , n60930 , n60562 );
and ( n60932 , n60929 , n60931 );
xor ( n60933 , n60590 , n60592 );
xor ( n60934 , n60933 , n60595 );
and ( n60935 , n60931 , n60934 );
and ( n60936 , n60929 , n60934 );
or ( n60937 , n60932 , n60935 , n60936 );
and ( n60938 , n60600 , n60937 );
and ( n60939 , n60598 , n60937 );
or ( n60940 , n60601 , n60938 , n60939 );
xor ( n60941 , n60210 , n60568 );
xor ( n60942 , n60941 , n60571 );
and ( n60943 , n60940 , n60942 );
xor ( n60944 , n60212 , n60214 );
xor ( n60945 , n60944 , n60565 );
xor ( n60946 , n60598 , n60600 );
xor ( n60947 , n60946 , n60937 );
and ( n60948 , n60945 , n60947 );
xor ( n60949 , n60582 , n60584 );
xor ( n60950 , n60949 , n60587 );
xor ( n60951 , n60484 , n60526 );
xor ( n60952 , n60951 , n60537 );
xor ( n60953 , n60551 , n60553 );
xor ( n60954 , n60953 , n60556 );
and ( n60955 , n60952 , n60954 );
xor ( n60956 , n60515 , n60517 );
xor ( n60957 , n60956 , n60520 );
xor ( n60958 , n60486 , n60488 );
xor ( n60959 , n60958 , n60491 );
xor ( n60960 , n60461 , n60465 );
xor ( n60961 , n60960 , n60469 );
xor ( n60962 , n60610 , n60611 );
and ( n60963 , n60961 , n60962 );
and ( n60964 , n47474 , n53357 );
and ( n60965 , n47351 , n53355 );
nor ( n60966 , n60964 , n60965 );
xnor ( n60967 , n60966 , n53060 );
and ( n60968 , n47778 , n52799 );
and ( n60969 , n47647 , n52797 );
nor ( n60970 , n60968 , n60969 );
xnor ( n60971 , n60970 , n52538 );
and ( n60972 , n60967 , n60971 );
and ( n60973 , n48384 , n51750 );
and ( n60974 , n48272 , n51748 );
nor ( n60975 , n60973 , n60974 );
xnor ( n60976 , n60975 , n51520 );
and ( n60977 , n60971 , n60976 );
and ( n60978 , n60967 , n60976 );
or ( n60979 , n60972 , n60977 , n60978 );
and ( n60980 , n49374 , n50338 );
and ( n60981 , n49115 , n50336 );
nor ( n60982 , n60980 , n60981 );
xnor ( n60983 , n60982 , n50111 );
and ( n60984 , n60979 , n60983 );
and ( n60985 , n49781 , n49896 );
and ( n60986 , n49570 , n49894 );
nor ( n60987 , n60985 , n60986 );
xnor ( n60988 , n60987 , n49711 );
and ( n60989 , n60983 , n60988 );
and ( n60990 , n60979 , n60988 );
or ( n60991 , n60984 , n60989 , n60990 );
and ( n60992 , n60962 , n60991 );
and ( n60993 , n60961 , n60991 );
or ( n60994 , n60963 , n60992 , n60993 );
and ( n60995 , n60959 , n60994 );
and ( n60996 , n58628 , n60372 );
not ( n60997 , n60996 );
and ( n60998 , n60376 , n58542 );
not ( n60999 , n60998 );
and ( n61000 , n60997 , n60999 );
not ( n61001 , n61000 );
and ( n61002 , n60376 , n58444 );
not ( n61003 , n61002 );
and ( n61004 , n61001 , n61003 );
buf ( n61005 , n61000 );
and ( n61006 , n61004 , n61005 );
buf ( n61007 , n20211 );
buf ( n61008 , n61007 );
and ( n61009 , n61008 , n58294 );
not ( n61010 , n61009 );
and ( n61011 , n59908 , n58911 );
not ( n61012 , n61011 );
or ( n61013 , n61010 , n61012 );
buf ( n61014 , n20211 );
buf ( n61015 , n61014 );
and ( n61016 , n57948 , n61015 );
not ( n61017 , n61016 );
and ( n61018 , n58915 , n59920 );
not ( n61019 , n61018 );
or ( n61020 , n61017 , n61019 );
and ( n61021 , n61013 , n61020 );
and ( n61022 , n61005 , n61021 );
and ( n61023 , n61004 , n61021 );
or ( n61024 , n61006 , n61022 , n61023 );
and ( n61025 , n60994 , n61024 );
and ( n61026 , n60959 , n61024 );
or ( n61027 , n60995 , n61025 , n61026 );
and ( n61028 , n60957 , n61027 );
xor ( n61029 , n60649 , n60653 );
xor ( n61030 , n61029 , n60658 );
xor ( n61031 , n60665 , n60669 );
xor ( n61032 , n61031 , n60674 );
and ( n61033 , n61030 , n61032 );
buf ( n61034 , n61033 );
xor ( n61035 , n60682 , n60686 );
xor ( n61036 , n61035 , n60691 );
xor ( n61037 , n60701 , n60705 );
xor ( n61038 , n61037 , n60467 );
and ( n61039 , n61036 , n61038 );
xor ( n61040 , n60713 , n60715 );
xor ( n61041 , n61040 , n60718 );
and ( n61042 , n61038 , n61041 );
and ( n61043 , n61036 , n61041 );
or ( n61044 , n61039 , n61042 , n61043 );
and ( n61045 , n61034 , n61044 );
xor ( n61046 , n60724 , n60726 );
xor ( n61047 , n61046 , n60729 );
and ( n61048 , n46530 , n55851 );
and ( n61049 , n46445 , n55849 );
nor ( n61050 , n61048 , n61049 );
xnor ( n61051 , n61050 , n55506 );
and ( n61052 , n47216 , n53928 );
and ( n61053 , n47090 , n53926 );
nor ( n61054 , n61052 , n61053 );
xnor ( n61055 , n61054 , n53652 );
and ( n61056 , n61051 , n61055 );
and ( n61057 , n48108 , n52269 );
and ( n61058 , n47962 , n52267 );
nor ( n61059 , n61057 , n61058 );
xnor ( n61060 , n61059 , n52008 );
and ( n61061 , n61055 , n61060 );
and ( n61062 , n61051 , n61060 );
or ( n61063 , n61056 , n61061 , n61062 );
and ( n61064 , n61047 , n61063 );
and ( n61065 , n46969 , n54535 );
and ( n61066 , n46843 , n54533 );
nor ( n61067 , n61065 , n61066 );
xnor ( n61068 , n61067 , n54237 );
and ( n61069 , n48709 , n51221 );
and ( n61070 , n48632 , n51219 );
nor ( n61071 , n61069 , n61070 );
xnor ( n61072 , n61071 , n51000 );
and ( n61073 , n61068 , n61072 );
and ( n61074 , n49115 , n50783 );
and ( n61075 , n48988 , n50781 );
nor ( n61076 , n61074 , n61075 );
xnor ( n61077 , n61076 , n50557 );
and ( n61078 , n61072 , n61077 );
and ( n61079 , n61068 , n61077 );
or ( n61080 , n61073 , n61078 , n61079 );
and ( n61081 , n61063 , n61080 );
and ( n61082 , n61047 , n61080 );
or ( n61083 , n61064 , n61081 , n61082 );
and ( n61084 , n61044 , n61083 );
and ( n61085 , n61034 , n61083 );
or ( n61086 , n61045 , n61084 , n61085 );
and ( n61087 , n52332 , n48042 );
and ( n61088 , n52082 , n48040 );
nor ( n61089 , n61087 , n61088 );
xnor ( n61090 , n61089 , n47921 );
and ( n61091 , n53328 , n47429 );
and ( n61092 , n53041 , n47427 );
nor ( n61093 , n61091 , n61092 );
xnor ( n61094 , n61093 , n47309 );
and ( n61095 , n61090 , n61094 );
and ( n61096 , n57063 , n46133 );
not ( n61097 , n61096 );
and ( n61098 , n61097 , n46067 );
and ( n61099 , n61094 , n61098 );
and ( n61100 , n61090 , n61098 );
or ( n61101 , n61095 , n61099 , n61100 );
and ( n61102 , n59365 , n59611 );
not ( n61103 , n61102 );
and ( n61104 , n59615 , n59207 );
not ( n61105 , n61104 );
and ( n61106 , n61103 , n61105 );
and ( n61107 , n61101 , n61106 );
and ( n61108 , n46169 , n57187 );
and ( n61109 , n46100 , n57184 );
nor ( n61110 , n61108 , n61109 );
xnor ( n61111 , n61110 , n56175 );
and ( n61112 , n46345 , n56503 );
and ( n61113 , n46264 , n56501 );
nor ( n61114 , n61112 , n61113 );
xnor ( n61115 , n61114 , n56178 );
and ( n61116 , n61111 , n61115 );
and ( n61117 , n46750 , n55159 );
and ( n61118 , n46577 , n55157 );
nor ( n61119 , n61117 , n61118 );
xnor ( n61120 , n61119 , n54864 );
and ( n61121 , n61115 , n61120 );
and ( n61122 , n61111 , n61120 );
or ( n61123 , n61116 , n61121 , n61122 );
and ( n61124 , n61106 , n61123 );
and ( n61125 , n61101 , n61123 );
or ( n61126 , n61107 , n61124 , n61125 );
and ( n61127 , n49976 , n49896 );
and ( n61128 , n49781 , n49894 );
nor ( n61129 , n61127 , n61128 );
xnor ( n61130 , n61129 , n49711 );
and ( n61131 , n50726 , n49121 );
and ( n61132 , n50625 , n49119 );
nor ( n61133 , n61131 , n61132 );
xnor ( n61134 , n61133 , n48932 );
and ( n61135 , n61130 , n61134 );
and ( n61136 , n51298 , n48740 );
and ( n61137 , n51077 , n48738 );
nor ( n61138 , n61136 , n61137 );
xnor ( n61139 , n61138 , n48571 );
and ( n61140 , n61134 , n61139 );
and ( n61141 , n61130 , n61139 );
or ( n61142 , n61135 , n61140 , n61141 );
and ( n61143 , n51734 , n48394 );
and ( n61144 , n51510 , n48392 );
nor ( n61145 , n61143 , n61144 );
xnor ( n61146 , n61145 , n48220 );
and ( n61147 , n52790 , n47734 );
and ( n61148 , n52612 , n47732 );
nor ( n61149 , n61147 , n61148 );
xnor ( n61150 , n61149 , n47606 );
and ( n61151 , n61146 , n61150 );
and ( n61152 , n53922 , n47178 );
and ( n61153 , n53639 , n47176 );
nor ( n61154 , n61152 , n61153 );
xnor ( n61155 , n61154 , n47039 );
and ( n61156 , n61150 , n61155 );
and ( n61157 , n61146 , n61155 );
or ( n61158 , n61151 , n61156 , n61157 );
and ( n61159 , n61142 , n61158 );
and ( n61160 , n54604 , n46911 );
and ( n61161 , n54227 , n46909 );
nor ( n61162 , n61160 , n61161 );
xnor ( n61163 , n61162 , n46802 );
and ( n61164 , n55143 , n46712 );
and ( n61165 , n54942 , n46710 );
nor ( n61166 , n61164 , n61165 );
xnor ( n61167 , n61166 , n46587 );
and ( n61168 , n61163 , n61167 );
and ( n61169 , n55756 , n46496 );
and ( n61170 , n55497 , n46494 );
nor ( n61171 , n61169 , n61170 );
xnor ( n61172 , n61171 , n46402 );
and ( n61173 , n61167 , n61172 );
and ( n61174 , n61163 , n61172 );
or ( n61175 , n61168 , n61173 , n61174 );
and ( n61176 , n61158 , n61175 );
and ( n61177 , n61142 , n61175 );
or ( n61178 , n61159 , n61176 , n61177 );
and ( n61179 , n61126 , n61178 );
xor ( n61180 , n39410 , n45569 );
buf ( n61181 , n61180 );
buf ( n61182 , n61181 );
buf ( n61183 , n61182 );
and ( n61184 , n60821 , n58444 );
not ( n61185 , n61184 );
and ( n61186 , n61183 , n61185 );
buf ( n61187 , n61186 );
xor ( n61188 , n60740 , n60744 );
xor ( n61189 , n61188 , n60749 );
and ( n61190 , n61187 , n61189 );
xor ( n61191 , n60756 , n60760 );
xor ( n61192 , n61191 , n60765 );
and ( n61193 , n61189 , n61192 );
and ( n61194 , n61187 , n61192 );
or ( n61195 , n61190 , n61193 , n61194 );
and ( n61196 , n61178 , n61195 );
and ( n61197 , n61126 , n61195 );
or ( n61198 , n61179 , n61196 , n61197 );
and ( n61199 , n61086 , n61198 );
xor ( n61200 , n60773 , n60777 );
xor ( n61201 , n61200 , n60782 );
xor ( n61202 , n60798 , n60802 );
xor ( n61203 , n61202 , n60807 );
and ( n61204 , n61201 , n61203 );
xor ( n61205 , n60814 , n60818 );
xor ( n61206 , n61205 , n60823 );
and ( n61207 , n61203 , n61206 );
and ( n61208 , n61201 , n61206 );
or ( n61209 , n61204 , n61207 , n61208 );
buf ( n61210 , n60619 );
xor ( n61211 , n61210 , n60621 );
and ( n61212 , n61209 , n61211 );
xor ( n61213 , n60625 , n60627 );
xor ( n61214 , n61213 , n60630 );
and ( n61215 , n61211 , n61214 );
and ( n61216 , n61209 , n61214 );
or ( n61217 , n61212 , n61215 , n61216 );
and ( n61218 , n61198 , n61217 );
and ( n61219 , n61086 , n61217 );
or ( n61220 , n61199 , n61218 , n61219 );
and ( n61221 , n61027 , n61220 );
and ( n61222 , n60957 , n61220 );
or ( n61223 , n61028 , n61221 , n61222 );
xor ( n61224 , n60635 , n60636 );
xor ( n61225 , n61224 , n60638 );
xor ( n61226 , n60661 , n60677 );
xor ( n61227 , n61226 , n60694 );
and ( n61228 , n61225 , n61227 );
xor ( n61229 , n60709 , n60721 );
xor ( n61230 , n61229 , n60732 );
and ( n61231 , n61227 , n61230 );
and ( n61232 , n61225 , n61230 );
or ( n61233 , n61228 , n61231 , n61232 );
xor ( n61234 , n60752 , n60768 );
xor ( n61235 , n61234 , n60785 );
xor ( n61236 , n60810 , n60826 );
xor ( n61237 , n61236 , n60829 );
and ( n61238 , n61235 , n61237 );
xor ( n61239 , n60834 , n60836 );
xor ( n61240 , n61239 , n60839 );
and ( n61241 , n61237 , n61240 );
and ( n61242 , n61235 , n61240 );
or ( n61243 , n61238 , n61241 , n61242 );
and ( n61244 , n61233 , n61243 );
xor ( n61245 , n60607 , n60608 );
xor ( n61246 , n61245 , n60612 );
and ( n61247 , n61243 , n61246 );
and ( n61248 , n61233 , n61246 );
or ( n61249 , n61244 , n61247 , n61248 );
xor ( n61250 , n60623 , n60633 );
xor ( n61251 , n61250 , n60641 );
xor ( n61252 , n60697 , n60735 );
xor ( n61253 , n61252 , n60788 );
and ( n61254 , n61251 , n61253 );
xor ( n61255 , n60832 , n60842 );
xor ( n61256 , n61255 , n60845 );
and ( n61257 , n61253 , n61256 );
and ( n61258 , n61251 , n61256 );
or ( n61259 , n61254 , n61257 , n61258 );
and ( n61260 , n61249 , n61259 );
xor ( n61261 , n60615 , n60644 );
xor ( n61262 , n61261 , n60791 );
and ( n61263 , n61259 , n61262 );
and ( n61264 , n61249 , n61262 );
or ( n61265 , n61260 , n61263 , n61264 );
and ( n61266 , n61223 , n61265 );
xor ( n61267 , n60848 , n60858 );
xor ( n61268 , n61267 , n60869 );
xor ( n61269 , n60875 , n60877 );
xor ( n61270 , n61269 , n60880 );
and ( n61271 , n61268 , n61270 );
xor ( n61272 , n60891 , n60893 );
xor ( n61273 , n61272 , n60896 );
and ( n61274 , n61270 , n61273 );
and ( n61275 , n61268 , n61273 );
or ( n61276 , n61271 , n61274 , n61275 );
and ( n61277 , n61265 , n61276 );
and ( n61278 , n61223 , n61276 );
or ( n61279 , n61266 , n61277 , n61278 );
and ( n61280 , n60954 , n61279 );
and ( n61281 , n60952 , n61279 );
or ( n61282 , n60955 , n61280 , n61281 );
and ( n61283 , n60950 , n61282 );
xor ( n61284 , n60794 , n60872 );
xor ( n61285 , n61284 , n60883 );
xor ( n61286 , n60899 , n60901 );
xor ( n61287 , n61286 , n60904 );
and ( n61288 , n61285 , n61287 );
xor ( n61289 , n60909 , n60911 );
xor ( n61290 , n61289 , n60914 );
and ( n61291 , n61287 , n61290 );
and ( n61292 , n61285 , n61290 );
or ( n61293 , n61288 , n61291 , n61292 );
xor ( n61294 , n60603 , n60605 );
xor ( n61295 , n61294 , n60886 );
and ( n61296 , n61293 , n61295 );
xor ( n61297 , n60907 , n60917 );
xor ( n61298 , n61297 , n60920 );
and ( n61299 , n61295 , n61298 );
and ( n61300 , n61293 , n61298 );
or ( n61301 , n61296 , n61299 , n61300 );
and ( n61302 , n61282 , n61301 );
and ( n61303 , n60950 , n61301 );
or ( n61304 , n61283 , n61302 , n61303 );
xor ( n61305 , n60929 , n60931 );
xor ( n61306 , n61305 , n60934 );
and ( n61307 , n61304 , n61306 );
xor ( n61308 , n60889 , n60923 );
xor ( n61309 , n61308 , n60926 );
xor ( n61310 , n60850 , n60852 );
xor ( n61311 , n61310 , n60855 );
xor ( n61312 , n60861 , n60863 );
xor ( n61313 , n61312 , n60866 );
and ( n61314 , n61311 , n61313 );
and ( n61315 , n48272 , n52269 );
and ( n61316 , n48108 , n52267 );
nor ( n61317 , n61315 , n61316 );
xnor ( n61318 , n61317 , n52008 );
and ( n61319 , n48632 , n51750 );
and ( n61320 , n48384 , n51748 );
nor ( n61321 , n61319 , n61320 );
xnor ( n61322 , n61321 , n51520 );
and ( n61323 , n61318 , n61322 );
and ( n61324 , n49374 , n50783 );
and ( n61325 , n49115 , n50781 );
nor ( n61326 , n61324 , n61325 );
xnor ( n61327 , n61326 , n50557 );
and ( n61328 , n61322 , n61327 );
and ( n61329 , n61318 , n61327 );
or ( n61330 , n61323 , n61328 , n61329 );
and ( n61331 , n46843 , n55159 );
and ( n61332 , n46750 , n55157 );
nor ( n61333 , n61331 , n61332 );
xnor ( n61334 , n61333 , n54864 );
and ( n61335 , n47090 , n54535 );
and ( n61336 , n46969 , n54533 );
nor ( n61337 , n61335 , n61336 );
xnor ( n61338 , n61337 , n54237 );
and ( n61339 , n61334 , n61338 );
and ( n61340 , n47351 , n53928 );
and ( n61341 , n47216 , n53926 );
nor ( n61342 , n61340 , n61341 );
xnor ( n61343 , n61342 , n53652 );
and ( n61344 , n61338 , n61343 );
and ( n61345 , n61334 , n61343 );
or ( n61346 , n61339 , n61344 , n61345 );
and ( n61347 , n61330 , n61346 );
and ( n61348 , n49570 , n50338 );
and ( n61349 , n49374 , n50336 );
nor ( n61350 , n61348 , n61349 );
xnor ( n61351 , n61350 , n50111 );
and ( n61352 , n61346 , n61351 );
and ( n61353 , n61330 , n61351 );
or ( n61354 , n61347 , n61352 , n61353 );
and ( n61355 , n46264 , n57187 );
and ( n61356 , n46169 , n57184 );
nor ( n61357 , n61355 , n61356 );
xnor ( n61358 , n61357 , n56175 );
and ( n61359 , n47647 , n53357 );
and ( n61360 , n47474 , n53355 );
nor ( n61361 , n61359 , n61360 );
xnor ( n61362 , n61361 , n53060 );
and ( n61363 , n61358 , n61362 );
and ( n61364 , n47962 , n52799 );
and ( n61365 , n47778 , n52797 );
nor ( n61366 , n61364 , n61365 );
xnor ( n61367 , n61366 , n52538 );
and ( n61368 , n61362 , n61367 );
and ( n61369 , n61358 , n61367 );
or ( n61370 , n61363 , n61368 , n61369 );
xor ( n61371 , n61051 , n61055 );
xor ( n61372 , n61371 , n61060 );
and ( n61373 , n61370 , n61372 );
xor ( n61374 , n61068 , n61072 );
xor ( n61375 , n61374 , n61077 );
and ( n61376 , n61372 , n61375 );
and ( n61377 , n61370 , n61375 );
or ( n61378 , n61373 , n61376 , n61377 );
and ( n61379 , n61354 , n61378 );
and ( n61380 , n50195 , n49513 );
and ( n61381 , n49976 , n49511 );
nor ( n61382 , n61380 , n61381 );
xnor ( n61383 , n61382 , n49310 );
and ( n61384 , n61378 , n61383 );
and ( n61385 , n61354 , n61383 );
or ( n61386 , n61379 , n61384 , n61385 );
xnor ( n61387 , n61010 , n61012 );
xnor ( n61388 , n61017 , n61019 );
and ( n61389 , n61387 , n61388 );
buf ( n61390 , n59365 );
not ( n61391 , n61390 );
or ( n61392 , n61389 , n61391 );
and ( n61393 , n61386 , n61392 );
xor ( n61394 , n60979 , n60983 );
xor ( n61395 , n61394 , n60988 );
xor ( n61396 , n61001 , n61003 );
and ( n61397 , n61395 , n61396 );
xor ( n61398 , n61013 , n61020 );
and ( n61399 , n61396 , n61398 );
and ( n61400 , n61395 , n61398 );
or ( n61401 , n61397 , n61399 , n61400 );
and ( n61402 , n61392 , n61401 );
and ( n61403 , n61386 , n61401 );
or ( n61404 , n61393 , n61402 , n61403 );
and ( n61405 , n61313 , n61404 );
and ( n61406 , n61311 , n61404 );
or ( n61407 , n61314 , n61405 , n61406 );
and ( n61408 , n52082 , n48394 );
and ( n61409 , n51734 , n48392 );
nor ( n61410 , n61408 , n61409 );
xnor ( n61411 , n61410 , n48220 );
and ( n61412 , n52612 , n48042 );
and ( n61413 , n52332 , n48040 );
nor ( n61414 , n61412 , n61413 );
xnor ( n61415 , n61414 , n47921 );
and ( n61416 , n61411 , n61415 );
and ( n61417 , n55497 , n46712 );
and ( n61418 , n55143 , n46710 );
nor ( n61419 , n61417 , n61418 );
xnor ( n61420 , n61419 , n46587 );
and ( n61421 , n61415 , n61420 );
and ( n61422 , n61411 , n61420 );
or ( n61423 , n61416 , n61421 , n61422 );
and ( n61424 , n56388 , n46306 );
and ( n61425 , n56255 , n46304 );
nor ( n61426 , n61424 , n61425 );
xnor ( n61427 , n61426 , n46228 );
and ( n61428 , n61423 , n61427 );
and ( n61429 , n57063 , n46135 );
and ( n61430 , n56915 , n46133 );
nor ( n61431 , n61429 , n61430 );
xnor ( n61432 , n61431 , n46067 );
and ( n61433 , n61427 , n61432 );
and ( n61434 , n61423 , n61432 );
or ( n61435 , n61428 , n61433 , n61434 );
and ( n61436 , n61008 , n58444 );
not ( n61437 , n61436 );
and ( n61438 , n58915 , n60372 );
not ( n61439 , n61438 );
and ( n61440 , n61437 , n61439 );
buf ( n61441 , n59615 );
not ( n61442 , n61441 );
and ( n61443 , n61439 , n61442 );
and ( n61444 , n61437 , n61442 );
or ( n61445 , n61440 , n61443 , n61444 );
and ( n61446 , n58292 , n60711 );
not ( n61447 , n61446 );
or ( n61448 , n61445 , n61447 );
and ( n61449 , n61435 , n61448 );
xor ( n61450 , n60967 , n60971 );
xor ( n61451 , n61450 , n60976 );
xor ( n61452 , n61090 , n61094 );
xor ( n61453 , n61452 , n61098 );
and ( n61454 , n61451 , n61453 );
xor ( n61455 , n60997 , n60999 );
and ( n61456 , n61453 , n61455 );
and ( n61457 , n61451 , n61455 );
or ( n61458 , n61454 , n61456 , n61457 );
and ( n61459 , n61448 , n61458 );
and ( n61460 , n61435 , n61458 );
or ( n61461 , n61449 , n61459 , n61460 );
xor ( n61462 , n61103 , n61105 );
and ( n61463 , n53639 , n47429 );
and ( n61464 , n53328 , n47427 );
nor ( n61465 , n61463 , n61464 );
xnor ( n61466 , n61465 , n47309 );
and ( n61467 , n54227 , n47178 );
and ( n61468 , n53922 , n47176 );
nor ( n61469 , n61467 , n61468 );
xnor ( n61470 , n61469 , n47039 );
and ( n61471 , n61466 , n61470 );
and ( n61472 , n54942 , n46911 );
and ( n61473 , n54604 , n46909 );
nor ( n61474 , n61472 , n61473 );
xnor ( n61475 , n61474 , n46802 );
and ( n61476 , n61470 , n61475 );
and ( n61477 , n61466 , n61475 );
or ( n61478 , n61471 , n61476 , n61477 );
and ( n61479 , n61462 , n61478 );
buf ( n61480 , n20214 );
buf ( n61481 , n61480 );
and ( n61482 , n57948 , n61481 );
not ( n61483 , n61482 );
and ( n61484 , n58292 , n61015 );
not ( n61485 , n61484 );
and ( n61486 , n61483 , n61485 );
and ( n61487 , n59365 , n59920 );
not ( n61488 , n61487 );
and ( n61489 , n61485 , n61488 );
and ( n61490 , n61483 , n61488 );
or ( n61491 , n61486 , n61489 , n61490 );
and ( n61492 , n61478 , n61491 );
and ( n61493 , n61462 , n61491 );
or ( n61494 , n61479 , n61492 , n61493 );
and ( n61495 , n46445 , n56503 );
and ( n61496 , n46345 , n56501 );
nor ( n61497 , n61495 , n61496 );
xnor ( n61498 , n61497 , n56178 );
and ( n61499 , n46577 , n55851 );
and ( n61500 , n46530 , n55849 );
nor ( n61501 , n61499 , n61500 );
xnor ( n61502 , n61501 , n55506 );
or ( n61503 , n61498 , n61502 );
buf ( n61504 , n20214 );
buf ( n61505 , n61504 );
and ( n61506 , n61505 , n58294 );
not ( n61507 , n61506 );
and ( n61508 , n59908 , n59207 );
not ( n61509 , n61508 );
and ( n61510 , n61507 , n61509 );
and ( n61511 , n61503 , n61510 );
and ( n61512 , n60821 , n58542 );
and ( n61513 , n60376 , n58911 );
not ( n61514 , n61513 );
and ( n61515 , n61512 , n61514 );
and ( n61516 , n61510 , n61515 );
and ( n61517 , n61503 , n61515 );
or ( n61518 , n61511 , n61516 , n61517 );
and ( n61519 , n61494 , n61518 );
not ( n61520 , n61512 );
buf ( n61521 , n61520 );
and ( n61522 , n48988 , n51221 );
and ( n61523 , n48709 , n51219 );
nor ( n61524 , n61522 , n61523 );
xnor ( n61525 , n61524 , n51000 );
and ( n61526 , n49781 , n50338 );
and ( n61527 , n49570 , n50336 );
nor ( n61528 , n61526 , n61527 );
xnor ( n61529 , n61528 , n50111 );
and ( n61530 , n61525 , n61529 );
and ( n61531 , n50195 , n49896 );
and ( n61532 , n49976 , n49894 );
nor ( n61533 , n61531 , n61532 );
xnor ( n61534 , n61533 , n49711 );
and ( n61535 , n61529 , n61534 );
and ( n61536 , n61525 , n61534 );
or ( n61537 , n61530 , n61535 , n61536 );
and ( n61538 , n61521 , n61537 );
and ( n61539 , n50625 , n49513 );
and ( n61540 , n50404 , n49511 );
nor ( n61541 , n61539 , n61540 );
xnor ( n61542 , n61541 , n49310 );
and ( n61543 , n51077 , n49121 );
and ( n61544 , n50726 , n49119 );
nor ( n61545 , n61543 , n61544 );
xnor ( n61546 , n61545 , n48932 );
and ( n61547 , n61542 , n61546 );
and ( n61548 , n51510 , n48740 );
and ( n61549 , n51298 , n48738 );
nor ( n61550 , n61548 , n61549 );
xnor ( n61551 , n61550 , n48571 );
and ( n61552 , n61546 , n61551 );
and ( n61553 , n61542 , n61551 );
or ( n61554 , n61547 , n61552 , n61553 );
and ( n61555 , n61537 , n61554 );
and ( n61556 , n61521 , n61554 );
or ( n61557 , n61538 , n61555 , n61556 );
and ( n61558 , n61518 , n61557 );
and ( n61559 , n61494 , n61557 );
or ( n61560 , n61519 , n61558 , n61559 );
and ( n61561 , n61461 , n61560 );
and ( n61562 , n53041 , n47734 );
and ( n61563 , n52790 , n47732 );
nor ( n61564 , n61562 , n61563 );
xnor ( n61565 , n61564 , n47606 );
and ( n61566 , n56255 , n46496 );
and ( n61567 , n55756 , n46494 );
nor ( n61568 , n61566 , n61567 );
xnor ( n61569 , n61568 , n46402 );
and ( n61570 , n61565 , n61569 );
and ( n61571 , n56915 , n46306 );
and ( n61572 , n56388 , n46304 );
nor ( n61573 , n61571 , n61572 );
xnor ( n61574 , n61573 , n46228 );
and ( n61575 , n61569 , n61574 );
and ( n61576 , n61565 , n61574 );
or ( n61577 , n61570 , n61575 , n61576 );
xor ( n61578 , n39412 , n45568 );
buf ( n61579 , n61578 );
buf ( n61580 , n61579 );
buf ( n61581 , n61580 );
and ( n61582 , n61096 , n61581 );
buf ( n61583 , n61582 );
and ( n61584 , n61577 , n61583 );
xor ( n61585 , n61111 , n61115 );
xor ( n61586 , n61585 , n61120 );
and ( n61587 , n61583 , n61586 );
and ( n61588 , n61577 , n61586 );
or ( n61589 , n61584 , n61587 , n61588 );
xor ( n61590 , n61130 , n61134 );
xor ( n61591 , n61590 , n61139 );
xor ( n61592 , n61146 , n61150 );
xor ( n61593 , n61592 , n61155 );
and ( n61594 , n61591 , n61593 );
xor ( n61595 , n61163 , n61167 );
xor ( n61596 , n61595 , n61172 );
and ( n61597 , n61593 , n61596 );
and ( n61598 , n61591 , n61596 );
or ( n61599 , n61594 , n61597 , n61598 );
and ( n61600 , n61589 , n61599 );
buf ( n61601 , n61030 );
xor ( n61602 , n61601 , n61032 );
and ( n61603 , n61599 , n61602 );
and ( n61604 , n61589 , n61602 );
or ( n61605 , n61600 , n61603 , n61604 );
and ( n61606 , n61560 , n61605 );
and ( n61607 , n61461 , n61605 );
or ( n61608 , n61561 , n61606 , n61607 );
xor ( n61609 , n61036 , n61038 );
xor ( n61610 , n61609 , n61041 );
xor ( n61611 , n61047 , n61063 );
xor ( n61612 , n61611 , n61080 );
and ( n61613 , n61610 , n61612 );
xor ( n61614 , n61101 , n61106 );
xor ( n61615 , n61614 , n61123 );
and ( n61616 , n61612 , n61615 );
and ( n61617 , n61610 , n61615 );
or ( n61618 , n61613 , n61616 , n61617 );
xor ( n61619 , n61142 , n61158 );
xor ( n61620 , n61619 , n61175 );
xor ( n61621 , n61187 , n61189 );
xor ( n61622 , n61621 , n61192 );
and ( n61623 , n61620 , n61622 );
xor ( n61624 , n61201 , n61203 );
xor ( n61625 , n61624 , n61206 );
and ( n61626 , n61622 , n61625 );
and ( n61627 , n61620 , n61625 );
or ( n61628 , n61623 , n61626 , n61627 );
and ( n61629 , n61618 , n61628 );
xor ( n61630 , n60961 , n60962 );
xor ( n61631 , n61630 , n60991 );
and ( n61632 , n61628 , n61631 );
and ( n61633 , n61618 , n61631 );
or ( n61634 , n61629 , n61632 , n61633 );
and ( n61635 , n61608 , n61634 );
xor ( n61636 , n61004 , n61005 );
xor ( n61637 , n61636 , n61021 );
xor ( n61638 , n61034 , n61044 );
xor ( n61639 , n61638 , n61083 );
and ( n61640 , n61637 , n61639 );
xor ( n61641 , n61126 , n61178 );
xor ( n61642 , n61641 , n61195 );
and ( n61643 , n61639 , n61642 );
and ( n61644 , n61637 , n61642 );
or ( n61645 , n61640 , n61643 , n61644 );
and ( n61646 , n61634 , n61645 );
and ( n61647 , n61608 , n61645 );
or ( n61648 , n61635 , n61646 , n61647 );
and ( n61649 , n61407 , n61648 );
xor ( n61650 , n61209 , n61211 );
xor ( n61651 , n61650 , n61214 );
xor ( n61652 , n61225 , n61227 );
xor ( n61653 , n61652 , n61230 );
and ( n61654 , n61651 , n61653 );
xor ( n61655 , n61235 , n61237 );
xor ( n61656 , n61655 , n61240 );
and ( n61657 , n61653 , n61656 );
and ( n61658 , n61651 , n61656 );
or ( n61659 , n61654 , n61657 , n61658 );
xor ( n61660 , n60959 , n60994 );
xor ( n61661 , n61660 , n61024 );
and ( n61662 , n61659 , n61661 );
xor ( n61663 , n61086 , n61198 );
xor ( n61664 , n61663 , n61217 );
and ( n61665 , n61661 , n61664 );
and ( n61666 , n61659 , n61664 );
or ( n61667 , n61662 , n61665 , n61666 );
and ( n61668 , n61648 , n61667 );
and ( n61669 , n61407 , n61667 );
or ( n61670 , n61649 , n61668 , n61669 );
xor ( n61671 , n60957 , n61027 );
xor ( n61672 , n61671 , n61220 );
xor ( n61673 , n61249 , n61259 );
xor ( n61674 , n61673 , n61262 );
and ( n61675 , n61672 , n61674 );
xor ( n61676 , n61268 , n61270 );
xor ( n61677 , n61676 , n61273 );
and ( n61678 , n61674 , n61677 );
and ( n61679 , n61672 , n61677 );
or ( n61680 , n61675 , n61678 , n61679 );
and ( n61681 , n61670 , n61680 );
xor ( n61682 , n61223 , n61265 );
xor ( n61683 , n61682 , n61276 );
and ( n61684 , n61680 , n61683 );
and ( n61685 , n61670 , n61683 );
or ( n61686 , n61681 , n61684 , n61685 );
xor ( n61687 , n60952 , n60954 );
xor ( n61688 , n61687 , n61279 );
and ( n61689 , n61686 , n61688 );
xor ( n61690 , n61293 , n61295 );
xor ( n61691 , n61690 , n61298 );
and ( n61692 , n61688 , n61691 );
and ( n61693 , n61686 , n61691 );
or ( n61694 , n61689 , n61692 , n61693 );
and ( n61695 , n61309 , n61694 );
xor ( n61696 , n60950 , n61282 );
xor ( n61697 , n61696 , n61301 );
and ( n61698 , n61694 , n61697 );
and ( n61699 , n61309 , n61697 );
or ( n61700 , n61695 , n61698 , n61699 );
and ( n61701 , n61306 , n61700 );
and ( n61702 , n61304 , n61700 );
or ( n61703 , n61307 , n61701 , n61702 );
and ( n61704 , n60947 , n61703 );
and ( n61705 , n60945 , n61703 );
or ( n61706 , n60948 , n61704 , n61705 );
and ( n61707 , n60942 , n61706 );
and ( n61708 , n60940 , n61706 );
or ( n61709 , n60943 , n61707 , n61708 );
or ( n61710 , n60580 , n61709 );
and ( n61711 , n60577 , n61710 );
and ( n61712 , n59856 , n61710 );
or ( n61713 , n60578 , n61711 , n61712 );
and ( n61714 , n59853 , n61713 );
and ( n61715 , n59851 , n61713 );
or ( n61716 , n59854 , n61714 , n61715 );
and ( n61717 , n59481 , n61716 );
xor ( n61718 , n59481 , n61716 );
xor ( n61719 , n59851 , n59853 );
xor ( n61720 , n61719 , n61713 );
xor ( n61721 , n59856 , n60577 );
xor ( n61722 , n61721 , n61710 );
not ( n61723 , n61722 );
xnor ( n61724 , n60580 , n61709 );
xor ( n61725 , n60940 , n60942 );
xor ( n61726 , n61725 , n61706 );
not ( n61727 , n61726 );
xor ( n61728 , n60945 , n60947 );
xor ( n61729 , n61728 , n61703 );
not ( n61730 , n61729 );
xor ( n61731 , n61304 , n61306 );
xor ( n61732 , n61731 , n61700 );
xor ( n61733 , n61309 , n61694 );
xor ( n61734 , n61733 , n61697 );
xor ( n61735 , n61285 , n61287 );
xor ( n61736 , n61735 , n61290 );
xor ( n61737 , n61233 , n61243 );
xor ( n61738 , n61737 , n61246 );
xor ( n61739 , n61251 , n61253 );
xor ( n61740 , n61739 , n61256 );
and ( n61741 , n61738 , n61740 );
xor ( n61742 , n61318 , n61322 );
xor ( n61743 , n61742 , n61327 );
xor ( n61744 , n61358 , n61362 );
xor ( n61745 , n61744 , n61367 );
and ( n61746 , n61743 , n61745 );
xor ( n61747 , n61334 , n61338 );
xor ( n61748 , n61747 , n61343 );
and ( n61749 , n61745 , n61748 );
and ( n61750 , n61743 , n61748 );
or ( n61751 , n61746 , n61749 , n61750 );
and ( n61752 , n50404 , n49513 );
and ( n61753 , n50195 , n49511 );
nor ( n61754 , n61752 , n61753 );
xnor ( n61755 , n61754 , n49310 );
and ( n61756 , n61751 , n61755 );
xor ( n61757 , n61330 , n61346 );
xor ( n61758 , n61757 , n61351 );
and ( n61759 , n61755 , n61758 );
and ( n61760 , n61751 , n61758 );
or ( n61761 , n61756 , n61759 , n61760 );
xor ( n61762 , n61354 , n61378 );
xor ( n61763 , n61762 , n61383 );
and ( n61764 , n61761 , n61763 );
xnor ( n61765 , n61389 , n61391 );
xor ( n61766 , n61183 , n61185 );
buf ( n61767 , n61766 );
xor ( n61768 , n61423 , n61427 );
xor ( n61769 , n61768 , n61432 );
and ( n61770 , n61767 , n61769 );
xor ( n61771 , n61370 , n61372 );
xor ( n61772 , n61771 , n61375 );
and ( n61773 , n61769 , n61772 );
and ( n61774 , n61767 , n61772 );
or ( n61775 , n61770 , n61773 , n61774 );
and ( n61776 , n61765 , n61775 );
xnor ( n61777 , n61445 , n61447 );
xor ( n61778 , n61387 , n61388 );
and ( n61779 , n61777 , n61778 );
and ( n61780 , n61505 , n58444 );
not ( n61781 , n61780 );
and ( n61782 , n61008 , n58542 );
not ( n61783 , n61782 );
and ( n61784 , n61781 , n61783 );
and ( n61785 , n60376 , n59207 );
not ( n61786 , n61785 );
and ( n61787 , n61783 , n61786 );
and ( n61788 , n61781 , n61786 );
or ( n61789 , n61784 , n61787 , n61788 );
and ( n61790 , n58628 , n60711 );
not ( n61791 , n61790 );
and ( n61792 , n61789 , n61791 );
xor ( n61793 , n61437 , n61439 );
xor ( n61794 , n61793 , n61442 );
and ( n61795 , n61791 , n61794 );
and ( n61796 , n61789 , n61794 );
or ( n61797 , n61792 , n61795 , n61796 );
and ( n61798 , n61778 , n61797 );
and ( n61799 , n61777 , n61797 );
or ( n61800 , n61779 , n61798 , n61799 );
and ( n61801 , n61775 , n61800 );
and ( n61802 , n61765 , n61800 );
or ( n61803 , n61776 , n61801 , n61802 );
and ( n61804 , n61764 , n61803 );
xor ( n61805 , n61411 , n61415 );
xor ( n61806 , n61805 , n61420 );
xor ( n61807 , n61466 , n61470 );
xor ( n61808 , n61807 , n61475 );
or ( n61809 , n61806 , n61808 );
xor ( n61810 , n61483 , n61485 );
xor ( n61811 , n61810 , n61488 );
xnor ( n61812 , n61498 , n61502 );
and ( n61813 , n61811 , n61812 );
xor ( n61814 , n61507 , n61509 );
and ( n61815 , n61812 , n61814 );
and ( n61816 , n61811 , n61814 );
or ( n61817 , n61813 , n61815 , n61816 );
and ( n61818 , n61809 , n61817 );
xor ( n61819 , n61512 , n61514 );
and ( n61820 , n48108 , n52799 );
and ( n61821 , n47962 , n52797 );
nor ( n61822 , n61820 , n61821 );
xnor ( n61823 , n61822 , n52538 );
and ( n61824 , n48384 , n52269 );
and ( n61825 , n48272 , n52267 );
nor ( n61826 , n61824 , n61825 );
xnor ( n61827 , n61826 , n52008 );
and ( n61828 , n61823 , n61827 );
and ( n61829 , n48709 , n51750 );
and ( n61830 , n48632 , n51748 );
nor ( n61831 , n61829 , n61830 );
xnor ( n61832 , n61831 , n51520 );
and ( n61833 , n61827 , n61832 );
and ( n61834 , n61823 , n61832 );
or ( n61835 , n61828 , n61833 , n61834 );
and ( n61836 , n61819 , n61835 );
and ( n61837 , n46345 , n57187 );
and ( n61838 , n46264 , n57184 );
nor ( n61839 , n61837 , n61838 );
xnor ( n61840 , n61839 , n56175 );
and ( n61841 , n46530 , n56503 );
and ( n61842 , n46445 , n56501 );
nor ( n61843 , n61841 , n61842 );
xnor ( n61844 , n61843 , n56178 );
and ( n61845 , n61840 , n61844 );
and ( n61846 , n46750 , n55851 );
and ( n61847 , n46577 , n55849 );
nor ( n61848 , n61846 , n61847 );
xnor ( n61849 , n61848 , n55506 );
and ( n61850 , n61844 , n61849 );
and ( n61851 , n61840 , n61849 );
or ( n61852 , n61845 , n61850 , n61851 );
and ( n61853 , n61835 , n61852 );
and ( n61854 , n61819 , n61852 );
or ( n61855 , n61836 , n61853 , n61854 );
and ( n61856 , n61817 , n61855 );
and ( n61857 , n61809 , n61855 );
or ( n61858 , n61818 , n61856 , n61857 );
and ( n61859 , n47216 , n54535 );
and ( n61860 , n47090 , n54533 );
nor ( n61861 , n61859 , n61860 );
xnor ( n61862 , n61861 , n54237 );
and ( n61863 , n47474 , n53928 );
and ( n61864 , n47351 , n53926 );
nor ( n61865 , n61863 , n61864 );
xnor ( n61866 , n61865 , n53652 );
and ( n61867 , n61862 , n61866 );
and ( n61868 , n47778 , n53357 );
and ( n61869 , n47647 , n53355 );
nor ( n61870 , n61868 , n61869 );
xnor ( n61871 , n61870 , n53060 );
and ( n61872 , n61866 , n61871 );
and ( n61873 , n61862 , n61871 );
or ( n61874 , n61867 , n61872 , n61873 );
and ( n61875 , n52790 , n48042 );
and ( n61876 , n52612 , n48040 );
nor ( n61877 , n61875 , n61876 );
xnor ( n61878 , n61877 , n47921 );
and ( n61879 , n54604 , n47178 );
and ( n61880 , n54227 , n47176 );
nor ( n61881 , n61879 , n61880 );
xnor ( n61882 , n61881 , n47039 );
and ( n61883 , n61878 , n61882 );
and ( n61884 , n55756 , n46712 );
and ( n61885 , n55497 , n46710 );
nor ( n61886 , n61884 , n61885 );
xnor ( n61887 , n61886 , n46587 );
and ( n61888 , n61882 , n61887 );
and ( n61889 , n61878 , n61887 );
or ( n61890 , n61883 , n61888 , n61889 );
and ( n61891 , n61874 , n61890 );
and ( n61892 , n58292 , n61481 );
not ( n61893 , n61892 );
and ( n61894 , n58628 , n61015 );
not ( n61895 , n61894 );
and ( n61896 , n61893 , n61895 );
and ( n61897 , n59615 , n59920 );
not ( n61898 , n61897 );
and ( n61899 , n61895 , n61898 );
and ( n61900 , n61893 , n61898 );
or ( n61901 , n61896 , n61899 , n61900 );
and ( n61902 , n61890 , n61901 );
and ( n61903 , n61874 , n61901 );
or ( n61904 , n61891 , n61902 , n61903 );
and ( n61905 , n53922 , n47429 );
and ( n61906 , n53639 , n47427 );
nor ( n61907 , n61905 , n61906 );
xnor ( n61908 , n61907 , n47309 );
and ( n61909 , n57063 , n46304 );
not ( n61910 , n61909 );
and ( n61911 , n61910 , n46228 );
or ( n61912 , n61908 , n61911 );
buf ( n61913 , n20217 );
buf ( n61914 , n61913 );
and ( n61915 , n57948 , n61914 );
not ( n61916 , n61915 );
buf ( n61917 , n20217 );
buf ( n61918 , n61917 );
and ( n61919 , n61918 , n58294 );
not ( n61920 , n61919 );
and ( n61921 , n61916 , n61920 );
and ( n61922 , n61912 , n61921 );
and ( n61923 , n58915 , n60711 );
not ( n61924 , n61923 );
and ( n61925 , n60821 , n58911 );
not ( n61926 , n61925 );
and ( n61927 , n61924 , n61926 );
and ( n61928 , n61921 , n61927 );
and ( n61929 , n61912 , n61927 );
or ( n61930 , n61922 , n61928 , n61929 );
and ( n61931 , n61904 , n61930 );
and ( n61932 , n46969 , n55159 );
and ( n61933 , n46843 , n55157 );
nor ( n61934 , n61932 , n61933 );
xnor ( n61935 , n61934 , n54864 );
and ( n61936 , n49115 , n51221 );
and ( n61937 , n48988 , n51219 );
nor ( n61938 , n61936 , n61937 );
xnor ( n61939 , n61938 , n51000 );
and ( n61940 , n61935 , n61939 );
and ( n61941 , n49570 , n50783 );
and ( n61942 , n49374 , n50781 );
nor ( n61943 , n61941 , n61942 );
xnor ( n61944 , n61943 , n50557 );
and ( n61945 , n61939 , n61944 );
and ( n61946 , n61935 , n61944 );
or ( n61947 , n61940 , n61945 , n61946 );
and ( n61948 , n49976 , n50338 );
and ( n61949 , n49781 , n50336 );
nor ( n61950 , n61948 , n61949 );
xnor ( n61951 , n61950 , n50111 );
and ( n61952 , n50404 , n49896 );
and ( n61953 , n50195 , n49894 );
nor ( n61954 , n61952 , n61953 );
xnor ( n61955 , n61954 , n49711 );
and ( n61956 , n61951 , n61955 );
and ( n61957 , n50726 , n49513 );
and ( n61958 , n50625 , n49511 );
nor ( n61959 , n61957 , n61958 );
xnor ( n61960 , n61959 , n49310 );
and ( n61961 , n61955 , n61960 );
and ( n61962 , n61951 , n61960 );
or ( n61963 , n61956 , n61961 , n61962 );
and ( n61964 , n61947 , n61963 );
and ( n61965 , n51298 , n49121 );
and ( n61966 , n51077 , n49119 );
nor ( n61967 , n61965 , n61966 );
xnor ( n61968 , n61967 , n48932 );
and ( n61969 , n51734 , n48740 );
and ( n61970 , n51510 , n48738 );
nor ( n61971 , n61969 , n61970 );
xnor ( n61972 , n61971 , n48571 );
and ( n61973 , n61968 , n61972 );
and ( n61974 , n52332 , n48394 );
and ( n61975 , n52082 , n48392 );
nor ( n61976 , n61974 , n61975 );
xnor ( n61977 , n61976 , n48220 );
and ( n61978 , n61972 , n61977 );
and ( n61979 , n61968 , n61977 );
or ( n61980 , n61973 , n61978 , n61979 );
and ( n61981 , n61963 , n61980 );
and ( n61982 , n61947 , n61980 );
or ( n61983 , n61964 , n61981 , n61982 );
and ( n61984 , n61930 , n61983 );
and ( n61985 , n61904 , n61983 );
or ( n61986 , n61931 , n61984 , n61985 );
and ( n61987 , n61858 , n61986 );
and ( n61988 , n53328 , n47734 );
and ( n61989 , n53041 , n47732 );
nor ( n61990 , n61988 , n61989 );
xnor ( n61991 , n61990 , n47606 );
and ( n61992 , n55143 , n46911 );
and ( n61993 , n54942 , n46909 );
nor ( n61994 , n61992 , n61993 );
xnor ( n61995 , n61994 , n46802 );
and ( n61996 , n61991 , n61995 );
and ( n61997 , n56388 , n46496 );
and ( n61998 , n56255 , n46494 );
nor ( n61999 , n61997 , n61998 );
xnor ( n62000 , n61999 , n46402 );
and ( n62001 , n61995 , n62000 );
and ( n62002 , n61991 , n62000 );
or ( n62003 , n61996 , n62001 , n62002 );
and ( n62004 , n57063 , n46306 );
and ( n62005 , n56915 , n46304 );
nor ( n62006 , n62004 , n62005 );
xnor ( n62007 , n62006 , n46228 );
xor ( n62008 , n39415 , n45566 );
buf ( n62009 , n62008 );
buf ( n62010 , n62009 );
buf ( n62011 , n62010 );
and ( n62012 , n62007 , n62011 );
and ( n62013 , n59908 , n59611 );
not ( n62014 , n62013 );
and ( n62015 , n62011 , n62014 );
and ( n62016 , n62007 , n62014 );
or ( n62017 , n62012 , n62015 , n62016 );
and ( n62018 , n62003 , n62017 );
xor ( n62019 , n61525 , n61529 );
xor ( n62020 , n62019 , n61534 );
and ( n62021 , n62017 , n62020 );
and ( n62022 , n62003 , n62020 );
or ( n62023 , n62018 , n62021 , n62022 );
xor ( n62024 , n61542 , n61546 );
xor ( n62025 , n62024 , n61551 );
xor ( n62026 , n61565 , n61569 );
xor ( n62027 , n62026 , n61574 );
and ( n62028 , n62025 , n62027 );
xor ( n62029 , n61096 , n61581 );
buf ( n62030 , n62029 );
and ( n62031 , n62027 , n62030 );
and ( n62032 , n62025 , n62030 );
or ( n62033 , n62028 , n62031 , n62032 );
and ( n62034 , n62023 , n62033 );
xor ( n62035 , n61451 , n61453 );
xor ( n62036 , n62035 , n61455 );
and ( n62037 , n62033 , n62036 );
and ( n62038 , n62023 , n62036 );
or ( n62039 , n62034 , n62037 , n62038 );
and ( n62040 , n61986 , n62039 );
and ( n62041 , n61858 , n62039 );
or ( n62042 , n61987 , n62040 , n62041 );
and ( n62043 , n61803 , n62042 );
and ( n62044 , n61764 , n62042 );
or ( n62045 , n61804 , n62043 , n62044 );
and ( n62046 , n61740 , n62045 );
and ( n62047 , n61738 , n62045 );
or ( n62048 , n61741 , n62046 , n62047 );
xor ( n62049 , n61462 , n61478 );
xor ( n62050 , n62049 , n61491 );
xor ( n62051 , n61503 , n61510 );
xor ( n62052 , n62051 , n61515 );
and ( n62053 , n62050 , n62052 );
xor ( n62054 , n61521 , n61537 );
xor ( n62055 , n62054 , n61554 );
and ( n62056 , n62052 , n62055 );
and ( n62057 , n62050 , n62055 );
or ( n62058 , n62053 , n62056 , n62057 );
xor ( n62059 , n61395 , n61396 );
xor ( n62060 , n62059 , n61398 );
and ( n62061 , n62058 , n62060 );
xor ( n62062 , n61435 , n61448 );
xor ( n62063 , n62062 , n61458 );
and ( n62064 , n62060 , n62063 );
and ( n62065 , n62058 , n62063 );
or ( n62066 , n62061 , n62064 , n62065 );
xor ( n62067 , n61494 , n61518 );
xor ( n62068 , n62067 , n61557 );
xor ( n62069 , n61589 , n61599 );
xor ( n62070 , n62069 , n61602 );
and ( n62071 , n62068 , n62070 );
xor ( n62072 , n61610 , n61612 );
xor ( n62073 , n62072 , n61615 );
and ( n62074 , n62070 , n62073 );
and ( n62075 , n62068 , n62073 );
or ( n62076 , n62071 , n62074 , n62075 );
and ( n62077 , n62066 , n62076 );
xor ( n62078 , n61386 , n61392 );
xor ( n62079 , n62078 , n61401 );
and ( n62080 , n62076 , n62079 );
and ( n62081 , n62066 , n62079 );
or ( n62082 , n62077 , n62080 , n62081 );
xor ( n62083 , n61461 , n61560 );
xor ( n62084 , n62083 , n61605 );
xor ( n62085 , n61618 , n61628 );
xor ( n62086 , n62085 , n61631 );
and ( n62087 , n62084 , n62086 );
xor ( n62088 , n61637 , n61639 );
xor ( n62089 , n62088 , n61642 );
and ( n62090 , n62086 , n62089 );
and ( n62091 , n62084 , n62089 );
or ( n62092 , n62087 , n62090 , n62091 );
and ( n62093 , n62082 , n62092 );
xor ( n62094 , n61311 , n61313 );
xor ( n62095 , n62094 , n61404 );
and ( n62096 , n62092 , n62095 );
and ( n62097 , n62082 , n62095 );
or ( n62098 , n62093 , n62096 , n62097 );
and ( n62099 , n62048 , n62098 );
xor ( n62100 , n61407 , n61648 );
xor ( n62101 , n62100 , n61667 );
and ( n62102 , n62098 , n62101 );
and ( n62103 , n62048 , n62101 );
or ( n62104 , n62099 , n62102 , n62103 );
and ( n62105 , n61736 , n62104 );
xor ( n62106 , n61670 , n61680 );
xor ( n62107 , n62106 , n61683 );
and ( n62108 , n62104 , n62107 );
and ( n62109 , n61736 , n62107 );
or ( n62110 , n62105 , n62108 , n62109 );
xor ( n62111 , n61686 , n61688 );
xor ( n62112 , n62111 , n61691 );
and ( n62113 , n62110 , n62112 );
xor ( n62114 , n61672 , n61674 );
xor ( n62115 , n62114 , n61677 );
xor ( n62116 , n61608 , n61634 );
xor ( n62117 , n62116 , n61645 );
xor ( n62118 , n61659 , n61661 );
xor ( n62119 , n62118 , n61664 );
and ( n62120 , n62117 , n62119 );
xor ( n62121 , n61651 , n61653 );
xor ( n62122 , n62121 , n61656 );
xor ( n62123 , n61620 , n61622 );
xor ( n62124 , n62123 , n61625 );
xor ( n62125 , n61761 , n61763 );
and ( n62126 , n62124 , n62125 );
xor ( n62127 , n61577 , n61583 );
xor ( n62128 , n62127 , n61586 );
xor ( n62129 , n61591 , n61593 );
xor ( n62130 , n62129 , n61596 );
and ( n62131 , n62128 , n62130 );
xor ( n62132 , n61751 , n61755 );
xor ( n62133 , n62132 , n61758 );
and ( n62134 , n62130 , n62133 );
and ( n62135 , n62128 , n62133 );
or ( n62136 , n62131 , n62134 , n62135 );
and ( n62137 , n62125 , n62136 );
and ( n62138 , n62124 , n62136 );
or ( n62139 , n62126 , n62137 , n62138 );
and ( n62140 , n62122 , n62139 );
xor ( n62141 , n61743 , n61745 );
xor ( n62142 , n62141 , n61748 );
xor ( n62143 , n61789 , n61791 );
xor ( n62144 , n62143 , n61794 );
and ( n62145 , n62142 , n62144 );
xnor ( n62146 , n61806 , n61808 );
and ( n62147 , n62144 , n62146 );
and ( n62148 , n62142 , n62146 );
or ( n62149 , n62145 , n62147 , n62148 );
buf ( n62150 , n20220 );
buf ( n62151 , n62150 );
and ( n62152 , n57948 , n62151 );
not ( n62153 , n62152 );
and ( n62154 , n58628 , n61481 );
not ( n62155 , n62154 );
and ( n62156 , n62153 , n62155 );
and ( n62157 , n59615 , n60372 );
not ( n62158 , n62157 );
and ( n62159 , n62155 , n62158 );
and ( n62160 , n62153 , n62158 );
or ( n62161 , n62156 , n62159 , n62160 );
and ( n62162 , n61918 , n58444 );
not ( n62163 , n62162 );
buf ( n62164 , n62163 );
and ( n62165 , n62161 , n62164 );
and ( n62166 , n59365 , n60372 );
not ( n62167 , n62166 );
and ( n62168 , n62164 , n62167 );
and ( n62169 , n62161 , n62167 );
or ( n62170 , n62165 , n62168 , n62169 );
and ( n62171 , n58292 , n61914 );
not ( n62172 , n62171 );
and ( n62173 , n61505 , n58542 );
not ( n62174 , n62173 );
and ( n62175 , n62172 , n62174 );
and ( n62176 , n58915 , n61015 );
not ( n62177 , n62176 );
and ( n62178 , n62174 , n62177 );
and ( n62179 , n62172 , n62177 );
or ( n62180 , n62175 , n62178 , n62179 );
xor ( n62181 , n61781 , n61783 );
xor ( n62182 , n62181 , n61786 );
and ( n62183 , n62180 , n62182 );
and ( n62184 , n62170 , n62183 );
xor ( n62185 , n61823 , n61827 );
xor ( n62186 , n62185 , n61832 );
xor ( n62187 , n61840 , n61844 );
xor ( n62188 , n62187 , n61849 );
and ( n62189 , n62186 , n62188 );
buf ( n62190 , n62189 );
and ( n62191 , n62183 , n62190 );
and ( n62192 , n62170 , n62190 );
or ( n62193 , n62184 , n62191 , n62192 );
and ( n62194 , n62149 , n62193 );
xor ( n62195 , n61862 , n61866 );
xor ( n62196 , n62195 , n61871 );
xor ( n62197 , n61878 , n61882 );
xor ( n62198 , n62197 , n61887 );
and ( n62199 , n62196 , n62198 );
xor ( n62200 , n61893 , n61895 );
xor ( n62201 , n62200 , n61898 );
and ( n62202 , n62198 , n62201 );
and ( n62203 , n62196 , n62201 );
or ( n62204 , n62199 , n62202 , n62203 );
xnor ( n62205 , n61908 , n61911 );
xor ( n62206 , n61916 , n61920 );
and ( n62207 , n62205 , n62206 );
xor ( n62208 , n61924 , n61926 );
and ( n62209 , n62206 , n62208 );
and ( n62210 , n62205 , n62208 );
or ( n62211 , n62207 , n62209 , n62210 );
and ( n62212 , n62204 , n62211 );
and ( n62213 , n47962 , n53357 );
and ( n62214 , n47778 , n53355 );
nor ( n62215 , n62213 , n62214 );
xnor ( n62216 , n62215 , n53060 );
and ( n62217 , n48272 , n52799 );
and ( n62218 , n48108 , n52797 );
nor ( n62219 , n62217 , n62218 );
xnor ( n62220 , n62219 , n52538 );
and ( n62221 , n62216 , n62220 );
and ( n62222 , n48632 , n52269 );
and ( n62223 , n48384 , n52267 );
nor ( n62224 , n62222 , n62223 );
xnor ( n62225 , n62224 , n52008 );
and ( n62226 , n62220 , n62225 );
and ( n62227 , n62216 , n62225 );
or ( n62228 , n62221 , n62226 , n62227 );
and ( n62229 , n52612 , n48394 );
and ( n62230 , n52332 , n48392 );
nor ( n62231 , n62229 , n62230 );
xnor ( n62232 , n62231 , n48220 );
and ( n62233 , n54227 , n47429 );
and ( n62234 , n53922 , n47427 );
nor ( n62235 , n62233 , n62234 );
xnor ( n62236 , n62235 , n47309 );
and ( n62237 , n62232 , n62236 );
and ( n62238 , n55497 , n46911 );
and ( n62239 , n55143 , n46909 );
nor ( n62240 , n62238 , n62239 );
xnor ( n62241 , n62240 , n46802 );
and ( n62242 , n62236 , n62241 );
and ( n62243 , n62232 , n62241 );
or ( n62244 , n62237 , n62242 , n62243 );
and ( n62245 , n62228 , n62244 );
and ( n62246 , n61008 , n58911 );
not ( n62247 , n62246 );
and ( n62248 , n62162 , n62247 );
and ( n62249 , n59365 , n60711 );
not ( n62250 , n62249 );
and ( n62251 , n62247 , n62250 );
and ( n62252 , n62162 , n62250 );
or ( n62253 , n62248 , n62251 , n62252 );
and ( n62254 , n62244 , n62253 );
and ( n62255 , n62228 , n62253 );
or ( n62256 , n62245 , n62254 , n62255 );
and ( n62257 , n62211 , n62256 );
and ( n62258 , n62204 , n62256 );
or ( n62259 , n62212 , n62257 , n62258 );
and ( n62260 , n62193 , n62259 );
and ( n62261 , n62149 , n62259 );
or ( n62262 , n62194 , n62260 , n62261 );
and ( n62263 , n46843 , n55851 );
and ( n62264 , n46750 , n55849 );
nor ( n62265 , n62263 , n62264 );
xnor ( n62266 , n62265 , n55506 );
and ( n62267 , n49781 , n50783 );
and ( n62268 , n49570 , n50781 );
nor ( n62269 , n62267 , n62268 );
xnor ( n62270 , n62269 , n50557 );
or ( n62271 , n62266 , n62270 );
and ( n62272 , n46445 , n57187 );
and ( n62273 , n46345 , n57184 );
nor ( n62274 , n62272 , n62273 );
xnor ( n62275 , n62274 , n56175 );
and ( n62276 , n46577 , n56503 );
and ( n62277 , n46530 , n56501 );
nor ( n62278 , n62276 , n62277 );
xnor ( n62279 , n62278 , n56178 );
or ( n62280 , n62275 , n62279 );
and ( n62281 , n62271 , n62280 );
and ( n62282 , n54942 , n47178 );
and ( n62283 , n54604 , n47176 );
nor ( n62284 , n62282 , n62283 );
xnor ( n62285 , n62284 , n47039 );
and ( n62286 , n62285 , n61909 );
and ( n62287 , n62280 , n62286 );
and ( n62288 , n62271 , n62286 );
or ( n62289 , n62281 , n62287 , n62288 );
and ( n62290 , n47090 , n55159 );
and ( n62291 , n46969 , n55157 );
nor ( n62292 , n62290 , n62291 );
xnor ( n62293 , n62292 , n54864 );
and ( n62294 , n47351 , n54535 );
and ( n62295 , n47216 , n54533 );
nor ( n62296 , n62294 , n62295 );
xnor ( n62297 , n62296 , n54237 );
and ( n62298 , n62293 , n62297 );
and ( n62299 , n47647 , n53928 );
and ( n62300 , n47474 , n53926 );
nor ( n62301 , n62299 , n62300 );
xnor ( n62302 , n62301 , n53652 );
and ( n62303 , n62297 , n62302 );
and ( n62304 , n62293 , n62302 );
or ( n62305 , n62298 , n62303 , n62304 );
and ( n62306 , n48988 , n51750 );
and ( n62307 , n48709 , n51748 );
nor ( n62308 , n62306 , n62307 );
xnor ( n62309 , n62308 , n51520 );
and ( n62310 , n49374 , n51221 );
and ( n62311 , n49115 , n51219 );
nor ( n62312 , n62310 , n62311 );
xnor ( n62313 , n62312 , n51000 );
and ( n62314 , n62309 , n62313 );
and ( n62315 , n50195 , n50338 );
and ( n62316 , n49976 , n50336 );
nor ( n62317 , n62315 , n62316 );
xnor ( n62318 , n62317 , n50111 );
and ( n62319 , n62313 , n62318 );
and ( n62320 , n62309 , n62318 );
or ( n62321 , n62314 , n62319 , n62320 );
and ( n62322 , n62305 , n62321 );
and ( n62323 , n50625 , n49896 );
and ( n62324 , n50404 , n49894 );
nor ( n62325 , n62323 , n62324 );
xnor ( n62326 , n62325 , n49711 );
and ( n62327 , n51077 , n49513 );
and ( n62328 , n50726 , n49511 );
nor ( n62329 , n62327 , n62328 );
xnor ( n62330 , n62329 , n49310 );
and ( n62331 , n62326 , n62330 );
and ( n62332 , n51510 , n49121 );
and ( n62333 , n51298 , n49119 );
nor ( n62334 , n62332 , n62333 );
xnor ( n62335 , n62334 , n48932 );
and ( n62336 , n62330 , n62335 );
and ( n62337 , n62326 , n62335 );
or ( n62338 , n62331 , n62336 , n62337 );
and ( n62339 , n62321 , n62338 );
and ( n62340 , n62305 , n62338 );
or ( n62341 , n62322 , n62339 , n62340 );
and ( n62342 , n62289 , n62341 );
and ( n62343 , n52082 , n48740 );
and ( n62344 , n51734 , n48738 );
nor ( n62345 , n62343 , n62344 );
xnor ( n62346 , n62345 , n48571 );
and ( n62347 , n53041 , n48042 );
and ( n62348 , n52790 , n48040 );
nor ( n62349 , n62347 , n62348 );
xnor ( n62350 , n62349 , n47921 );
and ( n62351 , n62346 , n62350 );
and ( n62352 , n53639 , n47734 );
and ( n62353 , n53328 , n47732 );
nor ( n62354 , n62352 , n62353 );
xnor ( n62355 , n62354 , n47606 );
and ( n62356 , n62350 , n62355 );
and ( n62357 , n62346 , n62355 );
or ( n62358 , n62351 , n62356 , n62357 );
and ( n62359 , n56255 , n46712 );
and ( n62360 , n55756 , n46710 );
nor ( n62361 , n62359 , n62360 );
xnor ( n62362 , n62361 , n46587 );
and ( n62363 , n56915 , n46496 );
and ( n62364 , n56388 , n46494 );
nor ( n62365 , n62363 , n62364 );
xnor ( n62366 , n62365 , n46402 );
and ( n62367 , n62362 , n62366 );
xor ( n62368 , n39418 , n45564 );
buf ( n62369 , n62368 );
buf ( n62370 , n62369 );
buf ( n62371 , n62370 );
and ( n62372 , n62366 , n62371 );
and ( n62373 , n62362 , n62371 );
or ( n62374 , n62367 , n62372 , n62373 );
and ( n62375 , n62358 , n62374 );
buf ( n62376 , n20220 );
buf ( n62377 , n62376 );
and ( n62378 , n62377 , n58294 );
not ( n62379 , n62378 );
and ( n62380 , n60821 , n59207 );
not ( n62381 , n62380 );
and ( n62382 , n62379 , n62381 );
and ( n62383 , n60376 , n59611 );
not ( n62384 , n62383 );
and ( n62385 , n62381 , n62384 );
and ( n62386 , n62379 , n62384 );
or ( n62387 , n62382 , n62385 , n62386 );
and ( n62388 , n62374 , n62387 );
and ( n62389 , n62358 , n62387 );
or ( n62390 , n62375 , n62388 , n62389 );
and ( n62391 , n62341 , n62390 );
and ( n62392 , n62289 , n62390 );
or ( n62393 , n62342 , n62391 , n62392 );
xor ( n62394 , n61935 , n61939 );
xor ( n62395 , n62394 , n61944 );
xor ( n62396 , n61951 , n61955 );
xor ( n62397 , n62396 , n61960 );
and ( n62398 , n62395 , n62397 );
xor ( n62399 , n61968 , n61972 );
xor ( n62400 , n62399 , n61977 );
and ( n62401 , n62397 , n62400 );
and ( n62402 , n62395 , n62400 );
or ( n62403 , n62398 , n62401 , n62402 );
xor ( n62404 , n61811 , n61812 );
xor ( n62405 , n62404 , n61814 );
and ( n62406 , n62403 , n62405 );
xor ( n62407 , n61819 , n61835 );
xor ( n62408 , n62407 , n61852 );
and ( n62409 , n62405 , n62408 );
and ( n62410 , n62403 , n62408 );
or ( n62411 , n62406 , n62409 , n62410 );
and ( n62412 , n62393 , n62411 );
xor ( n62413 , n61874 , n61890 );
xor ( n62414 , n62413 , n61901 );
xor ( n62415 , n61912 , n61921 );
xor ( n62416 , n62415 , n61927 );
and ( n62417 , n62414 , n62416 );
xor ( n62418 , n61947 , n61963 );
xor ( n62419 , n62418 , n61980 );
and ( n62420 , n62416 , n62419 );
and ( n62421 , n62414 , n62419 );
or ( n62422 , n62417 , n62420 , n62421 );
and ( n62423 , n62411 , n62422 );
and ( n62424 , n62393 , n62422 );
or ( n62425 , n62412 , n62423 , n62424 );
and ( n62426 , n62262 , n62425 );
xor ( n62427 , n61767 , n61769 );
xor ( n62428 , n62427 , n61772 );
xor ( n62429 , n61777 , n61778 );
xor ( n62430 , n62429 , n61797 );
and ( n62431 , n62428 , n62430 );
xor ( n62432 , n61809 , n61817 );
xor ( n62433 , n62432 , n61855 );
and ( n62434 , n62430 , n62433 );
and ( n62435 , n62428 , n62433 );
or ( n62436 , n62431 , n62434 , n62435 );
and ( n62437 , n62425 , n62436 );
and ( n62438 , n62262 , n62436 );
or ( n62439 , n62426 , n62437 , n62438 );
and ( n62440 , n62139 , n62439 );
and ( n62441 , n62122 , n62439 );
or ( n62442 , n62140 , n62440 , n62441 );
and ( n62443 , n62119 , n62442 );
and ( n62444 , n62117 , n62442 );
or ( n62445 , n62120 , n62443 , n62444 );
and ( n62446 , n62115 , n62445 );
xor ( n62447 , n61904 , n61930 );
xor ( n62448 , n62447 , n61983 );
xor ( n62449 , n62023 , n62033 );
xor ( n62450 , n62449 , n62036 );
and ( n62451 , n62448 , n62450 );
xor ( n62452 , n62050 , n62052 );
xor ( n62453 , n62452 , n62055 );
and ( n62454 , n62450 , n62453 );
and ( n62455 , n62448 , n62453 );
or ( n62456 , n62451 , n62454 , n62455 );
xor ( n62457 , n61765 , n61775 );
xor ( n62458 , n62457 , n61800 );
and ( n62459 , n62456 , n62458 );
xor ( n62460 , n61858 , n61986 );
xor ( n62461 , n62460 , n62039 );
and ( n62462 , n62458 , n62461 );
and ( n62463 , n62456 , n62461 );
or ( n62464 , n62459 , n62462 , n62463 );
xor ( n62465 , n61764 , n61803 );
xor ( n62466 , n62465 , n62042 );
and ( n62467 , n62464 , n62466 );
xor ( n62468 , n62066 , n62076 );
xor ( n62469 , n62468 , n62079 );
and ( n62470 , n62466 , n62469 );
and ( n62471 , n62464 , n62469 );
or ( n62472 , n62467 , n62470 , n62471 );
xor ( n62473 , n61738 , n61740 );
xor ( n62474 , n62473 , n62045 );
and ( n62475 , n62472 , n62474 );
xor ( n62476 , n62082 , n62092 );
xor ( n62477 , n62476 , n62095 );
and ( n62478 , n62474 , n62477 );
and ( n62479 , n62472 , n62477 );
or ( n62480 , n62475 , n62478 , n62479 );
and ( n62481 , n62445 , n62480 );
and ( n62482 , n62115 , n62480 );
or ( n62483 , n62446 , n62481 , n62482 );
xor ( n62484 , n61736 , n62104 );
xor ( n62485 , n62484 , n62107 );
and ( n62486 , n62483 , n62485 );
xor ( n62487 , n62048 , n62098 );
xor ( n62488 , n62487 , n62101 );
xor ( n62489 , n62084 , n62086 );
xor ( n62490 , n62489 , n62089 );
xor ( n62491 , n62058 , n62060 );
xor ( n62492 , n62491 , n62063 );
xor ( n62493 , n62068 , n62070 );
xor ( n62494 , n62493 , n62073 );
and ( n62495 , n62492 , n62494 );
xor ( n62496 , n62003 , n62017 );
xor ( n62497 , n62496 , n62020 );
xor ( n62498 , n62025 , n62027 );
xor ( n62499 , n62498 , n62030 );
and ( n62500 , n62497 , n62499 );
xor ( n62501 , n61991 , n61995 );
xor ( n62502 , n62501 , n62000 );
xor ( n62503 , n62007 , n62011 );
xor ( n62504 , n62503 , n62014 );
and ( n62505 , n62502 , n62504 );
xor ( n62506 , n62180 , n62182 );
and ( n62507 , n62504 , n62506 );
and ( n62508 , n62502 , n62506 );
or ( n62509 , n62505 , n62507 , n62508 );
and ( n62510 , n62499 , n62509 );
and ( n62511 , n62497 , n62509 );
or ( n62512 , n62500 , n62510 , n62511 );
xor ( n62513 , n62216 , n62220 );
xor ( n62514 , n62513 , n62225 );
xor ( n62515 , n62232 , n62236 );
xor ( n62516 , n62515 , n62241 );
and ( n62517 , n62514 , n62516 );
buf ( n62518 , n62517 );
xor ( n62519 , n62153 , n62155 );
xor ( n62520 , n62519 , n62158 );
xor ( n62521 , n62172 , n62174 );
xor ( n62522 , n62521 , n62177 );
and ( n62523 , n62520 , n62522 );
xor ( n62524 , n62162 , n62247 );
xor ( n62525 , n62524 , n62250 );
and ( n62526 , n62522 , n62525 );
and ( n62527 , n62520 , n62525 );
or ( n62528 , n62523 , n62526 , n62527 );
and ( n62529 , n62518 , n62528 );
xnor ( n62530 , n62266 , n62270 );
xnor ( n62531 , n62275 , n62279 );
and ( n62532 , n62530 , n62531 );
xor ( n62533 , n62285 , n61909 );
and ( n62534 , n62531 , n62533 );
and ( n62535 , n62530 , n62533 );
or ( n62536 , n62532 , n62534 , n62535 );
and ( n62537 , n62528 , n62536 );
and ( n62538 , n62518 , n62536 );
or ( n62539 , n62529 , n62537 , n62538 );
and ( n62540 , n47474 , n54535 );
and ( n62541 , n47351 , n54533 );
nor ( n62542 , n62540 , n62541 );
xnor ( n62543 , n62542 , n54237 );
and ( n62544 , n47778 , n53928 );
and ( n62545 , n47647 , n53926 );
nor ( n62546 , n62544 , n62545 );
xnor ( n62547 , n62546 , n53652 );
and ( n62548 , n62543 , n62547 );
and ( n62549 , n48108 , n53357 );
and ( n62550 , n47962 , n53355 );
nor ( n62551 , n62549 , n62550 );
xnor ( n62552 , n62551 , n53060 );
and ( n62553 , n62547 , n62552 );
and ( n62554 , n62543 , n62552 );
or ( n62555 , n62548 , n62553 , n62554 );
and ( n62556 , n46969 , n55851 );
and ( n62557 , n46843 , n55849 );
nor ( n62558 , n62556 , n62557 );
xnor ( n62559 , n62558 , n55506 );
and ( n62560 , n47216 , n55159 );
and ( n62561 , n47090 , n55157 );
nor ( n62562 , n62560 , n62561 );
xnor ( n62563 , n62562 , n54864 );
and ( n62564 , n62559 , n62563 );
and ( n62565 , n49976 , n50783 );
and ( n62566 , n49781 , n50781 );
nor ( n62567 , n62565 , n62566 );
xnor ( n62568 , n62567 , n50557 );
and ( n62569 , n62563 , n62568 );
and ( n62570 , n62559 , n62568 );
or ( n62571 , n62564 , n62569 , n62570 );
and ( n62572 , n62555 , n62571 );
and ( n62573 , n54604 , n47429 );
and ( n62574 , n54227 , n47427 );
nor ( n62575 , n62573 , n62574 );
xnor ( n62576 , n62575 , n47309 );
and ( n62577 , n55143 , n47178 );
and ( n62578 , n54942 , n47176 );
nor ( n62579 , n62577 , n62578 );
xnor ( n62580 , n62579 , n47039 );
and ( n62581 , n62576 , n62580 );
and ( n62582 , n55756 , n46911 );
and ( n62583 , n55497 , n46909 );
nor ( n62584 , n62582 , n62583 );
xnor ( n62585 , n62584 , n46802 );
and ( n62586 , n62580 , n62585 );
and ( n62587 , n62576 , n62585 );
or ( n62588 , n62581 , n62586 , n62587 );
and ( n62589 , n62571 , n62588 );
and ( n62590 , n62555 , n62588 );
or ( n62591 , n62572 , n62589 , n62590 );
buf ( n62592 , n20223 );
buf ( n62593 , n62592 );
and ( n62594 , n62593 , n58294 );
not ( n62595 , n62594 );
and ( n62596 , n58292 , n62151 );
not ( n62597 , n62596 );
and ( n62598 , n62595 , n62597 );
and ( n62599 , n58915 , n61481 );
not ( n62600 , n62599 );
and ( n62601 , n62597 , n62600 );
and ( n62602 , n62595 , n62600 );
or ( n62603 , n62598 , n62601 , n62602 );
and ( n62604 , n48384 , n52799 );
and ( n62605 , n48272 , n52797 );
nor ( n62606 , n62604 , n62605 );
xnor ( n62607 , n62606 , n52538 );
and ( n62608 , n48709 , n52269 );
and ( n62609 , n48632 , n52267 );
nor ( n62610 , n62608 , n62609 );
xnor ( n62611 , n62610 , n52008 );
or ( n62612 , n62607 , n62611 );
and ( n62613 , n62603 , n62612 );
and ( n62614 , n62377 , n58444 );
not ( n62615 , n62614 );
and ( n62616 , n61505 , n58911 );
not ( n62617 , n62616 );
or ( n62618 , n62615 , n62617 );
and ( n62619 , n62612 , n62618 );
and ( n62620 , n62603 , n62618 );
or ( n62621 , n62613 , n62619 , n62620 );
and ( n62622 , n62591 , n62621 );
and ( n62623 , n61918 , n58542 );
not ( n62624 , n62623 );
and ( n62625 , n60376 , n59920 );
not ( n62626 , n62625 );
or ( n62627 , n62624 , n62626 );
and ( n62628 , n52790 , n48394 );
and ( n62629 , n52612 , n48392 );
nor ( n62630 , n62628 , n62629 );
xnor ( n62631 , n62630 , n48220 );
and ( n62632 , n53328 , n48042 );
and ( n62633 , n53041 , n48040 );
nor ( n62634 , n62632 , n62633 );
xnor ( n62635 , n62634 , n47921 );
and ( n62636 , n62631 , n62635 );
and ( n62637 , n62627 , n62636 );
and ( n62638 , n46530 , n57187 );
and ( n62639 , n46445 , n57184 );
nor ( n62640 , n62638 , n62639 );
xnor ( n62641 , n62640 , n56175 );
and ( n62642 , n46750 , n56503 );
and ( n62643 , n46577 , n56501 );
nor ( n62644 , n62642 , n62643 );
xnor ( n62645 , n62644 , n56178 );
and ( n62646 , n62641 , n62645 );
and ( n62647 , n49115 , n51750 );
and ( n62648 , n48988 , n51748 );
nor ( n62649 , n62647 , n62648 );
xnor ( n62650 , n62649 , n51520 );
and ( n62651 , n62645 , n62650 );
and ( n62652 , n62641 , n62650 );
or ( n62653 , n62646 , n62651 , n62652 );
and ( n62654 , n62636 , n62653 );
and ( n62655 , n62627 , n62653 );
or ( n62656 , n62637 , n62654 , n62655 );
and ( n62657 , n62621 , n62656 );
and ( n62658 , n62591 , n62656 );
or ( n62659 , n62622 , n62657 , n62658 );
and ( n62660 , n62539 , n62659 );
and ( n62661 , n49570 , n51221 );
and ( n62662 , n49374 , n51219 );
nor ( n62663 , n62661 , n62662 );
xnor ( n62664 , n62663 , n51000 );
and ( n62665 , n51298 , n49513 );
and ( n62666 , n51077 , n49511 );
nor ( n62667 , n62665 , n62666 );
xnor ( n62668 , n62667 , n49310 );
and ( n62669 , n62664 , n62668 );
and ( n62670 , n51734 , n49121 );
and ( n62671 , n51510 , n49119 );
nor ( n62672 , n62670 , n62671 );
xnor ( n62673 , n62672 , n48932 );
and ( n62674 , n62668 , n62673 );
and ( n62675 , n62664 , n62673 );
or ( n62676 , n62669 , n62674 , n62675 );
and ( n62677 , n52332 , n48740 );
and ( n62678 , n52082 , n48738 );
nor ( n62679 , n62677 , n62678 );
xnor ( n62680 , n62679 , n48571 );
and ( n62681 , n53922 , n47734 );
and ( n62682 , n53639 , n47732 );
nor ( n62683 , n62681 , n62682 );
xnor ( n62684 , n62683 , n47606 );
and ( n62685 , n62680 , n62684 );
and ( n62686 , n56388 , n46712 );
and ( n62687 , n56255 , n46710 );
nor ( n62688 , n62686 , n62687 );
xnor ( n62689 , n62688 , n46587 );
and ( n62690 , n62684 , n62689 );
and ( n62691 , n62680 , n62689 );
or ( n62692 , n62685 , n62690 , n62691 );
and ( n62693 , n62676 , n62692 );
and ( n62694 , n57063 , n46496 );
and ( n62695 , n56915 , n46494 );
nor ( n62696 , n62694 , n62695 );
xnor ( n62697 , n62696 , n46402 );
and ( n62698 , n57063 , n46494 );
not ( n62699 , n62698 );
and ( n62700 , n62699 , n46402 );
and ( n62701 , n62697 , n62700 );
xor ( n62702 , n40494 , n45562 );
buf ( n62703 , n62702 );
buf ( n62704 , n62703 );
buf ( n62705 , n62704 );
and ( n62706 , n62700 , n62705 );
and ( n62707 , n62697 , n62705 );
or ( n62708 , n62701 , n62706 , n62707 );
and ( n62709 , n62692 , n62708 );
and ( n62710 , n62676 , n62708 );
or ( n62711 , n62693 , n62709 , n62710 );
xor ( n62712 , n62293 , n62297 );
xor ( n62713 , n62712 , n62302 );
xor ( n62714 , n62309 , n62313 );
xor ( n62715 , n62714 , n62318 );
and ( n62716 , n62713 , n62715 );
xor ( n62717 , n62326 , n62330 );
xor ( n62718 , n62717 , n62335 );
and ( n62719 , n62715 , n62718 );
and ( n62720 , n62713 , n62718 );
or ( n62721 , n62716 , n62719 , n62720 );
and ( n62722 , n62711 , n62721 );
xor ( n62723 , n62346 , n62350 );
xor ( n62724 , n62723 , n62355 );
xor ( n62725 , n62362 , n62366 );
xor ( n62726 , n62725 , n62371 );
and ( n62727 , n62724 , n62726 );
xor ( n62728 , n62379 , n62381 );
xor ( n62729 , n62728 , n62384 );
and ( n62730 , n62726 , n62729 );
and ( n62731 , n62724 , n62729 );
or ( n62732 , n62727 , n62730 , n62731 );
and ( n62733 , n62721 , n62732 );
and ( n62734 , n62711 , n62732 );
or ( n62735 , n62722 , n62733 , n62734 );
and ( n62736 , n62659 , n62735 );
and ( n62737 , n62539 , n62735 );
or ( n62738 , n62660 , n62736 , n62737 );
and ( n62739 , n62512 , n62738 );
buf ( n62740 , n62186 );
xor ( n62741 , n62740 , n62188 );
xor ( n62742 , n62196 , n62198 );
xor ( n62743 , n62742 , n62201 );
and ( n62744 , n62741 , n62743 );
xor ( n62745 , n62205 , n62206 );
xor ( n62746 , n62745 , n62208 );
and ( n62747 , n62743 , n62746 );
and ( n62748 , n62741 , n62746 );
or ( n62749 , n62744 , n62747 , n62748 );
xor ( n62750 , n62228 , n62244 );
xor ( n62751 , n62750 , n62253 );
xor ( n62752 , n62271 , n62280 );
xor ( n62753 , n62752 , n62286 );
and ( n62754 , n62751 , n62753 );
xor ( n62755 , n62305 , n62321 );
xor ( n62756 , n62755 , n62338 );
and ( n62757 , n62753 , n62756 );
and ( n62758 , n62751 , n62756 );
or ( n62759 , n62754 , n62757 , n62758 );
and ( n62760 , n62749 , n62759 );
xor ( n62761 , n62142 , n62144 );
xor ( n62762 , n62761 , n62146 );
and ( n62763 , n62759 , n62762 );
and ( n62764 , n62749 , n62762 );
or ( n62765 , n62760 , n62763 , n62764 );
and ( n62766 , n62738 , n62765 );
and ( n62767 , n62512 , n62765 );
or ( n62768 , n62739 , n62766 , n62767 );
and ( n62769 , n62494 , n62768 );
and ( n62770 , n62492 , n62768 );
or ( n62771 , n62495 , n62769 , n62770 );
and ( n62772 , n62490 , n62771 );
xor ( n62773 , n62170 , n62183 );
xor ( n62774 , n62773 , n62190 );
xor ( n62775 , n62204 , n62211 );
xor ( n62776 , n62775 , n62256 );
and ( n62777 , n62774 , n62776 );
xor ( n62778 , n62289 , n62341 );
xor ( n62779 , n62778 , n62390 );
and ( n62780 , n62776 , n62779 );
and ( n62781 , n62774 , n62779 );
or ( n62782 , n62777 , n62780 , n62781 );
xor ( n62783 , n62128 , n62130 );
xor ( n62784 , n62783 , n62133 );
and ( n62785 , n62782 , n62784 );
xor ( n62786 , n62149 , n62193 );
xor ( n62787 , n62786 , n62259 );
and ( n62788 , n62784 , n62787 );
and ( n62789 , n62782 , n62787 );
or ( n62790 , n62785 , n62788 , n62789 );
xor ( n62791 , n62393 , n62411 );
xor ( n62792 , n62791 , n62422 );
xor ( n62793 , n62428 , n62430 );
xor ( n62794 , n62793 , n62433 );
and ( n62795 , n62792 , n62794 );
xor ( n62796 , n62448 , n62450 );
xor ( n62797 , n62796 , n62453 );
and ( n62798 , n62794 , n62797 );
and ( n62799 , n62792 , n62797 );
or ( n62800 , n62795 , n62798 , n62799 );
and ( n62801 , n62790 , n62800 );
xor ( n62802 , n62124 , n62125 );
xor ( n62803 , n62802 , n62136 );
and ( n62804 , n62800 , n62803 );
and ( n62805 , n62790 , n62803 );
or ( n62806 , n62801 , n62804 , n62805 );
and ( n62807 , n62771 , n62806 );
and ( n62808 , n62490 , n62806 );
or ( n62809 , n62772 , n62807 , n62808 );
xor ( n62810 , n62117 , n62119 );
xor ( n62811 , n62810 , n62442 );
and ( n62812 , n62809 , n62811 );
xor ( n62813 , n62472 , n62474 );
xor ( n62814 , n62813 , n62477 );
and ( n62815 , n62811 , n62814 );
and ( n62816 , n62809 , n62814 );
or ( n62817 , n62812 , n62815 , n62816 );
and ( n62818 , n62488 , n62817 );
xor ( n62819 , n62115 , n62445 );
xor ( n62820 , n62819 , n62480 );
and ( n62821 , n62817 , n62820 );
and ( n62822 , n62488 , n62820 );
or ( n62823 , n62818 , n62821 , n62822 );
and ( n62824 , n62485 , n62823 );
and ( n62825 , n62483 , n62823 );
or ( n62826 , n62486 , n62824 , n62825 );
and ( n62827 , n62112 , n62826 );
and ( n62828 , n62110 , n62826 );
or ( n62829 , n62113 , n62827 , n62828 );
or ( n62830 , n61734 , n62829 );
and ( n62831 , n61732 , n62830 );
xor ( n62832 , n61732 , n62830 );
xnor ( n62833 , n61734 , n62829 );
xor ( n62834 , n62110 , n62112 );
xor ( n62835 , n62834 , n62826 );
not ( n62836 , n62835 );
xor ( n62837 , n62483 , n62485 );
xor ( n62838 , n62837 , n62823 );
xor ( n62839 , n62488 , n62817 );
xor ( n62840 , n62839 , n62820 );
xor ( n62841 , n62122 , n62139 );
xor ( n62842 , n62841 , n62439 );
xor ( n62843 , n62464 , n62466 );
xor ( n62844 , n62843 , n62469 );
and ( n62845 , n62842 , n62844 );
xor ( n62846 , n62262 , n62425 );
xor ( n62847 , n62846 , n62436 );
xor ( n62848 , n62456 , n62458 );
xor ( n62849 , n62848 , n62461 );
and ( n62850 , n62847 , n62849 );
xor ( n62851 , n62403 , n62405 );
xor ( n62852 , n62851 , n62408 );
xor ( n62853 , n62414 , n62416 );
xor ( n62854 , n62853 , n62419 );
and ( n62855 , n62852 , n62854 );
and ( n62856 , n58915 , n61914 );
not ( n62857 , n62856 );
buf ( n62858 , n62857 );
and ( n62859 , n59365 , n61015 );
not ( n62860 , n62859 );
and ( n62861 , n62858 , n62860 );
and ( n62862 , n59615 , n60711 );
not ( n62863 , n62862 );
and ( n62864 , n62860 , n62863 );
and ( n62865 , n62858 , n62863 );
or ( n62866 , n62861 , n62864 , n62865 );
buf ( n62867 , n20223 );
buf ( n62868 , n62867 );
and ( n62869 , n57948 , n62868 );
not ( n62870 , n62869 );
and ( n62871 , n58628 , n61914 );
not ( n62872 , n62871 );
and ( n62873 , n62870 , n62872 );
and ( n62874 , n59908 , n60372 );
not ( n62875 , n62874 );
and ( n62876 , n62872 , n62875 );
and ( n62877 , n62870 , n62875 );
or ( n62878 , n62873 , n62876 , n62877 );
and ( n62879 , n62866 , n62878 );
buf ( n62880 , n59908 );
not ( n62881 , n62880 );
and ( n62882 , n62878 , n62881 );
and ( n62883 , n62866 , n62881 );
or ( n62884 , n62879 , n62882 , n62883 );
xor ( n62885 , n62161 , n62164 );
xor ( n62886 , n62885 , n62167 );
or ( n62887 , n62884 , n62886 );
and ( n62888 , n62854 , n62887 );
and ( n62889 , n62852 , n62887 );
or ( n62890 , n62855 , n62888 , n62889 );
xor ( n62891 , n62358 , n62374 );
xor ( n62892 , n62891 , n62387 );
xor ( n62893 , n62395 , n62397 );
xor ( n62894 , n62893 , n62400 );
and ( n62895 , n62892 , n62894 );
and ( n62896 , n48632 , n52799 );
and ( n62897 , n48384 , n52797 );
nor ( n62898 , n62896 , n62897 );
xnor ( n62899 , n62898 , n52538 );
and ( n62900 , n48988 , n52269 );
and ( n62901 , n48709 , n52267 );
nor ( n62902 , n62900 , n62901 );
xnor ( n62903 , n62902 , n52008 );
and ( n62904 , n62899 , n62903 );
and ( n62905 , n50195 , n50783 );
and ( n62906 , n49976 , n50781 );
nor ( n62907 , n62905 , n62906 );
xnor ( n62908 , n62907 , n50557 );
and ( n62909 , n62903 , n62908 );
and ( n62910 , n62899 , n62908 );
or ( n62911 , n62904 , n62909 , n62910 );
and ( n62912 , n46843 , n56503 );
and ( n62913 , n46750 , n56501 );
nor ( n62914 , n62912 , n62913 );
xnor ( n62915 , n62914 , n56178 );
and ( n62916 , n47090 , n55851 );
and ( n62917 , n46969 , n55849 );
nor ( n62918 , n62916 , n62917 );
xnor ( n62919 , n62918 , n55506 );
and ( n62920 , n62915 , n62919 );
and ( n62921 , n47351 , n55159 );
and ( n62922 , n47216 , n55157 );
nor ( n62923 , n62921 , n62922 );
xnor ( n62924 , n62923 , n54864 );
and ( n62925 , n62919 , n62924 );
and ( n62926 , n62915 , n62924 );
or ( n62927 , n62920 , n62925 , n62926 );
and ( n62928 , n62911 , n62927 );
and ( n62929 , n50726 , n49896 );
and ( n62930 , n50625 , n49894 );
nor ( n62931 , n62929 , n62930 );
xnor ( n62932 , n62931 , n49711 );
and ( n62933 , n62927 , n62932 );
and ( n62934 , n62911 , n62932 );
or ( n62935 , n62928 , n62933 , n62934 );
and ( n62936 , n50404 , n50338 );
and ( n62937 , n50195 , n50336 );
nor ( n62938 , n62936 , n62937 );
xnor ( n62939 , n62938 , n50111 );
xor ( n62940 , n62543 , n62547 );
xor ( n62941 , n62940 , n62552 );
and ( n62942 , n62939 , n62941 );
and ( n62943 , n62935 , n62942 );
and ( n62944 , n60821 , n59611 );
not ( n62945 , n62944 );
xor ( n62946 , n62559 , n62563 );
xor ( n62947 , n62946 , n62568 );
and ( n62948 , n62945 , n62947 );
buf ( n62949 , n62948 );
and ( n62950 , n62942 , n62949 );
and ( n62951 , n62935 , n62949 );
or ( n62952 , n62943 , n62950 , n62951 );
and ( n62953 , n62894 , n62952 );
and ( n62954 , n62892 , n62952 );
or ( n62955 , n62895 , n62953 , n62954 );
xor ( n62956 , n62576 , n62580 );
xor ( n62957 , n62956 , n62585 );
xnor ( n62958 , n62607 , n62611 );
and ( n62959 , n62957 , n62958 );
xnor ( n62960 , n62615 , n62617 );
and ( n62961 , n62958 , n62960 );
and ( n62962 , n62957 , n62960 );
or ( n62963 , n62959 , n62961 , n62962 );
xnor ( n62964 , n62624 , n62626 );
xor ( n62965 , n62631 , n62635 );
and ( n62966 , n62964 , n62965 );
and ( n62967 , n53041 , n48394 );
and ( n62968 , n52790 , n48392 );
nor ( n62969 , n62967 , n62968 );
xnor ( n62970 , n62969 , n48220 );
and ( n62971 , n54942 , n47429 );
and ( n62972 , n54604 , n47427 );
nor ( n62973 , n62971 , n62972 );
xnor ( n62974 , n62973 , n47309 );
and ( n62975 , n62970 , n62974 );
and ( n62976 , n56915 , n46712 );
and ( n62977 , n56388 , n46710 );
nor ( n62978 , n62976 , n62977 );
xnor ( n62979 , n62978 , n46587 );
and ( n62980 , n62974 , n62979 );
and ( n62981 , n62970 , n62979 );
or ( n62982 , n62975 , n62980 , n62981 );
and ( n62983 , n62965 , n62982 );
and ( n62984 , n62964 , n62982 );
or ( n62985 , n62966 , n62983 , n62984 );
and ( n62986 , n62963 , n62985 );
and ( n62987 , n58292 , n62868 );
not ( n62988 , n62987 );
and ( n62989 , n59615 , n61015 );
not ( n62990 , n62989 );
and ( n62991 , n62988 , n62990 );
buf ( n62992 , n60376 );
not ( n62993 , n62992 );
and ( n62994 , n62990 , n62993 );
and ( n62995 , n62988 , n62993 );
or ( n62996 , n62991 , n62994 , n62995 );
buf ( n62997 , n20226 );
buf ( n62998 , n62997 );
and ( n62999 , n57948 , n62998 );
not ( n63000 , n62999 );
and ( n63001 , n62377 , n58542 );
not ( n63002 , n63001 );
and ( n63003 , n63000 , n63002 );
and ( n63004 , n63002 , n62856 );
and ( n63005 , n63000 , n62856 );
or ( n63006 , n63003 , n63004 , n63005 );
and ( n63007 , n62996 , n63006 );
and ( n63008 , n46577 , n57187 );
and ( n63009 , n46530 , n57184 );
nor ( n63010 , n63008 , n63009 );
xnor ( n63011 , n63010 , n56175 );
and ( n63012 , n48272 , n53357 );
and ( n63013 , n48108 , n53355 );
nor ( n63014 , n63012 , n63013 );
xnor ( n63015 , n63014 , n53060 );
and ( n63016 , n63011 , n63015 );
and ( n63017 , n63006 , n63016 );
and ( n63018 , n62996 , n63016 );
or ( n63019 , n63007 , n63017 , n63018 );
and ( n63020 , n62985 , n63019 );
and ( n63021 , n62963 , n63019 );
or ( n63022 , n62986 , n63020 , n63021 );
buf ( n63023 , n20226 );
buf ( n63024 , n63023 );
and ( n63025 , n63024 , n58294 );
not ( n63026 , n63025 );
and ( n63027 , n61505 , n59207 );
not ( n63028 , n63027 );
and ( n63029 , n63026 , n63028 );
and ( n63030 , n47647 , n54535 );
and ( n63031 , n47474 , n54533 );
nor ( n63032 , n63030 , n63031 );
xnor ( n63033 , n63032 , n54237 );
and ( n63034 , n47962 , n53928 );
and ( n63035 , n47778 , n53926 );
nor ( n63036 , n63034 , n63035 );
xnor ( n63037 , n63036 , n53652 );
and ( n63038 , n63033 , n63037 );
and ( n63039 , n49374 , n51750 );
and ( n63040 , n49115 , n51748 );
nor ( n63041 , n63039 , n63040 );
xnor ( n63042 , n63041 , n51520 );
and ( n63043 , n63037 , n63042 );
and ( n63044 , n63033 , n63042 );
or ( n63045 , n63038 , n63043 , n63044 );
and ( n63046 , n63029 , n63045 );
and ( n63047 , n49781 , n51221 );
and ( n63048 , n49570 , n51219 );
nor ( n63049 , n63047 , n63048 );
xnor ( n63050 , n63049 , n51000 );
and ( n63051 , n50625 , n50338 );
and ( n63052 , n50404 , n50336 );
nor ( n63053 , n63051 , n63052 );
xnor ( n63054 , n63053 , n50111 );
and ( n63055 , n63050 , n63054 );
and ( n63056 , n51510 , n49513 );
and ( n63057 , n51298 , n49511 );
nor ( n63058 , n63056 , n63057 );
xnor ( n63059 , n63058 , n49310 );
and ( n63060 , n63054 , n63059 );
and ( n63061 , n63050 , n63059 );
or ( n63062 , n63055 , n63060 , n63061 );
and ( n63063 , n63045 , n63062 );
and ( n63064 , n63029 , n63062 );
or ( n63065 , n63046 , n63063 , n63064 );
and ( n63066 , n52082 , n49121 );
and ( n63067 , n51734 , n49119 );
nor ( n63068 , n63066 , n63067 );
xnor ( n63069 , n63068 , n48932 );
and ( n63070 , n52612 , n48740 );
and ( n63071 , n52332 , n48738 );
nor ( n63072 , n63070 , n63071 );
xnor ( n63073 , n63072 , n48571 );
and ( n63074 , n63069 , n63073 );
and ( n63075 , n53639 , n48042 );
and ( n63076 , n53328 , n48040 );
nor ( n63077 , n63075 , n63076 );
xnor ( n63078 , n63077 , n47921 );
and ( n63079 , n63073 , n63078 );
and ( n63080 , n63069 , n63078 );
or ( n63081 , n63074 , n63079 , n63080 );
and ( n63082 , n54227 , n47734 );
and ( n63083 , n53922 , n47732 );
nor ( n63084 , n63082 , n63083 );
xnor ( n63085 , n63084 , n47606 );
and ( n63086 , n55497 , n47178 );
and ( n63087 , n55143 , n47176 );
nor ( n63088 , n63086 , n63087 );
xnor ( n63089 , n63088 , n47039 );
and ( n63090 , n63085 , n63089 );
and ( n63091 , n56255 , n46911 );
and ( n63092 , n55756 , n46909 );
nor ( n63093 , n63091 , n63092 );
xnor ( n63094 , n63093 , n46802 );
and ( n63095 , n63089 , n63094 );
and ( n63096 , n63085 , n63094 );
or ( n63097 , n63090 , n63095 , n63096 );
and ( n63098 , n63081 , n63097 );
xor ( n63099 , n40497 , n45560 );
buf ( n63100 , n63099 );
buf ( n63101 , n63100 );
buf ( n63102 , n63101 );
and ( n63103 , n62698 , n63102 );
and ( n63104 , n62593 , n58444 );
not ( n63105 , n63104 );
and ( n63106 , n63102 , n63105 );
and ( n63107 , n62698 , n63105 );
or ( n63108 , n63103 , n63106 , n63107 );
and ( n63109 , n63097 , n63108 );
and ( n63110 , n63081 , n63108 );
or ( n63111 , n63098 , n63109 , n63110 );
and ( n63112 , n63065 , n63111 );
xor ( n63113 , n62641 , n62645 );
xor ( n63114 , n63113 , n62650 );
xor ( n63115 , n62664 , n62668 );
xor ( n63116 , n63115 , n62673 );
and ( n63117 , n63114 , n63116 );
xor ( n63118 , n62680 , n62684 );
xor ( n63119 , n63118 , n62689 );
and ( n63120 , n63116 , n63119 );
and ( n63121 , n63114 , n63119 );
or ( n63122 , n63117 , n63120 , n63121 );
and ( n63123 , n63111 , n63122 );
and ( n63124 , n63065 , n63122 );
or ( n63125 , n63112 , n63123 , n63124 );
and ( n63126 , n63022 , n63125 );
buf ( n63127 , n62514 );
xor ( n63128 , n63127 , n62516 );
xor ( n63129 , n62520 , n62522 );
xor ( n63130 , n63129 , n62525 );
and ( n63131 , n63128 , n63130 );
xor ( n63132 , n62530 , n62531 );
xor ( n63133 , n63132 , n62533 );
and ( n63134 , n63130 , n63133 );
and ( n63135 , n63128 , n63133 );
or ( n63136 , n63131 , n63134 , n63135 );
and ( n63137 , n63125 , n63136 );
and ( n63138 , n63022 , n63136 );
or ( n63139 , n63126 , n63137 , n63138 );
and ( n63140 , n62955 , n63139 );
xor ( n63141 , n62555 , n62571 );
xor ( n63142 , n63141 , n62588 );
xor ( n63143 , n62603 , n62612 );
xor ( n63144 , n63143 , n62618 );
and ( n63145 , n63142 , n63144 );
xor ( n63146 , n62627 , n62636 );
xor ( n63147 , n63146 , n62653 );
and ( n63148 , n63144 , n63147 );
and ( n63149 , n63142 , n63147 );
or ( n63150 , n63145 , n63148 , n63149 );
xor ( n63151 , n62676 , n62692 );
xor ( n63152 , n63151 , n62708 );
xor ( n63153 , n62713 , n62715 );
xor ( n63154 , n63153 , n62718 );
and ( n63155 , n63152 , n63154 );
xor ( n63156 , n62724 , n62726 );
xor ( n63157 , n63156 , n62729 );
and ( n63158 , n63154 , n63157 );
and ( n63159 , n63152 , n63157 );
or ( n63160 , n63155 , n63158 , n63159 );
and ( n63161 , n63150 , n63160 );
xor ( n63162 , n62502 , n62504 );
xor ( n63163 , n63162 , n62506 );
and ( n63164 , n63160 , n63163 );
and ( n63165 , n63150 , n63163 );
or ( n63166 , n63161 , n63164 , n63165 );
and ( n63167 , n63139 , n63166 );
and ( n63168 , n62955 , n63166 );
or ( n63169 , n63140 , n63167 , n63168 );
and ( n63170 , n62890 , n63169 );
xor ( n63171 , n62518 , n62528 );
xor ( n63172 , n63171 , n62536 );
xor ( n63173 , n62591 , n62621 );
xor ( n63174 , n63173 , n62656 );
and ( n63175 , n63172 , n63174 );
xor ( n63176 , n62711 , n62721 );
xor ( n63177 , n63176 , n62732 );
and ( n63178 , n63174 , n63177 );
and ( n63179 , n63172 , n63177 );
or ( n63180 , n63175 , n63178 , n63179 );
xor ( n63181 , n62497 , n62499 );
xor ( n63182 , n63181 , n62509 );
and ( n63183 , n63180 , n63182 );
xor ( n63184 , n62539 , n62659 );
xor ( n63185 , n63184 , n62735 );
and ( n63186 , n63182 , n63185 );
and ( n63187 , n63180 , n63185 );
or ( n63188 , n63183 , n63186 , n63187 );
and ( n63189 , n63169 , n63188 );
and ( n63190 , n62890 , n63188 );
or ( n63191 , n63170 , n63189 , n63190 );
and ( n63192 , n62849 , n63191 );
and ( n63193 , n62847 , n63191 );
or ( n63194 , n62850 , n63192 , n63193 );
and ( n63195 , n62844 , n63194 );
and ( n63196 , n62842 , n63194 );
or ( n63197 , n62845 , n63195 , n63196 );
xor ( n63198 , n62809 , n62811 );
xor ( n63199 , n63198 , n62814 );
and ( n63200 , n63197 , n63199 );
xor ( n63201 , n62512 , n62738 );
xor ( n63202 , n63201 , n62765 );
xor ( n63203 , n62782 , n62784 );
xor ( n63204 , n63203 , n62787 );
and ( n63205 , n63202 , n63204 );
xor ( n63206 , n62792 , n62794 );
xor ( n63207 , n63206 , n62797 );
and ( n63208 , n63204 , n63207 );
and ( n63209 , n63202 , n63207 );
or ( n63210 , n63205 , n63208 , n63209 );
xor ( n63211 , n62492 , n62494 );
xor ( n63212 , n63211 , n62768 );
and ( n63213 , n63210 , n63212 );
xor ( n63214 , n62790 , n62800 );
xor ( n63215 , n63214 , n62803 );
and ( n63216 , n63212 , n63215 );
and ( n63217 , n63210 , n63215 );
or ( n63218 , n63213 , n63216 , n63217 );
xor ( n63219 , n62490 , n62771 );
xor ( n63220 , n63219 , n62806 );
and ( n63221 , n63218 , n63220 );
xor ( n63222 , n62749 , n62759 );
xor ( n63223 , n63222 , n62762 );
xor ( n63224 , n62774 , n62776 );
xor ( n63225 , n63224 , n62779 );
and ( n63226 , n63223 , n63225 );
xor ( n63227 , n62741 , n62743 );
xor ( n63228 , n63227 , n62746 );
xor ( n63229 , n62751 , n62753 );
xor ( n63230 , n63229 , n62756 );
and ( n63231 , n63228 , n63230 );
xnor ( n63232 , n62884 , n62886 );
and ( n63233 , n63230 , n63232 );
and ( n63234 , n63228 , n63232 );
or ( n63235 , n63231 , n63233 , n63234 );
and ( n63236 , n63225 , n63235 );
and ( n63237 , n63223 , n63235 );
or ( n63238 , n63226 , n63236 , n63237 );
xor ( n63239 , n62866 , n62878 );
xor ( n63240 , n63239 , n62881 );
and ( n63241 , n58292 , n62998 );
not ( n63242 , n63241 );
and ( n63243 , n58628 , n62868 );
not ( n63244 , n63243 );
and ( n63245 , n63242 , n63244 );
and ( n63246 , n59615 , n61481 );
not ( n63247 , n63246 );
and ( n63248 , n63244 , n63247 );
and ( n63249 , n63242 , n63247 );
or ( n63250 , n63245 , n63248 , n63249 );
and ( n63251 , n59365 , n61481 );
not ( n63252 , n63251 );
and ( n63253 , n63250 , n63252 );
and ( n63254 , n59908 , n60711 );
not ( n63255 , n63254 );
and ( n63256 , n63252 , n63255 );
and ( n63257 , n63250 , n63255 );
or ( n63258 , n63253 , n63256 , n63257 );
xor ( n63259 , n62858 , n62860 );
xor ( n63260 , n63259 , n62863 );
and ( n63261 , n63258 , n63260 );
xor ( n63262 , n62870 , n62872 );
xor ( n63263 , n63262 , n62875 );
and ( n63264 , n63260 , n63263 );
and ( n63265 , n63258 , n63263 );
or ( n63266 , n63261 , n63264 , n63265 );
and ( n63267 , n63240 , n63266 );
and ( n63268 , n63024 , n58444 );
not ( n63269 , n63268 );
and ( n63270 , n62593 , n58542 );
not ( n63271 , n63270 );
and ( n63272 , n63269 , n63271 );
and ( n63273 , n58628 , n62151 );
not ( n63274 , n63273 );
and ( n63275 , n63272 , n63274 );
and ( n63276 , n61008 , n59611 );
not ( n63277 , n63276 );
and ( n63278 , n63274 , n63277 );
and ( n63279 , n63272 , n63277 );
or ( n63280 , n63275 , n63278 , n63279 );
and ( n63281 , n61008 , n59207 );
not ( n63282 , n63281 );
and ( n63283 , n63280 , n63282 );
xor ( n63284 , n62595 , n62597 );
xor ( n63285 , n63284 , n62600 );
and ( n63286 , n63282 , n63285 );
and ( n63287 , n63280 , n63285 );
or ( n63288 , n63283 , n63286 , n63287 );
and ( n63289 , n63266 , n63288 );
and ( n63290 , n63240 , n63288 );
or ( n63291 , n63267 , n63289 , n63290 );
xor ( n63292 , n62697 , n62700 );
xor ( n63293 , n63292 , n62705 );
xor ( n63294 , n62911 , n62927 );
xor ( n63295 , n63294 , n62932 );
and ( n63296 , n63293 , n63295 );
xor ( n63297 , n62939 , n62941 );
and ( n63298 , n63295 , n63297 );
and ( n63299 , n63293 , n63297 );
or ( n63300 , n63296 , n63298 , n63299 );
and ( n63301 , n47778 , n54535 );
and ( n63302 , n47647 , n54533 );
nor ( n63303 , n63301 , n63302 );
xnor ( n63304 , n63303 , n54237 );
and ( n63305 , n48108 , n53928 );
and ( n63306 , n47962 , n53926 );
nor ( n63307 , n63305 , n63306 );
xnor ( n63308 , n63307 , n53652 );
and ( n63309 , n63304 , n63308 );
and ( n63310 , n48384 , n53357 );
and ( n63311 , n48272 , n53355 );
nor ( n63312 , n63310 , n63311 );
xnor ( n63313 , n63312 , n53060 );
and ( n63314 , n63308 , n63313 );
and ( n63315 , n63304 , n63313 );
or ( n63316 , n63309 , n63314 , n63315 );
and ( n63317 , n46969 , n56503 );
and ( n63318 , n46843 , n56501 );
nor ( n63319 , n63317 , n63318 );
xnor ( n63320 , n63319 , n56178 );
and ( n63321 , n47216 , n55851 );
and ( n63322 , n47090 , n55849 );
nor ( n63323 , n63321 , n63322 );
xnor ( n63324 , n63323 , n55506 );
and ( n63325 , n63320 , n63324 );
and ( n63326 , n47474 , n55159 );
and ( n63327 , n47351 , n55157 );
nor ( n63328 , n63326 , n63327 );
xnor ( n63329 , n63328 , n54864 );
and ( n63330 , n63324 , n63329 );
and ( n63331 , n63320 , n63329 );
or ( n63332 , n63325 , n63330 , n63331 );
and ( n63333 , n63316 , n63332 );
and ( n63334 , n51077 , n49896 );
and ( n63335 , n50726 , n49894 );
nor ( n63336 , n63334 , n63335 );
xnor ( n63337 , n63336 , n49711 );
and ( n63338 , n63332 , n63337 );
and ( n63339 , n63316 , n63337 );
or ( n63340 , n63333 , n63338 , n63339 );
and ( n63341 , n61918 , n58911 );
not ( n63342 , n63341 );
xor ( n63343 , n62899 , n62903 );
xor ( n63344 , n63343 , n62908 );
and ( n63345 , n63342 , n63344 );
buf ( n63346 , n63345 );
and ( n63347 , n63340 , n63346 );
xor ( n63348 , n62915 , n62919 );
xor ( n63349 , n63348 , n62924 );
xor ( n63350 , n62970 , n62974 );
xor ( n63351 , n63350 , n62979 );
and ( n63352 , n63349 , n63351 );
xor ( n63353 , n63000 , n63002 );
xor ( n63354 , n63353 , n62856 );
and ( n63355 , n63351 , n63354 );
and ( n63356 , n63349 , n63354 );
or ( n63357 , n63352 , n63355 , n63356 );
and ( n63358 , n63346 , n63357 );
and ( n63359 , n63340 , n63357 );
or ( n63360 , n63347 , n63358 , n63359 );
and ( n63361 , n63300 , n63360 );
xor ( n63362 , n63011 , n63015 );
xor ( n63363 , n63026 , n63028 );
and ( n63364 , n63362 , n63363 );
and ( n63365 , n53922 , n48042 );
and ( n63366 , n53639 , n48040 );
nor ( n63367 , n63365 , n63366 );
xnor ( n63368 , n63367 , n47921 );
and ( n63369 , n56388 , n46911 );
and ( n63370 , n56255 , n46909 );
nor ( n63371 , n63369 , n63370 );
xnor ( n63372 , n63371 , n46802 );
and ( n63373 , n63368 , n63372 );
and ( n63374 , n57063 , n46712 );
and ( n63375 , n56915 , n46710 );
nor ( n63376 , n63374 , n63375 );
xnor ( n63377 , n63376 , n46587 );
and ( n63378 , n63372 , n63377 );
and ( n63379 , n63368 , n63377 );
or ( n63380 , n63373 , n63378 , n63379 );
and ( n63381 , n63363 , n63380 );
and ( n63382 , n63362 , n63380 );
or ( n63383 , n63364 , n63381 , n63382 );
and ( n63384 , n59365 , n61914 );
not ( n63385 , n63384 );
and ( n63386 , n59908 , n61015 );
not ( n63387 , n63386 );
and ( n63388 , n63385 , n63387 );
and ( n63389 , n60376 , n60711 );
not ( n63390 , n63389 );
and ( n63391 , n63387 , n63390 );
and ( n63392 , n63385 , n63390 );
or ( n63393 , n63388 , n63391 , n63392 );
and ( n63394 , n48709 , n52799 );
and ( n63395 , n48632 , n52797 );
nor ( n63396 , n63394 , n63395 );
xnor ( n63397 , n63396 , n52538 );
and ( n63398 , n50404 , n50783 );
and ( n63399 , n50195 , n50781 );
nor ( n63400 , n63398 , n63399 );
xnor ( n63401 , n63400 , n50557 );
and ( n63402 , n63397 , n63401 );
and ( n63403 , n63393 , n63402 );
and ( n63404 , n46750 , n57187 );
and ( n63405 , n46577 , n57184 );
nor ( n63406 , n63404 , n63405 );
xnor ( n63407 , n63406 , n56175 );
and ( n63408 , n49115 , n52269 );
and ( n63409 , n48988 , n52267 );
nor ( n63410 , n63408 , n63409 );
xnor ( n63411 , n63410 , n52008 );
and ( n63412 , n63407 , n63411 );
and ( n63413 , n49570 , n51750 );
and ( n63414 , n49374 , n51748 );
nor ( n63415 , n63413 , n63414 );
xnor ( n63416 , n63415 , n51520 );
and ( n63417 , n63411 , n63416 );
and ( n63418 , n63407 , n63416 );
or ( n63419 , n63412 , n63417 , n63418 );
and ( n63420 , n63402 , n63419 );
and ( n63421 , n63393 , n63419 );
or ( n63422 , n63403 , n63420 , n63421 );
and ( n63423 , n63383 , n63422 );
and ( n63424 , n49976 , n51221 );
and ( n63425 , n49781 , n51219 );
nor ( n63426 , n63424 , n63425 );
xnor ( n63427 , n63426 , n51000 );
and ( n63428 , n50726 , n50338 );
and ( n63429 , n50625 , n50336 );
nor ( n63430 , n63428 , n63429 );
xnor ( n63431 , n63430 , n50111 );
and ( n63432 , n63427 , n63431 );
and ( n63433 , n51734 , n49513 );
and ( n63434 , n51510 , n49511 );
nor ( n63435 , n63433 , n63434 );
xnor ( n63436 , n63435 , n49310 );
and ( n63437 , n63431 , n63436 );
and ( n63438 , n63427 , n63436 );
or ( n63439 , n63432 , n63437 , n63438 );
and ( n63440 , n52332 , n49121 );
and ( n63441 , n52082 , n49119 );
nor ( n63442 , n63440 , n63441 );
xnor ( n63443 , n63442 , n48932 );
and ( n63444 , n52790 , n48740 );
and ( n63445 , n52612 , n48738 );
nor ( n63446 , n63444 , n63445 );
xnor ( n63447 , n63446 , n48571 );
and ( n63448 , n63443 , n63447 );
and ( n63449 , n53328 , n48394 );
and ( n63450 , n53041 , n48392 );
nor ( n63451 , n63449 , n63450 );
xnor ( n63452 , n63451 , n48220 );
and ( n63453 , n63447 , n63452 );
and ( n63454 , n63443 , n63452 );
or ( n63455 , n63448 , n63453 , n63454 );
and ( n63456 , n63439 , n63455 );
and ( n63457 , n54604 , n47734 );
and ( n63458 , n54227 , n47732 );
nor ( n63459 , n63457 , n63458 );
xnor ( n63460 , n63459 , n47606 );
and ( n63461 , n55143 , n47429 );
and ( n63462 , n54942 , n47427 );
nor ( n63463 , n63461 , n63462 );
xnor ( n63464 , n63463 , n47309 );
and ( n63465 , n63460 , n63464 );
and ( n63466 , n55756 , n47178 );
and ( n63467 , n55497 , n47176 );
nor ( n63468 , n63466 , n63467 );
xnor ( n63469 , n63468 , n47039 );
and ( n63470 , n63464 , n63469 );
and ( n63471 , n63460 , n63469 );
or ( n63472 , n63465 , n63470 , n63471 );
and ( n63473 , n63455 , n63472 );
and ( n63474 , n63439 , n63472 );
or ( n63475 , n63456 , n63473 , n63474 );
and ( n63476 , n63422 , n63475 );
and ( n63477 , n63383 , n63475 );
or ( n63478 , n63423 , n63476 , n63477 );
and ( n63479 , n63360 , n63478 );
and ( n63480 , n63300 , n63478 );
or ( n63481 , n63361 , n63479 , n63480 );
and ( n63482 , n63291 , n63481 );
and ( n63483 , n57063 , n46710 );
not ( n63484 , n63483 );
and ( n63485 , n63484 , n46587 );
xor ( n63486 , n40498 , n45559 );
buf ( n63487 , n63486 );
buf ( n63488 , n63487 );
buf ( n63489 , n63488 );
and ( n63490 , n63485 , n63489 );
buf ( n63491 , n20229 );
buf ( n63492 , n63491 );
and ( n63493 , n63492 , n58294 );
not ( n63494 , n63493 );
and ( n63495 , n63489 , n63494 );
and ( n63496 , n63485 , n63494 );
or ( n63497 , n63490 , n63495 , n63496 );
and ( n63498 , n62377 , n58911 );
not ( n63499 , n63498 );
and ( n63500 , n61918 , n59207 );
not ( n63501 , n63500 );
and ( n63502 , n63499 , n63501 );
and ( n63503 , n60821 , n60372 );
not ( n63504 , n63503 );
and ( n63505 , n63501 , n63504 );
and ( n63506 , n63499 , n63504 );
or ( n63507 , n63502 , n63505 , n63506 );
and ( n63508 , n63497 , n63507 );
xor ( n63509 , n63033 , n63037 );
xor ( n63510 , n63509 , n63042 );
and ( n63511 , n63507 , n63510 );
and ( n63512 , n63497 , n63510 );
or ( n63513 , n63508 , n63511 , n63512 );
xor ( n63514 , n63050 , n63054 );
xor ( n63515 , n63514 , n63059 );
xor ( n63516 , n63069 , n63073 );
xor ( n63517 , n63516 , n63078 );
and ( n63518 , n63515 , n63517 );
xor ( n63519 , n63085 , n63089 );
xor ( n63520 , n63519 , n63094 );
and ( n63521 , n63517 , n63520 );
and ( n63522 , n63515 , n63520 );
or ( n63523 , n63518 , n63521 , n63522 );
and ( n63524 , n63513 , n63523 );
buf ( n63525 , n62945 );
xor ( n63526 , n63525 , n62947 );
and ( n63527 , n63523 , n63526 );
and ( n63528 , n63513 , n63526 );
or ( n63529 , n63524 , n63527 , n63528 );
xor ( n63530 , n62957 , n62958 );
xor ( n63531 , n63530 , n62960 );
xor ( n63532 , n62964 , n62965 );
xor ( n63533 , n63532 , n62982 );
and ( n63534 , n63531 , n63533 );
xor ( n63535 , n62996 , n63006 );
xor ( n63536 , n63535 , n63016 );
and ( n63537 , n63533 , n63536 );
and ( n63538 , n63531 , n63536 );
or ( n63539 , n63534 , n63537 , n63538 );
and ( n63540 , n63529 , n63539 );
xor ( n63541 , n63029 , n63045 );
xor ( n63542 , n63541 , n63062 );
xor ( n63543 , n63081 , n63097 );
xor ( n63544 , n63543 , n63108 );
and ( n63545 , n63542 , n63544 );
xor ( n63546 , n63114 , n63116 );
xor ( n63547 , n63546 , n63119 );
and ( n63548 , n63544 , n63547 );
and ( n63549 , n63542 , n63547 );
or ( n63550 , n63545 , n63548 , n63549 );
and ( n63551 , n63539 , n63550 );
and ( n63552 , n63529 , n63550 );
or ( n63553 , n63540 , n63551 , n63552 );
and ( n63554 , n63481 , n63553 );
and ( n63555 , n63291 , n63553 );
or ( n63556 , n63482 , n63554 , n63555 );
xor ( n63557 , n62935 , n62942 );
xor ( n63558 , n63557 , n62949 );
xor ( n63559 , n62963 , n62985 );
xor ( n63560 , n63559 , n63019 );
and ( n63561 , n63558 , n63560 );
xor ( n63562 , n63065 , n63111 );
xor ( n63563 , n63562 , n63122 );
and ( n63564 , n63560 , n63563 );
and ( n63565 , n63558 , n63563 );
or ( n63566 , n63561 , n63564 , n63565 );
xor ( n63567 , n63128 , n63130 );
xor ( n63568 , n63567 , n63133 );
xor ( n63569 , n63142 , n63144 );
xor ( n63570 , n63569 , n63147 );
and ( n63571 , n63568 , n63570 );
xor ( n63572 , n63152 , n63154 );
xor ( n63573 , n63572 , n63157 );
and ( n63574 , n63570 , n63573 );
and ( n63575 , n63568 , n63573 );
or ( n63576 , n63571 , n63574 , n63575 );
and ( n63577 , n63566 , n63576 );
xor ( n63578 , n62892 , n62894 );
xor ( n63579 , n63578 , n62952 );
and ( n63580 , n63576 , n63579 );
and ( n63581 , n63566 , n63579 );
or ( n63582 , n63577 , n63580 , n63581 );
and ( n63583 , n63556 , n63582 );
xor ( n63584 , n63022 , n63125 );
xor ( n63585 , n63584 , n63136 );
xor ( n63586 , n63150 , n63160 );
xor ( n63587 , n63586 , n63163 );
and ( n63588 , n63585 , n63587 );
xor ( n63589 , n63172 , n63174 );
xor ( n63590 , n63589 , n63177 );
and ( n63591 , n63587 , n63590 );
and ( n63592 , n63585 , n63590 );
or ( n63593 , n63588 , n63591 , n63592 );
and ( n63594 , n63582 , n63593 );
and ( n63595 , n63556 , n63593 );
or ( n63596 , n63583 , n63594 , n63595 );
and ( n63597 , n63238 , n63596 );
xor ( n63598 , n62852 , n62854 );
xor ( n63599 , n63598 , n62887 );
xor ( n63600 , n62955 , n63139 );
xor ( n63601 , n63600 , n63166 );
and ( n63602 , n63599 , n63601 );
xor ( n63603 , n63180 , n63182 );
xor ( n63604 , n63603 , n63185 );
and ( n63605 , n63601 , n63604 );
and ( n63606 , n63599 , n63604 );
or ( n63607 , n63602 , n63605 , n63606 );
and ( n63608 , n63596 , n63607 );
and ( n63609 , n63238 , n63607 );
or ( n63610 , n63597 , n63608 , n63609 );
xor ( n63611 , n62847 , n62849 );
xor ( n63612 , n63611 , n63191 );
and ( n63613 , n63610 , n63612 );
xor ( n63614 , n63210 , n63212 );
xor ( n63615 , n63614 , n63215 );
and ( n63616 , n63612 , n63615 );
and ( n63617 , n63610 , n63615 );
or ( n63618 , n63613 , n63616 , n63617 );
and ( n63619 , n63220 , n63618 );
and ( n63620 , n63218 , n63618 );
or ( n63621 , n63221 , n63619 , n63620 );
and ( n63622 , n63199 , n63621 );
and ( n63623 , n63197 , n63621 );
or ( n63624 , n63200 , n63622 , n63623 );
and ( n63625 , n62840 , n63624 );
xor ( n63626 , n63197 , n63199 );
xor ( n63627 , n63626 , n63621 );
xor ( n63628 , n62842 , n62844 );
xor ( n63629 , n63628 , n63194 );
xor ( n63630 , n63218 , n63220 );
xor ( n63631 , n63630 , n63618 );
and ( n63632 , n63629 , n63631 );
xor ( n63633 , n62890 , n63169 );
xor ( n63634 , n63633 , n63188 );
xor ( n63635 , n63202 , n63204 );
xor ( n63636 , n63635 , n63207 );
and ( n63637 , n63634 , n63636 );
xor ( n63638 , n63258 , n63260 );
xor ( n63639 , n63638 , n63263 );
xor ( n63640 , n63280 , n63282 );
xor ( n63641 , n63640 , n63285 );
and ( n63642 , n63639 , n63641 );
xor ( n63643 , n63269 , n63271 );
and ( n63644 , n58915 , n62151 );
not ( n63645 , n63644 );
and ( n63646 , n63643 , n63645 );
and ( n63647 , n61008 , n59920 );
not ( n63648 , n63647 );
and ( n63649 , n63645 , n63648 );
and ( n63650 , n63643 , n63648 );
or ( n63651 , n63646 , n63649 , n63650 );
and ( n63652 , n60821 , n59920 );
not ( n63653 , n63652 );
and ( n63654 , n63651 , n63653 );
xor ( n63655 , n63272 , n63274 );
xor ( n63656 , n63655 , n63277 );
and ( n63657 , n63653 , n63656 );
and ( n63658 , n63651 , n63656 );
or ( n63659 , n63654 , n63657 , n63658 );
and ( n63660 , n63641 , n63659 );
and ( n63661 , n63639 , n63659 );
or ( n63662 , n63642 , n63660 , n63661 );
xor ( n63663 , n62698 , n63102 );
xor ( n63664 , n63663 , n63105 );
xor ( n63665 , n63316 , n63332 );
xor ( n63666 , n63665 , n63337 );
and ( n63667 , n63664 , n63666 );
and ( n63668 , n63492 , n58444 );
not ( n63669 , n63668 );
and ( n63670 , n63024 , n58542 );
not ( n63671 , n63670 );
and ( n63672 , n63669 , n63671 );
and ( n63673 , n58915 , n62868 );
not ( n63674 , n63673 );
and ( n63675 , n63671 , n63674 );
and ( n63676 , n63669 , n63674 );
or ( n63677 , n63672 , n63675 , n63676 );
buf ( n63678 , n20229 );
buf ( n63679 , n63678 );
and ( n63680 , n57948 , n63679 );
not ( n63681 , n63680 );
and ( n63682 , n63677 , n63681 );
and ( n63683 , n61505 , n59611 );
not ( n63684 , n63683 );
and ( n63685 , n63681 , n63684 );
and ( n63686 , n63677 , n63684 );
or ( n63687 , n63682 , n63685 , n63686 );
and ( n63688 , n63666 , n63687 );
and ( n63689 , n63664 , n63687 );
or ( n63690 , n63667 , n63688 , n63689 );
and ( n63691 , n46843 , n57187 );
and ( n63692 , n46750 , n57184 );
nor ( n63693 , n63691 , n63692 );
xnor ( n63694 , n63693 , n56175 );
and ( n63695 , n47090 , n56503 );
and ( n63696 , n46969 , n56501 );
nor ( n63697 , n63695 , n63696 );
xnor ( n63698 , n63697 , n56178 );
and ( n63699 , n63694 , n63698 );
and ( n63700 , n50625 , n50783 );
and ( n63701 , n50404 , n50781 );
nor ( n63702 , n63700 , n63701 );
xnor ( n63703 , n63702 , n50557 );
and ( n63704 , n63698 , n63703 );
and ( n63705 , n63694 , n63703 );
or ( n63706 , n63699 , n63704 , n63705 );
and ( n63707 , n51298 , n49896 );
and ( n63708 , n51077 , n49894 );
nor ( n63709 , n63707 , n63708 );
xnor ( n63710 , n63709 , n49711 );
and ( n63711 , n63706 , n63710 );
xor ( n63712 , n63304 , n63308 );
xor ( n63713 , n63712 , n63313 );
xor ( n63714 , n63320 , n63324 );
xor ( n63715 , n63714 , n63329 );
and ( n63716 , n63713 , n63715 );
buf ( n63717 , n63716 );
and ( n63718 , n63711 , n63717 );
xor ( n63719 , n63368 , n63372 );
xor ( n63720 , n63719 , n63377 );
xor ( n63721 , n63385 , n63387 );
xor ( n63722 , n63721 , n63390 );
and ( n63723 , n63720 , n63722 );
xor ( n63724 , n63397 , n63401 );
and ( n63725 , n63722 , n63724 );
and ( n63726 , n63720 , n63724 );
or ( n63727 , n63723 , n63725 , n63726 );
and ( n63728 , n63717 , n63727 );
and ( n63729 , n63711 , n63727 );
or ( n63730 , n63718 , n63728 , n63729 );
and ( n63731 , n63690 , n63730 );
and ( n63732 , n47962 , n54535 );
and ( n63733 , n47778 , n54533 );
nor ( n63734 , n63732 , n63733 );
xnor ( n63735 , n63734 , n54237 );
and ( n63736 , n48272 , n53928 );
and ( n63737 , n48108 , n53926 );
nor ( n63738 , n63736 , n63737 );
xnor ( n63739 , n63738 , n53652 );
and ( n63740 , n63735 , n63739 );
and ( n63741 , n48632 , n53357 );
and ( n63742 , n48384 , n53355 );
nor ( n63743 , n63741 , n63742 );
xnor ( n63744 , n63743 , n53060 );
and ( n63745 , n63739 , n63744 );
and ( n63746 , n63735 , n63744 );
or ( n63747 , n63740 , n63745 , n63746 );
and ( n63748 , n53639 , n48394 );
and ( n63749 , n53328 , n48392 );
nor ( n63750 , n63748 , n63749 );
xnor ( n63751 , n63750 , n48220 );
and ( n63752 , n56255 , n47178 );
and ( n63753 , n55756 , n47176 );
nor ( n63754 , n63752 , n63753 );
xnor ( n63755 , n63754 , n47039 );
and ( n63756 , n63751 , n63755 );
and ( n63757 , n56915 , n46911 );
and ( n63758 , n56388 , n46909 );
nor ( n63759 , n63757 , n63758 );
xnor ( n63760 , n63759 , n46802 );
and ( n63761 , n63755 , n63760 );
and ( n63762 , n63751 , n63760 );
or ( n63763 , n63756 , n63761 , n63762 );
and ( n63764 , n63747 , n63763 );
buf ( n63765 , n20232 );
buf ( n63766 , n63765 );
and ( n63767 , n57948 , n63766 );
not ( n63768 , n63767 );
and ( n63769 , n59615 , n61914 );
not ( n63770 , n63769 );
and ( n63771 , n63768 , n63770 );
and ( n63772 , n59908 , n61481 );
not ( n63773 , n63772 );
and ( n63774 , n63770 , n63773 );
and ( n63775 , n63768 , n63773 );
or ( n63776 , n63771 , n63774 , n63775 );
and ( n63777 , n63763 , n63776 );
and ( n63778 , n63747 , n63776 );
or ( n63779 , n63764 , n63777 , n63778 );
and ( n63780 , n47351 , n55851 );
and ( n63781 , n47216 , n55849 );
nor ( n63782 , n63780 , n63781 );
xnor ( n63783 , n63782 , n55506 );
and ( n63784 , n47647 , n55159 );
and ( n63785 , n47474 , n55157 );
nor ( n63786 , n63784 , n63785 );
xnor ( n63787 , n63786 , n54864 );
and ( n63788 , n63783 , n63787 );
and ( n63789 , n48988 , n52799 );
and ( n63790 , n48709 , n52797 );
nor ( n63791 , n63789 , n63790 );
xnor ( n63792 , n63791 , n52538 );
and ( n63793 , n63787 , n63792 );
and ( n63794 , n63783 , n63792 );
or ( n63795 , n63788 , n63793 , n63794 );
and ( n63796 , n49374 , n52269 );
and ( n63797 , n49115 , n52267 );
nor ( n63798 , n63796 , n63797 );
xnor ( n63799 , n63798 , n52008 );
and ( n63800 , n49781 , n51750 );
and ( n63801 , n49570 , n51748 );
nor ( n63802 , n63800 , n63801 );
xnor ( n63803 , n63802 , n51520 );
and ( n63804 , n63799 , n63803 );
and ( n63805 , n50195 , n51221 );
and ( n63806 , n49976 , n51219 );
nor ( n63807 , n63805 , n63806 );
xnor ( n63808 , n63807 , n51000 );
and ( n63809 , n63803 , n63808 );
and ( n63810 , n63799 , n63808 );
or ( n63811 , n63804 , n63809 , n63810 );
and ( n63812 , n63795 , n63811 );
and ( n63813 , n52082 , n49513 );
and ( n63814 , n51734 , n49511 );
nor ( n63815 , n63813 , n63814 );
xnor ( n63816 , n63815 , n49310 );
and ( n63817 , n52612 , n49121 );
and ( n63818 , n52332 , n49119 );
nor ( n63819 , n63817 , n63818 );
xnor ( n63820 , n63819 , n48932 );
and ( n63821 , n63816 , n63820 );
and ( n63822 , n53041 , n48740 );
and ( n63823 , n52790 , n48738 );
nor ( n63824 , n63822 , n63823 );
xnor ( n63825 , n63824 , n48571 );
and ( n63826 , n63820 , n63825 );
and ( n63827 , n63816 , n63825 );
or ( n63828 , n63821 , n63826 , n63827 );
and ( n63829 , n63811 , n63828 );
and ( n63830 , n63795 , n63828 );
or ( n63831 , n63812 , n63829 , n63830 );
and ( n63832 , n63779 , n63831 );
and ( n63833 , n54227 , n48042 );
and ( n63834 , n53922 , n48040 );
nor ( n63835 , n63833 , n63834 );
xnor ( n63836 , n63835 , n47921 );
and ( n63837 , n54942 , n47734 );
and ( n63838 , n54604 , n47732 );
nor ( n63839 , n63837 , n63838 );
xnor ( n63840 , n63839 , n47606 );
and ( n63841 , n63836 , n63840 );
and ( n63842 , n55497 , n47429 );
and ( n63843 , n55143 , n47427 );
nor ( n63844 , n63842 , n63843 );
xnor ( n63845 , n63844 , n47309 );
and ( n63846 , n63840 , n63845 );
and ( n63847 , n63836 , n63845 );
or ( n63848 , n63841 , n63846 , n63847 );
xor ( n63849 , n40500 , n45558 );
buf ( n63850 , n63849 );
buf ( n63851 , n63850 );
buf ( n63852 , n63851 );
and ( n63853 , n63483 , n63852 );
buf ( n63854 , n63853 );
and ( n63855 , n63848 , n63854 );
xor ( n63856 , n63407 , n63411 );
xor ( n63857 , n63856 , n63416 );
and ( n63858 , n63854 , n63857 );
and ( n63859 , n63848 , n63857 );
or ( n63860 , n63855 , n63858 , n63859 );
and ( n63861 , n63831 , n63860 );
and ( n63862 , n63779 , n63860 );
or ( n63863 , n63832 , n63861 , n63862 );
and ( n63864 , n63730 , n63863 );
and ( n63865 , n63690 , n63863 );
or ( n63866 , n63731 , n63864 , n63865 );
and ( n63867 , n63662 , n63866 );
xor ( n63868 , n63427 , n63431 );
xor ( n63869 , n63868 , n63436 );
xor ( n63870 , n63443 , n63447 );
xor ( n63871 , n63870 , n63452 );
and ( n63872 , n63869 , n63871 );
xor ( n63873 , n63460 , n63464 );
xor ( n63874 , n63873 , n63469 );
and ( n63875 , n63871 , n63874 );
and ( n63876 , n63869 , n63874 );
or ( n63877 , n63872 , n63875 , n63876 );
buf ( n63878 , n63342 );
xor ( n63879 , n63878 , n63344 );
and ( n63880 , n63877 , n63879 );
xor ( n63881 , n63349 , n63351 );
xor ( n63882 , n63881 , n63354 );
and ( n63883 , n63879 , n63882 );
and ( n63884 , n63877 , n63882 );
or ( n63885 , n63880 , n63883 , n63884 );
xor ( n63886 , n63362 , n63363 );
xor ( n63887 , n63886 , n63380 );
xor ( n63888 , n63393 , n63402 );
xor ( n63889 , n63888 , n63419 );
and ( n63890 , n63887 , n63889 );
xor ( n63891 , n63439 , n63455 );
xor ( n63892 , n63891 , n63472 );
and ( n63893 , n63889 , n63892 );
and ( n63894 , n63887 , n63892 );
or ( n63895 , n63890 , n63893 , n63894 );
and ( n63896 , n63885 , n63895 );
xor ( n63897 , n63293 , n63295 );
xor ( n63898 , n63897 , n63297 );
and ( n63899 , n63895 , n63898 );
and ( n63900 , n63885 , n63898 );
or ( n63901 , n63896 , n63899 , n63900 );
and ( n63902 , n63866 , n63901 );
and ( n63903 , n63662 , n63901 );
or ( n63904 , n63867 , n63902 , n63903 );
xor ( n63905 , n63340 , n63346 );
xor ( n63906 , n63905 , n63357 );
xor ( n63907 , n63383 , n63422 );
xor ( n63908 , n63907 , n63475 );
and ( n63909 , n63906 , n63908 );
xor ( n63910 , n63513 , n63523 );
xor ( n63911 , n63910 , n63526 );
and ( n63912 , n63908 , n63911 );
and ( n63913 , n63906 , n63911 );
or ( n63914 , n63909 , n63912 , n63913 );
xor ( n63915 , n63240 , n63266 );
xor ( n63916 , n63915 , n63288 );
and ( n63917 , n63914 , n63916 );
xor ( n63918 , n63300 , n63360 );
xor ( n63919 , n63918 , n63478 );
and ( n63920 , n63916 , n63919 );
and ( n63921 , n63914 , n63919 );
or ( n63922 , n63917 , n63920 , n63921 );
and ( n63923 , n63904 , n63922 );
xor ( n63924 , n63529 , n63539 );
xor ( n63925 , n63924 , n63550 );
xor ( n63926 , n63558 , n63560 );
xor ( n63927 , n63926 , n63563 );
and ( n63928 , n63925 , n63927 );
xor ( n63929 , n63568 , n63570 );
xor ( n63930 , n63929 , n63573 );
and ( n63931 , n63927 , n63930 );
and ( n63932 , n63925 , n63930 );
or ( n63933 , n63928 , n63931 , n63932 );
and ( n63934 , n63922 , n63933 );
and ( n63935 , n63904 , n63933 );
or ( n63936 , n63923 , n63934 , n63935 );
xor ( n63937 , n63228 , n63230 );
xor ( n63938 , n63937 , n63232 );
xor ( n63939 , n63291 , n63481 );
xor ( n63940 , n63939 , n63553 );
and ( n63941 , n63938 , n63940 );
xor ( n63942 , n63566 , n63576 );
xor ( n63943 , n63942 , n63579 );
and ( n63944 , n63940 , n63943 );
and ( n63945 , n63938 , n63943 );
or ( n63946 , n63941 , n63944 , n63945 );
and ( n63947 , n63936 , n63946 );
xor ( n63948 , n63223 , n63225 );
xor ( n63949 , n63948 , n63235 );
and ( n63950 , n63946 , n63949 );
and ( n63951 , n63936 , n63949 );
or ( n63952 , n63947 , n63950 , n63951 );
and ( n63953 , n63636 , n63952 );
and ( n63954 , n63634 , n63952 );
or ( n63955 , n63637 , n63953 , n63954 );
xor ( n63956 , n63610 , n63612 );
xor ( n63957 , n63956 , n63615 );
and ( n63958 , n63955 , n63957 );
xor ( n63959 , n63238 , n63596 );
xor ( n63960 , n63959 , n63607 );
xor ( n63961 , n63556 , n63582 );
xor ( n63962 , n63961 , n63593 );
xor ( n63963 , n63599 , n63601 );
xor ( n63964 , n63963 , n63604 );
and ( n63965 , n63962 , n63964 );
xor ( n63966 , n63585 , n63587 );
xor ( n63967 , n63966 , n63590 );
xor ( n63968 , n63531 , n63533 );
xor ( n63969 , n63968 , n63536 );
xor ( n63970 , n63542 , n63544 );
xor ( n63971 , n63970 , n63547 );
and ( n63972 , n63969 , n63971 );
xor ( n63973 , n63497 , n63507 );
xor ( n63974 , n63973 , n63510 );
xor ( n63975 , n63515 , n63517 );
xor ( n63976 , n63975 , n63520 );
and ( n63977 , n63974 , n63976 );
xor ( n63978 , n63651 , n63653 );
xor ( n63979 , n63978 , n63656 );
and ( n63980 , n63976 , n63979 );
and ( n63981 , n63974 , n63979 );
or ( n63982 , n63977 , n63980 , n63981 );
and ( n63983 , n63971 , n63982 );
and ( n63984 , n63969 , n63982 );
or ( n63985 , n63972 , n63983 , n63984 );
buf ( n63986 , n20232 );
buf ( n63987 , n63986 );
and ( n63988 , n63987 , n58294 );
not ( n63989 , n63988 );
and ( n63990 , n61918 , n59611 );
not ( n63991 , n63990 );
and ( n63992 , n63989 , n63991 );
buf ( n63993 , n60821 );
not ( n63994 , n63993 );
and ( n63995 , n63991 , n63994 );
and ( n63996 , n63989 , n63994 );
or ( n63997 , n63992 , n63995 , n63996 );
xor ( n63998 , n63677 , n63681 );
xor ( n63999 , n63998 , n63684 );
and ( n64000 , n63997 , n63999 );
xor ( n64001 , n63643 , n63645 );
xor ( n64002 , n64001 , n63648 );
and ( n64003 , n63999 , n64002 );
and ( n64004 , n63997 , n64002 );
or ( n64005 , n64000 , n64003 , n64004 );
xor ( n64006 , n63485 , n63489 );
xor ( n64007 , n64006 , n63494 );
xor ( n64008 , n63499 , n63501 );
xor ( n64009 , n64008 , n63504 );
and ( n64010 , n64007 , n64009 );
xor ( n64011 , n63706 , n63710 );
and ( n64012 , n64009 , n64011 );
and ( n64013 , n64007 , n64011 );
or ( n64014 , n64010 , n64012 , n64013 );
and ( n64015 , n64005 , n64014 );
and ( n64016 , n46969 , n57187 );
and ( n64017 , n46843 , n57184 );
nor ( n64018 , n64016 , n64017 );
xnor ( n64019 , n64018 , n56175 );
and ( n64020 , n47216 , n56503 );
and ( n64021 , n47090 , n56501 );
nor ( n64022 , n64020 , n64021 );
xnor ( n64023 , n64022 , n56178 );
and ( n64024 , n64019 , n64023 );
and ( n64025 , n48384 , n53928 );
and ( n64026 , n48272 , n53926 );
nor ( n64027 , n64025 , n64026 );
xnor ( n64028 , n64027 , n53652 );
and ( n64029 , n64023 , n64028 );
and ( n64030 , n64019 , n64028 );
or ( n64031 , n64024 , n64029 , n64030 );
and ( n64032 , n51077 , n50338 );
and ( n64033 , n50726 , n50336 );
nor ( n64034 , n64032 , n64033 );
xnor ( n64035 , n64034 , n50111 );
and ( n64036 , n64031 , n64035 );
and ( n64037 , n51510 , n49896 );
and ( n64038 , n51298 , n49894 );
nor ( n64039 , n64037 , n64038 );
xnor ( n64040 , n64039 , n49711 );
and ( n64041 , n64035 , n64040 );
and ( n64042 , n64031 , n64040 );
or ( n64043 , n64036 , n64041 , n64042 );
and ( n64044 , n63492 , n58542 );
not ( n64045 , n64044 );
and ( n64046 , n63024 , n58911 );
not ( n64047 , n64046 );
and ( n64048 , n64045 , n64047 );
and ( n64049 , n61505 , n59920 );
not ( n64050 , n64049 );
and ( n64051 , n64048 , n64050 );
and ( n64052 , n61008 , n60372 );
not ( n64053 , n64052 );
and ( n64054 , n64050 , n64053 );
and ( n64055 , n64048 , n64053 );
or ( n64056 , n64051 , n64054 , n64055 );
and ( n64057 , n64043 , n64056 );
and ( n64058 , n58292 , n63766 );
not ( n64059 , n64058 );
and ( n64060 , n58628 , n63679 );
not ( n64061 , n64060 );
and ( n64062 , n64059 , n64061 );
and ( n64063 , n59908 , n61914 );
not ( n64064 , n64063 );
and ( n64065 , n64061 , n64064 );
and ( n64066 , n64059 , n64064 );
or ( n64067 , n64062 , n64065 , n64066 );
and ( n64068 , n58292 , n63679 );
not ( n64069 , n64068 );
and ( n64070 , n58628 , n62998 );
not ( n64071 , n64070 );
xor ( n64072 , n64069 , n64071 );
and ( n64073 , n60376 , n61015 );
not ( n64074 , n64073 );
xor ( n64075 , n64072 , n64074 );
or ( n64076 , n64067 , n64075 );
and ( n64077 , n64056 , n64076 );
and ( n64078 , n64043 , n64076 );
or ( n64079 , n64057 , n64077 , n64078 );
and ( n64080 , n64014 , n64079 );
and ( n64081 , n64005 , n64079 );
or ( n64082 , n64015 , n64080 , n64081 );
xor ( n64083 , n63694 , n63698 );
xor ( n64084 , n64083 , n63703 );
xor ( n64085 , n63735 , n63739 );
xor ( n64086 , n64085 , n63744 );
and ( n64087 , n64084 , n64086 );
xor ( n64088 , n63751 , n63755 );
xor ( n64089 , n64088 , n63760 );
and ( n64090 , n64086 , n64089 );
and ( n64091 , n64084 , n64089 );
or ( n64092 , n64087 , n64090 , n64091 );
and ( n64093 , n47778 , n55159 );
and ( n64094 , n47647 , n55157 );
nor ( n64095 , n64093 , n64094 );
xnor ( n64096 , n64095 , n54864 );
and ( n64097 , n48709 , n53357 );
and ( n64098 , n48632 , n53355 );
nor ( n64099 , n64097 , n64098 );
xnor ( n64100 , n64099 , n53060 );
and ( n64101 , n64096 , n64100 );
and ( n64102 , n50726 , n50783 );
and ( n64103 , n50625 , n50781 );
nor ( n64104 , n64102 , n64103 );
xnor ( n64105 , n64104 , n50557 );
and ( n64106 , n64100 , n64105 );
and ( n64107 , n64096 , n64105 );
or ( n64108 , n64101 , n64106 , n64107 );
and ( n64109 , n53922 , n48394 );
and ( n64110 , n53639 , n48392 );
nor ( n64111 , n64109 , n64110 );
xnor ( n64112 , n64111 , n48220 );
and ( n64113 , n54604 , n48042 );
and ( n64114 , n54227 , n48040 );
nor ( n64115 , n64113 , n64114 );
xnor ( n64116 , n64115 , n47921 );
and ( n64117 , n64112 , n64116 );
and ( n64118 , n57063 , n46911 );
and ( n64119 , n56915 , n46909 );
nor ( n64120 , n64118 , n64119 );
xnor ( n64121 , n64120 , n46802 );
and ( n64122 , n64116 , n64121 );
and ( n64123 , n64112 , n64121 );
or ( n64124 , n64117 , n64122 , n64123 );
and ( n64125 , n64108 , n64124 );
and ( n64126 , n47474 , n55851 );
and ( n64127 , n47351 , n55849 );
nor ( n64128 , n64126 , n64127 );
xnor ( n64129 , n64128 , n55506 );
and ( n64130 , n48108 , n54535 );
and ( n64131 , n47962 , n54533 );
nor ( n64132 , n64130 , n64131 );
xnor ( n64133 , n64132 , n54237 );
and ( n64134 , n64129 , n64133 );
and ( n64135 , n49115 , n52799 );
and ( n64136 , n48988 , n52797 );
nor ( n64137 , n64135 , n64136 );
xnor ( n64138 , n64137 , n52538 );
and ( n64139 , n64133 , n64138 );
and ( n64140 , n64129 , n64138 );
or ( n64141 , n64134 , n64139 , n64140 );
and ( n64142 , n64124 , n64141 );
and ( n64143 , n64108 , n64141 );
or ( n64144 , n64125 , n64142 , n64143 );
and ( n64145 , n64092 , n64144 );
and ( n64146 , n49570 , n52269 );
and ( n64147 , n49374 , n52267 );
nor ( n64148 , n64146 , n64147 );
xnor ( n64149 , n64148 , n52008 );
and ( n64150 , n49976 , n51750 );
and ( n64151 , n49781 , n51748 );
nor ( n64152 , n64150 , n64151 );
xnor ( n64153 , n64152 , n51520 );
and ( n64154 , n64149 , n64153 );
and ( n64155 , n50404 , n51221 );
and ( n64156 , n50195 , n51219 );
nor ( n64157 , n64155 , n64156 );
xnor ( n64158 , n64157 , n51000 );
and ( n64159 , n64153 , n64158 );
and ( n64160 , n64149 , n64158 );
or ( n64161 , n64154 , n64159 , n64160 );
and ( n64162 , n51298 , n50338 );
and ( n64163 , n51077 , n50336 );
nor ( n64164 , n64162 , n64163 );
xnor ( n64165 , n64164 , n50111 );
and ( n64166 , n51734 , n49896 );
and ( n64167 , n51510 , n49894 );
nor ( n64168 , n64166 , n64167 );
xnor ( n64169 , n64168 , n49711 );
and ( n64170 , n64165 , n64169 );
and ( n64171 , n52332 , n49513 );
and ( n64172 , n52082 , n49511 );
nor ( n64173 , n64171 , n64172 );
xnor ( n64174 , n64173 , n49310 );
and ( n64175 , n64169 , n64174 );
and ( n64176 , n64165 , n64174 );
or ( n64177 , n64170 , n64175 , n64176 );
and ( n64178 , n64161 , n64177 );
and ( n64179 , n52790 , n49121 );
and ( n64180 , n52612 , n49119 );
nor ( n64181 , n64179 , n64180 );
xnor ( n64182 , n64181 , n48932 );
and ( n64183 , n53328 , n48740 );
and ( n64184 , n53041 , n48738 );
nor ( n64185 , n64183 , n64184 );
xnor ( n64186 , n64185 , n48571 );
and ( n64187 , n64182 , n64186 );
and ( n64188 , n55143 , n47734 );
and ( n64189 , n54942 , n47732 );
nor ( n64190 , n64188 , n64189 );
xnor ( n64191 , n64190 , n47606 );
and ( n64192 , n64186 , n64191 );
and ( n64193 , n64182 , n64191 );
or ( n64194 , n64187 , n64192 , n64193 );
and ( n64195 , n64177 , n64194 );
and ( n64196 , n64161 , n64194 );
or ( n64197 , n64178 , n64195 , n64196 );
and ( n64198 , n64144 , n64197 );
and ( n64199 , n64092 , n64197 );
or ( n64200 , n64145 , n64198 , n64199 );
and ( n64201 , n55756 , n47429 );
and ( n64202 , n55497 , n47427 );
nor ( n64203 , n64201 , n64202 );
xnor ( n64204 , n64203 , n47309 );
and ( n64205 , n56388 , n47178 );
and ( n64206 , n56255 , n47176 );
nor ( n64207 , n64205 , n64206 );
xnor ( n64208 , n64207 , n47039 );
and ( n64209 , n64204 , n64208 );
and ( n64210 , n57063 , n46909 );
not ( n64211 , n64210 );
and ( n64212 , n64211 , n46802 );
and ( n64213 , n64208 , n64212 );
and ( n64214 , n64204 , n64212 );
or ( n64215 , n64209 , n64213 , n64214 );
xor ( n64216 , n40503 , n45556 );
buf ( n64217 , n64216 );
buf ( n64218 , n64217 );
buf ( n64219 , n64218 );
buf ( n64220 , n20235 );
buf ( n64221 , n64220 );
and ( n64222 , n64221 , n58294 );
not ( n64223 , n64222 );
and ( n64224 , n64219 , n64223 );
and ( n64225 , n62593 , n59207 );
not ( n64226 , n64225 );
and ( n64227 , n64223 , n64226 );
and ( n64228 , n64219 , n64226 );
or ( n64229 , n64224 , n64227 , n64228 );
and ( n64230 , n64215 , n64229 );
and ( n64231 , n62377 , n59611 );
not ( n64232 , n64231 );
and ( n64233 , n61008 , n60711 );
not ( n64234 , n64233 );
and ( n64235 , n64232 , n64234 );
buf ( n64236 , n64235 );
and ( n64237 , n64229 , n64236 );
and ( n64238 , n64215 , n64236 );
or ( n64239 , n64230 , n64237 , n64238 );
xor ( n64240 , n63783 , n63787 );
xor ( n64241 , n64240 , n63792 );
xor ( n64242 , n63799 , n63803 );
xor ( n64243 , n64242 , n63808 );
and ( n64244 , n64241 , n64243 );
xor ( n64245 , n63816 , n63820 );
xor ( n64246 , n64245 , n63825 );
and ( n64247 , n64243 , n64246 );
and ( n64248 , n64241 , n64246 );
or ( n64249 , n64244 , n64247 , n64248 );
and ( n64250 , n64239 , n64249 );
buf ( n64251 , n63713 );
xor ( n64252 , n64251 , n63715 );
and ( n64253 , n64249 , n64252 );
and ( n64254 , n64239 , n64252 );
or ( n64255 , n64250 , n64253 , n64254 );
and ( n64256 , n64200 , n64255 );
xor ( n64257 , n63720 , n63722 );
xor ( n64258 , n64257 , n63724 );
xor ( n64259 , n63747 , n63763 );
xor ( n64260 , n64259 , n63776 );
and ( n64261 , n64258 , n64260 );
xor ( n64262 , n63795 , n63811 );
xor ( n64263 , n64262 , n63828 );
and ( n64264 , n64260 , n64263 );
and ( n64265 , n64258 , n64263 );
or ( n64266 , n64261 , n64264 , n64265 );
and ( n64267 , n64255 , n64266 );
and ( n64268 , n64200 , n64266 );
or ( n64269 , n64256 , n64267 , n64268 );
and ( n64270 , n64082 , n64269 );
xor ( n64271 , n63664 , n63666 );
xor ( n64272 , n64271 , n63687 );
xor ( n64273 , n63711 , n63717 );
xor ( n64274 , n64273 , n63727 );
and ( n64275 , n64272 , n64274 );
xor ( n64276 , n63779 , n63831 );
xor ( n64277 , n64276 , n63860 );
and ( n64278 , n64274 , n64277 );
and ( n64279 , n64272 , n64277 );
or ( n64280 , n64275 , n64278 , n64279 );
and ( n64281 , n64269 , n64280 );
and ( n64282 , n64082 , n64280 );
or ( n64283 , n64270 , n64281 , n64282 );
and ( n64284 , n63985 , n64283 );
xor ( n64285 , n63639 , n63641 );
xor ( n64286 , n64285 , n63659 );
xor ( n64287 , n63690 , n63730 );
xor ( n64288 , n64287 , n63863 );
and ( n64289 , n64286 , n64288 );
xor ( n64290 , n63885 , n63895 );
xor ( n64291 , n64290 , n63898 );
and ( n64292 , n64288 , n64291 );
and ( n64293 , n64286 , n64291 );
or ( n64294 , n64289 , n64292 , n64293 );
and ( n64295 , n64283 , n64294 );
and ( n64296 , n63985 , n64294 );
or ( n64297 , n64284 , n64295 , n64296 );
and ( n64298 , n63967 , n64297 );
xor ( n64299 , n63662 , n63866 );
xor ( n64300 , n64299 , n63901 );
xor ( n64301 , n63914 , n63916 );
xor ( n64302 , n64301 , n63919 );
and ( n64303 , n64300 , n64302 );
xor ( n64304 , n63925 , n63927 );
xor ( n64305 , n64304 , n63930 );
and ( n64306 , n64302 , n64305 );
and ( n64307 , n64300 , n64305 );
or ( n64308 , n64303 , n64306 , n64307 );
and ( n64309 , n64297 , n64308 );
and ( n64310 , n63967 , n64308 );
or ( n64311 , n64298 , n64309 , n64310 );
and ( n64312 , n63964 , n64311 );
and ( n64313 , n63962 , n64311 );
or ( n64314 , n63965 , n64312 , n64313 );
and ( n64315 , n63960 , n64314 );
xor ( n64316 , n63634 , n63636 );
xor ( n64317 , n64316 , n63952 );
and ( n64318 , n64314 , n64317 );
and ( n64319 , n63960 , n64317 );
or ( n64320 , n64315 , n64318 , n64319 );
and ( n64321 , n63957 , n64320 );
and ( n64322 , n63955 , n64320 );
or ( n64323 , n63958 , n64321 , n64322 );
and ( n64324 , n63631 , n64323 );
and ( n64325 , n63629 , n64323 );
or ( n64326 , n63632 , n64324 , n64325 );
and ( n64327 , n63627 , n64326 );
xor ( n64328 , n63629 , n63631 );
xor ( n64329 , n64328 , n64323 );
xor ( n64330 , n63955 , n63957 );
xor ( n64331 , n64330 , n64320 );
xor ( n64332 , n63936 , n63946 );
xor ( n64333 , n64332 , n63949 );
xor ( n64334 , n63904 , n63922 );
xor ( n64335 , n64334 , n63933 );
xor ( n64336 , n63938 , n63940 );
xor ( n64337 , n64336 , n63943 );
and ( n64338 , n64335 , n64337 );
xor ( n64339 , n63906 , n63908 );
xor ( n64340 , n64339 , n63911 );
and ( n64341 , n64069 , n64071 );
and ( n64342 , n64071 , n64074 );
and ( n64343 , n64069 , n64074 );
or ( n64344 , n64341 , n64342 , n64343 );
and ( n64345 , n62593 , n58911 );
not ( n64346 , n64345 );
buf ( n64347 , n64346 );
and ( n64348 , n64344 , n64347 );
xor ( n64349 , n63242 , n63244 );
xor ( n64350 , n64349 , n63247 );
and ( n64351 , n64347 , n64350 );
and ( n64352 , n64344 , n64350 );
or ( n64353 , n64348 , n64351 , n64352 );
xor ( n64354 , n62988 , n62990 );
xor ( n64355 , n64354 , n62993 );
and ( n64356 , n64353 , n64355 );
xor ( n64357 , n63250 , n63252 );
xor ( n64358 , n64357 , n63255 );
and ( n64359 , n64355 , n64358 );
and ( n64360 , n64353 , n64358 );
or ( n64361 , n64356 , n64359 , n64360 );
and ( n64362 , n64340 , n64361 );
xor ( n64363 , n63877 , n63879 );
xor ( n64364 , n64363 , n63882 );
xor ( n64365 , n63887 , n63889 );
xor ( n64366 , n64365 , n63892 );
and ( n64367 , n64364 , n64366 );
xor ( n64368 , n63848 , n63854 );
xor ( n64369 , n64368 , n63857 );
xor ( n64370 , n63869 , n63871 );
xor ( n64371 , n64370 , n63874 );
and ( n64372 , n64369 , n64371 );
xor ( n64373 , n63997 , n63999 );
xor ( n64374 , n64373 , n64002 );
and ( n64375 , n64371 , n64374 );
and ( n64376 , n64369 , n64374 );
or ( n64377 , n64372 , n64375 , n64376 );
and ( n64378 , n64366 , n64377 );
and ( n64379 , n64364 , n64377 );
or ( n64380 , n64367 , n64378 , n64379 );
and ( n64381 , n64361 , n64380 );
and ( n64382 , n64340 , n64380 );
or ( n64383 , n64362 , n64381 , n64382 );
and ( n64384 , n58915 , n62998 );
not ( n64385 , n64384 );
buf ( n64386 , n64385 );
and ( n64387 , n64386 , n64345 );
and ( n64388 , n59365 , n62151 );
not ( n64389 , n64388 );
and ( n64390 , n64345 , n64389 );
and ( n64391 , n64386 , n64389 );
or ( n64392 , n64387 , n64390 , n64391 );
xor ( n64393 , n64045 , n64047 );
and ( n64394 , n63987 , n58444 );
not ( n64395 , n64394 );
and ( n64396 , n64393 , n64395 );
and ( n64397 , n61505 , n60372 );
not ( n64398 , n64397 );
and ( n64399 , n64395 , n64398 );
and ( n64400 , n64393 , n64398 );
or ( n64401 , n64396 , n64399 , n64400 );
and ( n64402 , n62377 , n59207 );
not ( n64403 , n64402 );
and ( n64404 , n64401 , n64403 );
xor ( n64405 , n63669 , n63671 );
xor ( n64406 , n64405 , n63674 );
and ( n64407 , n64403 , n64406 );
and ( n64408 , n64401 , n64406 );
or ( n64409 , n64404 , n64407 , n64408 );
and ( n64410 , n64392 , n64409 );
buf ( n64411 , n20235 );
buf ( n64412 , n64411 );
and ( n64413 , n57948 , n64412 );
not ( n64414 , n64413 );
and ( n64415 , n59615 , n62151 );
not ( n64416 , n64415 );
and ( n64417 , n64414 , n64416 );
and ( n64418 , n61918 , n59920 );
not ( n64419 , n64418 );
and ( n64420 , n64416 , n64419 );
and ( n64421 , n64414 , n64419 );
or ( n64422 , n64417 , n64420 , n64421 );
xor ( n64423 , n63989 , n63991 );
xor ( n64424 , n64423 , n63994 );
and ( n64425 , n64422 , n64424 );
xor ( n64426 , n64048 , n64050 );
xor ( n64427 , n64426 , n64053 );
and ( n64428 , n64424 , n64427 );
and ( n64429 , n64422 , n64427 );
or ( n64430 , n64425 , n64428 , n64429 );
and ( n64431 , n64409 , n64430 );
and ( n64432 , n64392 , n64430 );
or ( n64433 , n64410 , n64431 , n64432 );
xor ( n64434 , n63836 , n63840 );
xor ( n64435 , n64434 , n63845 );
xor ( n64436 , n63483 , n63852 );
buf ( n64437 , n64436 );
and ( n64438 , n64435 , n64437 );
xor ( n64439 , n64031 , n64035 );
xor ( n64440 , n64439 , n64040 );
and ( n64441 , n64437 , n64440 );
and ( n64442 , n64435 , n64440 );
or ( n64443 , n64438 , n64441 , n64442 );
xnor ( n64444 , n64067 , n64075 );
and ( n64445 , n58292 , n64412 );
not ( n64446 , n64445 );
and ( n64447 , n58628 , n63766 );
not ( n64448 , n64447 );
and ( n64449 , n64446 , n64448 );
and ( n64450 , n60376 , n61914 );
not ( n64451 , n64450 );
and ( n64452 , n64448 , n64451 );
and ( n64453 , n64446 , n64451 );
or ( n64454 , n64449 , n64452 , n64453 );
and ( n64455 , n64454 , n64384 );
and ( n64456 , n59365 , n62868 );
not ( n64457 , n64456 );
and ( n64458 , n64384 , n64457 );
and ( n64459 , n64454 , n64457 );
or ( n64460 , n64455 , n64458 , n64459 );
and ( n64461 , n64444 , n64460 );
xor ( n64462 , n64096 , n64100 );
xor ( n64463 , n64462 , n64105 );
xor ( n64464 , n64019 , n64023 );
xor ( n64465 , n64464 , n64028 );
and ( n64466 , n64463 , n64465 );
xor ( n64467 , n64112 , n64116 );
xor ( n64468 , n64467 , n64121 );
and ( n64469 , n64465 , n64468 );
and ( n64470 , n64463 , n64468 );
or ( n64471 , n64466 , n64469 , n64470 );
and ( n64472 , n64460 , n64471 );
and ( n64473 , n64444 , n64471 );
or ( n64474 , n64461 , n64472 , n64473 );
and ( n64475 , n64443 , n64474 );
xor ( n64476 , n64059 , n64061 );
xor ( n64477 , n64476 , n64064 );
xor ( n64478 , n64414 , n64416 );
xor ( n64479 , n64478 , n64419 );
and ( n64480 , n64477 , n64479 );
and ( n64481 , n47647 , n55851 );
and ( n64482 , n47474 , n55849 );
nor ( n64483 , n64481 , n64482 );
xnor ( n64484 , n64483 , n55506 );
and ( n64485 , n48272 , n54535 );
and ( n64486 , n48108 , n54533 );
nor ( n64487 , n64485 , n64486 );
xnor ( n64488 , n64487 , n54237 );
and ( n64489 , n64484 , n64488 );
and ( n64490 , n48632 , n53928 );
and ( n64491 , n48384 , n53926 );
nor ( n64492 , n64490 , n64491 );
xnor ( n64493 , n64492 , n53652 );
and ( n64494 , n64488 , n64493 );
and ( n64495 , n64484 , n64493 );
or ( n64496 , n64489 , n64494 , n64495 );
and ( n64497 , n64479 , n64496 );
and ( n64498 , n64477 , n64496 );
or ( n64499 , n64480 , n64497 , n64498 );
and ( n64500 , n47351 , n56503 );
and ( n64501 , n47216 , n56501 );
nor ( n64502 , n64500 , n64501 );
xnor ( n64503 , n64502 , n56178 );
and ( n64504 , n47962 , n55159 );
and ( n64505 , n47778 , n55157 );
nor ( n64506 , n64504 , n64505 );
xnor ( n64507 , n64506 , n54864 );
and ( n64508 , n64503 , n64507 );
and ( n64509 , n51077 , n50783 );
and ( n64510 , n50726 , n50781 );
nor ( n64511 , n64509 , n64510 );
xnor ( n64512 , n64511 , n50557 );
and ( n64513 , n64507 , n64512 );
and ( n64514 , n64503 , n64512 );
or ( n64515 , n64508 , n64513 , n64514 );
and ( n64516 , n54227 , n48394 );
and ( n64517 , n53922 , n48392 );
nor ( n64518 , n64516 , n64517 );
xnor ( n64519 , n64518 , n48220 );
and ( n64520 , n54942 , n48042 );
and ( n64521 , n54604 , n48040 );
nor ( n64522 , n64520 , n64521 );
xnor ( n64523 , n64522 , n47921 );
and ( n64524 , n64519 , n64523 );
and ( n64525 , n56915 , n47178 );
and ( n64526 , n56388 , n47176 );
nor ( n64527 , n64525 , n64526 );
xnor ( n64528 , n64527 , n47039 );
and ( n64529 , n64523 , n64528 );
and ( n64530 , n64519 , n64528 );
or ( n64531 , n64524 , n64529 , n64530 );
and ( n64532 , n64515 , n64531 );
and ( n64533 , n63987 , n58542 );
not ( n64534 , n64533 );
and ( n64535 , n58915 , n63679 );
not ( n64536 , n64535 );
and ( n64537 , n64534 , n64536 );
and ( n64538 , n61918 , n60372 );
not ( n64539 , n64538 );
and ( n64540 , n64536 , n64539 );
and ( n64541 , n64534 , n64539 );
or ( n64542 , n64537 , n64540 , n64541 );
and ( n64543 , n64531 , n64542 );
and ( n64544 , n64515 , n64542 );
or ( n64545 , n64532 , n64543 , n64544 );
and ( n64546 , n64499 , n64545 );
buf ( n64547 , n20238 );
buf ( n64548 , n64547 );
and ( n64549 , n64548 , n58294 );
not ( n64550 , n64549 );
and ( n64551 , n63492 , n58911 );
and ( n64552 , n64550 , n64551 );
and ( n64553 , n62593 , n59611 );
not ( n64554 , n64553 );
and ( n64555 , n64551 , n64554 );
and ( n64556 , n64550 , n64554 );
or ( n64557 , n64552 , n64555 , n64556 );
and ( n64558 , n47090 , n57187 );
and ( n64559 , n46969 , n57184 );
nor ( n64560 , n64558 , n64559 );
xnor ( n64561 , n64560 , n56175 );
and ( n64562 , n48988 , n53357 );
and ( n64563 , n48709 , n53355 );
nor ( n64564 , n64562 , n64563 );
xnor ( n64565 , n64564 , n53060 );
and ( n64566 , n64561 , n64565 );
and ( n64567 , n49374 , n52799 );
and ( n64568 , n49115 , n52797 );
nor ( n64569 , n64567 , n64568 );
xnor ( n64570 , n64569 , n52538 );
and ( n64571 , n64565 , n64570 );
and ( n64572 , n64561 , n64570 );
or ( n64573 , n64566 , n64571 , n64572 );
and ( n64574 , n64557 , n64573 );
and ( n64575 , n49781 , n52269 );
and ( n64576 , n49570 , n52267 );
nor ( n64577 , n64575 , n64576 );
xnor ( n64578 , n64577 , n52008 );
and ( n64579 , n50195 , n51750 );
and ( n64580 , n49976 , n51748 );
nor ( n64581 , n64579 , n64580 );
xnor ( n64582 , n64581 , n51520 );
and ( n64583 , n64578 , n64582 );
and ( n64584 , n50625 , n51221 );
and ( n64585 , n50404 , n51219 );
nor ( n64586 , n64584 , n64585 );
xnor ( n64587 , n64586 , n51000 );
and ( n64588 , n64582 , n64587 );
and ( n64589 , n64578 , n64587 );
or ( n64590 , n64583 , n64588 , n64589 );
and ( n64591 , n64573 , n64590 );
and ( n64592 , n64557 , n64590 );
or ( n64593 , n64574 , n64591 , n64592 );
and ( n64594 , n64545 , n64593 );
and ( n64595 , n64499 , n64593 );
or ( n64596 , n64546 , n64594 , n64595 );
and ( n64597 , n64474 , n64596 );
and ( n64598 , n64443 , n64596 );
or ( n64599 , n64475 , n64597 , n64598 );
and ( n64600 , n64433 , n64599 );
and ( n64601 , n51510 , n50338 );
and ( n64602 , n51298 , n50336 );
nor ( n64603 , n64601 , n64602 );
xnor ( n64604 , n64603 , n50111 );
and ( n64605 , n52082 , n49896 );
and ( n64606 , n51734 , n49894 );
nor ( n64607 , n64605 , n64606 );
xnor ( n64608 , n64607 , n49711 );
and ( n64609 , n64604 , n64608 );
and ( n64610 , n52612 , n49513 );
and ( n64611 , n52332 , n49511 );
nor ( n64612 , n64610 , n64611 );
xnor ( n64613 , n64612 , n49310 );
and ( n64614 , n64608 , n64613 );
and ( n64615 , n64604 , n64613 );
or ( n64616 , n64609 , n64614 , n64615 );
and ( n64617 , n53041 , n49121 );
and ( n64618 , n52790 , n49119 );
nor ( n64619 , n64617 , n64618 );
xnor ( n64620 , n64619 , n48932 );
and ( n64621 , n53639 , n48740 );
and ( n64622 , n53328 , n48738 );
nor ( n64623 , n64621 , n64622 );
xnor ( n64624 , n64623 , n48571 );
and ( n64625 , n64620 , n64624 );
and ( n64626 , n55497 , n47734 );
and ( n64627 , n55143 , n47732 );
nor ( n64628 , n64626 , n64627 );
xnor ( n64629 , n64628 , n47606 );
and ( n64630 , n64624 , n64629 );
and ( n64631 , n64620 , n64629 );
or ( n64632 , n64625 , n64630 , n64631 );
and ( n64633 , n64616 , n64632 );
and ( n64634 , n56255 , n47429 );
and ( n64635 , n55756 , n47427 );
nor ( n64636 , n64634 , n64635 );
xnor ( n64637 , n64636 , n47309 );
and ( n64638 , n64637 , n64210 );
xor ( n64639 , n41787 , n45554 );
buf ( n64640 , n64639 );
buf ( n64641 , n64640 );
buf ( n64642 , n64641 );
and ( n64643 , n64210 , n64642 );
and ( n64644 , n64637 , n64642 );
or ( n64645 , n64638 , n64643 , n64644 );
and ( n64646 , n64632 , n64645 );
and ( n64647 , n64616 , n64645 );
or ( n64648 , n64633 , n64646 , n64647 );
xor ( n64649 , n64129 , n64133 );
xor ( n64650 , n64649 , n64138 );
xor ( n64651 , n64149 , n64153 );
xor ( n64652 , n64651 , n64158 );
and ( n64653 , n64650 , n64652 );
xor ( n64654 , n64165 , n64169 );
xor ( n64655 , n64654 , n64174 );
and ( n64656 , n64652 , n64655 );
and ( n64657 , n64650 , n64655 );
or ( n64658 , n64653 , n64656 , n64657 );
and ( n64659 , n64648 , n64658 );
xor ( n64660 , n64182 , n64186 );
xor ( n64661 , n64660 , n64191 );
xor ( n64662 , n64204 , n64208 );
xor ( n64663 , n64662 , n64212 );
and ( n64664 , n64661 , n64663 );
xor ( n64665 , n64219 , n64223 );
xor ( n64666 , n64665 , n64226 );
and ( n64667 , n64663 , n64666 );
and ( n64668 , n64661 , n64666 );
or ( n64669 , n64664 , n64667 , n64668 );
and ( n64670 , n64658 , n64669 );
and ( n64671 , n64648 , n64669 );
or ( n64672 , n64659 , n64670 , n64671 );
xor ( n64673 , n64084 , n64086 );
xor ( n64674 , n64673 , n64089 );
xor ( n64675 , n64108 , n64124 );
xor ( n64676 , n64675 , n64141 );
and ( n64677 , n64674 , n64676 );
xor ( n64678 , n64161 , n64177 );
xor ( n64679 , n64678 , n64194 );
and ( n64680 , n64676 , n64679 );
and ( n64681 , n64674 , n64679 );
or ( n64682 , n64677 , n64680 , n64681 );
and ( n64683 , n64672 , n64682 );
xor ( n64684 , n64007 , n64009 );
xor ( n64685 , n64684 , n64011 );
and ( n64686 , n64682 , n64685 );
and ( n64687 , n64672 , n64685 );
or ( n64688 , n64683 , n64686 , n64687 );
and ( n64689 , n64599 , n64688 );
and ( n64690 , n64433 , n64688 );
or ( n64691 , n64600 , n64689 , n64690 );
xor ( n64692 , n64043 , n64056 );
xor ( n64693 , n64692 , n64076 );
xor ( n64694 , n64092 , n64144 );
xor ( n64695 , n64694 , n64197 );
and ( n64696 , n64693 , n64695 );
xor ( n64697 , n64239 , n64249 );
xor ( n64698 , n64697 , n64252 );
and ( n64699 , n64695 , n64698 );
and ( n64700 , n64693 , n64698 );
or ( n64701 , n64696 , n64699 , n64700 );
xor ( n64702 , n63974 , n63976 );
xor ( n64703 , n64702 , n63979 );
and ( n64704 , n64701 , n64703 );
xor ( n64705 , n64005 , n64014 );
xor ( n64706 , n64705 , n64079 );
and ( n64707 , n64703 , n64706 );
and ( n64708 , n64701 , n64706 );
or ( n64709 , n64704 , n64707 , n64708 );
and ( n64710 , n64691 , n64709 );
xor ( n64711 , n63969 , n63971 );
xor ( n64712 , n64711 , n63982 );
and ( n64713 , n64709 , n64712 );
and ( n64714 , n64691 , n64712 );
or ( n64715 , n64710 , n64713 , n64714 );
and ( n64716 , n64383 , n64715 );
xor ( n64717 , n63985 , n64283 );
xor ( n64718 , n64717 , n64294 );
and ( n64719 , n64715 , n64718 );
and ( n64720 , n64383 , n64718 );
or ( n64721 , n64716 , n64719 , n64720 );
and ( n64722 , n64337 , n64721 );
and ( n64723 , n64335 , n64721 );
or ( n64724 , n64338 , n64722 , n64723 );
and ( n64725 , n64333 , n64724 );
xor ( n64726 , n63962 , n63964 );
xor ( n64727 , n64726 , n64311 );
and ( n64728 , n64724 , n64727 );
and ( n64729 , n64333 , n64727 );
or ( n64730 , n64725 , n64728 , n64729 );
xor ( n64731 , n63960 , n64314 );
xor ( n64732 , n64731 , n64317 );
and ( n64733 , n64730 , n64732 );
xor ( n64734 , n63967 , n64297 );
xor ( n64735 , n64734 , n64308 );
xor ( n64736 , n64300 , n64302 );
xor ( n64737 , n64736 , n64305 );
xor ( n64738 , n64082 , n64269 );
xor ( n64739 , n64738 , n64280 );
xor ( n64740 , n64286 , n64288 );
xor ( n64741 , n64740 , n64291 );
and ( n64742 , n64739 , n64741 );
xor ( n64743 , n64200 , n64255 );
xor ( n64744 , n64743 , n64266 );
xor ( n64745 , n64272 , n64274 );
xor ( n64746 , n64745 , n64277 );
and ( n64747 , n64744 , n64746 );
xor ( n64748 , n64353 , n64355 );
xor ( n64749 , n64748 , n64358 );
and ( n64750 , n64746 , n64749 );
and ( n64751 , n64744 , n64749 );
or ( n64752 , n64747 , n64750 , n64751 );
and ( n64753 , n64741 , n64752 );
and ( n64754 , n64739 , n64752 );
or ( n64755 , n64742 , n64753 , n64754 );
and ( n64756 , n64737 , n64755 );
xor ( n64757 , n64258 , n64260 );
xor ( n64758 , n64757 , n64263 );
xor ( n64759 , n64344 , n64347 );
xor ( n64760 , n64759 , n64350 );
and ( n64761 , n64758 , n64760 );
not ( n64762 , n64551 );
buf ( n64763 , n64762 );
and ( n64764 , n60376 , n61481 );
not ( n64765 , n64764 );
and ( n64766 , n64763 , n64765 );
and ( n64767 , n60821 , n61015 );
not ( n64768 , n64767 );
and ( n64769 , n64765 , n64768 );
and ( n64770 , n64763 , n64768 );
or ( n64771 , n64766 , n64769 , n64770 );
xor ( n64772 , n63768 , n63770 );
xor ( n64773 , n64772 , n63773 );
and ( n64774 , n64771 , n64773 );
xor ( n64775 , n64386 , n64345 );
xor ( n64776 , n64775 , n64389 );
and ( n64777 , n64773 , n64776 );
and ( n64778 , n64771 , n64776 );
or ( n64779 , n64774 , n64777 , n64778 );
and ( n64780 , n64760 , n64779 );
and ( n64781 , n64758 , n64779 );
or ( n64782 , n64761 , n64780 , n64781 );
xor ( n64783 , n64215 , n64229 );
xor ( n64784 , n64783 , n64236 );
xor ( n64785 , n64241 , n64243 );
xor ( n64786 , n64785 , n64246 );
and ( n64787 , n64784 , n64786 );
xor ( n64788 , n64401 , n64403 );
xor ( n64789 , n64788 , n64406 );
and ( n64790 , n64786 , n64789 );
and ( n64791 , n64784 , n64789 );
or ( n64792 , n64787 , n64790 , n64791 );
xor ( n64793 , n64422 , n64424 );
xor ( n64794 , n64793 , n64427 );
and ( n64795 , n64221 , n58444 );
not ( n64796 , n64795 );
and ( n64797 , n59615 , n62868 );
not ( n64798 , n64797 );
and ( n64799 , n64796 , n64798 );
buf ( n64800 , n61008 );
not ( n64801 , n64800 );
and ( n64802 , n64798 , n64801 );
and ( n64803 , n64796 , n64801 );
or ( n64804 , n64799 , n64802 , n64803 );
and ( n64805 , n58628 , n64412 );
not ( n64806 , n64805 );
and ( n64807 , n63987 , n58911 );
not ( n64808 , n64807 );
and ( n64809 , n64806 , n64808 );
buf ( n64810 , n20238 );
buf ( n64811 , n64810 );
and ( n64812 , n57948 , n64811 );
not ( n64813 , n64812 );
and ( n64814 , n64809 , n64813 );
and ( n64815 , n62377 , n59920 );
not ( n64816 , n64815 );
and ( n64817 , n64813 , n64816 );
and ( n64818 , n64809 , n64816 );
or ( n64819 , n64814 , n64817 , n64818 );
and ( n64820 , n64804 , n64819 );
xor ( n64821 , n64393 , n64395 );
xor ( n64822 , n64821 , n64398 );
and ( n64823 , n64819 , n64822 );
and ( n64824 , n64804 , n64822 );
or ( n64825 , n64820 , n64823 , n64824 );
and ( n64826 , n64794 , n64825 );
xor ( n64827 , n64232 , n64234 );
buf ( n64828 , n64827 );
and ( n64829 , n63024 , n59207 );
not ( n64830 , n64829 );
and ( n64831 , n61505 , n60711 );
not ( n64832 , n64831 );
and ( n64833 , n64830 , n64832 );
xor ( n64834 , n64534 , n64536 );
xor ( n64835 , n64834 , n64539 );
and ( n64836 , n64832 , n64835 );
and ( n64837 , n64830 , n64835 );
or ( n64838 , n64833 , n64836 , n64837 );
and ( n64839 , n64828 , n64838 );
and ( n64840 , n58915 , n63766 );
and ( n64841 , n59365 , n63679 );
not ( n64842 , n64841 );
and ( n64843 , n64840 , n64842 );
and ( n64844 , n61918 , n60711 );
not ( n64845 , n64844 );
and ( n64846 , n64842 , n64845 );
and ( n64847 , n64840 , n64845 );
or ( n64848 , n64843 , n64846 , n64847 );
and ( n64849 , n59365 , n62998 );
not ( n64850 , n64849 );
and ( n64851 , n59908 , n62151 );
not ( n64852 , n64851 );
xor ( n64853 , n64850 , n64852 );
and ( n64854 , n60821 , n61481 );
not ( n64855 , n64854 );
xor ( n64856 , n64853 , n64855 );
or ( n64857 , n64848 , n64856 );
and ( n64858 , n64838 , n64857 );
and ( n64859 , n64828 , n64857 );
or ( n64860 , n64839 , n64858 , n64859 );
and ( n64861 , n64825 , n64860 );
and ( n64862 , n64794 , n64860 );
or ( n64863 , n64826 , n64861 , n64862 );
and ( n64864 , n64792 , n64863 );
xor ( n64865 , n64484 , n64488 );
xor ( n64866 , n64865 , n64493 );
xor ( n64867 , n64503 , n64507 );
xor ( n64868 , n64867 , n64512 );
and ( n64869 , n64866 , n64868 );
xor ( n64870 , n64519 , n64523 );
xor ( n64871 , n64870 , n64528 );
xor ( n64872 , n64446 , n64448 );
xor ( n64873 , n64872 , n64451 );
and ( n64874 , n64871 , n64873 );
buf ( n64875 , n64874 );
and ( n64876 , n64869 , n64875 );
and ( n64877 , n48108 , n55159 );
and ( n64878 , n47962 , n55157 );
nor ( n64879 , n64877 , n64878 );
xnor ( n64880 , n64879 , n54864 );
and ( n64881 , n48384 , n54535 );
and ( n64882 , n48272 , n54533 );
nor ( n64883 , n64881 , n64882 );
xnor ( n64884 , n64883 , n54237 );
and ( n64885 , n64880 , n64884 );
and ( n64886 , n51298 , n50783 );
and ( n64887 , n51077 , n50781 );
nor ( n64888 , n64886 , n64887 );
xnor ( n64889 , n64888 , n50557 );
and ( n64890 , n64884 , n64889 );
and ( n64891 , n64880 , n64889 );
or ( n64892 , n64885 , n64890 , n64891 );
not ( n64893 , n64840 );
buf ( n64894 , n64893 );
and ( n64895 , n64892 , n64894 );
and ( n64896 , n64548 , n58444 );
not ( n64897 , n64896 );
and ( n64898 , n64221 , n58542 );
not ( n64899 , n64898 );
or ( n64900 , n64897 , n64899 );
and ( n64901 , n64894 , n64900 );
and ( n64902 , n64892 , n64900 );
or ( n64903 , n64895 , n64901 , n64902 );
and ( n64904 , n64875 , n64903 );
and ( n64905 , n64869 , n64903 );
or ( n64906 , n64876 , n64904 , n64905 );
and ( n64907 , n47216 , n57187 );
and ( n64908 , n47090 , n57184 );
nor ( n64909 , n64907 , n64908 );
xnor ( n64910 , n64909 , n56175 );
and ( n64911 , n47474 , n56503 );
and ( n64912 , n47351 , n56501 );
nor ( n64913 , n64911 , n64912 );
xnor ( n64914 , n64913 , n56178 );
and ( n64915 , n64910 , n64914 );
and ( n64916 , n47778 , n55851 );
and ( n64917 , n47647 , n55849 );
nor ( n64918 , n64916 , n64917 );
xnor ( n64919 , n64918 , n55506 );
and ( n64920 , n64914 , n64919 );
and ( n64921 , n64910 , n64919 );
or ( n64922 , n64915 , n64920 , n64921 );
and ( n64923 , n48709 , n53928 );
and ( n64924 , n48632 , n53926 );
nor ( n64925 , n64923 , n64924 );
xnor ( n64926 , n64925 , n53652 );
and ( n64927 , n49115 , n53357 );
and ( n64928 , n48988 , n53355 );
nor ( n64929 , n64927 , n64928 );
xnor ( n64930 , n64929 , n53060 );
and ( n64931 , n64926 , n64930 );
and ( n64932 , n49570 , n52799 );
and ( n64933 , n49374 , n52797 );
nor ( n64934 , n64932 , n64933 );
xnor ( n64935 , n64934 , n52538 );
and ( n64936 , n64930 , n64935 );
and ( n64937 , n64926 , n64935 );
or ( n64938 , n64931 , n64936 , n64937 );
and ( n64939 , n64922 , n64938 );
and ( n64940 , n49976 , n52269 );
and ( n64941 , n49781 , n52267 );
nor ( n64942 , n64940 , n64941 );
xnor ( n64943 , n64942 , n52008 );
and ( n64944 , n50404 , n51750 );
and ( n64945 , n50195 , n51748 );
nor ( n64946 , n64944 , n64945 );
xnor ( n64947 , n64946 , n51520 );
and ( n64948 , n64943 , n64947 );
and ( n64949 , n50726 , n51221 );
and ( n64950 , n50625 , n51219 );
nor ( n64951 , n64949 , n64950 );
xnor ( n64952 , n64951 , n51000 );
and ( n64953 , n64947 , n64952 );
and ( n64954 , n64943 , n64952 );
or ( n64955 , n64948 , n64953 , n64954 );
and ( n64956 , n64938 , n64955 );
and ( n64957 , n64922 , n64955 );
or ( n64958 , n64939 , n64956 , n64957 );
and ( n64959 , n51734 , n50338 );
and ( n64960 , n51510 , n50336 );
nor ( n64961 , n64959 , n64960 );
xnor ( n64962 , n64961 , n50111 );
and ( n64963 , n52332 , n49896 );
and ( n64964 , n52082 , n49894 );
nor ( n64965 , n64963 , n64964 );
xnor ( n64966 , n64965 , n49711 );
and ( n64967 , n64962 , n64966 );
and ( n64968 , n52790 , n49513 );
and ( n64969 , n52612 , n49511 );
nor ( n64970 , n64968 , n64969 );
xnor ( n64971 , n64970 , n49310 );
and ( n64972 , n64966 , n64971 );
and ( n64973 , n64962 , n64971 );
or ( n64974 , n64967 , n64972 , n64973 );
and ( n64975 , n53328 , n49121 );
and ( n64976 , n53041 , n49119 );
nor ( n64977 , n64975 , n64976 );
xnor ( n64978 , n64977 , n48932 );
and ( n64979 , n53922 , n48740 );
and ( n64980 , n53639 , n48738 );
nor ( n64981 , n64979 , n64980 );
xnor ( n64982 , n64981 , n48571 );
and ( n64983 , n64978 , n64982 );
and ( n64984 , n54604 , n48394 );
and ( n64985 , n54227 , n48392 );
nor ( n64986 , n64984 , n64985 );
xnor ( n64987 , n64986 , n48220 );
and ( n64988 , n64982 , n64987 );
and ( n64989 , n64978 , n64987 );
or ( n64990 , n64983 , n64988 , n64989 );
and ( n64991 , n64974 , n64990 );
and ( n64992 , n55143 , n48042 );
and ( n64993 , n54942 , n48040 );
nor ( n64994 , n64992 , n64993 );
xnor ( n64995 , n64994 , n47921 );
and ( n64996 , n55756 , n47734 );
and ( n64997 , n55497 , n47732 );
nor ( n64998 , n64996 , n64997 );
xnor ( n64999 , n64998 , n47606 );
and ( n65000 , n64995 , n64999 );
and ( n65001 , n56388 , n47429 );
and ( n65002 , n56255 , n47427 );
nor ( n65003 , n65001 , n65002 );
xnor ( n65004 , n65003 , n47309 );
and ( n65005 , n64999 , n65004 );
and ( n65006 , n64995 , n65004 );
or ( n65007 , n65000 , n65005 , n65006 );
and ( n65008 , n64990 , n65007 );
and ( n65009 , n64974 , n65007 );
or ( n65010 , n64991 , n65008 , n65009 );
and ( n65011 , n64958 , n65010 );
and ( n65012 , n57063 , n47178 );
and ( n65013 , n56915 , n47176 );
nor ( n65014 , n65012 , n65013 );
xnor ( n65015 , n65014 , n47039 );
and ( n65016 , n57063 , n47176 );
not ( n65017 , n65016 );
and ( n65018 , n65017 , n47039 );
and ( n65019 , n65015 , n65018 );
xor ( n65020 , n41790 , n45552 );
buf ( n65021 , n65020 );
buf ( n65022 , n65021 );
buf ( n65023 , n65022 );
and ( n65024 , n65018 , n65023 );
and ( n65025 , n65015 , n65023 );
or ( n65026 , n65019 , n65024 , n65025 );
and ( n65027 , n63492 , n59207 );
not ( n65028 , n65027 );
and ( n65029 , n61505 , n61015 );
not ( n65030 , n65029 );
and ( n65031 , n65028 , n65030 );
buf ( n65032 , n65031 );
and ( n65033 , n65026 , n65032 );
xor ( n65034 , n64561 , n64565 );
xor ( n65035 , n65034 , n64570 );
and ( n65036 , n65032 , n65035 );
and ( n65037 , n65026 , n65035 );
or ( n65038 , n65033 , n65036 , n65037 );
and ( n65039 , n65010 , n65038 );
and ( n65040 , n64958 , n65038 );
or ( n65041 , n65011 , n65039 , n65040 );
and ( n65042 , n64906 , n65041 );
xor ( n65043 , n64578 , n64582 );
xor ( n65044 , n65043 , n64587 );
xor ( n65045 , n64604 , n64608 );
xor ( n65046 , n65045 , n64613 );
and ( n65047 , n65044 , n65046 );
xor ( n65048 , n64620 , n64624 );
xor ( n65049 , n65048 , n64629 );
and ( n65050 , n65046 , n65049 );
and ( n65051 , n65044 , n65049 );
or ( n65052 , n65047 , n65050 , n65051 );
xor ( n65053 , n64463 , n64465 );
xor ( n65054 , n65053 , n64468 );
and ( n65055 , n65052 , n65054 );
xor ( n65056 , n64477 , n64479 );
xor ( n65057 , n65056 , n64496 );
and ( n65058 , n65054 , n65057 );
and ( n65059 , n65052 , n65057 );
or ( n65060 , n65055 , n65058 , n65059 );
and ( n65061 , n65041 , n65060 );
and ( n65062 , n64906 , n65060 );
or ( n65063 , n65042 , n65061 , n65062 );
and ( n65064 , n64863 , n65063 );
and ( n65065 , n64792 , n65063 );
or ( n65066 , n64864 , n65064 , n65065 );
and ( n65067 , n64782 , n65066 );
xor ( n65068 , n64515 , n64531 );
xor ( n65069 , n65068 , n64542 );
xor ( n65070 , n64557 , n64573 );
xor ( n65071 , n65070 , n64590 );
and ( n65072 , n65069 , n65071 );
xor ( n65073 , n64616 , n64632 );
xor ( n65074 , n65073 , n64645 );
and ( n65075 , n65071 , n65074 );
and ( n65076 , n65069 , n65074 );
or ( n65077 , n65072 , n65075 , n65076 );
xor ( n65078 , n64435 , n64437 );
xor ( n65079 , n65078 , n64440 );
and ( n65080 , n65077 , n65079 );
xor ( n65081 , n64444 , n64460 );
xor ( n65082 , n65081 , n64471 );
and ( n65083 , n65079 , n65082 );
and ( n65084 , n65077 , n65082 );
or ( n65085 , n65080 , n65083 , n65084 );
xor ( n65086 , n64499 , n64545 );
xor ( n65087 , n65086 , n64593 );
xor ( n65088 , n64648 , n64658 );
xor ( n65089 , n65088 , n64669 );
and ( n65090 , n65087 , n65089 );
xor ( n65091 , n64674 , n64676 );
xor ( n65092 , n65091 , n64679 );
and ( n65093 , n65089 , n65092 );
and ( n65094 , n65087 , n65092 );
or ( n65095 , n65090 , n65093 , n65094 );
and ( n65096 , n65085 , n65095 );
xor ( n65097 , n64369 , n64371 );
xor ( n65098 , n65097 , n64374 );
and ( n65099 , n65095 , n65098 );
and ( n65100 , n65085 , n65098 );
or ( n65101 , n65096 , n65099 , n65100 );
and ( n65102 , n65066 , n65101 );
and ( n65103 , n64782 , n65101 );
or ( n65104 , n65067 , n65102 , n65103 );
xor ( n65105 , n64392 , n64409 );
xor ( n65106 , n65105 , n64430 );
xor ( n65107 , n64443 , n64474 );
xor ( n65108 , n65107 , n64596 );
and ( n65109 , n65106 , n65108 );
xor ( n65110 , n64672 , n64682 );
xor ( n65111 , n65110 , n64685 );
and ( n65112 , n65108 , n65111 );
and ( n65113 , n65106 , n65111 );
or ( n65114 , n65109 , n65112 , n65113 );
xor ( n65115 , n64364 , n64366 );
xor ( n65116 , n65115 , n64377 );
and ( n65117 , n65114 , n65116 );
xor ( n65118 , n64433 , n64599 );
xor ( n65119 , n65118 , n64688 );
and ( n65120 , n65116 , n65119 );
and ( n65121 , n65114 , n65119 );
or ( n65122 , n65117 , n65120 , n65121 );
and ( n65123 , n65104 , n65122 );
xor ( n65124 , n64340 , n64361 );
xor ( n65125 , n65124 , n64380 );
and ( n65126 , n65122 , n65125 );
and ( n65127 , n65104 , n65125 );
or ( n65128 , n65123 , n65126 , n65127 );
and ( n65129 , n64755 , n65128 );
and ( n65130 , n64737 , n65128 );
or ( n65131 , n64756 , n65129 , n65130 );
and ( n65132 , n64735 , n65131 );
xor ( n65133 , n64335 , n64337 );
xor ( n65134 , n65133 , n64721 );
and ( n65135 , n65131 , n65134 );
and ( n65136 , n64735 , n65134 );
or ( n65137 , n65132 , n65135 , n65136 );
xor ( n65138 , n64333 , n64724 );
xor ( n65139 , n65138 , n64727 );
and ( n65140 , n65137 , n65139 );
xor ( n65141 , n64383 , n64715 );
xor ( n65142 , n65141 , n64718 );
xor ( n65143 , n64691 , n64709 );
xor ( n65144 , n65143 , n64712 );
xor ( n65145 , n64701 , n64703 );
xor ( n65146 , n65145 , n64706 );
xor ( n65147 , n64693 , n64695 );
xor ( n65148 , n65147 , n64698 );
and ( n65149 , n64850 , n64852 );
and ( n65150 , n64852 , n64855 );
and ( n65151 , n64850 , n64855 );
or ( n65152 , n65149 , n65150 , n65151 );
xor ( n65153 , n64763 , n64765 );
xor ( n65154 , n65153 , n64768 );
and ( n65155 , n65152 , n65154 );
xor ( n65156 , n64454 , n64384 );
xor ( n65157 , n65156 , n64457 );
and ( n65158 , n65154 , n65157 );
and ( n65159 , n65152 , n65157 );
or ( n65160 , n65155 , n65158 , n65159 );
xor ( n65161 , n64771 , n64773 );
xor ( n65162 , n65161 , n64776 );
or ( n65163 , n65160 , n65162 );
and ( n65164 , n65148 , n65163 );
and ( n65165 , n58292 , n64811 );
not ( n65166 , n65165 );
and ( n65167 , n63024 , n59611 );
not ( n65168 , n65167 );
and ( n65169 , n65166 , n65168 );
and ( n65170 , n62377 , n60372 );
not ( n65171 , n65170 );
and ( n65172 , n65168 , n65171 );
and ( n65173 , n65166 , n65171 );
or ( n65174 , n65169 , n65172 , n65173 );
xor ( n65175 , n64806 , n64808 );
buf ( n65176 , n20241 );
buf ( n65177 , n65176 );
and ( n65178 , n65177 , n58294 );
not ( n65179 , n65178 );
and ( n65180 , n65175 , n65179 );
and ( n65181 , n62593 , n59920 );
not ( n65182 , n65181 );
and ( n65183 , n65179 , n65182 );
and ( n65184 , n65175 , n65182 );
or ( n65185 , n65180 , n65183 , n65184 );
and ( n65186 , n65174 , n65185 );
xor ( n65187 , n64796 , n64798 );
xor ( n65188 , n65187 , n64801 );
and ( n65189 , n65185 , n65188 );
and ( n65190 , n65174 , n65188 );
or ( n65191 , n65186 , n65189 , n65190 );
xor ( n65192 , n64804 , n64819 );
xor ( n65193 , n65192 , n64822 );
and ( n65194 , n65191 , n65193 );
xor ( n65195 , n64650 , n64652 );
xor ( n65196 , n65195 , n64655 );
xor ( n65197 , n64661 , n64663 );
xor ( n65198 , n65197 , n64666 );
and ( n65199 , n65196 , n65198 );
xor ( n65200 , n65152 , n65154 );
xor ( n65201 , n65200 , n65157 );
and ( n65202 , n65198 , n65201 );
and ( n65203 , n65196 , n65201 );
or ( n65204 , n65199 , n65202 , n65203 );
and ( n65205 , n65194 , n65204 );
and ( n65206 , n64221 , n58911 );
not ( n65207 , n65206 );
buf ( n65208 , n65207 );
buf ( n65209 , n20241 );
buf ( n65210 , n65209 );
and ( n65211 , n57948 , n65210 );
not ( n65212 , n65211 );
and ( n65213 , n65208 , n65212 );
and ( n65214 , n59615 , n62998 );
not ( n65215 , n65214 );
and ( n65216 , n65212 , n65215 );
and ( n65217 , n65208 , n65215 );
or ( n65218 , n65213 , n65216 , n65217 );
and ( n65219 , n59908 , n62868 );
not ( n65220 , n65219 );
and ( n65221 , n60376 , n62151 );
not ( n65222 , n65221 );
and ( n65223 , n65220 , n65222 );
and ( n65224 , n61008 , n61481 );
not ( n65225 , n65224 );
and ( n65226 , n65222 , n65225 );
and ( n65227 , n65220 , n65225 );
or ( n65228 , n65223 , n65226 , n65227 );
and ( n65229 , n65218 , n65228 );
xor ( n65230 , n64550 , n64551 );
xor ( n65231 , n65230 , n64554 );
and ( n65232 , n65228 , n65231 );
and ( n65233 , n65218 , n65231 );
or ( n65234 , n65229 , n65232 , n65233 );
xor ( n65235 , n64637 , n64210 );
xor ( n65236 , n65235 , n64642 );
xor ( n65237 , n64809 , n64813 );
xor ( n65238 , n65237 , n64816 );
and ( n65239 , n65236 , n65238 );
xor ( n65240 , n64830 , n64832 );
xor ( n65241 , n65240 , n64835 );
and ( n65242 , n65238 , n65241 );
and ( n65243 , n65236 , n65241 );
or ( n65244 , n65239 , n65242 , n65243 );
and ( n65245 , n65234 , n65244 );
xnor ( n65246 , n64848 , n64856 );
xor ( n65247 , n64866 , n64868 );
and ( n65248 , n65246 , n65247 );
xor ( n65249 , n64880 , n64884 );
xor ( n65250 , n65249 , n64889 );
xor ( n65251 , n64840 , n64842 );
xor ( n65252 , n65251 , n64845 );
and ( n65253 , n65250 , n65252 );
xnor ( n65254 , n64897 , n64899 );
and ( n65255 , n65252 , n65254 );
and ( n65256 , n65250 , n65254 );
or ( n65257 , n65253 , n65255 , n65256 );
and ( n65258 , n65247 , n65257 );
and ( n65259 , n65246 , n65257 );
or ( n65260 , n65248 , n65258 , n65259 );
and ( n65261 , n65244 , n65260 );
and ( n65262 , n65234 , n65260 );
or ( n65263 , n65245 , n65261 , n65262 );
and ( n65264 , n65204 , n65263 );
and ( n65265 , n65194 , n65263 );
or ( n65266 , n65205 , n65264 , n65265 );
and ( n65267 , n65163 , n65266 );
and ( n65268 , n65148 , n65266 );
or ( n65269 , n65164 , n65267 , n65268 );
and ( n65270 , n65146 , n65269 );
and ( n65271 , n58292 , n65210 );
not ( n65272 , n65271 );
and ( n65273 , n58628 , n64811 );
not ( n65274 , n65273 );
and ( n65275 , n65272 , n65274 );
and ( n65276 , n60376 , n62868 );
not ( n65277 , n65276 );
and ( n65278 , n65274 , n65277 );
and ( n65279 , n65272 , n65277 );
or ( n65280 , n65275 , n65278 , n65279 );
and ( n65281 , n64548 , n58542 );
not ( n65282 , n65281 );
and ( n65283 , n58915 , n64412 );
not ( n65284 , n65283 );
and ( n65285 , n65282 , n65284 );
and ( n65286 , n62593 , n60372 );
not ( n65287 , n65286 );
and ( n65288 , n65284 , n65287 );
and ( n65289 , n65282 , n65287 );
or ( n65290 , n65285 , n65288 , n65289 );
and ( n65291 , n65280 , n65290 );
and ( n65292 , n47351 , n57187 );
and ( n65293 , n47216 , n57184 );
nor ( n65294 , n65292 , n65293 );
xnor ( n65295 , n65294 , n56175 );
and ( n65296 , n51510 , n50783 );
and ( n65297 , n51298 , n50781 );
nor ( n65298 , n65296 , n65297 );
xnor ( n65299 , n65298 , n50557 );
or ( n65300 , n65295 , n65299 );
and ( n65301 , n65290 , n65300 );
and ( n65302 , n65280 , n65300 );
or ( n65303 , n65291 , n65301 , n65302 );
and ( n65304 , n47647 , n56503 );
and ( n65305 , n47474 , n56501 );
nor ( n65306 , n65304 , n65305 );
xnor ( n65307 , n65306 , n56178 );
and ( n65308 , n48632 , n54535 );
and ( n65309 , n48384 , n54533 );
nor ( n65310 , n65308 , n65309 );
xnor ( n65311 , n65310 , n54237 );
or ( n65312 , n65307 , n65311 );
and ( n65313 , n48272 , n55159 );
and ( n65314 , n48108 , n55157 );
nor ( n65315 , n65313 , n65314 );
xnor ( n65316 , n65315 , n54864 );
and ( n65317 , n48988 , n53928 );
and ( n65318 , n48709 , n53926 );
nor ( n65319 , n65317 , n65318 );
xnor ( n65320 , n65319 , n53652 );
or ( n65321 , n65316 , n65320 );
and ( n65322 , n65312 , n65321 );
and ( n65323 , n50195 , n52269 );
and ( n65324 , n49976 , n52267 );
nor ( n65325 , n65323 , n65324 );
xnor ( n65326 , n65325 , n52008 );
and ( n65327 , n50625 , n51750 );
and ( n65328 , n50404 , n51748 );
nor ( n65329 , n65327 , n65328 );
xnor ( n65330 , n65329 , n51520 );
and ( n65331 , n65326 , n65330 );
and ( n65332 , n65321 , n65331 );
and ( n65333 , n65312 , n65331 );
or ( n65334 , n65322 , n65332 , n65333 );
and ( n65335 , n65303 , n65334 );
and ( n65336 , n52082 , n50338 );
and ( n65337 , n51734 , n50336 );
nor ( n65338 , n65336 , n65337 );
xnor ( n65339 , n65338 , n50111 );
and ( n65340 , n52612 , n49896 );
and ( n65341 , n52332 , n49894 );
nor ( n65342 , n65340 , n65341 );
xnor ( n65343 , n65342 , n49711 );
and ( n65344 , n65339 , n65343 );
and ( n65345 , n47962 , n55851 );
and ( n65346 , n47778 , n55849 );
nor ( n65347 , n65345 , n65346 );
xnor ( n65348 , n65347 , n55506 );
and ( n65349 , n49374 , n53357 );
and ( n65350 , n49115 , n53355 );
nor ( n65351 , n65349 , n65350 );
xnor ( n65352 , n65351 , n53060 );
and ( n65353 , n65348 , n65352 );
and ( n65354 , n49781 , n52799 );
and ( n65355 , n49570 , n52797 );
nor ( n65356 , n65354 , n65355 );
xnor ( n65357 , n65356 , n52538 );
and ( n65358 , n65352 , n65357 );
and ( n65359 , n65348 , n65357 );
or ( n65360 , n65353 , n65358 , n65359 );
and ( n65361 , n65344 , n65360 );
and ( n65362 , n51077 , n51221 );
and ( n65363 , n50726 , n51219 );
nor ( n65364 , n65362 , n65363 );
xnor ( n65365 , n65364 , n51000 );
and ( n65366 , n53041 , n49513 );
and ( n65367 , n52790 , n49511 );
nor ( n65368 , n65366 , n65367 );
xnor ( n65369 , n65368 , n49310 );
and ( n65370 , n65365 , n65369 );
and ( n65371 , n53639 , n49121 );
and ( n65372 , n53328 , n49119 );
nor ( n65373 , n65371 , n65372 );
xnor ( n65374 , n65373 , n48932 );
and ( n65375 , n65369 , n65374 );
and ( n65376 , n65365 , n65374 );
or ( n65377 , n65370 , n65375 , n65376 );
and ( n65378 , n65360 , n65377 );
and ( n65379 , n65344 , n65377 );
or ( n65380 , n65361 , n65378 , n65379 );
and ( n65381 , n65334 , n65380 );
and ( n65382 , n65303 , n65380 );
or ( n65383 , n65335 , n65381 , n65382 );
and ( n65384 , n54227 , n48740 );
and ( n65385 , n53922 , n48738 );
nor ( n65386 , n65384 , n65385 );
xnor ( n65387 , n65386 , n48571 );
and ( n65388 , n54942 , n48394 );
and ( n65389 , n54604 , n48392 );
nor ( n65390 , n65388 , n65389 );
xnor ( n65391 , n65390 , n48220 );
and ( n65392 , n65387 , n65391 );
and ( n65393 , n55497 , n48042 );
and ( n65394 , n55143 , n48040 );
nor ( n65395 , n65393 , n65394 );
xnor ( n65396 , n65395 , n47921 );
and ( n65397 , n65391 , n65396 );
and ( n65398 , n65387 , n65396 );
or ( n65399 , n65392 , n65397 , n65398 );
and ( n65400 , n56255 , n47734 );
and ( n65401 , n55756 , n47732 );
nor ( n65402 , n65400 , n65401 );
xnor ( n65403 , n65402 , n47606 );
and ( n65404 , n56915 , n47429 );
and ( n65405 , n56388 , n47427 );
nor ( n65406 , n65404 , n65405 );
xnor ( n65407 , n65406 , n47309 );
and ( n65408 , n65403 , n65407 );
and ( n65409 , n65407 , n65016 );
and ( n65410 , n65403 , n65016 );
or ( n65411 , n65408 , n65409 , n65410 );
and ( n65412 , n65399 , n65411 );
xor ( n65413 , n41793 , n45550 );
buf ( n65414 , n65413 );
buf ( n65415 , n65414 );
buf ( n65416 , n65415 );
and ( n65417 , n63987 , n59207 );
not ( n65418 , n65417 );
and ( n65419 , n65416 , n65418 );
and ( n65420 , n62377 , n60711 );
not ( n65421 , n65420 );
and ( n65422 , n65418 , n65421 );
and ( n65423 , n65416 , n65421 );
or ( n65424 , n65419 , n65422 , n65423 );
and ( n65425 , n65411 , n65424 );
and ( n65426 , n65399 , n65424 );
or ( n65427 , n65412 , n65425 , n65426 );
xor ( n65428 , n64910 , n64914 );
xor ( n65429 , n65428 , n64919 );
xor ( n65430 , n64926 , n64930 );
xor ( n65431 , n65430 , n64935 );
and ( n65432 , n65429 , n65431 );
xor ( n65433 , n64943 , n64947 );
xor ( n65434 , n65433 , n64952 );
and ( n65435 , n65431 , n65434 );
and ( n65436 , n65429 , n65434 );
or ( n65437 , n65432 , n65435 , n65436 );
and ( n65438 , n65427 , n65437 );
xor ( n65439 , n64962 , n64966 );
xor ( n65440 , n65439 , n64971 );
xor ( n65441 , n64978 , n64982 );
xor ( n65442 , n65441 , n64987 );
and ( n65443 , n65440 , n65442 );
xor ( n65444 , n64995 , n64999 );
xor ( n65445 , n65444 , n65004 );
and ( n65446 , n65442 , n65445 );
and ( n65447 , n65440 , n65445 );
or ( n65448 , n65443 , n65446 , n65447 );
and ( n65449 , n65437 , n65448 );
and ( n65450 , n65427 , n65448 );
or ( n65451 , n65438 , n65449 , n65450 );
and ( n65452 , n65383 , n65451 );
buf ( n65453 , n64871 );
xor ( n65454 , n65453 , n64873 );
xor ( n65455 , n64892 , n64894 );
xor ( n65456 , n65455 , n64900 );
and ( n65457 , n65454 , n65456 );
xor ( n65458 , n64922 , n64938 );
xor ( n65459 , n65458 , n64955 );
and ( n65460 , n65456 , n65459 );
and ( n65461 , n65454 , n65459 );
or ( n65462 , n65457 , n65460 , n65461 );
and ( n65463 , n65451 , n65462 );
and ( n65464 , n65383 , n65462 );
or ( n65465 , n65452 , n65463 , n65464 );
xor ( n65466 , n64974 , n64990 );
xor ( n65467 , n65466 , n65007 );
xor ( n65468 , n65026 , n65032 );
xor ( n65469 , n65468 , n65035 );
and ( n65470 , n65467 , n65469 );
xor ( n65471 , n65044 , n65046 );
xor ( n65472 , n65471 , n65049 );
and ( n65473 , n65469 , n65472 );
and ( n65474 , n65467 , n65472 );
or ( n65475 , n65470 , n65473 , n65474 );
xor ( n65476 , n64828 , n64838 );
xor ( n65477 , n65476 , n64857 );
and ( n65478 , n65475 , n65477 );
xor ( n65479 , n64869 , n64875 );
xor ( n65480 , n65479 , n64903 );
and ( n65481 , n65477 , n65480 );
and ( n65482 , n65475 , n65480 );
or ( n65483 , n65478 , n65481 , n65482 );
and ( n65484 , n65465 , n65483 );
xor ( n65485 , n64958 , n65010 );
xor ( n65486 , n65485 , n65038 );
xor ( n65487 , n65052 , n65054 );
xor ( n65488 , n65487 , n65057 );
and ( n65489 , n65486 , n65488 );
xor ( n65490 , n65069 , n65071 );
xor ( n65491 , n65490 , n65074 );
and ( n65492 , n65488 , n65491 );
and ( n65493 , n65486 , n65491 );
or ( n65494 , n65489 , n65492 , n65493 );
and ( n65495 , n65483 , n65494 );
and ( n65496 , n65465 , n65494 );
or ( n65497 , n65484 , n65495 , n65496 );
xor ( n65498 , n64784 , n64786 );
xor ( n65499 , n65498 , n64789 );
xor ( n65500 , n64794 , n64825 );
xor ( n65501 , n65500 , n64860 );
and ( n65502 , n65499 , n65501 );
xor ( n65503 , n64906 , n65041 );
xor ( n65504 , n65503 , n65060 );
and ( n65505 , n65501 , n65504 );
and ( n65506 , n65499 , n65504 );
or ( n65507 , n65502 , n65505 , n65506 );
and ( n65508 , n65497 , n65507 );
xor ( n65509 , n64758 , n64760 );
xor ( n65510 , n65509 , n64779 );
and ( n65511 , n65507 , n65510 );
and ( n65512 , n65497 , n65510 );
or ( n65513 , n65508 , n65511 , n65512 );
and ( n65514 , n65269 , n65513 );
and ( n65515 , n65146 , n65513 );
or ( n65516 , n65270 , n65514 , n65515 );
and ( n65517 , n65144 , n65516 );
xor ( n65518 , n64792 , n64863 );
xor ( n65519 , n65518 , n65063 );
xor ( n65520 , n65085 , n65095 );
xor ( n65521 , n65520 , n65098 );
and ( n65522 , n65519 , n65521 );
xor ( n65523 , n65106 , n65108 );
xor ( n65524 , n65523 , n65111 );
and ( n65525 , n65521 , n65524 );
and ( n65526 , n65519 , n65524 );
or ( n65527 , n65522 , n65525 , n65526 );
xor ( n65528 , n64744 , n64746 );
xor ( n65529 , n65528 , n64749 );
and ( n65530 , n65527 , n65529 );
xor ( n65531 , n64782 , n65066 );
xor ( n65532 , n65531 , n65101 );
and ( n65533 , n65529 , n65532 );
and ( n65534 , n65527 , n65532 );
or ( n65535 , n65530 , n65533 , n65534 );
and ( n65536 , n65516 , n65535 );
and ( n65537 , n65144 , n65535 );
or ( n65538 , n65517 , n65536 , n65537 );
and ( n65539 , n65142 , n65538 );
xor ( n65540 , n64737 , n64755 );
xor ( n65541 , n65540 , n65128 );
and ( n65542 , n65538 , n65541 );
and ( n65543 , n65142 , n65541 );
or ( n65544 , n65539 , n65542 , n65543 );
xor ( n65545 , n64735 , n65131 );
xor ( n65546 , n65545 , n65134 );
and ( n65547 , n65544 , n65546 );
xor ( n65548 , n64739 , n64741 );
xor ( n65549 , n65548 , n64752 );
xor ( n65550 , n65104 , n65122 );
xor ( n65551 , n65550 , n65125 );
and ( n65552 , n65549 , n65551 );
xor ( n65553 , n65114 , n65116 );
xor ( n65554 , n65553 , n65119 );
xor ( n65555 , n65077 , n65079 );
xor ( n65556 , n65555 , n65082 );
xor ( n65557 , n65087 , n65089 );
xor ( n65558 , n65557 , n65092 );
and ( n65559 , n65556 , n65558 );
xnor ( n65560 , n65160 , n65162 );
and ( n65561 , n65558 , n65560 );
and ( n65562 , n65556 , n65560 );
or ( n65563 , n65559 , n65561 , n65562 );
xor ( n65564 , n65191 , n65193 );
xor ( n65565 , n65218 , n65228 );
xor ( n65566 , n65565 , n65231 );
xor ( n65567 , n65174 , n65185 );
xor ( n65568 , n65567 , n65188 );
and ( n65569 , n65566 , n65568 );
and ( n65570 , n65177 , n58444 );
not ( n65571 , n65570 );
and ( n65572 , n59908 , n62998 );
not ( n65573 , n65572 );
and ( n65574 , n65571 , n65573 );
buf ( n65575 , n61505 );
not ( n65576 , n65575 );
and ( n65577 , n65573 , n65576 );
and ( n65578 , n65571 , n65576 );
or ( n65579 , n65574 , n65577 , n65578 );
and ( n65580 , n64548 , n58911 );
not ( n65581 , n65580 );
and ( n65582 , n60376 , n62998 );
not ( n65583 , n65582 );
and ( n65584 , n65581 , n65583 );
buf ( n65585 , n20244 );
buf ( n65586 , n65585 );
and ( n65587 , n57948 , n65586 );
not ( n65588 , n65587 );
and ( n65589 , n65584 , n65588 );
and ( n65590 , n63492 , n59611 );
not ( n65591 , n65590 );
and ( n65592 , n65588 , n65591 );
and ( n65593 , n65584 , n65591 );
or ( n65594 , n65589 , n65592 , n65593 );
and ( n65595 , n65579 , n65594 );
and ( n65596 , n60821 , n61914 );
not ( n65597 , n65596 );
and ( n65598 , n65594 , n65597 );
and ( n65599 , n65579 , n65597 );
or ( n65600 , n65595 , n65598 , n65599 );
and ( n65601 , n65568 , n65600 );
and ( n65602 , n65566 , n65600 );
or ( n65603 , n65569 , n65601 , n65602 );
and ( n65604 , n65564 , n65603 );
buf ( n65605 , n20244 );
buf ( n65606 , n65605 );
and ( n65607 , n65606 , n58294 );
not ( n65608 , n65607 );
and ( n65609 , n65608 , n65206 );
and ( n65610 , n63024 , n59920 );
not ( n65611 , n65610 );
and ( n65612 , n65206 , n65611 );
and ( n65613 , n65608 , n65611 );
or ( n65614 , n65609 , n65612 , n65613 );
xor ( n65615 , n65208 , n65212 );
xor ( n65616 , n65615 , n65215 );
and ( n65617 , n65614 , n65616 );
xor ( n65618 , n65220 , n65222 );
xor ( n65619 , n65618 , n65225 );
and ( n65620 , n65616 , n65619 );
and ( n65621 , n65614 , n65619 );
or ( n65622 , n65617 , n65620 , n65621 );
and ( n65623 , n59365 , n63766 );
not ( n65624 , n65623 );
and ( n65625 , n61918 , n61015 );
not ( n65626 , n65625 );
and ( n65627 , n65624 , n65626 );
xor ( n65628 , n65282 , n65284 );
xor ( n65629 , n65628 , n65287 );
and ( n65630 , n65626 , n65629 );
and ( n65631 , n65624 , n65629 );
or ( n65632 , n65627 , n65630 , n65631 );
xor ( n65633 , n65166 , n65168 );
xor ( n65634 , n65633 , n65171 );
and ( n65635 , n65632 , n65634 );
xor ( n65636 , n65175 , n65179 );
xor ( n65637 , n65636 , n65182 );
and ( n65638 , n65634 , n65637 );
and ( n65639 , n65632 , n65637 );
or ( n65640 , n65635 , n65638 , n65639 );
and ( n65641 , n65622 , n65640 );
xor ( n65642 , n65015 , n65018 );
xor ( n65643 , n65642 , n65023 );
xor ( n65644 , n65028 , n65030 );
buf ( n65645 , n65644 );
and ( n65646 , n65643 , n65645 );
and ( n65647 , n58915 , n64811 );
not ( n65648 , n65647 );
buf ( n65649 , n65648 );
and ( n65650 , n59615 , n63679 );
not ( n65651 , n65650 );
and ( n65652 , n65649 , n65651 );
and ( n65653 , n61008 , n61914 );
not ( n65654 , n65653 );
and ( n65655 , n65651 , n65654 );
and ( n65656 , n65649 , n65654 );
or ( n65657 , n65652 , n65655 , n65656 );
and ( n65658 , n65645 , n65657 );
and ( n65659 , n65643 , n65657 );
or ( n65660 , n65646 , n65658 , n65659 );
and ( n65661 , n65640 , n65660 );
and ( n65662 , n65622 , n65660 );
or ( n65663 , n65641 , n65661 , n65662 );
and ( n65664 , n65603 , n65663 );
and ( n65665 , n65564 , n65663 );
or ( n65666 , n65604 , n65664 , n65665 );
and ( n65667 , n58292 , n65586 );
not ( n65668 , n65667 );
and ( n65669 , n61008 , n62151 );
not ( n65670 , n65669 );
and ( n65671 , n65668 , n65670 );
and ( n65672 , n61505 , n61914 );
not ( n65673 , n65672 );
and ( n65674 , n65670 , n65673 );
and ( n65675 , n65668 , n65673 );
or ( n65676 , n65671 , n65674 , n65675 );
buf ( n65677 , n20247 );
buf ( n65678 , n65677 );
and ( n65679 , n65678 , n58294 );
not ( n65680 , n65679 );
and ( n65681 , n65680 , n65647 );
and ( n65682 , n59908 , n63679 );
not ( n65683 , n65682 );
and ( n65684 , n65647 , n65683 );
and ( n65685 , n65680 , n65683 );
or ( n65686 , n65681 , n65684 , n65685 );
and ( n65687 , n65676 , n65686 );
xor ( n65688 , n65272 , n65274 );
xor ( n65689 , n65688 , n65277 );
and ( n65690 , n65686 , n65689 );
and ( n65691 , n65676 , n65689 );
or ( n65692 , n65687 , n65690 , n65691 );
xnor ( n65693 , n65295 , n65299 );
xnor ( n65694 , n65307 , n65311 );
and ( n65695 , n65693 , n65694 );
buf ( n65696 , n65695 );
and ( n65697 , n65692 , n65696 );
xnor ( n65698 , n65316 , n65320 );
xor ( n65699 , n65326 , n65330 );
and ( n65700 , n65698 , n65699 );
xor ( n65701 , n65339 , n65343 );
and ( n65702 , n65699 , n65701 );
and ( n65703 , n65698 , n65701 );
or ( n65704 , n65700 , n65702 , n65703 );
and ( n65705 , n65696 , n65704 );
and ( n65706 , n65692 , n65704 );
or ( n65707 , n65697 , n65705 , n65706 );
and ( n65708 , n47778 , n56503 );
and ( n65709 , n47647 , n56501 );
nor ( n65710 , n65708 , n65709 );
xnor ( n65711 , n65710 , n56178 );
and ( n65712 , n48384 , n55159 );
and ( n65713 , n48272 , n55157 );
nor ( n65714 , n65712 , n65713 );
xnor ( n65715 , n65714 , n54864 );
and ( n65716 , n65711 , n65715 );
and ( n65717 , n48709 , n54535 );
and ( n65718 , n48632 , n54533 );
nor ( n65719 , n65717 , n65718 );
xnor ( n65720 , n65719 , n54237 );
and ( n65721 , n65715 , n65720 );
and ( n65722 , n65711 , n65720 );
or ( n65723 , n65716 , n65721 , n65722 );
and ( n65724 , n54604 , n48740 );
and ( n65725 , n54227 , n48738 );
nor ( n65726 , n65724 , n65725 );
xnor ( n65727 , n65726 , n48571 );
and ( n65728 , n56388 , n47734 );
and ( n65729 , n56255 , n47732 );
nor ( n65730 , n65728 , n65729 );
xnor ( n65731 , n65730 , n47606 );
and ( n65732 , n65727 , n65731 );
and ( n65733 , n57063 , n47427 );
not ( n65734 , n65733 );
and ( n65735 , n65734 , n47309 );
and ( n65736 , n65731 , n65735 );
and ( n65737 , n65727 , n65735 );
or ( n65738 , n65732 , n65736 , n65737 );
and ( n65739 , n65723 , n65738 );
and ( n65740 , n47474 , n57187 );
and ( n65741 , n47351 , n57184 );
nor ( n65742 , n65740 , n65741 );
xnor ( n65743 , n65742 , n56175 );
and ( n65744 , n51734 , n50783 );
and ( n65745 , n51510 , n50781 );
nor ( n65746 , n65744 , n65745 );
xnor ( n65747 , n65746 , n50557 );
or ( n65748 , n65743 , n65747 );
and ( n65749 , n65738 , n65748 );
and ( n65750 , n65723 , n65748 );
or ( n65751 , n65739 , n65749 , n65750 );
and ( n65752 , n65177 , n58542 );
not ( n65753 , n65752 );
and ( n65754 , n63024 , n60372 );
not ( n65755 , n65754 );
or ( n65756 , n65753 , n65755 );
and ( n65757 , n48108 , n55851 );
and ( n65758 , n47962 , n55849 );
nor ( n65759 , n65757 , n65758 );
xnor ( n65760 , n65759 , n55506 );
and ( n65761 , n49115 , n53928 );
and ( n65762 , n48988 , n53926 );
nor ( n65763 , n65761 , n65762 );
xnor ( n65764 , n65763 , n53652 );
and ( n65765 , n65760 , n65764 );
and ( n65766 , n49570 , n53357 );
and ( n65767 , n49374 , n53355 );
nor ( n65768 , n65766 , n65767 );
xnor ( n65769 , n65768 , n53060 );
and ( n65770 , n65764 , n65769 );
and ( n65771 , n65760 , n65769 );
or ( n65772 , n65765 , n65770 , n65771 );
and ( n65773 , n65756 , n65772 );
and ( n65774 , n49976 , n52799 );
and ( n65775 , n49781 , n52797 );
nor ( n65776 , n65774 , n65775 );
xnor ( n65777 , n65776 , n52538 );
and ( n65778 , n50404 , n52269 );
and ( n65779 , n50195 , n52267 );
nor ( n65780 , n65778 , n65779 );
xnor ( n65781 , n65780 , n52008 );
and ( n65782 , n65777 , n65781 );
and ( n65783 , n50726 , n51750 );
and ( n65784 , n50625 , n51748 );
nor ( n65785 , n65783 , n65784 );
xnor ( n65786 , n65785 , n51520 );
and ( n65787 , n65781 , n65786 );
and ( n65788 , n65777 , n65786 );
or ( n65789 , n65782 , n65787 , n65788 );
and ( n65790 , n65772 , n65789 );
and ( n65791 , n65756 , n65789 );
or ( n65792 , n65773 , n65790 , n65791 );
and ( n65793 , n65751 , n65792 );
and ( n65794 , n51298 , n51221 );
and ( n65795 , n51077 , n51219 );
nor ( n65796 , n65794 , n65795 );
xnor ( n65797 , n65796 , n51000 );
and ( n65798 , n52790 , n49896 );
and ( n65799 , n52612 , n49894 );
nor ( n65800 , n65798 , n65799 );
xnor ( n65801 , n65800 , n49711 );
and ( n65802 , n65797 , n65801 );
and ( n65803 , n53328 , n49513 );
and ( n65804 , n53041 , n49511 );
nor ( n65805 , n65803 , n65804 );
xnor ( n65806 , n65805 , n49310 );
and ( n65807 , n65801 , n65806 );
and ( n65808 , n65797 , n65806 );
or ( n65809 , n65802 , n65807 , n65808 );
and ( n65810 , n53922 , n49121 );
and ( n65811 , n53639 , n49119 );
nor ( n65812 , n65810 , n65811 );
xnor ( n65813 , n65812 , n48932 );
and ( n65814 , n55143 , n48394 );
and ( n65815 , n54942 , n48392 );
nor ( n65816 , n65814 , n65815 );
xnor ( n65817 , n65816 , n48220 );
and ( n65818 , n65813 , n65817 );
and ( n65819 , n55756 , n48042 );
and ( n65820 , n55497 , n48040 );
nor ( n65821 , n65819 , n65820 );
xnor ( n65822 , n65821 , n47921 );
and ( n65823 , n65817 , n65822 );
and ( n65824 , n65813 , n65822 );
or ( n65825 , n65818 , n65823 , n65824 );
and ( n65826 , n65809 , n65825 );
and ( n65827 , n57063 , n47429 );
and ( n65828 , n56915 , n47427 );
nor ( n65829 , n65827 , n65828 );
xnor ( n65830 , n65829 , n47309 );
xor ( n65831 , n41796 , n45548 );
buf ( n65832 , n65831 );
buf ( n65833 , n65832 );
buf ( n65834 , n65833 );
and ( n65835 , n65830 , n65834 );
and ( n65836 , n63492 , n59920 );
not ( n65837 , n65836 );
and ( n65838 , n65834 , n65837 );
and ( n65839 , n65830 , n65837 );
or ( n65840 , n65835 , n65838 , n65839 );
and ( n65841 , n65825 , n65840 );
and ( n65842 , n65809 , n65840 );
or ( n65843 , n65826 , n65841 , n65842 );
and ( n65844 , n65792 , n65843 );
and ( n65845 , n65751 , n65843 );
or ( n65846 , n65793 , n65844 , n65845 );
and ( n65847 , n65707 , n65846 );
xor ( n65848 , n65348 , n65352 );
xor ( n65849 , n65848 , n65357 );
xor ( n65850 , n65365 , n65369 );
xor ( n65851 , n65850 , n65374 );
and ( n65852 , n65849 , n65851 );
xor ( n65853 , n65387 , n65391 );
xor ( n65854 , n65853 , n65396 );
and ( n65855 , n65851 , n65854 );
and ( n65856 , n65849 , n65854 );
or ( n65857 , n65852 , n65855 , n65856 );
xor ( n65858 , n65250 , n65252 );
xor ( n65859 , n65858 , n65254 );
and ( n65860 , n65857 , n65859 );
xor ( n65861 , n65280 , n65290 );
xor ( n65862 , n65861 , n65300 );
and ( n65863 , n65859 , n65862 );
and ( n65864 , n65857 , n65862 );
or ( n65865 , n65860 , n65863 , n65864 );
and ( n65866 , n65846 , n65865 );
and ( n65867 , n65707 , n65865 );
or ( n65868 , n65847 , n65866 , n65867 );
xor ( n65869 , n65312 , n65321 );
xor ( n65870 , n65869 , n65331 );
xor ( n65871 , n65344 , n65360 );
xor ( n65872 , n65871 , n65377 );
and ( n65873 , n65870 , n65872 );
xor ( n65874 , n65399 , n65411 );
xor ( n65875 , n65874 , n65424 );
and ( n65876 , n65872 , n65875 );
and ( n65877 , n65870 , n65875 );
or ( n65878 , n65873 , n65876 , n65877 );
xor ( n65879 , n65236 , n65238 );
xor ( n65880 , n65879 , n65241 );
and ( n65881 , n65878 , n65880 );
xor ( n65882 , n65246 , n65247 );
xor ( n65883 , n65882 , n65257 );
and ( n65884 , n65880 , n65883 );
and ( n65885 , n65878 , n65883 );
or ( n65886 , n65881 , n65884 , n65885 );
and ( n65887 , n65868 , n65886 );
xor ( n65888 , n65303 , n65334 );
xor ( n65889 , n65888 , n65380 );
xor ( n65890 , n65427 , n65437 );
xor ( n65891 , n65890 , n65448 );
and ( n65892 , n65889 , n65891 );
xor ( n65893 , n65454 , n65456 );
xor ( n65894 , n65893 , n65459 );
and ( n65895 , n65891 , n65894 );
and ( n65896 , n65889 , n65894 );
or ( n65897 , n65892 , n65895 , n65896 );
and ( n65898 , n65886 , n65897 );
and ( n65899 , n65868 , n65897 );
or ( n65900 , n65887 , n65898 , n65899 );
and ( n65901 , n65666 , n65900 );
xor ( n65902 , n65196 , n65198 );
xor ( n65903 , n65902 , n65201 );
xor ( n65904 , n65234 , n65244 );
xor ( n65905 , n65904 , n65260 );
and ( n65906 , n65903 , n65905 );
xor ( n65907 , n65383 , n65451 );
xor ( n65908 , n65907 , n65462 );
and ( n65909 , n65905 , n65908 );
and ( n65910 , n65903 , n65908 );
or ( n65911 , n65906 , n65909 , n65910 );
and ( n65912 , n65900 , n65911 );
and ( n65913 , n65666 , n65911 );
or ( n65914 , n65901 , n65912 , n65913 );
and ( n65915 , n65563 , n65914 );
xor ( n65916 , n65194 , n65204 );
xor ( n65917 , n65916 , n65263 );
xor ( n65918 , n65465 , n65483 );
xor ( n65919 , n65918 , n65494 );
and ( n65920 , n65917 , n65919 );
xor ( n65921 , n65499 , n65501 );
xor ( n65922 , n65921 , n65504 );
and ( n65923 , n65919 , n65922 );
and ( n65924 , n65917 , n65922 );
or ( n65925 , n65920 , n65923 , n65924 );
and ( n65926 , n65914 , n65925 );
and ( n65927 , n65563 , n65925 );
or ( n65928 , n65915 , n65926 , n65927 );
and ( n65929 , n65554 , n65928 );
xor ( n65930 , n65148 , n65163 );
xor ( n65931 , n65930 , n65266 );
xor ( n65932 , n65497 , n65507 );
xor ( n65933 , n65932 , n65510 );
and ( n65934 , n65931 , n65933 );
xor ( n65935 , n65519 , n65521 );
xor ( n65936 , n65935 , n65524 );
and ( n65937 , n65933 , n65936 );
and ( n65938 , n65931 , n65936 );
or ( n65939 , n65934 , n65937 , n65938 );
and ( n65940 , n65928 , n65939 );
and ( n65941 , n65554 , n65939 );
or ( n65942 , n65929 , n65940 , n65941 );
and ( n65943 , n65551 , n65942 );
and ( n65944 , n65549 , n65942 );
or ( n65945 , n65552 , n65943 , n65944 );
xor ( n65946 , n65142 , n65538 );
xor ( n65947 , n65946 , n65541 );
and ( n65948 , n65945 , n65947 );
xor ( n65949 , n65144 , n65516 );
xor ( n65950 , n65949 , n65535 );
xor ( n65951 , n65146 , n65269 );
xor ( n65952 , n65951 , n65513 );
xor ( n65953 , n65527 , n65529 );
xor ( n65954 , n65953 , n65532 );
and ( n65955 , n65952 , n65954 );
xor ( n65956 , n65475 , n65477 );
xor ( n65957 , n65956 , n65480 );
xor ( n65958 , n65486 , n65488 );
xor ( n65959 , n65958 , n65491 );
and ( n65960 , n65957 , n65959 );
xor ( n65961 , n65467 , n65469 );
xor ( n65962 , n65961 , n65472 );
and ( n65963 , n65177 , n58911 );
not ( n65964 , n65963 );
buf ( n65965 , n65964 );
and ( n65966 , n59365 , n64412 );
not ( n65967 , n65966 );
and ( n65968 , n65965 , n65967 );
and ( n65969 , n59615 , n63766 );
not ( n65970 , n65969 );
and ( n65971 , n65967 , n65970 );
and ( n65972 , n65965 , n65970 );
or ( n65973 , n65968 , n65971 , n65972 );
xor ( n65974 , n65649 , n65651 );
xor ( n65975 , n65974 , n65654 );
and ( n65976 , n65973 , n65975 );
xor ( n65977 , n65608 , n65206 );
xor ( n65978 , n65977 , n65611 );
and ( n65979 , n65975 , n65978 );
and ( n65980 , n65973 , n65978 );
or ( n65981 , n65976 , n65979 , n65980 );
xor ( n65982 , n65614 , n65616 );
xor ( n65983 , n65982 , n65619 );
or ( n65984 , n65981 , n65983 );
and ( n65985 , n65962 , n65984 );
xor ( n65986 , n65429 , n65431 );
xor ( n65987 , n65986 , n65434 );
xor ( n65988 , n65440 , n65442 );
xor ( n65989 , n65988 , n65445 );
and ( n65990 , n65987 , n65989 );
xor ( n65991 , n65579 , n65594 );
xor ( n65992 , n65991 , n65597 );
and ( n65993 , n65989 , n65992 );
and ( n65994 , n65987 , n65992 );
or ( n65995 , n65990 , n65993 , n65994 );
and ( n65996 , n65984 , n65995 );
and ( n65997 , n65962 , n65995 );
or ( n65998 , n65985 , n65996 , n65997 );
and ( n65999 , n65959 , n65998 );
and ( n66000 , n65957 , n65998 );
or ( n66001 , n65960 , n65999 , n66000 );
xor ( n66002 , n65632 , n65634 );
xor ( n66003 , n66002 , n65637 );
buf ( n66004 , n20247 );
buf ( n66005 , n66004 );
and ( n66006 , n57948 , n66005 );
not ( n66007 , n66006 );
and ( n66008 , n65606 , n58444 );
not ( n66009 , n66008 );
and ( n66010 , n66007 , n66009 );
and ( n66011 , n58628 , n65210 );
not ( n66012 , n66011 );
and ( n66013 , n66009 , n66012 );
and ( n66014 , n66007 , n66012 );
or ( n66015 , n66010 , n66013 , n66014 );
xor ( n66016 , n65581 , n65583 );
and ( n66017 , n63987 , n59611 );
not ( n66018 , n66017 );
and ( n66019 , n66016 , n66018 );
and ( n66020 , n62377 , n61015 );
not ( n66021 , n66020 );
and ( n66022 , n66018 , n66021 );
and ( n66023 , n66016 , n66021 );
or ( n66024 , n66019 , n66022 , n66023 );
and ( n66025 , n66015 , n66024 );
and ( n66026 , n60821 , n62151 );
not ( n66027 , n66026 );
and ( n66028 , n66024 , n66027 );
and ( n66029 , n66015 , n66027 );
or ( n66030 , n66025 , n66028 , n66029 );
and ( n66031 , n66003 , n66030 );
xor ( n66032 , n65571 , n65573 );
xor ( n66033 , n66032 , n65576 );
xor ( n66034 , n65584 , n65588 );
xor ( n66035 , n66034 , n65591 );
or ( n66036 , n66033 , n66035 );
and ( n66037 , n66030 , n66036 );
and ( n66038 , n66003 , n66036 );
or ( n66039 , n66031 , n66037 , n66038 );
xor ( n66040 , n65403 , n65407 );
xor ( n66041 , n66040 , n65016 );
xor ( n66042 , n65416 , n65418 );
xor ( n66043 , n66042 , n65421 );
and ( n66044 , n66041 , n66043 );
xor ( n66045 , n65676 , n65686 );
xor ( n66046 , n66045 , n65689 );
and ( n66047 , n66043 , n66046 );
and ( n66048 , n66041 , n66046 );
or ( n66049 , n66044 , n66047 , n66048 );
and ( n66050 , n59365 , n64811 );
not ( n66051 , n66050 );
and ( n66052 , n65963 , n66051 );
and ( n66053 , n60821 , n62998 );
not ( n66054 , n66053 );
and ( n66055 , n66051 , n66054 );
and ( n66056 , n65963 , n66054 );
or ( n66057 , n66052 , n66055 , n66056 );
xor ( n66058 , n65668 , n65670 );
xor ( n66059 , n66058 , n65673 );
and ( n66060 , n66057 , n66059 );
xor ( n66061 , n65680 , n65647 );
xor ( n66062 , n66061 , n65683 );
and ( n66063 , n66059 , n66062 );
and ( n66064 , n66057 , n66062 );
or ( n66065 , n66060 , n66063 , n66064 );
and ( n66066 , n47962 , n56503 );
and ( n66067 , n47778 , n56501 );
nor ( n66068 , n66066 , n66067 );
xnor ( n66069 , n66068 , n56178 );
and ( n66070 , n48632 , n55159 );
and ( n66071 , n48384 , n55157 );
nor ( n66072 , n66070 , n66071 );
xnor ( n66073 , n66072 , n54864 );
and ( n66074 , n66069 , n66073 );
and ( n66075 , n52082 , n50783 );
and ( n66076 , n51734 , n50781 );
nor ( n66077 , n66075 , n66076 );
xnor ( n66078 , n66077 , n50557 );
and ( n66079 , n66073 , n66078 );
and ( n66080 , n66069 , n66078 );
or ( n66081 , n66074 , n66079 , n66080 );
and ( n66082 , n52332 , n50338 );
and ( n66083 , n52082 , n50336 );
nor ( n66084 , n66082 , n66083 );
xnor ( n66085 , n66084 , n50111 );
or ( n66086 , n66081 , n66085 );
and ( n66087 , n66065 , n66086 );
and ( n66088 , n61918 , n61481 );
not ( n66089 , n66088 );
xor ( n66090 , n65711 , n65715 );
xor ( n66091 , n66090 , n65720 );
and ( n66092 , n66089 , n66091 );
buf ( n66093 , n66092 );
and ( n66094 , n66086 , n66093 );
and ( n66095 , n66065 , n66093 );
or ( n66096 , n66087 , n66094 , n66095 );
and ( n66097 , n66049 , n66096 );
xor ( n66098 , n65727 , n65731 );
xor ( n66099 , n66098 , n65735 );
xnor ( n66100 , n65743 , n65747 );
and ( n66101 , n66099 , n66100 );
xnor ( n66102 , n65753 , n65755 );
and ( n66103 , n66100 , n66102 );
and ( n66104 , n66099 , n66102 );
or ( n66105 , n66101 , n66103 , n66104 );
and ( n66106 , n59908 , n63766 );
not ( n66107 , n66106 );
and ( n66108 , n61008 , n62868 );
not ( n66109 , n66108 );
and ( n66110 , n66107 , n66109 );
and ( n66111 , n61505 , n62151 );
not ( n66112 , n66111 );
and ( n66113 , n66109 , n66112 );
and ( n66114 , n66107 , n66112 );
or ( n66115 , n66110 , n66113 , n66114 );
and ( n66116 , n65606 , n58542 );
not ( n66117 , n66116 );
and ( n66118 , n58915 , n65210 );
not ( n66119 , n66118 );
and ( n66120 , n66117 , n66119 );
and ( n66121 , n63492 , n60372 );
not ( n66122 , n66121 );
and ( n66123 , n66119 , n66122 );
and ( n66124 , n66117 , n66122 );
or ( n66125 , n66120 , n66123 , n66124 );
and ( n66126 , n66115 , n66125 );
and ( n66127 , n64548 , n59207 );
not ( n66128 , n66127 );
and ( n66129 , n63024 , n60711 );
not ( n66130 , n66129 );
or ( n66131 , n66128 , n66130 );
and ( n66132 , n66125 , n66131 );
and ( n66133 , n66115 , n66131 );
or ( n66134 , n66126 , n66132 , n66133 );
and ( n66135 , n66105 , n66134 );
and ( n66136 , n47647 , n57187 );
and ( n66137 , n47474 , n57184 );
nor ( n66138 , n66136 , n66137 );
xnor ( n66139 , n66138 , n56175 );
and ( n66140 , n48272 , n55851 );
and ( n66141 , n48108 , n55849 );
nor ( n66142 , n66140 , n66141 );
xnor ( n66143 , n66142 , n55506 );
and ( n66144 , n66139 , n66143 );
and ( n66145 , n48988 , n54535 );
and ( n66146 , n48709 , n54533 );
nor ( n66147 , n66145 , n66146 );
xnor ( n66148 , n66147 , n54237 );
and ( n66149 , n66143 , n66148 );
and ( n66150 , n66139 , n66148 );
or ( n66151 , n66144 , n66149 , n66150 );
and ( n66152 , n49374 , n53928 );
and ( n66153 , n49115 , n53926 );
nor ( n66154 , n66152 , n66153 );
xnor ( n66155 , n66154 , n53652 );
and ( n66156 , n49781 , n53357 );
and ( n66157 , n49570 , n53355 );
nor ( n66158 , n66156 , n66157 );
xnor ( n66159 , n66158 , n53060 );
and ( n66160 , n66155 , n66159 );
and ( n66161 , n50195 , n52799 );
and ( n66162 , n49976 , n52797 );
nor ( n66163 , n66161 , n66162 );
xnor ( n66164 , n66163 , n52538 );
and ( n66165 , n66159 , n66164 );
and ( n66166 , n66155 , n66164 );
or ( n66167 , n66160 , n66165 , n66166 );
and ( n66168 , n66151 , n66167 );
and ( n66169 , n50625 , n52269 );
and ( n66170 , n50404 , n52267 );
nor ( n66171 , n66169 , n66170 );
xnor ( n66172 , n66171 , n52008 );
and ( n66173 , n51077 , n51750 );
and ( n66174 , n50726 , n51748 );
nor ( n66175 , n66173 , n66174 );
xnor ( n66176 , n66175 , n51520 );
and ( n66177 , n66172 , n66176 );
and ( n66178 , n51510 , n51221 );
and ( n66179 , n51298 , n51219 );
nor ( n66180 , n66178 , n66179 );
xnor ( n66181 , n66180 , n51000 );
and ( n66182 , n66176 , n66181 );
and ( n66183 , n66172 , n66181 );
or ( n66184 , n66177 , n66182 , n66183 );
and ( n66185 , n66167 , n66184 );
and ( n66186 , n66151 , n66184 );
or ( n66187 , n66168 , n66185 , n66186 );
and ( n66188 , n66134 , n66187 );
and ( n66189 , n66105 , n66187 );
or ( n66190 , n66135 , n66188 , n66189 );
and ( n66191 , n66096 , n66190 );
and ( n66192 , n66049 , n66190 );
or ( n66193 , n66097 , n66191 , n66192 );
and ( n66194 , n66039 , n66193 );
and ( n66195 , n53639 , n49513 );
and ( n66196 , n53328 , n49511 );
nor ( n66197 , n66195 , n66196 );
xnor ( n66198 , n66197 , n49310 );
and ( n66199 , n54227 , n49121 );
and ( n66200 , n53922 , n49119 );
nor ( n66201 , n66199 , n66200 );
xnor ( n66202 , n66201 , n48932 );
and ( n66203 , n66198 , n66202 );
and ( n66204 , n54942 , n48740 );
and ( n66205 , n54604 , n48738 );
nor ( n66206 , n66204 , n66205 );
xnor ( n66207 , n66206 , n48571 );
and ( n66208 , n66202 , n66207 );
and ( n66209 , n66198 , n66207 );
or ( n66210 , n66203 , n66208 , n66209 );
and ( n66211 , n55497 , n48394 );
and ( n66212 , n55143 , n48392 );
nor ( n66213 , n66211 , n66212 );
xnor ( n66214 , n66213 , n48220 );
and ( n66215 , n56255 , n48042 );
and ( n66216 , n55756 , n48040 );
nor ( n66217 , n66215 , n66216 );
xnor ( n66218 , n66217 , n47921 );
and ( n66219 , n66214 , n66218 );
and ( n66220 , n56915 , n47734 );
and ( n66221 , n56388 , n47732 );
nor ( n66222 , n66220 , n66221 );
xnor ( n66223 , n66222 , n47606 );
and ( n66224 , n66218 , n66223 );
and ( n66225 , n66214 , n66223 );
or ( n66226 , n66219 , n66224 , n66225 );
and ( n66227 , n66210 , n66226 );
xor ( n66228 , n42762 , n45546 );
buf ( n66229 , n66228 );
buf ( n66230 , n66229 );
buf ( n66231 , n66230 );
and ( n66232 , n65733 , n66231 );
and ( n66233 , n63987 , n59920 );
not ( n66234 , n66233 );
and ( n66235 , n66231 , n66234 );
and ( n66236 , n65733 , n66234 );
or ( n66237 , n66232 , n66235 , n66236 );
and ( n66238 , n66226 , n66237 );
and ( n66239 , n66210 , n66237 );
or ( n66240 , n66227 , n66238 , n66239 );
xor ( n66241 , n65760 , n65764 );
xor ( n66242 , n66241 , n65769 );
xor ( n66243 , n65777 , n65781 );
xor ( n66244 , n66243 , n65786 );
and ( n66245 , n66242 , n66244 );
xor ( n66246 , n65797 , n65801 );
xor ( n66247 , n66246 , n65806 );
and ( n66248 , n66244 , n66247 );
and ( n66249 , n66242 , n66247 );
or ( n66250 , n66245 , n66248 , n66249 );
and ( n66251 , n66240 , n66250 );
buf ( n66252 , n65693 );
xor ( n66253 , n66252 , n65694 );
and ( n66254 , n66250 , n66253 );
and ( n66255 , n66240 , n66253 );
or ( n66256 , n66251 , n66254 , n66255 );
xor ( n66257 , n65698 , n65699 );
xor ( n66258 , n66257 , n65701 );
xor ( n66259 , n65723 , n65738 );
xor ( n66260 , n66259 , n65748 );
and ( n66261 , n66258 , n66260 );
xor ( n66262 , n65756 , n65772 );
xor ( n66263 , n66262 , n65789 );
and ( n66264 , n66260 , n66263 );
and ( n66265 , n66258 , n66263 );
or ( n66266 , n66261 , n66264 , n66265 );
and ( n66267 , n66256 , n66266 );
xor ( n66268 , n65643 , n65645 );
xor ( n66269 , n66268 , n65657 );
and ( n66270 , n66266 , n66269 );
and ( n66271 , n66256 , n66269 );
or ( n66272 , n66267 , n66270 , n66271 );
and ( n66273 , n66193 , n66272 );
and ( n66274 , n66039 , n66272 );
or ( n66275 , n66194 , n66273 , n66274 );
xor ( n66276 , n65692 , n65696 );
xor ( n66277 , n66276 , n65704 );
xor ( n66278 , n65751 , n65792 );
xor ( n66279 , n66278 , n65843 );
and ( n66280 , n66277 , n66279 );
xor ( n66281 , n65857 , n65859 );
xor ( n66282 , n66281 , n65862 );
and ( n66283 , n66279 , n66282 );
and ( n66284 , n66277 , n66282 );
or ( n66285 , n66280 , n66283 , n66284 );
xor ( n66286 , n65566 , n65568 );
xor ( n66287 , n66286 , n65600 );
and ( n66288 , n66285 , n66287 );
xor ( n66289 , n65622 , n65640 );
xor ( n66290 , n66289 , n65660 );
and ( n66291 , n66287 , n66290 );
and ( n66292 , n66285 , n66290 );
or ( n66293 , n66288 , n66291 , n66292 );
and ( n66294 , n66275 , n66293 );
xor ( n66295 , n65707 , n65846 );
xor ( n66296 , n66295 , n65865 );
xor ( n66297 , n65878 , n65880 );
xor ( n66298 , n66297 , n65883 );
and ( n66299 , n66296 , n66298 );
xor ( n66300 , n65889 , n65891 );
xor ( n66301 , n66300 , n65894 );
and ( n66302 , n66298 , n66301 );
and ( n66303 , n66296 , n66301 );
or ( n66304 , n66299 , n66302 , n66303 );
and ( n66305 , n66293 , n66304 );
and ( n66306 , n66275 , n66304 );
or ( n66307 , n66294 , n66305 , n66306 );
and ( n66308 , n66001 , n66307 );
xor ( n66309 , n65564 , n65603 );
xor ( n66310 , n66309 , n65663 );
xor ( n66311 , n65868 , n65886 );
xor ( n66312 , n66311 , n65897 );
and ( n66313 , n66310 , n66312 );
xor ( n66314 , n65903 , n65905 );
xor ( n66315 , n66314 , n65908 );
and ( n66316 , n66312 , n66315 );
and ( n66317 , n66310 , n66315 );
or ( n66318 , n66313 , n66316 , n66317 );
and ( n66319 , n66307 , n66318 );
and ( n66320 , n66001 , n66318 );
or ( n66321 , n66308 , n66319 , n66320 );
xor ( n66322 , n65556 , n65558 );
xor ( n66323 , n66322 , n65560 );
xor ( n66324 , n65666 , n65900 );
xor ( n66325 , n66324 , n65911 );
and ( n66326 , n66323 , n66325 );
xor ( n66327 , n65917 , n65919 );
xor ( n66328 , n66327 , n65922 );
and ( n66329 , n66325 , n66328 );
and ( n66330 , n66323 , n66328 );
or ( n66331 , n66326 , n66329 , n66330 );
and ( n66332 , n66321 , n66331 );
xor ( n66333 , n65563 , n65914 );
xor ( n66334 , n66333 , n65925 );
and ( n66335 , n66331 , n66334 );
and ( n66336 , n66321 , n66334 );
or ( n66337 , n66332 , n66335 , n66336 );
and ( n66338 , n65954 , n66337 );
and ( n66339 , n65952 , n66337 );
or ( n66340 , n65955 , n66338 , n66339 );
and ( n66341 , n65950 , n66340 );
xor ( n66342 , n65549 , n65551 );
xor ( n66343 , n66342 , n65942 );
and ( n66344 , n66340 , n66343 );
and ( n66345 , n65950 , n66343 );
or ( n66346 , n66341 , n66344 , n66345 );
and ( n66347 , n65947 , n66346 );
and ( n66348 , n65945 , n66346 );
or ( n66349 , n65948 , n66347 , n66348 );
and ( n66350 , n65546 , n66349 );
and ( n66351 , n65544 , n66349 );
or ( n66352 , n65547 , n66350 , n66351 );
and ( n66353 , n65139 , n66352 );
and ( n66354 , n65137 , n66352 );
or ( n66355 , n65140 , n66353 , n66354 );
and ( n66356 , n64732 , n66355 );
and ( n66357 , n64730 , n66355 );
or ( n66358 , n64733 , n66356 , n66357 );
or ( n66359 , n64331 , n66358 );
or ( n66360 , n64329 , n66359 );
and ( n66361 , n64326 , n66360 );
and ( n66362 , n63627 , n66360 );
or ( n66363 , n64327 , n66361 , n66362 );
and ( n66364 , n63624 , n66363 );
and ( n66365 , n62840 , n66363 );
or ( n66366 , n63625 , n66364 , n66365 );
and ( n66367 , n62838 , n66366 );
xor ( n66368 , n62838 , n66366 );
xor ( n66369 , n62840 , n63624 );
xor ( n66370 , n66369 , n66363 );
not ( n66371 , n66370 );
xor ( n66372 , n63627 , n64326 );
xor ( n66373 , n66372 , n66360 );
not ( n66374 , n66373 );
xnor ( n66375 , n64329 , n66359 );
xnor ( n66376 , n64331 , n66358 );
xor ( n66377 , n64730 , n64732 );
xor ( n66378 , n66377 , n66355 );
xor ( n66379 , n65137 , n65139 );
xor ( n66380 , n66379 , n66352 );
xor ( n66381 , n65544 , n65546 );
xor ( n66382 , n66381 , n66349 );
not ( n66383 , n66382 );
xor ( n66384 , n65945 , n65947 );
xor ( n66385 , n66384 , n66346 );
xor ( n66386 , n65554 , n65928 );
xor ( n66387 , n66386 , n65939 );
xor ( n66388 , n65931 , n65933 );
xor ( n66389 , n66388 , n65936 );
xor ( n66390 , n65870 , n65872 );
xor ( n66391 , n66390 , n65875 );
xnor ( n66392 , n65981 , n65983 );
and ( n66393 , n66391 , n66392 );
and ( n66394 , n64221 , n59207 );
not ( n66395 , n66394 );
and ( n66396 , n62593 , n60711 );
not ( n66397 , n66396 );
and ( n66398 , n66395 , n66397 );
xor ( n66399 , n66007 , n66009 );
xor ( n66400 , n66399 , n66012 );
and ( n66401 , n66397 , n66400 );
and ( n66402 , n66395 , n66400 );
or ( n66403 , n66398 , n66401 , n66402 );
and ( n66404 , n65678 , n58444 );
not ( n66405 , n66404 );
and ( n66406 , n64221 , n59611 );
not ( n66407 , n66406 );
and ( n66408 , n66405 , n66407 );
buf ( n66409 , n61918 );
not ( n66410 , n66409 );
and ( n66411 , n66407 , n66410 );
and ( n66412 , n66405 , n66410 );
or ( n66413 , n66408 , n66411 , n66412 );
buf ( n66414 , n20252 );
buf ( n66415 , n66414 );
and ( n66416 , n66415 , n58294 );
not ( n66417 , n66416 );
and ( n66418 , n62593 , n61015 );
not ( n66419 , n66418 );
and ( n66420 , n66417 , n66419 );
and ( n66421 , n62377 , n61481 );
not ( n66422 , n66421 );
and ( n66423 , n66419 , n66422 );
and ( n66424 , n66417 , n66422 );
or ( n66425 , n66420 , n66423 , n66424 );
and ( n66426 , n66413 , n66425 );
xor ( n66427 , n66016 , n66018 );
xor ( n66428 , n66427 , n66021 );
and ( n66429 , n66425 , n66428 );
and ( n66430 , n66413 , n66428 );
or ( n66431 , n66426 , n66429 , n66430 );
and ( n66432 , n66403 , n66431 );
xor ( n66433 , n65624 , n65626 );
xor ( n66434 , n66433 , n65629 );
and ( n66435 , n66431 , n66434 );
and ( n66436 , n66403 , n66434 );
or ( n66437 , n66432 , n66435 , n66436 );
and ( n66438 , n66392 , n66437 );
and ( n66439 , n66391 , n66437 );
or ( n66440 , n66393 , n66438 , n66439 );
xor ( n66441 , n65809 , n65825 );
xor ( n66442 , n66441 , n65840 );
xor ( n66443 , n65849 , n65851 );
xor ( n66444 , n66443 , n65854 );
and ( n66445 , n66442 , n66444 );
xor ( n66446 , n66015 , n66024 );
xor ( n66447 , n66446 , n66027 );
and ( n66448 , n66444 , n66447 );
and ( n66449 , n66442 , n66447 );
or ( n66450 , n66445 , n66448 , n66449 );
xor ( n66451 , n65973 , n65975 );
xor ( n66452 , n66451 , n65978 );
xnor ( n66453 , n66033 , n66035 );
and ( n66454 , n66452 , n66453 );
and ( n66455 , n58292 , n66005 );
not ( n66456 , n66455 );
and ( n66457 , n58628 , n65586 );
not ( n66458 , n66457 );
and ( n66459 , n66456 , n66458 );
and ( n66460 , n60376 , n63679 );
not ( n66461 , n66460 );
and ( n66462 , n66458 , n66461 );
and ( n66463 , n66456 , n66461 );
or ( n66464 , n66459 , n66462 , n66463 );
and ( n66465 , n65606 , n58911 );
not ( n66466 , n66465 );
buf ( n66467 , n66466 );
buf ( n66468 , n20252 );
buf ( n66469 , n66468 );
and ( n66470 , n57948 , n66469 );
not ( n66471 , n66470 );
and ( n66472 , n66467 , n66471 );
and ( n66473 , n59615 , n64412 );
not ( n66474 , n66473 );
and ( n66475 , n66471 , n66474 );
and ( n66476 , n66467 , n66474 );
or ( n66477 , n66472 , n66475 , n66476 );
and ( n66478 , n66464 , n66477 );
and ( n66479 , n60821 , n62868 );
not ( n66480 , n66479 );
and ( n66481 , n66477 , n66480 );
and ( n66482 , n66464 , n66480 );
or ( n66483 , n66478 , n66481 , n66482 );
and ( n66484 , n66453 , n66483 );
and ( n66485 , n66452 , n66483 );
or ( n66486 , n66454 , n66484 , n66485 );
and ( n66487 , n66450 , n66486 );
xor ( n66488 , n65813 , n65817 );
xor ( n66489 , n66488 , n65822 );
xor ( n66490 , n65830 , n65834 );
xor ( n66491 , n66490 , n65837 );
and ( n66492 , n66489 , n66491 );
xor ( n66493 , n65965 , n65967 );
xor ( n66494 , n66493 , n65970 );
and ( n66495 , n66491 , n66494 );
and ( n66496 , n66489 , n66494 );
or ( n66497 , n66492 , n66495 , n66496 );
xor ( n66498 , n66057 , n66059 );
xor ( n66499 , n66498 , n66062 );
xor ( n66500 , n66395 , n66397 );
xor ( n66501 , n66500 , n66400 );
and ( n66502 , n66499 , n66501 );
xnor ( n66503 , n66081 , n66085 );
and ( n66504 , n66501 , n66503 );
and ( n66505 , n66499 , n66503 );
or ( n66506 , n66502 , n66504 , n66505 );
and ( n66507 , n66497 , n66506 );
and ( n66508 , n47778 , n57187 );
and ( n66509 , n47647 , n57184 );
nor ( n66510 , n66508 , n66509 );
xnor ( n66511 , n66510 , n56175 );
and ( n66512 , n48709 , n55159 );
and ( n66513 , n48632 , n55157 );
nor ( n66514 , n66512 , n66513 );
xnor ( n66515 , n66514 , n54864 );
and ( n66516 , n66511 , n66515 );
and ( n66517 , n52332 , n50783 );
and ( n66518 , n52082 , n50781 );
nor ( n66519 , n66517 , n66518 );
xnor ( n66520 , n66519 , n50557 );
and ( n66521 , n66515 , n66520 );
and ( n66522 , n66511 , n66520 );
or ( n66523 , n66516 , n66521 , n66522 );
and ( n66524 , n52612 , n50338 );
and ( n66525 , n52332 , n50336 );
nor ( n66526 , n66524 , n66525 );
xnor ( n66527 , n66526 , n50111 );
and ( n66528 , n66523 , n66527 );
and ( n66529 , n53041 , n49896 );
and ( n66530 , n52790 , n49894 );
nor ( n66531 , n66529 , n66530 );
xnor ( n66532 , n66531 , n49711 );
and ( n66533 , n66527 , n66532 );
and ( n66534 , n66523 , n66532 );
or ( n66535 , n66528 , n66533 , n66534 );
and ( n66536 , n66415 , n58444 );
and ( n66537 , n65678 , n58542 );
not ( n66538 , n66537 );
and ( n66539 , n66536 , n66538 );
and ( n66540 , n58292 , n66469 );
and ( n66541 , n58628 , n66005 );
not ( n66542 , n66541 );
and ( n66543 , n66540 , n66542 );
and ( n66544 , n66539 , n66543 );
and ( n66545 , n66535 , n66544 );
not ( n66546 , n66536 );
buf ( n66547 , n66546 );
not ( n66548 , n66540 );
buf ( n66549 , n66548 );
and ( n66550 , n66547 , n66549 );
and ( n66551 , n66544 , n66550 );
and ( n66552 , n66535 , n66550 );
or ( n66553 , n66545 , n66551 , n66552 );
and ( n66554 , n66506 , n66553 );
and ( n66555 , n66497 , n66553 );
or ( n66556 , n66507 , n66554 , n66555 );
and ( n66557 , n66486 , n66556 );
and ( n66558 , n66450 , n66556 );
or ( n66559 , n66487 , n66557 , n66558 );
and ( n66560 , n66440 , n66559 );
xor ( n66561 , n66069 , n66073 );
xor ( n66562 , n66561 , n66078 );
xor ( n66563 , n66405 , n66407 );
xor ( n66564 , n66563 , n66410 );
and ( n66565 , n66562 , n66564 );
buf ( n66566 , n66565 );
xor ( n66567 , n66117 , n66119 );
xor ( n66568 , n66567 , n66122 );
xnor ( n66569 , n66128 , n66130 );
and ( n66570 , n66568 , n66569 );
and ( n66571 , n59615 , n64811 );
not ( n66572 , n66571 );
and ( n66573 , n61505 , n62868 );
not ( n66574 , n66573 );
and ( n66575 , n66572 , n66574 );
and ( n66576 , n61918 , n62151 );
not ( n66577 , n66576 );
and ( n66578 , n66574 , n66577 );
and ( n66579 , n66572 , n66577 );
or ( n66580 , n66575 , n66578 , n66579 );
and ( n66581 , n66569 , n66580 );
and ( n66582 , n66568 , n66580 );
or ( n66583 , n66570 , n66581 , n66582 );
and ( n66584 , n66566 , n66583 );
and ( n66585 , n64548 , n59611 );
not ( n66586 , n66585 );
and ( n66587 , n64221 , n59920 );
not ( n66588 , n66587 );
and ( n66589 , n66586 , n66588 );
and ( n66590 , n62593 , n61481 );
not ( n66591 , n66590 );
and ( n66592 , n66588 , n66591 );
and ( n66593 , n66586 , n66591 );
or ( n66594 , n66589 , n66592 , n66593 );
and ( n66595 , n58915 , n65586 );
and ( n66596 , n60376 , n63766 );
not ( n66597 , n66596 );
and ( n66598 , n66595 , n66597 );
and ( n66599 , n61008 , n62998 );
not ( n66600 , n66599 );
and ( n66601 , n66597 , n66600 );
and ( n66602 , n66595 , n66600 );
or ( n66603 , n66598 , n66601 , n66602 );
and ( n66604 , n66594 , n66603 );
not ( n66605 , n66595 );
buf ( n66606 , n66605 );
and ( n66607 , n66603 , n66606 );
and ( n66608 , n66594 , n66606 );
or ( n66609 , n66604 , n66607 , n66608 );
and ( n66610 , n66583 , n66609 );
and ( n66611 , n66566 , n66609 );
or ( n66612 , n66584 , n66610 , n66611 );
and ( n66613 , n49115 , n54535 );
and ( n66614 , n48988 , n54533 );
nor ( n66615 , n66613 , n66614 );
xnor ( n66616 , n66615 , n54237 );
and ( n66617 , n51734 , n51221 );
and ( n66618 , n51510 , n51219 );
nor ( n66619 , n66617 , n66618 );
xnor ( n66620 , n66619 , n51000 );
or ( n66621 , n66616 , n66620 );
and ( n66622 , n48108 , n56503 );
and ( n66623 , n47962 , n56501 );
nor ( n66624 , n66622 , n66623 );
xnor ( n66625 , n66624 , n56178 );
and ( n66626 , n48384 , n55851 );
and ( n66627 , n48272 , n55849 );
nor ( n66628 , n66626 , n66627 );
xnor ( n66629 , n66628 , n55506 );
and ( n66630 , n66625 , n66629 );
and ( n66631 , n49570 , n53928 );
and ( n66632 , n49374 , n53926 );
nor ( n66633 , n66631 , n66632 );
xnor ( n66634 , n66633 , n53652 );
and ( n66635 , n66629 , n66634 );
and ( n66636 , n66625 , n66634 );
or ( n66637 , n66630 , n66635 , n66636 );
and ( n66638 , n66621 , n66637 );
and ( n66639 , n49976 , n53357 );
and ( n66640 , n49781 , n53355 );
nor ( n66641 , n66639 , n66640 );
xnor ( n66642 , n66641 , n53060 );
and ( n66643 , n50404 , n52799 );
and ( n66644 , n50195 , n52797 );
nor ( n66645 , n66643 , n66644 );
xnor ( n66646 , n66645 , n52538 );
and ( n66647 , n66642 , n66646 );
and ( n66648 , n50726 , n52269 );
and ( n66649 , n50625 , n52267 );
nor ( n66650 , n66648 , n66649 );
xnor ( n66651 , n66650 , n52008 );
and ( n66652 , n66646 , n66651 );
and ( n66653 , n66642 , n66651 );
or ( n66654 , n66647 , n66652 , n66653 );
and ( n66655 , n66637 , n66654 );
and ( n66656 , n66621 , n66654 );
or ( n66657 , n66638 , n66655 , n66656 );
and ( n66658 , n51298 , n51750 );
and ( n66659 , n51077 , n51748 );
nor ( n66660 , n66658 , n66659 );
xnor ( n66661 , n66660 , n51520 );
and ( n66662 , n52790 , n50338 );
and ( n66663 , n52612 , n50336 );
nor ( n66664 , n66662 , n66663 );
xnor ( n66665 , n66664 , n50111 );
and ( n66666 , n66661 , n66665 );
and ( n66667 , n53328 , n49896 );
and ( n66668 , n53041 , n49894 );
nor ( n66669 , n66667 , n66668 );
xnor ( n66670 , n66669 , n49711 );
and ( n66671 , n66665 , n66670 );
and ( n66672 , n66661 , n66670 );
or ( n66673 , n66666 , n66671 , n66672 );
and ( n66674 , n53922 , n49513 );
and ( n66675 , n53639 , n49511 );
nor ( n66676 , n66674 , n66675 );
xnor ( n66677 , n66676 , n49310 );
and ( n66678 , n54604 , n49121 );
and ( n66679 , n54227 , n49119 );
nor ( n66680 , n66678 , n66679 );
xnor ( n66681 , n66680 , n48932 );
and ( n66682 , n66677 , n66681 );
and ( n66683 , n55143 , n48740 );
and ( n66684 , n54942 , n48738 );
nor ( n66685 , n66683 , n66684 );
xnor ( n66686 , n66685 , n48571 );
and ( n66687 , n66681 , n66686 );
and ( n66688 , n66677 , n66686 );
or ( n66689 , n66682 , n66687 , n66688 );
and ( n66690 , n66673 , n66689 );
and ( n66691 , n55756 , n48394 );
and ( n66692 , n55497 , n48392 );
nor ( n66693 , n66691 , n66692 );
xnor ( n66694 , n66693 , n48220 );
and ( n66695 , n56388 , n48042 );
and ( n66696 , n56255 , n48040 );
nor ( n66697 , n66695 , n66696 );
xnor ( n66698 , n66697 , n47921 );
and ( n66699 , n66694 , n66698 );
and ( n66700 , n57063 , n47734 );
and ( n66701 , n56915 , n47732 );
nor ( n66702 , n66700 , n66701 );
xnor ( n66703 , n66702 , n47606 );
and ( n66704 , n66698 , n66703 );
and ( n66705 , n66694 , n66703 );
or ( n66706 , n66699 , n66704 , n66705 );
and ( n66707 , n66689 , n66706 );
and ( n66708 , n66673 , n66706 );
or ( n66709 , n66690 , n66707 , n66708 );
and ( n66710 , n66657 , n66709 );
and ( n66711 , n57063 , n47732 );
not ( n66712 , n66711 );
and ( n66713 , n66712 , n47606 );
xor ( n66714 , n42763 , n45545 );
buf ( n66715 , n66714 );
buf ( n66716 , n66715 );
buf ( n66717 , n66716 );
and ( n66718 , n66713 , n66717 );
buf ( n66719 , n20257 );
buf ( n66720 , n66719 );
and ( n66721 , n66720 , n58294 );
not ( n66722 , n66721 );
and ( n66723 , n66717 , n66722 );
and ( n66724 , n66713 , n66722 );
or ( n66725 , n66718 , n66723 , n66724 );
xor ( n66726 , n66139 , n66143 );
xor ( n66727 , n66726 , n66148 );
and ( n66728 , n66725 , n66727 );
xor ( n66729 , n66155 , n66159 );
xor ( n66730 , n66729 , n66164 );
and ( n66731 , n66727 , n66730 );
and ( n66732 , n66725 , n66730 );
or ( n66733 , n66728 , n66731 , n66732 );
and ( n66734 , n66709 , n66733 );
and ( n66735 , n66657 , n66733 );
or ( n66736 , n66710 , n66734 , n66735 );
and ( n66737 , n66612 , n66736 );
xor ( n66738 , n66172 , n66176 );
xor ( n66739 , n66738 , n66181 );
xor ( n66740 , n66198 , n66202 );
xor ( n66741 , n66740 , n66207 );
and ( n66742 , n66739 , n66741 );
xor ( n66743 , n66214 , n66218 );
xor ( n66744 , n66743 , n66223 );
and ( n66745 , n66741 , n66744 );
and ( n66746 , n66739 , n66744 );
or ( n66747 , n66742 , n66745 , n66746 );
buf ( n66748 , n66089 );
xor ( n66749 , n66748 , n66091 );
and ( n66750 , n66747 , n66749 );
xor ( n66751 , n66099 , n66100 );
xor ( n66752 , n66751 , n66102 );
and ( n66753 , n66749 , n66752 );
and ( n66754 , n66747 , n66752 );
or ( n66755 , n66750 , n66753 , n66754 );
and ( n66756 , n66736 , n66755 );
and ( n66757 , n66612 , n66755 );
or ( n66758 , n66737 , n66756 , n66757 );
xor ( n66759 , n66115 , n66125 );
xor ( n66760 , n66759 , n66131 );
xor ( n66761 , n66151 , n66167 );
xor ( n66762 , n66761 , n66184 );
and ( n66763 , n66760 , n66762 );
xor ( n66764 , n66210 , n66226 );
xor ( n66765 , n66764 , n66237 );
and ( n66766 , n66762 , n66765 );
and ( n66767 , n66760 , n66765 );
or ( n66768 , n66763 , n66766 , n66767 );
xor ( n66769 , n66041 , n66043 );
xor ( n66770 , n66769 , n66046 );
and ( n66771 , n66768 , n66770 );
xor ( n66772 , n66065 , n66086 );
xor ( n66773 , n66772 , n66093 );
and ( n66774 , n66770 , n66773 );
and ( n66775 , n66768 , n66773 );
or ( n66776 , n66771 , n66774 , n66775 );
and ( n66777 , n66758 , n66776 );
xor ( n66778 , n66105 , n66134 );
xor ( n66779 , n66778 , n66187 );
xor ( n66780 , n66240 , n66250 );
xor ( n66781 , n66780 , n66253 );
and ( n66782 , n66779 , n66781 );
xor ( n66783 , n66258 , n66260 );
xor ( n66784 , n66783 , n66263 );
and ( n66785 , n66781 , n66784 );
and ( n66786 , n66779 , n66784 );
or ( n66787 , n66782 , n66785 , n66786 );
and ( n66788 , n66776 , n66787 );
and ( n66789 , n66758 , n66787 );
or ( n66790 , n66777 , n66788 , n66789 );
and ( n66791 , n66559 , n66790 );
and ( n66792 , n66440 , n66790 );
or ( n66793 , n66560 , n66791 , n66792 );
xor ( n66794 , n65987 , n65989 );
xor ( n66795 , n66794 , n65992 );
xor ( n66796 , n66003 , n66030 );
xor ( n66797 , n66796 , n66036 );
and ( n66798 , n66795 , n66797 );
xor ( n66799 , n66049 , n66096 );
xor ( n66800 , n66799 , n66190 );
and ( n66801 , n66797 , n66800 );
and ( n66802 , n66795 , n66800 );
or ( n66803 , n66798 , n66801 , n66802 );
xor ( n66804 , n65962 , n65984 );
xor ( n66805 , n66804 , n65995 );
and ( n66806 , n66803 , n66805 );
xor ( n66807 , n66039 , n66193 );
xor ( n66808 , n66807 , n66272 );
and ( n66809 , n66805 , n66808 );
and ( n66810 , n66803 , n66808 );
or ( n66811 , n66806 , n66809 , n66810 );
and ( n66812 , n66793 , n66811 );
xor ( n66813 , n65957 , n65959 );
xor ( n66814 , n66813 , n65998 );
and ( n66815 , n66811 , n66814 );
and ( n66816 , n66793 , n66814 );
or ( n66817 , n66812 , n66815 , n66816 );
xor ( n66818 , n66001 , n66307 );
xor ( n66819 , n66818 , n66318 );
and ( n66820 , n66817 , n66819 );
xor ( n66821 , n66323 , n66325 );
xor ( n66822 , n66821 , n66328 );
and ( n66823 , n66819 , n66822 );
and ( n66824 , n66817 , n66822 );
or ( n66825 , n66820 , n66823 , n66824 );
and ( n66826 , n66389 , n66825 );
xor ( n66827 , n66321 , n66331 );
xor ( n66828 , n66827 , n66334 );
and ( n66829 , n66825 , n66828 );
and ( n66830 , n66389 , n66828 );
or ( n66831 , n66826 , n66829 , n66830 );
and ( n66832 , n66387 , n66831 );
xor ( n66833 , n65952 , n65954 );
xor ( n66834 , n66833 , n66337 );
and ( n66835 , n66831 , n66834 );
and ( n66836 , n66387 , n66834 );
or ( n66837 , n66832 , n66835 , n66836 );
xor ( n66838 , n65950 , n66340 );
xor ( n66839 , n66838 , n66343 );
and ( n66840 , n66837 , n66839 );
xor ( n66841 , n66387 , n66831 );
xor ( n66842 , n66841 , n66834 );
xor ( n66843 , n66389 , n66825 );
xor ( n66844 , n66843 , n66828 );
xor ( n66845 , n66275 , n66293 );
xor ( n66846 , n66845 , n66304 );
xor ( n66847 , n66310 , n66312 );
xor ( n66848 , n66847 , n66315 );
and ( n66849 , n66846 , n66848 );
xor ( n66850 , n66285 , n66287 );
xor ( n66851 , n66850 , n66290 );
xor ( n66852 , n66296 , n66298 );
xor ( n66853 , n66852 , n66301 );
and ( n66854 , n66851 , n66853 );
xor ( n66855 , n66256 , n66266 );
xor ( n66856 , n66855 , n66269 );
xor ( n66857 , n66277 , n66279 );
xor ( n66858 , n66857 , n66282 );
and ( n66859 , n66856 , n66858 );
xor ( n66860 , n66403 , n66431 );
xor ( n66861 , n66860 , n66434 );
xor ( n66862 , n66242 , n66244 );
xor ( n66863 , n66862 , n66247 );
xor ( n66864 , n66464 , n66477 );
xor ( n66865 , n66864 , n66480 );
and ( n66866 , n66863 , n66865 );
xor ( n66867 , n66413 , n66425 );
xor ( n66868 , n66867 , n66428 );
and ( n66869 , n66865 , n66868 );
and ( n66870 , n66863 , n66868 );
or ( n66871 , n66866 , n66869 , n66870 );
and ( n66872 , n66861 , n66871 );
and ( n66873 , n63987 , n60372 );
not ( n66874 , n66873 );
and ( n66875 , n66465 , n66874 );
and ( n66876 , n63024 , n61015 );
not ( n66877 , n66876 );
and ( n66878 , n66874 , n66877 );
and ( n66879 , n66465 , n66877 );
or ( n66880 , n66875 , n66878 , n66879 );
xor ( n66881 , n66456 , n66458 );
xor ( n66882 , n66881 , n66461 );
and ( n66883 , n66880 , n66882 );
xor ( n66884 , n66467 , n66471 );
xor ( n66885 , n66884 , n66474 );
and ( n66886 , n66882 , n66885 );
and ( n66887 , n66880 , n66885 );
or ( n66888 , n66883 , n66886 , n66887 );
and ( n66889 , n58628 , n66469 );
not ( n66890 , n66889 );
and ( n66891 , n60376 , n64412 );
not ( n66892 , n66891 );
and ( n66893 , n66890 , n66892 );
and ( n66894 , n61918 , n62868 );
not ( n66895 , n66894 );
and ( n66896 , n66892 , n66895 );
and ( n66897 , n66890 , n66895 );
or ( n66898 , n66893 , n66896 , n66897 );
and ( n66899 , n59365 , n65210 );
not ( n66900 , n66899 );
and ( n66901 , n66898 , n66900 );
and ( n66902 , n60821 , n63679 );
not ( n66903 , n66902 );
and ( n66904 , n66900 , n66903 );
and ( n66905 , n66898 , n66903 );
or ( n66906 , n66901 , n66904 , n66905 );
xor ( n66907 , n66107 , n66109 );
xor ( n66908 , n66907 , n66112 );
and ( n66909 , n66906 , n66908 );
xor ( n66910 , n65963 , n66051 );
xor ( n66911 , n66910 , n66054 );
and ( n66912 , n66908 , n66911 );
and ( n66913 , n66906 , n66911 );
or ( n66914 , n66909 , n66912 , n66913 );
and ( n66915 , n66888 , n66914 );
buf ( n66916 , n20257 );
buf ( n66917 , n66916 );
and ( n66918 , n58292 , n66917 );
not ( n66919 , n66918 );
and ( n66920 , n58915 , n66005 );
not ( n66921 , n66920 );
and ( n66922 , n66919 , n66921 );
and ( n66923 , n62593 , n61914 );
not ( n66924 , n66923 );
and ( n66925 , n66921 , n66924 );
and ( n66926 , n66919 , n66924 );
or ( n66927 , n66922 , n66925 , n66926 );
and ( n66928 , n65177 , n59207 );
not ( n66929 , n66928 );
and ( n66930 , n66927 , n66929 );
and ( n66931 , n63492 , n60711 );
not ( n66932 , n66931 );
and ( n66933 , n66929 , n66932 );
and ( n66934 , n66927 , n66932 );
or ( n66935 , n66930 , n66933 , n66934 );
xor ( n66936 , n66417 , n66419 );
xor ( n66937 , n66936 , n66422 );
or ( n66938 , n66935 , n66937 );
and ( n66939 , n66914 , n66938 );
and ( n66940 , n66888 , n66938 );
or ( n66941 , n66915 , n66939 , n66940 );
and ( n66942 , n66871 , n66941 );
and ( n66943 , n66861 , n66941 );
or ( n66944 , n66872 , n66942 , n66943 );
and ( n66945 , n66858 , n66944 );
and ( n66946 , n66856 , n66944 );
or ( n66947 , n66859 , n66945 , n66946 );
and ( n66948 , n66853 , n66947 );
and ( n66949 , n66851 , n66947 );
or ( n66950 , n66854 , n66948 , n66949 );
and ( n66951 , n66848 , n66950 );
and ( n66952 , n66846 , n66950 );
or ( n66953 , n66849 , n66951 , n66952 );
xor ( n66954 , n66817 , n66819 );
xor ( n66955 , n66954 , n66822 );
and ( n66956 , n66953 , n66955 );
xor ( n66957 , n65733 , n66231 );
xor ( n66958 , n66957 , n66234 );
xor ( n66959 , n66523 , n66527 );
xor ( n66960 , n66959 , n66532 );
and ( n66961 , n66958 , n66960 );
xor ( n66962 , n66539 , n66543 );
and ( n66963 , n66960 , n66962 );
and ( n66964 , n66958 , n66962 );
or ( n66965 , n66961 , n66963 , n66964 );
xor ( n66966 , n66547 , n66549 );
and ( n66967 , n65678 , n58911 );
not ( n66968 , n66967 );
buf ( n66969 , n66968 );
and ( n66970 , n57948 , n66917 );
not ( n66971 , n66970 );
and ( n66972 , n66969 , n66971 );
and ( n66973 , n59908 , n64412 );
not ( n66974 , n66973 );
and ( n66975 , n66971 , n66974 );
and ( n66976 , n66969 , n66974 );
or ( n66977 , n66972 , n66975 , n66976 );
and ( n66978 , n66966 , n66977 );
buf ( n66979 , n20262 );
buf ( n66980 , n66979 );
and ( n66981 , n66980 , n58294 );
not ( n66982 , n66981 );
and ( n66983 , n64548 , n59920 );
not ( n66984 , n66983 );
and ( n66985 , n66982 , n66984 );
buf ( n66986 , n62377 );
not ( n66987 , n66986 );
and ( n66988 , n66984 , n66987 );
and ( n66989 , n66982 , n66987 );
or ( n66990 , n66985 , n66988 , n66989 );
xor ( n66991 , n66586 , n66588 );
xor ( n66992 , n66991 , n66591 );
or ( n66993 , n66990 , n66992 );
and ( n66994 , n66977 , n66993 );
and ( n66995 , n66966 , n66993 );
or ( n66996 , n66978 , n66994 , n66995 );
and ( n66997 , n66965 , n66996 );
xor ( n66998 , n66536 , n66538 );
xor ( n66999 , n66540 , n66542 );
and ( n67000 , n66998 , n66999 );
and ( n67001 , n62377 , n61914 );
not ( n67002 , n67001 );
xor ( n67003 , n66511 , n66515 );
xor ( n67004 , n67003 , n66520 );
and ( n67005 , n67002 , n67004 );
buf ( n67006 , n67005 );
and ( n67007 , n67000 , n67006 );
xor ( n67008 , n66465 , n66874 );
xor ( n67009 , n67008 , n66877 );
xnor ( n67010 , n66616 , n66620 );
and ( n67011 , n67009 , n67010 );
buf ( n67012 , n20262 );
buf ( n67013 , n67012 );
and ( n67014 , n57948 , n67013 );
not ( n67015 , n67014 );
and ( n67016 , n59908 , n64811 );
not ( n67017 , n67016 );
and ( n67018 , n67015 , n67017 );
and ( n67019 , n61008 , n63679 );
not ( n67020 , n67019 );
and ( n67021 , n67017 , n67020 );
and ( n67022 , n67015 , n67020 );
or ( n67023 , n67018 , n67021 , n67022 );
and ( n67024 , n67010 , n67023 );
and ( n67025 , n67009 , n67023 );
or ( n67026 , n67011 , n67024 , n67025 );
and ( n67027 , n67006 , n67026 );
and ( n67028 , n67000 , n67026 );
or ( n67029 , n67007 , n67027 , n67028 );
and ( n67030 , n66996 , n67029 );
and ( n67031 , n66965 , n67029 );
or ( n67032 , n66997 , n67030 , n67031 );
and ( n67033 , n65177 , n59611 );
not ( n67034 , n67033 );
and ( n67035 , n63492 , n61015 );
not ( n67036 , n67035 );
and ( n67037 , n67034 , n67036 );
and ( n67038 , n61505 , n62998 );
not ( n67039 , n67038 );
and ( n67040 , n67036 , n67039 );
and ( n67041 , n67034 , n67039 );
or ( n67042 , n67037 , n67040 , n67041 );
and ( n67043 , n66720 , n58444 );
not ( n67044 , n67043 );
and ( n67045 , n67044 , n66967 );
and ( n67046 , n63024 , n61481 );
not ( n67047 , n67046 );
and ( n67048 , n66967 , n67047 );
and ( n67049 , n67044 , n67047 );
or ( n67050 , n67045 , n67048 , n67049 );
and ( n67051 , n67042 , n67050 );
and ( n67052 , n66415 , n58542 );
not ( n67053 , n67052 );
and ( n67054 , n64221 , n60372 );
not ( n67055 , n67054 );
or ( n67056 , n67053 , n67055 );
and ( n67057 , n67050 , n67056 );
and ( n67058 , n67042 , n67056 );
or ( n67059 , n67051 , n67057 , n67058 );
and ( n67060 , n60821 , n63766 );
not ( n67061 , n67060 );
and ( n67062 , n63987 , n60711 );
not ( n67063 , n67062 );
and ( n67064 , n67061 , n67063 );
and ( n67065 , n47962 , n57187 );
and ( n67066 , n47778 , n57184 );
nor ( n67067 , n67065 , n67066 );
xnor ( n67068 , n67067 , n56175 );
and ( n67069 , n48272 , n56503 );
and ( n67070 , n48108 , n56501 );
nor ( n67071 , n67069 , n67070 );
xnor ( n67072 , n67071 , n56178 );
and ( n67073 , n67068 , n67072 );
and ( n67074 , n48632 , n55851 );
and ( n67075 , n48384 , n55849 );
nor ( n67076 , n67074 , n67075 );
xnor ( n67077 , n67076 , n55506 );
and ( n67078 , n67072 , n67077 );
and ( n67079 , n67068 , n67077 );
or ( n67080 , n67073 , n67078 , n67079 );
and ( n67081 , n67064 , n67080 );
and ( n67082 , n48988 , n55159 );
and ( n67083 , n48709 , n55157 );
nor ( n67084 , n67082 , n67083 );
xnor ( n67085 , n67084 , n54864 );
and ( n67086 , n49374 , n54535 );
and ( n67087 , n49115 , n54533 );
nor ( n67088 , n67086 , n67087 );
xnor ( n67089 , n67088 , n54237 );
and ( n67090 , n67085 , n67089 );
and ( n67091 , n49781 , n53928 );
and ( n67092 , n49570 , n53926 );
nor ( n67093 , n67091 , n67092 );
xnor ( n67094 , n67093 , n53652 );
and ( n67095 , n67089 , n67094 );
and ( n67096 , n67085 , n67094 );
or ( n67097 , n67090 , n67095 , n67096 );
and ( n67098 , n67080 , n67097 );
and ( n67099 , n67064 , n67097 );
or ( n67100 , n67081 , n67098 , n67099 );
and ( n67101 , n67059 , n67100 );
and ( n67102 , n50195 , n53357 );
and ( n67103 , n49976 , n53355 );
nor ( n67104 , n67102 , n67103 );
xnor ( n67105 , n67104 , n53060 );
and ( n67106 , n50625 , n52799 );
and ( n67107 , n50404 , n52797 );
nor ( n67108 , n67106 , n67107 );
xnor ( n67109 , n67108 , n52538 );
and ( n67110 , n67105 , n67109 );
and ( n67111 , n51077 , n52269 );
and ( n67112 , n50726 , n52267 );
nor ( n67113 , n67111 , n67112 );
xnor ( n67114 , n67113 , n52008 );
and ( n67115 , n67109 , n67114 );
and ( n67116 , n67105 , n67114 );
or ( n67117 , n67110 , n67115 , n67116 );
and ( n67118 , n51510 , n51750 );
and ( n67119 , n51298 , n51748 );
nor ( n67120 , n67118 , n67119 );
xnor ( n67121 , n67120 , n51520 );
and ( n67122 , n52082 , n51221 );
and ( n67123 , n51734 , n51219 );
nor ( n67124 , n67122 , n67123 );
xnor ( n67125 , n67124 , n51000 );
and ( n67126 , n67121 , n67125 );
and ( n67127 , n52612 , n50783 );
and ( n67128 , n52332 , n50781 );
nor ( n67129 , n67127 , n67128 );
xnor ( n67130 , n67129 , n50557 );
and ( n67131 , n67125 , n67130 );
and ( n67132 , n67121 , n67130 );
or ( n67133 , n67126 , n67131 , n67132 );
and ( n67134 , n67117 , n67133 );
and ( n67135 , n53041 , n50338 );
and ( n67136 , n52790 , n50336 );
nor ( n67137 , n67135 , n67136 );
xnor ( n67138 , n67137 , n50111 );
and ( n67139 , n53639 , n49896 );
and ( n67140 , n53328 , n49894 );
nor ( n67141 , n67139 , n67140 );
xnor ( n67142 , n67141 , n49711 );
and ( n67143 , n67138 , n67142 );
and ( n67144 , n54227 , n49513 );
and ( n67145 , n53922 , n49511 );
nor ( n67146 , n67144 , n67145 );
xnor ( n67147 , n67146 , n49310 );
and ( n67148 , n67142 , n67147 );
and ( n67149 , n67138 , n67147 );
or ( n67150 , n67143 , n67148 , n67149 );
and ( n67151 , n67133 , n67150 );
and ( n67152 , n67117 , n67150 );
or ( n67153 , n67134 , n67151 , n67152 );
and ( n67154 , n67100 , n67153 );
and ( n67155 , n67059 , n67153 );
or ( n67156 , n67101 , n67154 , n67155 );
and ( n67157 , n54942 , n49121 );
and ( n67158 , n54604 , n49119 );
nor ( n67159 , n67157 , n67158 );
xnor ( n67160 , n67159 , n48932 );
and ( n67161 , n55497 , n48740 );
and ( n67162 , n55143 , n48738 );
nor ( n67163 , n67161 , n67162 );
xnor ( n67164 , n67163 , n48571 );
and ( n67165 , n67160 , n67164 );
and ( n67166 , n56255 , n48394 );
and ( n67167 , n55756 , n48392 );
nor ( n67168 , n67166 , n67167 );
xnor ( n67169 , n67168 , n48220 );
and ( n67170 , n67164 , n67169 );
and ( n67171 , n67160 , n67169 );
or ( n67172 , n67165 , n67170 , n67171 );
and ( n67173 , n56915 , n48042 );
and ( n67174 , n56388 , n48040 );
nor ( n67175 , n67173 , n67174 );
xnor ( n67176 , n67175 , n47921 );
and ( n67177 , n67176 , n66711 );
xor ( n67178 , n42764 , n45544 );
buf ( n67179 , n67178 );
buf ( n67180 , n67179 );
buf ( n67181 , n67180 );
and ( n67182 , n66711 , n67181 );
and ( n67183 , n67176 , n67181 );
or ( n67184 , n67177 , n67182 , n67183 );
and ( n67185 , n67172 , n67184 );
xor ( n67186 , n66625 , n66629 );
xor ( n67187 , n67186 , n66634 );
and ( n67188 , n67184 , n67187 );
and ( n67189 , n67172 , n67187 );
or ( n67190 , n67185 , n67188 , n67189 );
xor ( n67191 , n66642 , n66646 );
xor ( n67192 , n67191 , n66651 );
xor ( n67193 , n66661 , n66665 );
xor ( n67194 , n67193 , n66670 );
and ( n67195 , n67192 , n67194 );
xor ( n67196 , n66677 , n66681 );
xor ( n67197 , n67196 , n66686 );
and ( n67198 , n67194 , n67197 );
and ( n67199 , n67192 , n67197 );
or ( n67200 , n67195 , n67198 , n67199 );
and ( n67201 , n67190 , n67200 );
buf ( n67202 , n66562 );
xor ( n67203 , n67202 , n66564 );
and ( n67204 , n67200 , n67203 );
and ( n67205 , n67190 , n67203 );
or ( n67206 , n67201 , n67204 , n67205 );
and ( n67207 , n67156 , n67206 );
xor ( n67208 , n66568 , n66569 );
xor ( n67209 , n67208 , n66580 );
xor ( n67210 , n66594 , n66603 );
xor ( n67211 , n67210 , n66606 );
and ( n67212 , n67209 , n67211 );
xor ( n67213 , n66621 , n66637 );
xor ( n67214 , n67213 , n66654 );
and ( n67215 , n67211 , n67214 );
and ( n67216 , n67209 , n67214 );
or ( n67217 , n67212 , n67215 , n67216 );
and ( n67218 , n67206 , n67217 );
and ( n67219 , n67156 , n67217 );
or ( n67220 , n67207 , n67218 , n67219 );
and ( n67221 , n67032 , n67220 );
xor ( n67222 , n66673 , n66689 );
xor ( n67223 , n67222 , n66706 );
xor ( n67224 , n66725 , n66727 );
xor ( n67225 , n67224 , n66730 );
and ( n67226 , n67223 , n67225 );
xor ( n67227 , n66739 , n66741 );
xor ( n67228 , n67227 , n66744 );
and ( n67229 , n67225 , n67228 );
and ( n67230 , n67223 , n67228 );
or ( n67231 , n67226 , n67229 , n67230 );
xor ( n67232 , n66489 , n66491 );
xor ( n67233 , n67232 , n66494 );
and ( n67234 , n67231 , n67233 );
xor ( n67235 , n66499 , n66501 );
xor ( n67236 , n67235 , n66503 );
and ( n67237 , n67233 , n67236 );
and ( n67238 , n67231 , n67236 );
or ( n67239 , n67234 , n67237 , n67238 );
and ( n67240 , n67220 , n67239 );
and ( n67241 , n67032 , n67239 );
or ( n67242 , n67221 , n67240 , n67241 );
xor ( n67243 , n66535 , n66544 );
xor ( n67244 , n67243 , n66550 );
xor ( n67245 , n66566 , n66583 );
xor ( n67246 , n67245 , n66609 );
and ( n67247 , n67244 , n67246 );
xor ( n67248 , n66657 , n66709 );
xor ( n67249 , n67248 , n66733 );
and ( n67250 , n67246 , n67249 );
and ( n67251 , n67244 , n67249 );
or ( n67252 , n67247 , n67250 , n67251 );
xor ( n67253 , n66442 , n66444 );
xor ( n67254 , n67253 , n66447 );
and ( n67255 , n67252 , n67254 );
xor ( n67256 , n66452 , n66453 );
xor ( n67257 , n67256 , n66483 );
and ( n67258 , n67254 , n67257 );
and ( n67259 , n67252 , n67257 );
or ( n67260 , n67255 , n67258 , n67259 );
and ( n67261 , n67242 , n67260 );
xor ( n67262 , n66497 , n66506 );
xor ( n67263 , n67262 , n66553 );
xor ( n67264 , n66612 , n66736 );
xor ( n67265 , n67264 , n66755 );
and ( n67266 , n67263 , n67265 );
xor ( n67267 , n66768 , n66770 );
xor ( n67268 , n67267 , n66773 );
and ( n67269 , n67265 , n67268 );
and ( n67270 , n67263 , n67268 );
or ( n67271 , n67266 , n67269 , n67270 );
and ( n67272 , n67260 , n67271 );
and ( n67273 , n67242 , n67271 );
or ( n67274 , n67261 , n67272 , n67273 );
xor ( n67275 , n66391 , n66392 );
xor ( n67276 , n67275 , n66437 );
xor ( n67277 , n66450 , n66486 );
xor ( n67278 , n67277 , n66556 );
and ( n67279 , n67276 , n67278 );
xor ( n67280 , n66758 , n66776 );
xor ( n67281 , n67280 , n66787 );
and ( n67282 , n67278 , n67281 );
and ( n67283 , n67276 , n67281 );
or ( n67284 , n67279 , n67282 , n67283 );
and ( n67285 , n67274 , n67284 );
xor ( n67286 , n66440 , n66559 );
xor ( n67287 , n67286 , n66790 );
and ( n67288 , n67284 , n67287 );
and ( n67289 , n67274 , n67287 );
or ( n67290 , n67285 , n67288 , n67289 );
xor ( n67291 , n66793 , n66811 );
xor ( n67292 , n67291 , n66814 );
and ( n67293 , n67290 , n67292 );
xor ( n67294 , n66803 , n66805 );
xor ( n67295 , n67294 , n66808 );
xor ( n67296 , n66795 , n66797 );
xor ( n67297 , n67296 , n66800 );
xor ( n67298 , n66779 , n66781 );
xor ( n67299 , n67298 , n66784 );
xor ( n67300 , n66747 , n66749 );
xor ( n67301 , n67300 , n66752 );
xor ( n67302 , n66760 , n66762 );
xor ( n67303 , n67302 , n66765 );
and ( n67304 , n67301 , n67303 );
xor ( n67305 , n66880 , n66882 );
xor ( n67306 , n67305 , n66885 );
xor ( n67307 , n66906 , n66908 );
xor ( n67308 , n67307 , n66911 );
and ( n67309 , n67306 , n67308 );
xnor ( n67310 , n66935 , n66937 );
and ( n67311 , n67308 , n67310 );
and ( n67312 , n67306 , n67310 );
or ( n67313 , n67309 , n67311 , n67312 );
and ( n67314 , n67303 , n67313 );
and ( n67315 , n67301 , n67313 );
or ( n67316 , n67304 , n67314 , n67315 );
and ( n67317 , n67299 , n67316 );
xor ( n67318 , n66969 , n66971 );
xor ( n67319 , n67318 , n66974 );
xor ( n67320 , n66572 , n66574 );
xor ( n67321 , n67320 , n66577 );
and ( n67322 , n67319 , n67321 );
xor ( n67323 , n66595 , n66597 );
xor ( n67324 , n67323 , n66600 );
and ( n67325 , n67321 , n67324 );
and ( n67326 , n67319 , n67324 );
or ( n67327 , n67322 , n67325 , n67326 );
xor ( n67328 , n66694 , n66698 );
xor ( n67329 , n67328 , n66703 );
xor ( n67330 , n66713 , n66717 );
xor ( n67331 , n67330 , n66722 );
and ( n67332 , n67329 , n67331 );
xor ( n67333 , n66927 , n66929 );
xor ( n67334 , n67333 , n66932 );
and ( n67335 , n67331 , n67334 );
and ( n67336 , n67329 , n67334 );
or ( n67337 , n67332 , n67335 , n67336 );
and ( n67338 , n67327 , n67337 );
xnor ( n67339 , n66990 , n66992 );
xor ( n67340 , n66998 , n66999 );
and ( n67341 , n67339 , n67340 );
buf ( n67342 , n20267 );
buf ( n67343 , n67342 );
and ( n67344 , n67343 , n58294 );
not ( n67345 , n67344 );
and ( n67346 , n65678 , n59207 );
not ( n67347 , n67346 );
and ( n67348 , n67345 , n67347 );
and ( n67349 , n64221 , n60711 );
not ( n67350 , n67349 );
and ( n67351 , n67347 , n67350 );
and ( n67352 , n67345 , n67350 );
or ( n67353 , n67348 , n67351 , n67352 );
xor ( n67354 , n67015 , n67017 );
xor ( n67355 , n67354 , n67020 );
and ( n67356 , n67353 , n67355 );
xor ( n67357 , n67044 , n66967 );
xor ( n67358 , n67357 , n67047 );
and ( n67359 , n67355 , n67358 );
and ( n67360 , n67353 , n67358 );
or ( n67361 , n67356 , n67359 , n67360 );
and ( n67362 , n67340 , n67361 );
and ( n67363 , n67339 , n67361 );
or ( n67364 , n67341 , n67362 , n67363 );
and ( n67365 , n67337 , n67364 );
and ( n67366 , n67327 , n67364 );
or ( n67367 , n67338 , n67365 , n67366 );
and ( n67368 , n58292 , n67013 );
not ( n67369 , n67368 );
and ( n67370 , n58628 , n66917 );
not ( n67371 , n67370 );
and ( n67372 , n67369 , n67371 );
and ( n67373 , n63024 , n61914 );
not ( n67374 , n67373 );
and ( n67375 , n67371 , n67374 );
and ( n67376 , n67369 , n67374 );
or ( n67377 , n67372 , n67375 , n67376 );
and ( n67378 , n65606 , n59207 );
not ( n67379 , n67378 );
and ( n67380 , n67377 , n67379 );
xor ( n67381 , n66919 , n66921 );
xor ( n67382 , n67381 , n66924 );
and ( n67383 , n67379 , n67382 );
and ( n67384 , n67377 , n67382 );
or ( n67385 , n67380 , n67383 , n67384 );
xor ( n67386 , n67034 , n67036 );
xor ( n67387 , n67386 , n67039 );
xnor ( n67388 , n67053 , n67055 );
and ( n67389 , n67387 , n67388 );
buf ( n67390 , n67389 );
and ( n67391 , n67385 , n67390 );
xor ( n67392 , n67061 , n67063 );
and ( n67393 , n48108 , n57187 );
and ( n67394 , n47962 , n57184 );
nor ( n67395 , n67393 , n67394 );
xnor ( n67396 , n67395 , n56175 );
and ( n67397 , n48384 , n56503 );
and ( n67398 , n48272 , n56501 );
nor ( n67399 , n67397 , n67398 );
xnor ( n67400 , n67399 , n56178 );
and ( n67401 , n67396 , n67400 );
and ( n67402 , n52790 , n50783 );
and ( n67403 , n52612 , n50781 );
nor ( n67404 , n67402 , n67403 );
xnor ( n67405 , n67404 , n50557 );
and ( n67406 , n67400 , n67405 );
and ( n67407 , n67396 , n67405 );
or ( n67408 , n67401 , n67406 , n67407 );
and ( n67409 , n67392 , n67408 );
buf ( n67410 , n20267 );
buf ( n67411 , n67410 );
and ( n67412 , n57948 , n67411 );
not ( n67413 , n67412 );
and ( n67414 , n59365 , n66005 );
not ( n67415 , n67414 );
and ( n67416 , n67413 , n67415 );
and ( n67417 , n60821 , n64412 );
not ( n67418 , n67417 );
and ( n67419 , n67415 , n67418 );
and ( n67420 , n67413 , n67418 );
or ( n67421 , n67416 , n67419 , n67420 );
and ( n67422 , n67408 , n67421 );
and ( n67423 , n67392 , n67421 );
or ( n67424 , n67409 , n67422 , n67423 );
and ( n67425 , n67390 , n67424 );
and ( n67426 , n67385 , n67424 );
or ( n67427 , n67391 , n67425 , n67426 );
and ( n67428 , n60376 , n64811 );
not ( n67429 , n67428 );
and ( n67430 , n61505 , n63679 );
not ( n67431 , n67430 );
and ( n67432 , n67429 , n67431 );
and ( n67433 , n61918 , n62998 );
not ( n67434 , n67433 );
and ( n67435 , n67431 , n67434 );
and ( n67436 , n67429 , n67434 );
or ( n67437 , n67432 , n67435 , n67436 );
and ( n67438 , n66415 , n58911 );
not ( n67439 , n67438 );
and ( n67440 , n64548 , n60372 );
not ( n67441 , n67440 );
and ( n67442 , n67439 , n67441 );
and ( n67443 , n67437 , n67442 );
and ( n67444 , n66980 , n58444 );
not ( n67445 , n67444 );
and ( n67446 , n66720 , n58542 );
not ( n67447 , n67446 );
or ( n67448 , n67445 , n67447 );
and ( n67449 , n67442 , n67448 );
and ( n67450 , n67437 , n67448 );
or ( n67451 , n67443 , n67449 , n67450 );
and ( n67452 , n53328 , n50338 );
and ( n67453 , n53041 , n50336 );
nor ( n67454 , n67452 , n67453 );
xnor ( n67455 , n67454 , n50111 );
and ( n67456 , n53922 , n49896 );
and ( n67457 , n53639 , n49894 );
nor ( n67458 , n67456 , n67457 );
xnor ( n67459 , n67458 , n49711 );
and ( n67460 , n67455 , n67459 );
and ( n67461 , n48709 , n55851 );
and ( n67462 , n48632 , n55849 );
nor ( n67463 , n67461 , n67462 );
xnor ( n67464 , n67463 , n55506 );
and ( n67465 , n49115 , n55159 );
and ( n67466 , n48988 , n55157 );
nor ( n67467 , n67465 , n67466 );
xnor ( n67468 , n67467 , n54864 );
and ( n67469 , n67464 , n67468 );
and ( n67470 , n49570 , n54535 );
and ( n67471 , n49374 , n54533 );
nor ( n67472 , n67470 , n67471 );
xnor ( n67473 , n67472 , n54237 );
and ( n67474 , n67468 , n67473 );
and ( n67475 , n67464 , n67473 );
or ( n67476 , n67469 , n67474 , n67475 );
and ( n67477 , n67460 , n67476 );
and ( n67478 , n49976 , n53928 );
and ( n67479 , n49781 , n53926 );
nor ( n67480 , n67478 , n67479 );
xnor ( n67481 , n67480 , n53652 );
and ( n67482 , n50404 , n53357 );
and ( n67483 , n50195 , n53355 );
nor ( n67484 , n67482 , n67483 );
xnor ( n67485 , n67484 , n53060 );
and ( n67486 , n67481 , n67485 );
and ( n67487 , n50726 , n52799 );
and ( n67488 , n50625 , n52797 );
nor ( n67489 , n67487 , n67488 );
xnor ( n67490 , n67489 , n52538 );
and ( n67491 , n67485 , n67490 );
and ( n67492 , n67481 , n67490 );
or ( n67493 , n67486 , n67491 , n67492 );
and ( n67494 , n67476 , n67493 );
and ( n67495 , n67460 , n67493 );
or ( n67496 , n67477 , n67494 , n67495 );
and ( n67497 , n67451 , n67496 );
and ( n67498 , n51298 , n52269 );
and ( n67499 , n51077 , n52267 );
nor ( n67500 , n67498 , n67499 );
xnor ( n67501 , n67500 , n52008 );
and ( n67502 , n51734 , n51750 );
and ( n67503 , n51510 , n51748 );
nor ( n67504 , n67502 , n67503 );
xnor ( n67505 , n67504 , n51520 );
and ( n67506 , n67501 , n67505 );
and ( n67507 , n52332 , n51221 );
and ( n67508 , n52082 , n51219 );
nor ( n67509 , n67507 , n67508 );
xnor ( n67510 , n67509 , n51000 );
and ( n67511 , n67505 , n67510 );
and ( n67512 , n67501 , n67510 );
or ( n67513 , n67506 , n67511 , n67512 );
and ( n67514 , n54604 , n49513 );
and ( n67515 , n54227 , n49511 );
nor ( n67516 , n67514 , n67515 );
xnor ( n67517 , n67516 , n49310 );
and ( n67518 , n55143 , n49121 );
and ( n67519 , n54942 , n49119 );
nor ( n67520 , n67518 , n67519 );
xnor ( n67521 , n67520 , n48932 );
and ( n67522 , n67517 , n67521 );
and ( n67523 , n55756 , n48740 );
and ( n67524 , n55497 , n48738 );
nor ( n67525 , n67523 , n67524 );
xnor ( n67526 , n67525 , n48571 );
and ( n67527 , n67521 , n67526 );
and ( n67528 , n67517 , n67526 );
or ( n67529 , n67522 , n67527 , n67528 );
and ( n67530 , n67513 , n67529 );
and ( n67531 , n56388 , n48394 );
and ( n67532 , n56255 , n48392 );
nor ( n67533 , n67531 , n67532 );
xnor ( n67534 , n67533 , n48220 );
and ( n67535 , n57063 , n48042 );
and ( n67536 , n56915 , n48040 );
nor ( n67537 , n67535 , n67536 );
xnor ( n67538 , n67537 , n47921 );
and ( n67539 , n67534 , n67538 );
and ( n67540 , n57063 , n48040 );
not ( n67541 , n67540 );
and ( n67542 , n67541 , n47921 );
and ( n67543 , n67538 , n67542 );
and ( n67544 , n67534 , n67542 );
or ( n67545 , n67539 , n67543 , n67544 );
and ( n67546 , n67529 , n67545 );
and ( n67547 , n67513 , n67545 );
or ( n67548 , n67530 , n67546 , n67547 );
and ( n67549 , n67496 , n67548 );
and ( n67550 , n67451 , n67548 );
or ( n67551 , n67497 , n67549 , n67550 );
and ( n67552 , n67427 , n67551 );
xor ( n67553 , n42765 , n45543 );
buf ( n67554 , n67553 );
buf ( n67555 , n67554 );
buf ( n67556 , n67555 );
and ( n67557 , n65177 , n59920 );
not ( n67558 , n67557 );
and ( n67559 , n67556 , n67558 );
and ( n67560 , n63987 , n61015 );
not ( n67561 , n67560 );
and ( n67562 , n67558 , n67561 );
and ( n67563 , n67556 , n67561 );
or ( n67564 , n67559 , n67562 , n67563 );
xor ( n67565 , n67068 , n67072 );
xor ( n67566 , n67565 , n67077 );
and ( n67567 , n67564 , n67566 );
xor ( n67568 , n67085 , n67089 );
xor ( n67569 , n67568 , n67094 );
and ( n67570 , n67566 , n67569 );
and ( n67571 , n67564 , n67569 );
or ( n67572 , n67567 , n67570 , n67571 );
xor ( n67573 , n67105 , n67109 );
xor ( n67574 , n67573 , n67114 );
xor ( n67575 , n67121 , n67125 );
xor ( n67576 , n67575 , n67130 );
and ( n67577 , n67574 , n67576 );
xor ( n67578 , n67138 , n67142 );
xor ( n67579 , n67578 , n67147 );
and ( n67580 , n67576 , n67579 );
and ( n67581 , n67574 , n67579 );
or ( n67582 , n67577 , n67580 , n67581 );
and ( n67583 , n67572 , n67582 );
buf ( n67584 , n67002 );
xor ( n67585 , n67584 , n67004 );
and ( n67586 , n67582 , n67585 );
and ( n67587 , n67572 , n67585 );
or ( n67588 , n67583 , n67586 , n67587 );
and ( n67589 , n67551 , n67588 );
and ( n67590 , n67427 , n67588 );
or ( n67591 , n67552 , n67589 , n67590 );
and ( n67592 , n67367 , n67591 );
xor ( n67593 , n67009 , n67010 );
xor ( n67594 , n67593 , n67023 );
xor ( n67595 , n67042 , n67050 );
xor ( n67596 , n67595 , n67056 );
and ( n67597 , n67594 , n67596 );
xor ( n67598 , n67064 , n67080 );
xor ( n67599 , n67598 , n67097 );
and ( n67600 , n67596 , n67599 );
and ( n67601 , n67594 , n67599 );
or ( n67602 , n67597 , n67600 , n67601 );
xor ( n67603 , n67117 , n67133 );
xor ( n67604 , n67603 , n67150 );
xor ( n67605 , n67172 , n67184 );
xor ( n67606 , n67605 , n67187 );
and ( n67607 , n67604 , n67606 );
xor ( n67608 , n67192 , n67194 );
xor ( n67609 , n67608 , n67197 );
and ( n67610 , n67606 , n67609 );
and ( n67611 , n67604 , n67609 );
or ( n67612 , n67607 , n67610 , n67611 );
and ( n67613 , n67602 , n67612 );
xor ( n67614 , n66958 , n66960 );
xor ( n67615 , n67614 , n66962 );
and ( n67616 , n67612 , n67615 );
and ( n67617 , n67602 , n67615 );
or ( n67618 , n67613 , n67616 , n67617 );
and ( n67619 , n67591 , n67618 );
and ( n67620 , n67367 , n67618 );
or ( n67621 , n67592 , n67619 , n67620 );
and ( n67622 , n67316 , n67621 );
and ( n67623 , n67299 , n67621 );
or ( n67624 , n67317 , n67622 , n67623 );
and ( n67625 , n67297 , n67624 );
xor ( n67626 , n66966 , n66977 );
xor ( n67627 , n67626 , n66993 );
xor ( n67628 , n67000 , n67006 );
xor ( n67629 , n67628 , n67026 );
and ( n67630 , n67627 , n67629 );
xor ( n67631 , n67059 , n67100 );
xor ( n67632 , n67631 , n67153 );
and ( n67633 , n67629 , n67632 );
and ( n67634 , n67627 , n67632 );
or ( n67635 , n67630 , n67633 , n67634 );
xor ( n67636 , n67190 , n67200 );
xor ( n67637 , n67636 , n67203 );
xor ( n67638 , n67209 , n67211 );
xor ( n67639 , n67638 , n67214 );
and ( n67640 , n67637 , n67639 );
xor ( n67641 , n67223 , n67225 );
xor ( n67642 , n67641 , n67228 );
and ( n67643 , n67639 , n67642 );
and ( n67644 , n67637 , n67642 );
or ( n67645 , n67640 , n67643 , n67644 );
and ( n67646 , n67635 , n67645 );
xor ( n67647 , n66863 , n66865 );
xor ( n67648 , n67647 , n66868 );
and ( n67649 , n67645 , n67648 );
and ( n67650 , n67635 , n67648 );
or ( n67651 , n67646 , n67649 , n67650 );
xor ( n67652 , n66888 , n66914 );
xor ( n67653 , n67652 , n66938 );
xor ( n67654 , n66965 , n66996 );
xor ( n67655 , n67654 , n67029 );
and ( n67656 , n67653 , n67655 );
xor ( n67657 , n67156 , n67206 );
xor ( n67658 , n67657 , n67217 );
and ( n67659 , n67655 , n67658 );
and ( n67660 , n67653 , n67658 );
or ( n67661 , n67656 , n67659 , n67660 );
and ( n67662 , n67651 , n67661 );
xor ( n67663 , n66861 , n66871 );
xor ( n67664 , n67663 , n66941 );
and ( n67665 , n67661 , n67664 );
and ( n67666 , n67651 , n67664 );
or ( n67667 , n67662 , n67665 , n67666 );
and ( n67668 , n67624 , n67667 );
and ( n67669 , n67297 , n67667 );
or ( n67670 , n67625 , n67668 , n67669 );
and ( n67671 , n67295 , n67670 );
xor ( n67672 , n67032 , n67220 );
xor ( n67673 , n67672 , n67239 );
xor ( n67674 , n67252 , n67254 );
xor ( n67675 , n67674 , n67257 );
and ( n67676 , n67673 , n67675 );
xor ( n67677 , n67263 , n67265 );
xor ( n67678 , n67677 , n67268 );
and ( n67679 , n67675 , n67678 );
and ( n67680 , n67673 , n67678 );
or ( n67681 , n67676 , n67679 , n67680 );
xor ( n67682 , n66856 , n66858 );
xor ( n67683 , n67682 , n66944 );
and ( n67684 , n67681 , n67683 );
xor ( n67685 , n67242 , n67260 );
xor ( n67686 , n67685 , n67271 );
and ( n67687 , n67683 , n67686 );
and ( n67688 , n67681 , n67686 );
or ( n67689 , n67684 , n67687 , n67688 );
and ( n67690 , n67670 , n67689 );
and ( n67691 , n67295 , n67689 );
or ( n67692 , n67671 , n67690 , n67691 );
and ( n67693 , n67292 , n67692 );
and ( n67694 , n67290 , n67692 );
or ( n67695 , n67293 , n67693 , n67694 );
and ( n67696 , n66955 , n67695 );
and ( n67697 , n66953 , n67695 );
or ( n67698 , n66956 , n67696 , n67697 );
and ( n67699 , n66844 , n67698 );
xor ( n67700 , n66846 , n66848 );
xor ( n67701 , n67700 , n66950 );
xor ( n67702 , n66851 , n66853 );
xor ( n67703 , n67702 , n66947 );
xor ( n67704 , n67274 , n67284 );
xor ( n67705 , n67704 , n67287 );
and ( n67706 , n67703 , n67705 );
xor ( n67707 , n67276 , n67278 );
xor ( n67708 , n67707 , n67281 );
xor ( n67709 , n67231 , n67233 );
xor ( n67710 , n67709 , n67236 );
xor ( n67711 , n67244 , n67246 );
xor ( n67712 , n67711 , n67249 );
and ( n67713 , n67710 , n67712 );
and ( n67714 , n58915 , n66469 );
not ( n67715 , n67714 );
buf ( n67716 , n67715 );
and ( n67717 , n59365 , n65586 );
not ( n67718 , n67717 );
and ( n67719 , n67716 , n67718 );
and ( n67720 , n59615 , n65210 );
not ( n67721 , n67720 );
and ( n67722 , n67718 , n67721 );
and ( n67723 , n67716 , n67721 );
or ( n67724 , n67719 , n67722 , n67723 );
and ( n67725 , n66720 , n58911 );
not ( n67726 , n67725 );
buf ( n67727 , n67726 );
and ( n67728 , n59615 , n65586 );
not ( n67729 , n67728 );
and ( n67730 , n67727 , n67729 );
and ( n67731 , n59908 , n65210 );
not ( n67732 , n67731 );
and ( n67733 , n67729 , n67732 );
and ( n67734 , n67727 , n67732 );
or ( n67735 , n67730 , n67733 , n67734 );
and ( n67736 , n61008 , n63766 );
not ( n67737 , n67736 );
and ( n67738 , n67714 , n67737 );
and ( n67739 , n62377 , n62868 );
not ( n67740 , n67739 );
and ( n67741 , n67737 , n67740 );
and ( n67742 , n67714 , n67740 );
or ( n67743 , n67738 , n67741 , n67742 );
and ( n67744 , n67735 , n67743 );
xor ( n67745 , n66890 , n66892 );
xor ( n67746 , n67745 , n66895 );
and ( n67747 , n67743 , n67746 );
and ( n67748 , n67735 , n67746 );
or ( n67749 , n67744 , n67747 , n67748 );
and ( n67750 , n67724 , n67749 );
xor ( n67751 , n66898 , n66900 );
xor ( n67752 , n67751 , n66903 );
and ( n67753 , n67749 , n67752 );
and ( n67754 , n67724 , n67752 );
or ( n67755 , n67750 , n67753 , n67754 );
xor ( n67756 , n67439 , n67441 );
and ( n67757 , n65606 , n59611 );
not ( n67758 , n67757 );
and ( n67759 , n67756 , n67758 );
and ( n67760 , n63492 , n61481 );
not ( n67761 , n67760 );
and ( n67762 , n67758 , n67761 );
and ( n67763 , n67756 , n67761 );
or ( n67764 , n67759 , n67762 , n67763 );
xor ( n67765 , n66982 , n66984 );
xor ( n67766 , n67765 , n66987 );
or ( n67767 , n67764 , n67766 );
xor ( n67768 , n67160 , n67164 );
xor ( n67769 , n67768 , n67169 );
xor ( n67770 , n67176 , n66711 );
xor ( n67771 , n67770 , n67181 );
and ( n67772 , n67769 , n67771 );
xor ( n67773 , n67716 , n67718 );
xor ( n67774 , n67773 , n67721 );
and ( n67775 , n67771 , n67774 );
and ( n67776 , n67769 , n67774 );
or ( n67777 , n67772 , n67775 , n67776 );
and ( n67778 , n67767 , n67777 );
xor ( n67779 , n67353 , n67355 );
xor ( n67780 , n67779 , n67358 );
xor ( n67781 , n67377 , n67379 );
xor ( n67782 , n67781 , n67382 );
and ( n67783 , n67780 , n67782 );
and ( n67784 , n58292 , n67411 );
not ( n67785 , n67784 );
and ( n67786 , n58628 , n67013 );
not ( n67787 , n67786 );
and ( n67788 , n67785 , n67787 );
and ( n67789 , n61918 , n63679 );
not ( n67790 , n67789 );
and ( n67791 , n67787 , n67790 );
and ( n67792 , n67785 , n67790 );
or ( n67793 , n67788 , n67791 , n67792 );
and ( n67794 , n59615 , n66005 );
not ( n67795 , n67794 );
and ( n67796 , n61505 , n63766 );
not ( n67797 , n67796 );
and ( n67798 , n67795 , n67797 );
and ( n67799 , n62377 , n62998 );
not ( n67800 , n67799 );
and ( n67801 , n67797 , n67800 );
and ( n67802 , n67795 , n67800 );
or ( n67803 , n67798 , n67801 , n67802 );
and ( n67804 , n67793 , n67803 );
and ( n67805 , n65177 , n60372 );
not ( n67806 , n67805 );
and ( n67807 , n67725 , n67806 );
and ( n67808 , n61008 , n64412 );
not ( n67809 , n67808 );
and ( n67810 , n67806 , n67809 );
and ( n67811 , n67725 , n67809 );
or ( n67812 , n67807 , n67810 , n67811 );
and ( n67813 , n67803 , n67812 );
and ( n67814 , n67793 , n67812 );
or ( n67815 , n67804 , n67813 , n67814 );
and ( n67816 , n67782 , n67815 );
and ( n67817 , n67780 , n67815 );
or ( n67818 , n67783 , n67816 , n67817 );
and ( n67819 , n67777 , n67818 );
and ( n67820 , n67767 , n67818 );
or ( n67821 , n67778 , n67819 , n67820 );
and ( n67822 , n67755 , n67821 );
and ( n67823 , n62593 , n62151 );
not ( n67824 , n67823 );
xor ( n67825 , n67396 , n67400 );
xor ( n67826 , n67825 , n67405 );
and ( n67827 , n67824 , n67826 );
buf ( n67828 , n67827 );
xor ( n67829 , n67429 , n67431 );
xor ( n67830 , n67829 , n67434 );
xor ( n67831 , n67369 , n67371 );
xor ( n67832 , n67831 , n67374 );
and ( n67833 , n67830 , n67832 );
xor ( n67834 , n67345 , n67347 );
xor ( n67835 , n67834 , n67350 );
and ( n67836 , n67832 , n67835 );
and ( n67837 , n67830 , n67835 );
or ( n67838 , n67833 , n67836 , n67837 );
and ( n67839 , n67828 , n67838 );
xnor ( n67840 , n67445 , n67447 );
xor ( n67841 , n67455 , n67459 );
and ( n67842 , n67840 , n67841 );
buf ( n67843 , n20270 );
buf ( n67844 , n67843 );
and ( n67845 , n57948 , n67844 );
not ( n67846 , n67845 );
and ( n67847 , n59908 , n65586 );
not ( n67848 , n67847 );
and ( n67849 , n67846 , n67848 );
buf ( n67850 , n62593 );
not ( n67851 , n67850 );
and ( n67852 , n67848 , n67851 );
and ( n67853 , n67846 , n67851 );
or ( n67854 , n67849 , n67852 , n67853 );
and ( n67855 , n67841 , n67854 );
and ( n67856 , n67840 , n67854 );
or ( n67857 , n67842 , n67855 , n67856 );
and ( n67858 , n67838 , n67857 );
and ( n67859 , n67828 , n67857 );
or ( n67860 , n67839 , n67858 , n67859 );
and ( n67861 , n67343 , n58444 );
not ( n67862 , n67861 );
and ( n67863 , n58915 , n66917 );
not ( n67864 , n67863 );
and ( n67865 , n67862 , n67864 );
and ( n67866 , n60376 , n65210 );
not ( n67867 , n67866 );
and ( n67868 , n67864 , n67867 );
and ( n67869 , n67862 , n67867 );
or ( n67870 , n67865 , n67868 , n67869 );
and ( n67871 , n65606 , n59920 );
not ( n67872 , n67871 );
and ( n67873 , n63987 , n61481 );
not ( n67874 , n67873 );
and ( n67875 , n67872 , n67874 );
and ( n67876 , n63024 , n62151 );
not ( n67877 , n67876 );
and ( n67878 , n67874 , n67877 );
and ( n67879 , n67872 , n67877 );
or ( n67880 , n67875 , n67878 , n67879 );
and ( n67881 , n67870 , n67880 );
and ( n67882 , n49781 , n54535 );
and ( n67883 , n49570 , n54533 );
nor ( n67884 , n67882 , n67883 );
xnor ( n67885 , n67884 , n54237 );
and ( n67886 , n50195 , n53928 );
and ( n67887 , n49976 , n53926 );
nor ( n67888 , n67886 , n67887 );
xnor ( n67889 , n67888 , n53652 );
or ( n67890 , n67885 , n67889 );
and ( n67891 , n67880 , n67890 );
and ( n67892 , n67870 , n67890 );
or ( n67893 , n67881 , n67891 , n67892 );
and ( n67894 , n48632 , n56503 );
and ( n67895 , n48384 , n56501 );
nor ( n67896 , n67894 , n67895 );
xnor ( n67897 , n67896 , n56178 );
and ( n67898 , n53041 , n50783 );
and ( n67899 , n52790 , n50781 );
nor ( n67900 , n67898 , n67899 );
xnor ( n67901 , n67900 , n50557 );
and ( n67902 , n67897 , n67901 );
and ( n67903 , n48272 , n57187 );
and ( n67904 , n48108 , n57184 );
nor ( n67905 , n67903 , n67904 );
xnor ( n67906 , n67905 , n56175 );
and ( n67907 , n48988 , n55851 );
and ( n67908 , n48709 , n55849 );
nor ( n67909 , n67907 , n67908 );
xnor ( n67910 , n67909 , n55506 );
and ( n67911 , n67906 , n67910 );
and ( n67912 , n49374 , n55159 );
and ( n67913 , n49115 , n55157 );
nor ( n67914 , n67912 , n67913 );
xnor ( n67915 , n67914 , n54864 );
and ( n67916 , n67910 , n67915 );
and ( n67917 , n67906 , n67915 );
or ( n67918 , n67911 , n67916 , n67917 );
and ( n67919 , n67902 , n67918 );
and ( n67920 , n50625 , n53357 );
and ( n67921 , n50404 , n53355 );
nor ( n67922 , n67920 , n67921 );
xnor ( n67923 , n67922 , n53060 );
and ( n67924 , n51077 , n52799 );
and ( n67925 , n50726 , n52797 );
nor ( n67926 , n67924 , n67925 );
xnor ( n67927 , n67926 , n52538 );
and ( n67928 , n67923 , n67927 );
and ( n67929 , n51510 , n52269 );
and ( n67930 , n51298 , n52267 );
nor ( n67931 , n67929 , n67930 );
xnor ( n67932 , n67931 , n52008 );
and ( n67933 , n67927 , n67932 );
and ( n67934 , n67923 , n67932 );
or ( n67935 , n67928 , n67933 , n67934 );
and ( n67936 , n67918 , n67935 );
and ( n67937 , n67902 , n67935 );
or ( n67938 , n67919 , n67936 , n67937 );
and ( n67939 , n67893 , n67938 );
and ( n67940 , n52082 , n51750 );
and ( n67941 , n51734 , n51748 );
nor ( n67942 , n67940 , n67941 );
xnor ( n67943 , n67942 , n51520 );
and ( n67944 , n52612 , n51221 );
and ( n67945 , n52332 , n51219 );
nor ( n67946 , n67944 , n67945 );
xnor ( n67947 , n67946 , n51000 );
and ( n67948 , n67943 , n67947 );
and ( n67949 , n53639 , n50338 );
and ( n67950 , n53328 , n50336 );
nor ( n67951 , n67949 , n67950 );
xnor ( n67952 , n67951 , n50111 );
and ( n67953 , n67947 , n67952 );
and ( n67954 , n67943 , n67952 );
or ( n67955 , n67948 , n67953 , n67954 );
and ( n67956 , n54227 , n49896 );
and ( n67957 , n53922 , n49894 );
nor ( n67958 , n67956 , n67957 );
xnor ( n67959 , n67958 , n49711 );
and ( n67960 , n54942 , n49513 );
and ( n67961 , n54604 , n49511 );
nor ( n67962 , n67960 , n67961 );
xnor ( n67963 , n67962 , n49310 );
and ( n67964 , n67959 , n67963 );
and ( n67965 , n55497 , n49121 );
and ( n67966 , n55143 , n49119 );
nor ( n67967 , n67965 , n67966 );
xnor ( n67968 , n67967 , n48932 );
and ( n67969 , n67963 , n67968 );
and ( n67970 , n67959 , n67968 );
or ( n67971 , n67964 , n67969 , n67970 );
and ( n67972 , n67955 , n67971 );
and ( n67973 , n56255 , n48740 );
and ( n67974 , n55756 , n48738 );
nor ( n67975 , n67973 , n67974 );
xnor ( n67976 , n67975 , n48571 );
and ( n67977 , n56915 , n48394 );
and ( n67978 , n56388 , n48392 );
nor ( n67979 , n67977 , n67978 );
xnor ( n67980 , n67979 , n48220 );
and ( n67981 , n67976 , n67980 );
and ( n67982 , n67980 , n67540 );
and ( n67983 , n67976 , n67540 );
or ( n67984 , n67981 , n67982 , n67983 );
and ( n67985 , n67971 , n67984 );
and ( n67986 , n67955 , n67984 );
or ( n67987 , n67972 , n67985 , n67986 );
and ( n67988 , n67938 , n67987 );
and ( n67989 , n67893 , n67987 );
or ( n67990 , n67939 , n67988 , n67989 );
and ( n67991 , n67860 , n67990 );
xor ( n67992 , n42767 , n45542 );
buf ( n67993 , n67992 );
buf ( n67994 , n67993 );
buf ( n67995 , n67994 );
buf ( n67996 , n20270 );
buf ( n67997 , n67996 );
and ( n67998 , n67997 , n58294 );
not ( n67999 , n67998 );
and ( n68000 , n67995 , n67999 );
and ( n68001 , n66980 , n58542 );
not ( n68002 , n68001 );
and ( n68003 , n67999 , n68002 );
and ( n68004 , n67995 , n68002 );
or ( n68005 , n68000 , n68003 , n68004 );
and ( n68006 , n66415 , n59207 );
not ( n68007 , n68006 );
and ( n68008 , n64548 , n60711 );
not ( n68009 , n68008 );
and ( n68010 , n68007 , n68009 );
and ( n68011 , n64221 , n61015 );
not ( n68012 , n68011 );
and ( n68013 , n68009 , n68012 );
and ( n68014 , n68007 , n68012 );
or ( n68015 , n68010 , n68013 , n68014 );
and ( n68016 , n68005 , n68015 );
xor ( n68017 , n67464 , n67468 );
xor ( n68018 , n68017 , n67473 );
and ( n68019 , n68015 , n68018 );
and ( n68020 , n68005 , n68018 );
or ( n68021 , n68016 , n68019 , n68020 );
xor ( n68022 , n67481 , n67485 );
xor ( n68023 , n68022 , n67490 );
xor ( n68024 , n67501 , n67505 );
xor ( n68025 , n68024 , n67510 );
and ( n68026 , n68023 , n68025 );
xor ( n68027 , n67517 , n67521 );
xor ( n68028 , n68027 , n67526 );
and ( n68029 , n68025 , n68028 );
and ( n68030 , n68023 , n68028 );
or ( n68031 , n68026 , n68029 , n68030 );
and ( n68032 , n68021 , n68031 );
buf ( n68033 , n67387 );
xor ( n68034 , n68033 , n67388 );
and ( n68035 , n68031 , n68034 );
and ( n68036 , n68021 , n68034 );
or ( n68037 , n68032 , n68035 , n68036 );
and ( n68038 , n67990 , n68037 );
and ( n68039 , n67860 , n68037 );
or ( n68040 , n67991 , n68038 , n68039 );
and ( n68041 , n67821 , n68040 );
and ( n68042 , n67755 , n68040 );
or ( n68043 , n67822 , n68041 , n68042 );
and ( n68044 , n67712 , n68043 );
and ( n68045 , n67710 , n68043 );
or ( n68046 , n67713 , n68044 , n68045 );
xor ( n68047 , n67392 , n67408 );
xor ( n68048 , n68047 , n67421 );
xor ( n68049 , n67437 , n67442 );
xor ( n68050 , n68049 , n67448 );
and ( n68051 , n68048 , n68050 );
xor ( n68052 , n67460 , n67476 );
xor ( n68053 , n68052 , n67493 );
and ( n68054 , n68050 , n68053 );
and ( n68055 , n68048 , n68053 );
or ( n68056 , n68051 , n68054 , n68055 );
xor ( n68057 , n67513 , n67529 );
xor ( n68058 , n68057 , n67545 );
xor ( n68059 , n67564 , n67566 );
xor ( n68060 , n68059 , n67569 );
and ( n68061 , n68058 , n68060 );
xor ( n68062 , n67574 , n67576 );
xor ( n68063 , n68062 , n67579 );
and ( n68064 , n68060 , n68063 );
and ( n68065 , n68058 , n68063 );
or ( n68066 , n68061 , n68064 , n68065 );
and ( n68067 , n68056 , n68066 );
xor ( n68068 , n67329 , n67331 );
xor ( n68069 , n68068 , n67334 );
and ( n68070 , n68066 , n68069 );
and ( n68071 , n68056 , n68069 );
or ( n68072 , n68067 , n68070 , n68071 );
xor ( n68073 , n67339 , n67340 );
xor ( n68074 , n68073 , n67361 );
xor ( n68075 , n67385 , n67390 );
xor ( n68076 , n68075 , n67424 );
and ( n68077 , n68074 , n68076 );
xor ( n68078 , n67451 , n67496 );
xor ( n68079 , n68078 , n67548 );
and ( n68080 , n68076 , n68079 );
and ( n68081 , n68074 , n68079 );
or ( n68082 , n68077 , n68080 , n68081 );
and ( n68083 , n68072 , n68082 );
xor ( n68084 , n67572 , n67582 );
xor ( n68085 , n68084 , n67585 );
xor ( n68086 , n67594 , n67596 );
xor ( n68087 , n68086 , n67599 );
and ( n68088 , n68085 , n68087 );
xor ( n68089 , n67604 , n67606 );
xor ( n68090 , n68089 , n67609 );
and ( n68091 , n68087 , n68090 );
and ( n68092 , n68085 , n68090 );
or ( n68093 , n68088 , n68091 , n68092 );
and ( n68094 , n68082 , n68093 );
and ( n68095 , n68072 , n68093 );
or ( n68096 , n68083 , n68094 , n68095 );
xor ( n68097 , n67306 , n67308 );
xor ( n68098 , n68097 , n67310 );
xor ( n68099 , n67327 , n67337 );
xor ( n68100 , n68099 , n67364 );
and ( n68101 , n68098 , n68100 );
xor ( n68102 , n67427 , n67551 );
xor ( n68103 , n68102 , n67588 );
and ( n68104 , n68100 , n68103 );
and ( n68105 , n68098 , n68103 );
or ( n68106 , n68101 , n68104 , n68105 );
and ( n68107 , n68096 , n68106 );
xor ( n68108 , n67602 , n67612 );
xor ( n68109 , n68108 , n67615 );
xor ( n68110 , n67627 , n67629 );
xor ( n68111 , n68110 , n67632 );
and ( n68112 , n68109 , n68111 );
xor ( n68113 , n67637 , n67639 );
xor ( n68114 , n68113 , n67642 );
and ( n68115 , n68111 , n68114 );
and ( n68116 , n68109 , n68114 );
or ( n68117 , n68112 , n68115 , n68116 );
and ( n68118 , n68106 , n68117 );
and ( n68119 , n68096 , n68117 );
or ( n68120 , n68107 , n68118 , n68119 );
and ( n68121 , n68046 , n68120 );
xor ( n68122 , n67301 , n67303 );
xor ( n68123 , n68122 , n67313 );
xor ( n68124 , n67367 , n67591 );
xor ( n68125 , n68124 , n67618 );
and ( n68126 , n68123 , n68125 );
xor ( n68127 , n67635 , n67645 );
xor ( n68128 , n68127 , n67648 );
and ( n68129 , n68125 , n68128 );
and ( n68130 , n68123 , n68128 );
or ( n68131 , n68126 , n68129 , n68130 );
and ( n68132 , n68120 , n68131 );
and ( n68133 , n68046 , n68131 );
or ( n68134 , n68121 , n68132 , n68133 );
and ( n68135 , n67708 , n68134 );
xor ( n68136 , n67299 , n67316 );
xor ( n68137 , n68136 , n67621 );
xor ( n68138 , n67651 , n67661 );
xor ( n68139 , n68138 , n67664 );
and ( n68140 , n68137 , n68139 );
xor ( n68141 , n67673 , n67675 );
xor ( n68142 , n68141 , n67678 );
and ( n68143 , n68139 , n68142 );
and ( n68144 , n68137 , n68142 );
or ( n68145 , n68140 , n68143 , n68144 );
and ( n68146 , n68134 , n68145 );
and ( n68147 , n67708 , n68145 );
or ( n68148 , n68135 , n68146 , n68147 );
and ( n68149 , n67705 , n68148 );
and ( n68150 , n67703 , n68148 );
or ( n68151 , n67706 , n68149 , n68150 );
and ( n68152 , n67701 , n68151 );
xor ( n68153 , n67290 , n67292 );
xor ( n68154 , n68153 , n67692 );
and ( n68155 , n68151 , n68154 );
and ( n68156 , n67701 , n68154 );
or ( n68157 , n68152 , n68155 , n68156 );
xor ( n68158 , n66953 , n66955 );
xor ( n68159 , n68158 , n67695 );
or ( n68160 , n68157 , n68159 );
and ( n68161 , n67698 , n68160 );
and ( n68162 , n66844 , n68160 );
or ( n68163 , n67699 , n68161 , n68162 );
or ( n68164 , n66842 , n68163 );
and ( n68165 , n66839 , n68164 );
and ( n68166 , n66837 , n68164 );
or ( n68167 , n66840 , n68165 , n68166 );
and ( n68168 , n66385 , n68167 );
xor ( n68169 , n66385 , n68167 );
xor ( n68170 , n66837 , n66839 );
xor ( n68171 , n68170 , n68164 );
not ( n68172 , n68171 );
xnor ( n68173 , n66842 , n68163 );
xor ( n68174 , n66844 , n67698 );
xor ( n68175 , n68174 , n68160 );
not ( n68176 , n68175 );
xnor ( n68177 , n68157 , n68159 );
xor ( n68178 , n67295 , n67670 );
xor ( n68179 , n68178 , n67689 );
xor ( n68180 , n67297 , n67624 );
xor ( n68181 , n68180 , n67667 );
xor ( n68182 , n67681 , n67683 );
xor ( n68183 , n68182 , n67686 );
and ( n68184 , n68181 , n68183 );
xor ( n68185 , n67653 , n67655 );
xor ( n68186 , n68185 , n67658 );
xor ( n68187 , n67319 , n67321 );
xor ( n68188 , n68187 , n67324 );
xor ( n68189 , n67724 , n67749 );
xor ( n68190 , n68189 , n67752 );
or ( n68191 , n68188 , n68190 );
xor ( n68192 , n67735 , n67743 );
xor ( n68193 , n68192 , n67746 );
xnor ( n68194 , n67764 , n67766 );
and ( n68195 , n68193 , n68194 );
xor ( n68196 , n67727 , n67729 );
xor ( n68197 , n68196 , n67732 );
xor ( n68198 , n67413 , n67415 );
xor ( n68199 , n68198 , n67418 );
and ( n68200 , n68197 , n68199 );
xor ( n68201 , n67714 , n67737 );
xor ( n68202 , n68201 , n67740 );
and ( n68203 , n68199 , n68202 );
and ( n68204 , n68197 , n68202 );
or ( n68205 , n68200 , n68203 , n68204 );
and ( n68206 , n68194 , n68205 );
and ( n68207 , n68193 , n68205 );
or ( n68208 , n68195 , n68206 , n68207 );
xor ( n68209 , n67534 , n67538 );
xor ( n68210 , n68209 , n67542 );
xor ( n68211 , n67556 , n67558 );
xor ( n68212 , n68211 , n67561 );
and ( n68213 , n68210 , n68212 );
xor ( n68214 , n67756 , n67758 );
xor ( n68215 , n68214 , n67761 );
and ( n68216 , n68212 , n68215 );
and ( n68217 , n68210 , n68215 );
or ( n68218 , n68213 , n68216 , n68217 );
and ( n68219 , n58915 , n67013 );
not ( n68220 , n68219 );
and ( n68221 , n61918 , n63766 );
not ( n68222 , n68221 );
and ( n68223 , n68220 , n68222 );
and ( n68224 , n62593 , n62998 );
not ( n68225 , n68224 );
and ( n68226 , n68222 , n68225 );
and ( n68227 , n68220 , n68225 );
or ( n68228 , n68223 , n68226 , n68227 );
and ( n68229 , n59365 , n66469 );
not ( n68230 , n68229 );
and ( n68231 , n68228 , n68230 );
and ( n68232 , n60821 , n64811 );
not ( n68233 , n68232 );
and ( n68234 , n68230 , n68233 );
and ( n68235 , n68228 , n68233 );
or ( n68236 , n68231 , n68234 , n68235 );
and ( n68237 , n67997 , n58444 );
not ( n68238 , n68237 );
and ( n68239 , n65606 , n60372 );
not ( n68240 , n68239 );
and ( n68241 , n68238 , n68240 );
and ( n68242 , n63987 , n61914 );
not ( n68243 , n68242 );
and ( n68244 , n68240 , n68243 );
and ( n68245 , n68238 , n68243 );
or ( n68246 , n68241 , n68244 , n68245 );
and ( n68247 , n65678 , n59611 );
not ( n68248 , n68247 );
and ( n68249 , n68246 , n68248 );
xor ( n68250 , n67862 , n67864 );
xor ( n68251 , n68250 , n67867 );
and ( n68252 , n68248 , n68251 );
and ( n68253 , n68246 , n68251 );
or ( n68254 , n68249 , n68252 , n68253 );
and ( n68255 , n68236 , n68254 );
and ( n68256 , n63492 , n61914 );
not ( n68257 , n68256 );
xnor ( n68258 , n67885 , n67889 );
and ( n68259 , n68257 , n68258 );
buf ( n68260 , n68259 );
and ( n68261 , n68254 , n68260 );
and ( n68262 , n68236 , n68260 );
or ( n68263 , n68255 , n68261 , n68262 );
and ( n68264 , n68218 , n68263 );
xor ( n68265 , n67897 , n67901 );
and ( n68266 , n59615 , n66469 );
not ( n68267 , n68266 );
and ( n68268 , n61008 , n64811 );
not ( n68269 , n68268 );
and ( n68270 , n68267 , n68269 );
and ( n68271 , n61505 , n64412 );
not ( n68272 , n68271 );
and ( n68273 , n68269 , n68272 );
and ( n68274 , n68267 , n68272 );
or ( n68275 , n68270 , n68273 , n68274 );
and ( n68276 , n68265 , n68275 );
and ( n68277 , n58292 , n67844 );
not ( n68278 , n68277 );
and ( n68279 , n58628 , n67411 );
not ( n68280 , n68279 );
and ( n68281 , n68278 , n68280 );
and ( n68282 , n60376 , n65586 );
not ( n68283 , n68282 );
and ( n68284 , n68280 , n68283 );
and ( n68285 , n68278 , n68283 );
or ( n68286 , n68281 , n68284 , n68285 );
and ( n68287 , n68275 , n68286 );
and ( n68288 , n68265 , n68286 );
or ( n68289 , n68276 , n68287 , n68288 );
and ( n68290 , n66415 , n59611 );
not ( n68291 , n68290 );
and ( n68292 , n59908 , n66005 );
not ( n68293 , n68292 );
and ( n68294 , n68291 , n68293 );
and ( n68295 , n63492 , n62151 );
not ( n68296 , n68295 );
and ( n68297 , n68293 , n68296 );
and ( n68298 , n68291 , n68296 );
or ( n68299 , n68294 , n68297 , n68298 );
and ( n68300 , n66980 , n58911 );
not ( n68301 , n68300 );
and ( n68302 , n63024 , n62868 );
not ( n68303 , n68302 );
or ( n68304 , n68301 , n68303 );
and ( n68305 , n68299 , n68304 );
buf ( n68306 , n20273 );
buf ( n68307 , n68306 );
and ( n68308 , n68307 , n58294 );
not ( n68309 , n68308 );
and ( n68310 , n67343 , n58542 );
not ( n68311 , n68310 );
and ( n68312 , n68309 , n68311 );
and ( n68313 , n68304 , n68312 );
and ( n68314 , n68299 , n68312 );
or ( n68315 , n68305 , n68313 , n68314 );
and ( n68316 , n68289 , n68315 );
and ( n68317 , n48384 , n57187 );
and ( n68318 , n48272 , n57184 );
nor ( n68319 , n68317 , n68318 );
xnor ( n68320 , n68319 , n56175 );
and ( n68321 , n48709 , n56503 );
and ( n68322 , n48632 , n56501 );
nor ( n68323 , n68321 , n68322 );
xnor ( n68324 , n68323 , n56178 );
and ( n68325 , n68320 , n68324 );
and ( n68326 , n49115 , n55851 );
and ( n68327 , n48988 , n55849 );
nor ( n68328 , n68326 , n68327 );
xnor ( n68329 , n68328 , n55506 );
and ( n68330 , n68324 , n68329 );
and ( n68331 , n68320 , n68329 );
or ( n68332 , n68325 , n68330 , n68331 );
and ( n68333 , n49570 , n55159 );
and ( n68334 , n49374 , n55157 );
nor ( n68335 , n68333 , n68334 );
xnor ( n68336 , n68335 , n54864 );
and ( n68337 , n49976 , n54535 );
and ( n68338 , n49781 , n54533 );
nor ( n68339 , n68337 , n68338 );
xnor ( n68340 , n68339 , n54237 );
and ( n68341 , n68336 , n68340 );
and ( n68342 , n50404 , n53928 );
and ( n68343 , n50195 , n53926 );
nor ( n68344 , n68342 , n68343 );
xnor ( n68345 , n68344 , n53652 );
and ( n68346 , n68340 , n68345 );
and ( n68347 , n68336 , n68345 );
or ( n68348 , n68341 , n68346 , n68347 );
and ( n68349 , n68332 , n68348 );
and ( n68350 , n50726 , n53357 );
and ( n68351 , n50625 , n53355 );
nor ( n68352 , n68350 , n68351 );
xnor ( n68353 , n68352 , n53060 );
and ( n68354 , n51298 , n52799 );
and ( n68355 , n51077 , n52797 );
nor ( n68356 , n68354 , n68355 );
xnor ( n68357 , n68356 , n52538 );
and ( n68358 , n68353 , n68357 );
and ( n68359 , n51734 , n52269 );
and ( n68360 , n51510 , n52267 );
nor ( n68361 , n68359 , n68360 );
xnor ( n68362 , n68361 , n52008 );
and ( n68363 , n68357 , n68362 );
and ( n68364 , n68353 , n68362 );
or ( n68365 , n68358 , n68363 , n68364 );
and ( n68366 , n68348 , n68365 );
and ( n68367 , n68332 , n68365 );
or ( n68368 , n68349 , n68366 , n68367 );
and ( n68369 , n68315 , n68368 );
and ( n68370 , n68289 , n68368 );
or ( n68371 , n68316 , n68369 , n68370 );
and ( n68372 , n68263 , n68371 );
and ( n68373 , n68218 , n68371 );
or ( n68374 , n68264 , n68372 , n68373 );
and ( n68375 , n68208 , n68374 );
and ( n68376 , n52332 , n51750 );
and ( n68377 , n52082 , n51748 );
nor ( n68378 , n68376 , n68377 );
xnor ( n68379 , n68378 , n51520 );
and ( n68380 , n52790 , n51221 );
and ( n68381 , n52612 , n51219 );
nor ( n68382 , n68380 , n68381 );
xnor ( n68383 , n68382 , n51000 );
and ( n68384 , n68379 , n68383 );
and ( n68385 , n53328 , n50783 );
and ( n68386 , n53041 , n50781 );
nor ( n68387 , n68385 , n68386 );
xnor ( n68388 , n68387 , n50557 );
and ( n68389 , n68383 , n68388 );
and ( n68390 , n68379 , n68388 );
or ( n68391 , n68384 , n68389 , n68390 );
and ( n68392 , n53922 , n50338 );
and ( n68393 , n53639 , n50336 );
nor ( n68394 , n68392 , n68393 );
xnor ( n68395 , n68394 , n50111 );
and ( n68396 , n54604 , n49896 );
and ( n68397 , n54227 , n49894 );
nor ( n68398 , n68396 , n68397 );
xnor ( n68399 , n68398 , n49711 );
and ( n68400 , n68395 , n68399 );
and ( n68401 , n55143 , n49513 );
and ( n68402 , n54942 , n49511 );
nor ( n68403 , n68401 , n68402 );
xnor ( n68404 , n68403 , n49310 );
and ( n68405 , n68399 , n68404 );
and ( n68406 , n68395 , n68404 );
or ( n68407 , n68400 , n68405 , n68406 );
and ( n68408 , n68391 , n68407 );
and ( n68409 , n55756 , n49121 );
and ( n68410 , n55497 , n49119 );
nor ( n68411 , n68409 , n68410 );
xnor ( n68412 , n68411 , n48932 );
and ( n68413 , n56388 , n48740 );
and ( n68414 , n56255 , n48738 );
nor ( n68415 , n68413 , n68414 );
xnor ( n68416 , n68415 , n48571 );
and ( n68417 , n68412 , n68416 );
and ( n68418 , n57063 , n48394 );
and ( n68419 , n56915 , n48392 );
nor ( n68420 , n68418 , n68419 );
xnor ( n68421 , n68420 , n48220 );
and ( n68422 , n68416 , n68421 );
and ( n68423 , n68412 , n68421 );
or ( n68424 , n68417 , n68422 , n68423 );
and ( n68425 , n68407 , n68424 );
and ( n68426 , n68391 , n68424 );
or ( n68427 , n68408 , n68425 , n68426 );
and ( n68428 , n57063 , n48392 );
not ( n68429 , n68428 );
and ( n68430 , n68429 , n48220 );
xor ( n68431 , n42770 , n45540 );
buf ( n68432 , n68431 );
buf ( n68433 , n68432 );
buf ( n68434 , n68433 );
and ( n68435 , n68430 , n68434 );
and ( n68436 , n66720 , n59207 );
not ( n68437 , n68436 );
and ( n68438 , n68434 , n68437 );
and ( n68439 , n68430 , n68437 );
or ( n68440 , n68435 , n68438 , n68439 );
and ( n68441 , n65678 , n59920 );
not ( n68442 , n68441 );
and ( n68443 , n65177 , n60711 );
not ( n68444 , n68443 );
and ( n68445 , n68442 , n68444 );
buf ( n68446 , n68445 );
and ( n68447 , n68440 , n68446 );
xor ( n68448 , n67906 , n67910 );
xor ( n68449 , n68448 , n67915 );
and ( n68450 , n68446 , n68449 );
and ( n68451 , n68440 , n68449 );
or ( n68452 , n68447 , n68450 , n68451 );
and ( n68453 , n68427 , n68452 );
xor ( n68454 , n67923 , n67927 );
xor ( n68455 , n68454 , n67932 );
xor ( n68456 , n67943 , n67947 );
xor ( n68457 , n68456 , n67952 );
and ( n68458 , n68455 , n68457 );
xor ( n68459 , n67959 , n67963 );
xor ( n68460 , n68459 , n67968 );
and ( n68461 , n68457 , n68460 );
and ( n68462 , n68455 , n68460 );
or ( n68463 , n68458 , n68461 , n68462 );
and ( n68464 , n68452 , n68463 );
and ( n68465 , n68427 , n68463 );
or ( n68466 , n68453 , n68464 , n68465 );
xor ( n68467 , n67976 , n67980 );
xor ( n68468 , n68467 , n67540 );
xor ( n68469 , n67995 , n67999 );
xor ( n68470 , n68469 , n68002 );
and ( n68471 , n68468 , n68470 );
xor ( n68472 , n68007 , n68009 );
xor ( n68473 , n68472 , n68012 );
and ( n68474 , n68470 , n68473 );
and ( n68475 , n68468 , n68473 );
or ( n68476 , n68471 , n68474 , n68475 );
buf ( n68477 , n67824 );
xor ( n68478 , n68477 , n67826 );
and ( n68479 , n68476 , n68478 );
xor ( n68480 , n67830 , n67832 );
xor ( n68481 , n68480 , n67835 );
and ( n68482 , n68478 , n68481 );
and ( n68483 , n68476 , n68481 );
or ( n68484 , n68479 , n68482 , n68483 );
and ( n68485 , n68466 , n68484 );
xor ( n68486 , n67840 , n67841 );
xor ( n68487 , n68486 , n67854 );
xor ( n68488 , n67870 , n67880 );
xor ( n68489 , n68488 , n67890 );
and ( n68490 , n68487 , n68489 );
xor ( n68491 , n67902 , n67918 );
xor ( n68492 , n68491 , n67935 );
and ( n68493 , n68489 , n68492 );
and ( n68494 , n68487 , n68492 );
or ( n68495 , n68490 , n68493 , n68494 );
and ( n68496 , n68484 , n68495 );
and ( n68497 , n68466 , n68495 );
or ( n68498 , n68485 , n68496 , n68497 );
and ( n68499 , n68374 , n68498 );
and ( n68500 , n68208 , n68498 );
or ( n68501 , n68375 , n68499 , n68500 );
and ( n68502 , n68191 , n68501 );
xor ( n68503 , n67955 , n67971 );
xor ( n68504 , n68503 , n67984 );
xor ( n68505 , n68005 , n68015 );
xor ( n68506 , n68505 , n68018 );
and ( n68507 , n68504 , n68506 );
xor ( n68508 , n68023 , n68025 );
xor ( n68509 , n68508 , n68028 );
and ( n68510 , n68506 , n68509 );
and ( n68511 , n68504 , n68509 );
or ( n68512 , n68507 , n68510 , n68511 );
xor ( n68513 , n67769 , n67771 );
xor ( n68514 , n68513 , n67774 );
and ( n68515 , n68512 , n68514 );
xor ( n68516 , n67780 , n67782 );
xor ( n68517 , n68516 , n67815 );
and ( n68518 , n68514 , n68517 );
and ( n68519 , n68512 , n68517 );
or ( n68520 , n68515 , n68518 , n68519 );
xor ( n68521 , n67828 , n67838 );
xor ( n68522 , n68521 , n67857 );
xor ( n68523 , n67893 , n67938 );
xor ( n68524 , n68523 , n67987 );
and ( n68525 , n68522 , n68524 );
xor ( n68526 , n68021 , n68031 );
xor ( n68527 , n68526 , n68034 );
and ( n68528 , n68524 , n68527 );
and ( n68529 , n68522 , n68527 );
or ( n68530 , n68525 , n68528 , n68529 );
and ( n68531 , n68520 , n68530 );
xor ( n68532 , n67767 , n67777 );
xor ( n68533 , n68532 , n67818 );
and ( n68534 , n68530 , n68533 );
and ( n68535 , n68520 , n68533 );
or ( n68536 , n68531 , n68534 , n68535 );
and ( n68537 , n68501 , n68536 );
and ( n68538 , n68191 , n68536 );
or ( n68539 , n68502 , n68537 , n68538 );
and ( n68540 , n68186 , n68539 );
xor ( n68541 , n67860 , n67990 );
xor ( n68542 , n68541 , n68037 );
xor ( n68543 , n68056 , n68066 );
xor ( n68544 , n68543 , n68069 );
and ( n68545 , n68542 , n68544 );
xor ( n68546 , n68074 , n68076 );
xor ( n68547 , n68546 , n68079 );
and ( n68548 , n68544 , n68547 );
and ( n68549 , n68542 , n68547 );
or ( n68550 , n68545 , n68548 , n68549 );
xor ( n68551 , n67755 , n67821 );
xor ( n68552 , n68551 , n68040 );
and ( n68553 , n68550 , n68552 );
xor ( n68554 , n68072 , n68082 );
xor ( n68555 , n68554 , n68093 );
and ( n68556 , n68552 , n68555 );
and ( n68557 , n68550 , n68555 );
or ( n68558 , n68553 , n68556 , n68557 );
and ( n68559 , n68539 , n68558 );
and ( n68560 , n68186 , n68558 );
or ( n68561 , n68540 , n68559 , n68560 );
xor ( n68562 , n67710 , n67712 );
xor ( n68563 , n68562 , n68043 );
xor ( n68564 , n68096 , n68106 );
xor ( n68565 , n68564 , n68117 );
and ( n68566 , n68563 , n68565 );
xor ( n68567 , n68123 , n68125 );
xor ( n68568 , n68567 , n68128 );
and ( n68569 , n68565 , n68568 );
and ( n68570 , n68563 , n68568 );
or ( n68571 , n68566 , n68569 , n68570 );
and ( n68572 , n68561 , n68571 );
xor ( n68573 , n68046 , n68120 );
xor ( n68574 , n68573 , n68131 );
and ( n68575 , n68571 , n68574 );
and ( n68576 , n68561 , n68574 );
or ( n68577 , n68572 , n68575 , n68576 );
and ( n68578 , n68183 , n68577 );
and ( n68579 , n68181 , n68577 );
or ( n68580 , n68184 , n68578 , n68579 );
and ( n68581 , n68179 , n68580 );
xor ( n68582 , n67703 , n67705 );
xor ( n68583 , n68582 , n68148 );
and ( n68584 , n68580 , n68583 );
and ( n68585 , n68179 , n68583 );
or ( n68586 , n68581 , n68584 , n68585 );
xor ( n68587 , n67701 , n68151 );
xor ( n68588 , n68587 , n68154 );
and ( n68589 , n68586 , n68588 );
xor ( n68590 , n68586 , n68588 );
xor ( n68591 , n67708 , n68134 );
xor ( n68592 , n68591 , n68145 );
xor ( n68593 , n68137 , n68139 );
xor ( n68594 , n68593 , n68142 );
xor ( n68595 , n68098 , n68100 );
xor ( n68596 , n68595 , n68103 );
xor ( n68597 , n68109 , n68111 );
xor ( n68598 , n68597 , n68114 );
and ( n68599 , n68596 , n68598 );
xor ( n68600 , n68085 , n68087 );
xor ( n68601 , n68600 , n68090 );
xnor ( n68602 , n68188 , n68190 );
and ( n68603 , n68601 , n68602 );
xor ( n68604 , n68048 , n68050 );
xor ( n68605 , n68604 , n68053 );
xor ( n68606 , n68058 , n68060 );
xor ( n68607 , n68606 , n68063 );
and ( n68608 , n68605 , n68607 );
buf ( n68609 , n20273 );
buf ( n68610 , n68609 );
and ( n68611 , n57948 , n68610 );
not ( n68612 , n68611 );
and ( n68613 , n59365 , n66917 );
not ( n68614 , n68613 );
and ( n68615 , n68612 , n68614 );
and ( n68616 , n62377 , n63679 );
not ( n68617 , n68616 );
and ( n68618 , n68614 , n68617 );
and ( n68619 , n68612 , n68617 );
or ( n68620 , n68615 , n68618 , n68619 );
xor ( n68621 , n67785 , n67787 );
xor ( n68622 , n68621 , n67790 );
and ( n68623 , n68620 , n68622 );
xor ( n68624 , n67846 , n67848 );
xor ( n68625 , n68624 , n67851 );
and ( n68626 , n68622 , n68625 );
and ( n68627 , n68620 , n68625 );
or ( n68628 , n68623 , n68626 , n68627 );
xor ( n68629 , n67795 , n67797 );
xor ( n68630 , n68629 , n67800 );
xor ( n68631 , n68228 , n68230 );
xor ( n68632 , n68631 , n68233 );
and ( n68633 , n68630 , n68632 );
xor ( n68634 , n67725 , n67806 );
xor ( n68635 , n68634 , n67809 );
and ( n68636 , n68632 , n68635 );
and ( n68637 , n68630 , n68635 );
or ( n68638 , n68633 , n68636 , n68637 );
and ( n68639 , n68628 , n68638 );
xor ( n68640 , n67793 , n67803 );
xor ( n68641 , n68640 , n67812 );
and ( n68642 , n68638 , n68641 );
and ( n68643 , n68628 , n68641 );
or ( n68644 , n68639 , n68642 , n68643 );
and ( n68645 , n68607 , n68644 );
and ( n68646 , n68605 , n68644 );
or ( n68647 , n68608 , n68645 , n68646 );
and ( n68648 , n68602 , n68647 );
and ( n68649 , n68601 , n68647 );
or ( n68650 , n68603 , n68648 , n68649 );
and ( n68651 , n68598 , n68650 );
and ( n68652 , n68596 , n68650 );
or ( n68653 , n68599 , n68651 , n68652 );
xor ( n68654 , n68197 , n68199 );
xor ( n68655 , n68654 , n68202 );
and ( n68656 , n67997 , n58542 );
not ( n68657 , n68656 );
and ( n68658 , n58915 , n67411 );
not ( n68659 , n68658 );
and ( n68660 , n68657 , n68659 );
and ( n68661 , n64221 , n61914 );
not ( n68662 , n68661 );
and ( n68663 , n68659 , n68662 );
and ( n68664 , n68657 , n68662 );
or ( n68665 , n68660 , n68663 , n68664 );
and ( n68666 , n64548 , n61015 );
not ( n68667 , n68666 );
and ( n68668 , n68665 , n68667 );
and ( n68669 , n64221 , n61481 );
not ( n68670 , n68669 );
and ( n68671 , n68667 , n68670 );
and ( n68672 , n68665 , n68670 );
or ( n68673 , n68668 , n68671 , n68672 );
xor ( n68674 , n67872 , n67874 );
xor ( n68675 , n68674 , n67877 );
and ( n68676 , n68673 , n68675 );
and ( n68677 , n68655 , n68676 );
xor ( n68678 , n68246 , n68248 );
xor ( n68679 , n68678 , n68251 );
and ( n68680 , n60376 , n66005 );
not ( n68681 , n68680 );
and ( n68682 , n61505 , n64811 );
not ( n68683 , n68682 );
and ( n68684 , n68681 , n68683 );
and ( n68685 , n61918 , n64412 );
not ( n68686 , n68685 );
and ( n68687 , n68683 , n68686 );
and ( n68688 , n68681 , n68686 );
or ( n68689 , n68684 , n68687 , n68688 );
and ( n68690 , n58292 , n68610 );
not ( n68691 , n68690 );
and ( n68692 , n58628 , n67844 );
not ( n68693 , n68692 );
and ( n68694 , n68691 , n68693 );
and ( n68695 , n62593 , n63679 );
not ( n68696 , n68695 );
and ( n68697 , n68693 , n68696 );
and ( n68698 , n68691 , n68696 );
or ( n68699 , n68694 , n68697 , n68698 );
and ( n68700 , n68689 , n68699 );
and ( n68701 , n60821 , n65210 );
not ( n68702 , n68701 );
and ( n68703 , n68699 , n68702 );
and ( n68704 , n68689 , n68702 );
or ( n68705 , n68700 , n68703 , n68704 );
and ( n68706 , n68679 , n68705 );
and ( n68707 , n59615 , n66917 );
not ( n68708 , n68707 );
and ( n68709 , n59908 , n66469 );
not ( n68710 , n68709 );
and ( n68711 , n68708 , n68710 );
buf ( n68712 , n63024 );
not ( n68713 , n68712 );
and ( n68714 , n68710 , n68713 );
and ( n68715 , n68708 , n68713 );
or ( n68716 , n68711 , n68714 , n68715 );
and ( n68717 , n67343 , n58911 );
and ( n68718 , n65177 , n61015 );
not ( n68719 , n68718 );
and ( n68720 , n68717 , n68719 );
and ( n68721 , n62377 , n63766 );
not ( n68722 , n68721 );
and ( n68723 , n68719 , n68722 );
and ( n68724 , n68717 , n68722 );
or ( n68725 , n68720 , n68723 , n68724 );
and ( n68726 , n68716 , n68725 );
xor ( n68727 , n68278 , n68280 );
xor ( n68728 , n68727 , n68283 );
and ( n68729 , n68725 , n68728 );
and ( n68730 , n68716 , n68728 );
or ( n68731 , n68726 , n68729 , n68730 );
and ( n68732 , n68705 , n68731 );
and ( n68733 , n68679 , n68731 );
or ( n68734 , n68706 , n68732 , n68733 );
and ( n68735 , n68676 , n68734 );
and ( n68736 , n68655 , n68734 );
or ( n68737 , n68677 , n68735 , n68736 );
xor ( n68738 , n68267 , n68269 );
xor ( n68739 , n68738 , n68272 );
xor ( n68740 , n68238 , n68240 );
xor ( n68741 , n68740 , n68243 );
and ( n68742 , n68739 , n68741 );
xor ( n68743 , n68291 , n68293 );
xor ( n68744 , n68743 , n68296 );
and ( n68745 , n68741 , n68744 );
and ( n68746 , n68739 , n68744 );
or ( n68747 , n68742 , n68745 , n68746 );
xnor ( n68748 , n68301 , n68303 );
xor ( n68749 , n68309 , n68311 );
and ( n68750 , n68748 , n68749 );
buf ( n68751 , n20276 );
buf ( n68752 , n68751 );
and ( n68753 , n57948 , n68752 );
not ( n68754 , n68753 );
and ( n68755 , n59365 , n67013 );
not ( n68756 , n68755 );
and ( n68757 , n68754 , n68756 );
and ( n68758 , n60821 , n65586 );
not ( n68759 , n68758 );
and ( n68760 , n68756 , n68759 );
and ( n68761 , n68754 , n68759 );
or ( n68762 , n68757 , n68760 , n68761 );
and ( n68763 , n68749 , n68762 );
and ( n68764 , n68748 , n68762 );
or ( n68765 , n68750 , n68763 , n68764 );
and ( n68766 , n68747 , n68765 );
and ( n68767 , n66720 , n59611 );
not ( n68768 , n68767 );
and ( n68769 , n61008 , n65210 );
not ( n68770 , n68769 );
and ( n68771 , n68768 , n68770 );
and ( n68772 , n64548 , n61481 );
not ( n68773 , n68772 );
and ( n68774 , n68770 , n68773 );
and ( n68775 , n68768 , n68773 );
or ( n68776 , n68771 , n68774 , n68775 );
not ( n68777 , n68717 );
buf ( n68778 , n68777 );
and ( n68779 , n68776 , n68778 );
and ( n68780 , n68307 , n58444 );
and ( n68781 , n63492 , n62868 );
not ( n68782 , n68781 );
and ( n68783 , n68780 , n68782 );
and ( n68784 , n68778 , n68783 );
and ( n68785 , n68776 , n68783 );
or ( n68786 , n68779 , n68784 , n68785 );
and ( n68787 , n68765 , n68786 );
and ( n68788 , n68747 , n68786 );
or ( n68789 , n68766 , n68787 , n68788 );
not ( n68790 , n68780 );
buf ( n68791 , n68790 );
and ( n68792 , n48632 , n57187 );
and ( n68793 , n48384 , n57184 );
nor ( n68794 , n68792 , n68793 );
xnor ( n68795 , n68794 , n56175 );
and ( n68796 , n48988 , n56503 );
and ( n68797 , n48709 , n56501 );
nor ( n68798 , n68796 , n68797 );
xnor ( n68799 , n68798 , n56178 );
and ( n68800 , n68795 , n68799 );
and ( n68801 , n49781 , n55159 );
and ( n68802 , n49570 , n55157 );
nor ( n68803 , n68801 , n68802 );
xnor ( n68804 , n68803 , n54864 );
and ( n68805 , n68799 , n68804 );
and ( n68806 , n68795 , n68804 );
or ( n68807 , n68800 , n68805 , n68806 );
and ( n68808 , n68791 , n68807 );
and ( n68809 , n50195 , n54535 );
and ( n68810 , n49976 , n54533 );
nor ( n68811 , n68809 , n68810 );
xnor ( n68812 , n68811 , n54237 );
and ( n68813 , n50625 , n53928 );
and ( n68814 , n50404 , n53926 );
nor ( n68815 , n68813 , n68814 );
xnor ( n68816 , n68815 , n53652 );
and ( n68817 , n68812 , n68816 );
and ( n68818 , n51077 , n53357 );
and ( n68819 , n50726 , n53355 );
nor ( n68820 , n68818 , n68819 );
xnor ( n68821 , n68820 , n53060 );
and ( n68822 , n68816 , n68821 );
and ( n68823 , n68812 , n68821 );
or ( n68824 , n68817 , n68822 , n68823 );
and ( n68825 , n68807 , n68824 );
and ( n68826 , n68791 , n68824 );
or ( n68827 , n68808 , n68825 , n68826 );
and ( n68828 , n51510 , n52799 );
and ( n68829 , n51298 , n52797 );
nor ( n68830 , n68828 , n68829 );
xnor ( n68831 , n68830 , n52538 );
and ( n68832 , n52082 , n52269 );
and ( n68833 , n51734 , n52267 );
nor ( n68834 , n68832 , n68833 );
xnor ( n68835 , n68834 , n52008 );
and ( n68836 , n68831 , n68835 );
and ( n68837 , n52612 , n51750 );
and ( n68838 , n52332 , n51748 );
nor ( n68839 , n68837 , n68838 );
xnor ( n68840 , n68839 , n51520 );
and ( n68841 , n68835 , n68840 );
and ( n68842 , n68831 , n68840 );
or ( n68843 , n68836 , n68841 , n68842 );
and ( n68844 , n53041 , n51221 );
and ( n68845 , n52790 , n51219 );
nor ( n68846 , n68844 , n68845 );
xnor ( n68847 , n68846 , n51000 );
and ( n68848 , n53639 , n50783 );
and ( n68849 , n53328 , n50781 );
nor ( n68850 , n68848 , n68849 );
xnor ( n68851 , n68850 , n50557 );
and ( n68852 , n68847 , n68851 );
and ( n68853 , n54227 , n50338 );
and ( n68854 , n53922 , n50336 );
nor ( n68855 , n68853 , n68854 );
xnor ( n68856 , n68855 , n50111 );
and ( n68857 , n68851 , n68856 );
and ( n68858 , n68847 , n68856 );
or ( n68859 , n68852 , n68857 , n68858 );
and ( n68860 , n68843 , n68859 );
and ( n68861 , n54942 , n49896 );
and ( n68862 , n54604 , n49894 );
nor ( n68863 , n68861 , n68862 );
xnor ( n68864 , n68863 , n49711 );
and ( n68865 , n55497 , n49513 );
and ( n68866 , n55143 , n49511 );
nor ( n68867 , n68865 , n68866 );
xnor ( n68868 , n68867 , n49310 );
and ( n68869 , n68864 , n68868 );
and ( n68870 , n56255 , n49121 );
and ( n68871 , n55756 , n49119 );
nor ( n68872 , n68870 , n68871 );
xnor ( n68873 , n68872 , n48932 );
and ( n68874 , n68868 , n68873 );
and ( n68875 , n68864 , n68873 );
or ( n68876 , n68869 , n68874 , n68875 );
and ( n68877 , n68859 , n68876 );
and ( n68878 , n68843 , n68876 );
or ( n68879 , n68860 , n68877 , n68878 );
and ( n68880 , n68827 , n68879 );
and ( n68881 , n56915 , n48740 );
and ( n68882 , n56388 , n48738 );
nor ( n68883 , n68881 , n68882 );
xnor ( n68884 , n68883 , n48571 );
and ( n68885 , n68884 , n68428 );
xor ( n68886 , n42773 , n45538 );
buf ( n68887 , n68886 );
buf ( n68888 , n68887 );
buf ( n68889 , n68888 );
and ( n68890 , n68428 , n68889 );
and ( n68891 , n68884 , n68889 );
or ( n68892 , n68885 , n68890 , n68891 );
and ( n68893 , n66415 , n59920 );
not ( n68894 , n68893 );
and ( n68895 , n65678 , n60372 );
not ( n68896 , n68895 );
and ( n68897 , n68894 , n68896 );
and ( n68898 , n63987 , n62151 );
not ( n68899 , n68898 );
and ( n68900 , n68896 , n68899 );
and ( n68901 , n68894 , n68899 );
or ( n68902 , n68897 , n68900 , n68901 );
and ( n68903 , n68892 , n68902 );
xor ( n68904 , n68320 , n68324 );
xor ( n68905 , n68904 , n68329 );
and ( n68906 , n68902 , n68905 );
and ( n68907 , n68892 , n68905 );
or ( n68908 , n68903 , n68906 , n68907 );
and ( n68909 , n68879 , n68908 );
and ( n68910 , n68827 , n68908 );
or ( n68911 , n68880 , n68909 , n68910 );
and ( n68912 , n68789 , n68911 );
xor ( n68913 , n68336 , n68340 );
xor ( n68914 , n68913 , n68345 );
xor ( n68915 , n68353 , n68357 );
xor ( n68916 , n68915 , n68362 );
and ( n68917 , n68914 , n68916 );
xor ( n68918 , n68379 , n68383 );
xor ( n68919 , n68918 , n68388 );
and ( n68920 , n68916 , n68919 );
and ( n68921 , n68914 , n68919 );
or ( n68922 , n68917 , n68920 , n68921 );
xor ( n68923 , n68395 , n68399 );
xor ( n68924 , n68923 , n68404 );
xor ( n68925 , n68412 , n68416 );
xor ( n68926 , n68925 , n68421 );
and ( n68927 , n68924 , n68926 );
xor ( n68928 , n68430 , n68434 );
xor ( n68929 , n68928 , n68437 );
and ( n68930 , n68926 , n68929 );
and ( n68931 , n68924 , n68929 );
or ( n68932 , n68927 , n68930 , n68931 );
and ( n68933 , n68922 , n68932 );
buf ( n68934 , n68257 );
xor ( n68935 , n68934 , n68258 );
and ( n68936 , n68932 , n68935 );
and ( n68937 , n68922 , n68935 );
or ( n68938 , n68933 , n68936 , n68937 );
and ( n68939 , n68911 , n68938 );
and ( n68940 , n68789 , n68938 );
or ( n68941 , n68912 , n68939 , n68940 );
and ( n68942 , n68737 , n68941 );
xor ( n68943 , n68265 , n68275 );
xor ( n68944 , n68943 , n68286 );
xor ( n68945 , n68299 , n68304 );
xor ( n68946 , n68945 , n68312 );
and ( n68947 , n68944 , n68946 );
xor ( n68948 , n68332 , n68348 );
xor ( n68949 , n68948 , n68365 );
and ( n68950 , n68946 , n68949 );
and ( n68951 , n68944 , n68949 );
or ( n68952 , n68947 , n68950 , n68951 );
xor ( n68953 , n68391 , n68407 );
xor ( n68954 , n68953 , n68424 );
xor ( n68955 , n68440 , n68446 );
xor ( n68956 , n68955 , n68449 );
and ( n68957 , n68954 , n68956 );
xor ( n68958 , n68455 , n68457 );
xor ( n68959 , n68958 , n68460 );
and ( n68960 , n68956 , n68959 );
and ( n68961 , n68954 , n68959 );
or ( n68962 , n68957 , n68960 , n68961 );
and ( n68963 , n68952 , n68962 );
xor ( n68964 , n68210 , n68212 );
xor ( n68965 , n68964 , n68215 );
and ( n68966 , n68962 , n68965 );
and ( n68967 , n68952 , n68965 );
or ( n68968 , n68963 , n68966 , n68967 );
and ( n68969 , n68941 , n68968 );
and ( n68970 , n68737 , n68968 );
or ( n68971 , n68942 , n68969 , n68970 );
xor ( n68972 , n68236 , n68254 );
xor ( n68973 , n68972 , n68260 );
xor ( n68974 , n68289 , n68315 );
xor ( n68975 , n68974 , n68368 );
and ( n68976 , n68973 , n68975 );
xor ( n68977 , n68427 , n68452 );
xor ( n68978 , n68977 , n68463 );
and ( n68979 , n68975 , n68978 );
and ( n68980 , n68973 , n68978 );
or ( n68981 , n68976 , n68979 , n68980 );
xor ( n68982 , n68476 , n68478 );
xor ( n68983 , n68982 , n68481 );
xor ( n68984 , n68487 , n68489 );
xor ( n68985 , n68984 , n68492 );
and ( n68986 , n68983 , n68985 );
xor ( n68987 , n68504 , n68506 );
xor ( n68988 , n68987 , n68509 );
and ( n68989 , n68985 , n68988 );
and ( n68990 , n68983 , n68988 );
or ( n68991 , n68986 , n68989 , n68990 );
and ( n68992 , n68981 , n68991 );
xor ( n68993 , n68193 , n68194 );
xor ( n68994 , n68993 , n68205 );
and ( n68995 , n68991 , n68994 );
and ( n68996 , n68981 , n68994 );
or ( n68997 , n68992 , n68995 , n68996 );
and ( n68998 , n68971 , n68997 );
xor ( n68999 , n68218 , n68263 );
xor ( n69000 , n68999 , n68371 );
xor ( n69001 , n68466 , n68484 );
xor ( n69002 , n69001 , n68495 );
and ( n69003 , n69000 , n69002 );
xor ( n69004 , n68512 , n68514 );
xor ( n69005 , n69004 , n68517 );
and ( n69006 , n69002 , n69005 );
and ( n69007 , n69000 , n69005 );
or ( n69008 , n69003 , n69006 , n69007 );
and ( n69009 , n68997 , n69008 );
and ( n69010 , n68971 , n69008 );
or ( n69011 , n68998 , n69009 , n69010 );
xor ( n69012 , n68208 , n68374 );
xor ( n69013 , n69012 , n68498 );
xor ( n69014 , n68520 , n68530 );
xor ( n69015 , n69014 , n68533 );
and ( n69016 , n69013 , n69015 );
xor ( n69017 , n68542 , n68544 );
xor ( n69018 , n69017 , n68547 );
and ( n69019 , n69015 , n69018 );
and ( n69020 , n69013 , n69018 );
or ( n69021 , n69016 , n69019 , n69020 );
and ( n69022 , n69011 , n69021 );
xor ( n69023 , n68191 , n68501 );
xor ( n69024 , n69023 , n68536 );
and ( n69025 , n69021 , n69024 );
and ( n69026 , n69011 , n69024 );
or ( n69027 , n69022 , n69025 , n69026 );
and ( n69028 , n68653 , n69027 );
xor ( n69029 , n68186 , n68539 );
xor ( n69030 , n69029 , n68558 );
and ( n69031 , n69027 , n69030 );
and ( n69032 , n68653 , n69030 );
or ( n69033 , n69028 , n69031 , n69032 );
and ( n69034 , n68594 , n69033 );
xor ( n69035 , n68561 , n68571 );
xor ( n69036 , n69035 , n68574 );
and ( n69037 , n69033 , n69036 );
and ( n69038 , n68594 , n69036 );
or ( n69039 , n69034 , n69037 , n69038 );
and ( n69040 , n68592 , n69039 );
xor ( n69041 , n68181 , n68183 );
xor ( n69042 , n69041 , n68577 );
and ( n69043 , n69039 , n69042 );
and ( n69044 , n68592 , n69042 );
or ( n69045 , n69040 , n69043 , n69044 );
xor ( n69046 , n68179 , n68580 );
xor ( n69047 , n69046 , n68583 );
and ( n69048 , n69045 , n69047 );
xor ( n69049 , n69045 , n69047 );
xor ( n69050 , n68592 , n69039 );
xor ( n69051 , n69050 , n69042 );
xor ( n69052 , n68563 , n68565 );
xor ( n69053 , n69052 , n68568 );
xor ( n69054 , n68550 , n68552 );
xor ( n69055 , n69054 , n68555 );
xor ( n69056 , n68522 , n68524 );
xor ( n69057 , n69056 , n68527 );
buf ( n69058 , n20276 );
buf ( n69059 , n69058 );
and ( n69060 , n69059 , n58294 );
not ( n69061 , n69060 );
and ( n69062 , n66980 , n59207 );
not ( n69063 , n69062 );
and ( n69064 , n69061 , n69063 );
and ( n69065 , n65606 , n60711 );
not ( n69066 , n69065 );
and ( n69067 , n69063 , n69066 );
and ( n69068 , n69061 , n69066 );
or ( n69069 , n69064 , n69067 , n69068 );
xor ( n69070 , n68220 , n68222 );
xor ( n69071 , n69070 , n68225 );
and ( n69072 , n69069 , n69071 );
xor ( n69073 , n68612 , n68614 );
xor ( n69074 , n69073 , n68617 );
and ( n69075 , n69071 , n69074 );
and ( n69076 , n69069 , n69074 );
or ( n69077 , n69072 , n69075 , n69076 );
xor ( n69078 , n68620 , n68622 );
xor ( n69079 , n69078 , n68625 );
and ( n69080 , n69077 , n69079 );
xor ( n69081 , n68630 , n68632 );
xor ( n69082 , n69081 , n68635 );
and ( n69083 , n69079 , n69082 );
and ( n69084 , n69077 , n69082 );
or ( n69085 , n69080 , n69083 , n69084 );
xor ( n69086 , n68628 , n68638 );
xor ( n69087 , n69086 , n68641 );
or ( n69088 , n69085 , n69087 );
and ( n69089 , n69057 , n69088 );
xor ( n69090 , n68468 , n68470 );
xor ( n69091 , n69090 , n68473 );
xor ( n69092 , n68673 , n68675 );
and ( n69093 , n69091 , n69092 );
xor ( n69094 , n68691 , n68693 );
xor ( n69095 , n69094 , n68696 );
xor ( n69096 , n68708 , n68710 );
xor ( n69097 , n69096 , n68713 );
and ( n69098 , n69095 , n69097 );
xor ( n69099 , n68717 , n68719 );
xor ( n69100 , n69099 , n68722 );
and ( n69101 , n69097 , n69100 );
and ( n69102 , n69095 , n69100 );
or ( n69103 , n69098 , n69101 , n69102 );
xor ( n69104 , n69069 , n69071 );
xor ( n69105 , n69104 , n69074 );
or ( n69106 , n69103 , n69105 );
and ( n69107 , n69092 , n69106 );
and ( n69108 , n69091 , n69106 );
or ( n69109 , n69093 , n69107 , n69108 );
xor ( n69110 , n68442 , n68444 );
buf ( n69111 , n69110 );
xor ( n69112 , n68689 , n68699 );
xor ( n69113 , n69112 , n68702 );
and ( n69114 , n69111 , n69113 );
xor ( n69115 , n68665 , n68667 );
xor ( n69116 , n69115 , n68670 );
and ( n69117 , n69113 , n69116 );
and ( n69118 , n69111 , n69116 );
or ( n69119 , n69114 , n69117 , n69118 );
xor ( n69120 , n68716 , n68725 );
xor ( n69121 , n69120 , n68728 );
and ( n69122 , n58915 , n67844 );
not ( n69123 , n69122 );
and ( n69124 , n60376 , n66469 );
not ( n69125 , n69124 );
and ( n69126 , n69123 , n69125 );
and ( n69127 , n63024 , n63679 );
not ( n69128 , n69127 );
and ( n69129 , n69125 , n69128 );
and ( n69130 , n69123 , n69128 );
or ( n69131 , n69126 , n69129 , n69130 );
and ( n69132 , n58628 , n68610 );
not ( n69133 , n69132 );
and ( n69134 , n61918 , n64811 );
not ( n69135 , n69134 );
and ( n69136 , n69133 , n69135 );
and ( n69137 , n62593 , n63766 );
not ( n69138 , n69137 );
and ( n69139 , n69135 , n69138 );
and ( n69140 , n69133 , n69138 );
or ( n69141 , n69136 , n69139 , n69140 );
or ( n69142 , n69131 , n69141 );
and ( n69143 , n69121 , n69142 );
and ( n69144 , n50726 , n53928 );
and ( n69145 , n50625 , n53926 );
nor ( n69146 , n69144 , n69145 );
xnor ( n69147 , n69146 , n53652 );
and ( n69148 , n51298 , n53357 );
and ( n69149 , n51077 , n53355 );
nor ( n69150 , n69148 , n69149 );
xnor ( n69151 , n69150 , n53060 );
and ( n69152 , n69147 , n69151 );
and ( n69153 , n51734 , n52799 );
and ( n69154 , n51510 , n52797 );
nor ( n69155 , n69153 , n69154 );
xnor ( n69156 , n69155 , n52538 );
and ( n69157 , n69151 , n69156 );
and ( n69158 , n69147 , n69156 );
or ( n69159 , n69152 , n69157 , n69158 );
and ( n69160 , n49374 , n55851 );
and ( n69161 , n49115 , n55849 );
nor ( n69162 , n69160 , n69161 );
xnor ( n69163 , n69162 , n55506 );
and ( n69164 , n69159 , n69163 );
and ( n69165 , n69142 , n69164 );
and ( n69166 , n69121 , n69164 );
or ( n69167 , n69143 , n69165 , n69166 );
and ( n69168 , n69119 , n69167 );
xor ( n69169 , n68754 , n68756 );
xor ( n69170 , n69169 , n68759 );
xor ( n69171 , n68657 , n68659 );
xor ( n69172 , n69171 , n68662 );
and ( n69173 , n69170 , n69172 );
buf ( n69174 , n69173 );
xor ( n69175 , n68768 , n68770 );
xor ( n69176 , n69175 , n68773 );
xor ( n69177 , n68780 , n68782 );
and ( n69178 , n69176 , n69177 );
and ( n69179 , n58292 , n68752 );
not ( n69180 , n69179 );
and ( n69181 , n64548 , n61914 );
not ( n69182 , n69181 );
and ( n69183 , n69180 , n69182 );
and ( n69184 , n63987 , n62868 );
not ( n69185 , n69184 );
and ( n69186 , n69182 , n69185 );
and ( n69187 , n69180 , n69185 );
or ( n69188 , n69183 , n69186 , n69187 );
and ( n69189 , n69177 , n69188 );
and ( n69190 , n69176 , n69188 );
or ( n69191 , n69178 , n69189 , n69190 );
and ( n69192 , n69174 , n69191 );
and ( n69193 , n68307 , n58542 );
not ( n69194 , n69193 );
and ( n69195 , n66415 , n60372 );
not ( n69196 , n69195 );
and ( n69197 , n69194 , n69196 );
and ( n69198 , n65177 , n61481 );
not ( n69199 , n69198 );
and ( n69200 , n69196 , n69199 );
and ( n69201 , n69194 , n69199 );
or ( n69202 , n69197 , n69200 , n69201 );
buf ( n69203 , n20279 );
buf ( n69204 , n69203 );
and ( n69205 , n57948 , n69204 );
not ( n69206 , n69205 );
and ( n69207 , n66980 , n59611 );
not ( n69208 , n69207 );
and ( n69209 , n69206 , n69208 );
and ( n69210 , n66720 , n59920 );
not ( n69211 , n69210 );
and ( n69212 , n69208 , n69211 );
and ( n69213 , n69206 , n69211 );
or ( n69214 , n69209 , n69212 , n69213 );
and ( n69215 , n69202 , n69214 );
and ( n69216 , n49976 , n55159 );
and ( n69217 , n49781 , n55157 );
nor ( n69218 , n69216 , n69217 );
xnor ( n69219 , n69218 , n54864 );
and ( n69220 , n50404 , n54535 );
and ( n69221 , n50195 , n54533 );
nor ( n69222 , n69220 , n69221 );
xnor ( n69223 , n69222 , n54237 );
and ( n69224 , n69219 , n69223 );
and ( n69225 , n69214 , n69224 );
and ( n69226 , n69202 , n69224 );
or ( n69227 , n69215 , n69225 , n69226 );
and ( n69228 , n69191 , n69227 );
and ( n69229 , n69174 , n69227 );
or ( n69230 , n69192 , n69228 , n69229 );
and ( n69231 , n69167 , n69230 );
and ( n69232 , n69119 , n69230 );
or ( n69233 , n69168 , n69231 , n69232 );
and ( n69234 , n69109 , n69233 );
and ( n69235 , n48709 , n57187 );
and ( n69236 , n48632 , n57184 );
nor ( n69237 , n69235 , n69236 );
xnor ( n69238 , n69237 , n56175 );
and ( n69239 , n49570 , n55851 );
and ( n69240 , n49374 , n55849 );
nor ( n69241 , n69239 , n69240 );
xnor ( n69242 , n69241 , n55506 );
and ( n69243 , n69238 , n69242 );
and ( n69244 , n52332 , n52269 );
and ( n69245 , n52082 , n52267 );
nor ( n69246 , n69244 , n69245 );
xnor ( n69247 , n69246 , n52008 );
and ( n69248 , n69242 , n69247 );
and ( n69249 , n69238 , n69247 );
or ( n69250 , n69243 , n69248 , n69249 );
and ( n69251 , n52790 , n51750 );
and ( n69252 , n52612 , n51748 );
nor ( n69253 , n69251 , n69252 );
xnor ( n69254 , n69253 , n51520 );
and ( n69255 , n53922 , n50783 );
and ( n69256 , n53639 , n50781 );
nor ( n69257 , n69255 , n69256 );
xnor ( n69258 , n69257 , n50557 );
and ( n69259 , n69254 , n69258 );
and ( n69260 , n54604 , n50338 );
and ( n69261 , n54227 , n50336 );
nor ( n69262 , n69260 , n69261 );
xnor ( n69263 , n69262 , n50111 );
and ( n69264 , n69258 , n69263 );
and ( n69265 , n69254 , n69263 );
or ( n69266 , n69259 , n69264 , n69265 );
and ( n69267 , n69250 , n69266 );
and ( n69268 , n55143 , n49896 );
and ( n69269 , n54942 , n49894 );
nor ( n69270 , n69268 , n69269 );
xnor ( n69271 , n69270 , n49711 );
and ( n69272 , n55756 , n49513 );
and ( n69273 , n55497 , n49511 );
nor ( n69274 , n69272 , n69273 );
xnor ( n69275 , n69274 , n49310 );
and ( n69276 , n69271 , n69275 );
and ( n69277 , n56388 , n49121 );
and ( n69278 , n56255 , n49119 );
nor ( n69279 , n69277 , n69278 );
xnor ( n69280 , n69279 , n48932 );
and ( n69281 , n69275 , n69280 );
and ( n69282 , n69271 , n69280 );
or ( n69283 , n69276 , n69281 , n69282 );
and ( n69284 , n69266 , n69283 );
and ( n69285 , n69250 , n69283 );
or ( n69286 , n69267 , n69284 , n69285 );
and ( n69287 , n57063 , n48740 );
and ( n69288 , n56915 , n48738 );
nor ( n69289 , n69287 , n69288 );
xnor ( n69290 , n69289 , n48571 );
and ( n69291 , n57063 , n48738 );
not ( n69292 , n69291 );
and ( n69293 , n69292 , n48571 );
and ( n69294 , n69290 , n69293 );
xor ( n69295 , n42776 , n45536 );
buf ( n69296 , n69295 );
buf ( n69297 , n69296 );
buf ( n69298 , n69297 );
and ( n69299 , n69293 , n69298 );
and ( n69300 , n69290 , n69298 );
or ( n69301 , n69294 , n69299 , n69300 );
buf ( n69302 , n20279 );
buf ( n69303 , n69302 );
and ( n69304 , n69303 , n58294 );
not ( n69305 , n69304 );
and ( n69306 , n69059 , n58444 );
not ( n69307 , n69306 );
and ( n69308 , n69305 , n69307 );
and ( n69309 , n67997 , n58911 );
not ( n69310 , n69309 );
and ( n69311 , n69307 , n69310 );
and ( n69312 , n69305 , n69310 );
or ( n69313 , n69308 , n69311 , n69312 );
and ( n69314 , n69301 , n69313 );
and ( n69315 , n65606 , n61015 );
not ( n69316 , n69315 );
and ( n69317 , n63492 , n62998 );
not ( n69318 , n69317 );
and ( n69319 , n69316 , n69318 );
buf ( n69320 , n69319 );
and ( n69321 , n69313 , n69320 );
and ( n69322 , n69301 , n69320 );
or ( n69323 , n69314 , n69321 , n69322 );
and ( n69324 , n69286 , n69323 );
xor ( n69325 , n68795 , n68799 );
xor ( n69326 , n69325 , n68804 );
xor ( n69327 , n68812 , n68816 );
xor ( n69328 , n69327 , n68821 );
and ( n69329 , n69326 , n69328 );
xor ( n69330 , n68831 , n68835 );
xor ( n69331 , n69330 , n68840 );
and ( n69332 , n69328 , n69331 );
and ( n69333 , n69326 , n69331 );
or ( n69334 , n69329 , n69332 , n69333 );
and ( n69335 , n69323 , n69334 );
and ( n69336 , n69286 , n69334 );
or ( n69337 , n69324 , n69335 , n69336 );
xor ( n69338 , n68847 , n68851 );
xor ( n69339 , n69338 , n68856 );
xor ( n69340 , n68864 , n68868 );
xor ( n69341 , n69340 , n68873 );
and ( n69342 , n69339 , n69341 );
xor ( n69343 , n68884 , n68428 );
xor ( n69344 , n69343 , n68889 );
and ( n69345 , n69341 , n69344 );
and ( n69346 , n69339 , n69344 );
or ( n69347 , n69342 , n69345 , n69346 );
xor ( n69348 , n68739 , n68741 );
xor ( n69349 , n69348 , n68744 );
and ( n69350 , n69347 , n69349 );
xor ( n69351 , n68748 , n68749 );
xor ( n69352 , n69351 , n68762 );
and ( n69353 , n69349 , n69352 );
and ( n69354 , n69347 , n69352 );
or ( n69355 , n69350 , n69353 , n69354 );
and ( n69356 , n69337 , n69355 );
xor ( n69357 , n68776 , n68778 );
xor ( n69358 , n69357 , n68783 );
xor ( n69359 , n68791 , n68807 );
xor ( n69360 , n69359 , n68824 );
and ( n69361 , n69358 , n69360 );
xor ( n69362 , n68843 , n68859 );
xor ( n69363 , n69362 , n68876 );
and ( n69364 , n69360 , n69363 );
and ( n69365 , n69358 , n69363 );
or ( n69366 , n69361 , n69364 , n69365 );
and ( n69367 , n69355 , n69366 );
and ( n69368 , n69337 , n69366 );
or ( n69369 , n69356 , n69367 , n69368 );
and ( n69370 , n69233 , n69369 );
and ( n69371 , n69109 , n69369 );
or ( n69372 , n69234 , n69370 , n69371 );
and ( n69373 , n69088 , n69372 );
and ( n69374 , n69057 , n69372 );
or ( n69375 , n69089 , n69373 , n69374 );
xor ( n69376 , n68892 , n68902 );
xor ( n69377 , n69376 , n68905 );
xor ( n69378 , n68914 , n68916 );
xor ( n69379 , n69378 , n68919 );
and ( n69380 , n69377 , n69379 );
xor ( n69381 , n68924 , n68926 );
xor ( n69382 , n69381 , n68929 );
and ( n69383 , n69379 , n69382 );
and ( n69384 , n69377 , n69382 );
or ( n69385 , n69380 , n69383 , n69384 );
xor ( n69386 , n68679 , n68705 );
xor ( n69387 , n69386 , n68731 );
and ( n69388 , n69385 , n69387 );
xor ( n69389 , n68747 , n68765 );
xor ( n69390 , n69389 , n68786 );
and ( n69391 , n69387 , n69390 );
and ( n69392 , n69385 , n69390 );
or ( n69393 , n69388 , n69391 , n69392 );
xor ( n69394 , n68827 , n68879 );
xor ( n69395 , n69394 , n68908 );
xor ( n69396 , n68922 , n68932 );
xor ( n69397 , n69396 , n68935 );
and ( n69398 , n69395 , n69397 );
xor ( n69399 , n68944 , n68946 );
xor ( n69400 , n69399 , n68949 );
and ( n69401 , n69397 , n69400 );
and ( n69402 , n69395 , n69400 );
or ( n69403 , n69398 , n69401 , n69402 );
and ( n69404 , n69393 , n69403 );
xor ( n69405 , n68655 , n68676 );
xor ( n69406 , n69405 , n68734 );
and ( n69407 , n69403 , n69406 );
and ( n69408 , n69393 , n69406 );
or ( n69409 , n69404 , n69407 , n69408 );
xor ( n69410 , n68789 , n68911 );
xor ( n69411 , n69410 , n68938 );
xor ( n69412 , n68952 , n68962 );
xor ( n69413 , n69412 , n68965 );
and ( n69414 , n69411 , n69413 );
xor ( n69415 , n68973 , n68975 );
xor ( n69416 , n69415 , n68978 );
and ( n69417 , n69413 , n69416 );
and ( n69418 , n69411 , n69416 );
or ( n69419 , n69414 , n69417 , n69418 );
and ( n69420 , n69409 , n69419 );
xor ( n69421 , n68605 , n68607 );
xor ( n69422 , n69421 , n68644 );
and ( n69423 , n69419 , n69422 );
and ( n69424 , n69409 , n69422 );
or ( n69425 , n69420 , n69423 , n69424 );
and ( n69426 , n69375 , n69425 );
xor ( n69427 , n68737 , n68941 );
xor ( n69428 , n69427 , n68968 );
xor ( n69429 , n68981 , n68991 );
xor ( n69430 , n69429 , n68994 );
and ( n69431 , n69428 , n69430 );
xor ( n69432 , n69000 , n69002 );
xor ( n69433 , n69432 , n69005 );
and ( n69434 , n69430 , n69433 );
and ( n69435 , n69428 , n69433 );
or ( n69436 , n69431 , n69434 , n69435 );
and ( n69437 , n69425 , n69436 );
and ( n69438 , n69375 , n69436 );
or ( n69439 , n69426 , n69437 , n69438 );
and ( n69440 , n69055 , n69439 );
xor ( n69441 , n68601 , n68602 );
xor ( n69442 , n69441 , n68647 );
xor ( n69443 , n68971 , n68997 );
xor ( n69444 , n69443 , n69008 );
and ( n69445 , n69442 , n69444 );
xor ( n69446 , n69013 , n69015 );
xor ( n69447 , n69446 , n69018 );
and ( n69448 , n69444 , n69447 );
and ( n69449 , n69442 , n69447 );
or ( n69450 , n69445 , n69448 , n69449 );
and ( n69451 , n69439 , n69450 );
and ( n69452 , n69055 , n69450 );
or ( n69453 , n69440 , n69451 , n69452 );
and ( n69454 , n69053 , n69453 );
xor ( n69455 , n68653 , n69027 );
xor ( n69456 , n69455 , n69030 );
and ( n69457 , n69453 , n69456 );
and ( n69458 , n69053 , n69456 );
or ( n69459 , n69454 , n69457 , n69458 );
xor ( n69460 , n68594 , n69033 );
xor ( n69461 , n69460 , n69036 );
and ( n69462 , n69459 , n69461 );
xor ( n69463 , n68596 , n68598 );
xor ( n69464 , n69463 , n68650 );
xor ( n69465 , n69011 , n69021 );
xor ( n69466 , n69465 , n69024 );
and ( n69467 , n69464 , n69466 );
xor ( n69468 , n68983 , n68985 );
xor ( n69469 , n69468 , n68988 );
xnor ( n69470 , n69085 , n69087 );
and ( n69471 , n69469 , n69470 );
xor ( n69472 , n68954 , n68956 );
xor ( n69473 , n69472 , n68959 );
xor ( n69474 , n69077 , n69079 );
xor ( n69475 , n69474 , n69082 );
and ( n69476 , n69473 , n69475 );
xnor ( n69477 , n69103 , n69105 );
and ( n69478 , n58915 , n68610 );
not ( n69479 , n69478 );
buf ( n69480 , n69479 );
and ( n69481 , n59908 , n66917 );
not ( n69482 , n69481 );
and ( n69483 , n69480 , n69482 );
and ( n69484 , n62377 , n64412 );
not ( n69485 , n69484 );
and ( n69486 , n69482 , n69485 );
and ( n69487 , n69480 , n69485 );
or ( n69488 , n69483 , n69486 , n69487 );
and ( n69489 , n59615 , n67013 );
not ( n69490 , n69489 );
and ( n69491 , n61008 , n65586 );
not ( n69492 , n69491 );
and ( n69493 , n69490 , n69492 );
and ( n69494 , n61505 , n65210 );
not ( n69495 , n69494 );
and ( n69496 , n69492 , n69495 );
and ( n69497 , n69490 , n69495 );
or ( n69498 , n69493 , n69496 , n69497 );
and ( n69499 , n69488 , n69498 );
xor ( n69500 , n68681 , n68683 );
xor ( n69501 , n69500 , n68686 );
and ( n69502 , n69498 , n69501 );
and ( n69503 , n69488 , n69501 );
or ( n69504 , n69499 , n69502 , n69503 );
and ( n69505 , n69477 , n69504 );
buf ( n69506 , n10629 );
buf ( n69507 , n69506 );
and ( n69508 , n57948 , n69507 );
not ( n69509 , n69508 );
and ( n69510 , n59365 , n67844 );
not ( n69511 , n69510 );
and ( n69512 , n69509 , n69511 );
and ( n69513 , n62377 , n64811 );
not ( n69514 , n69513 );
and ( n69515 , n69511 , n69514 );
and ( n69516 , n69509 , n69514 );
or ( n69517 , n69512 , n69515 , n69516 );
xor ( n69518 , n69123 , n69125 );
xor ( n69519 , n69518 , n69128 );
and ( n69520 , n69517 , n69519 );
xor ( n69521 , n69133 , n69135 );
xor ( n69522 , n69521 , n69138 );
and ( n69523 , n69519 , n69522 );
and ( n69524 , n69517 , n69522 );
or ( n69525 , n69520 , n69523 , n69524 );
xor ( n69526 , n69095 , n69097 );
xor ( n69527 , n69526 , n69100 );
or ( n69528 , n69525 , n69527 );
and ( n69529 , n69504 , n69528 );
and ( n69530 , n69477 , n69528 );
or ( n69531 , n69505 , n69529 , n69530 );
and ( n69532 , n69475 , n69531 );
and ( n69533 , n69473 , n69531 );
or ( n69534 , n69476 , n69532 , n69533 );
and ( n69535 , n69470 , n69534 );
and ( n69536 , n69469 , n69534 );
or ( n69537 , n69471 , n69535 , n69536 );
and ( n69538 , n60376 , n66917 );
not ( n69539 , n69538 );
and ( n69540 , n61918 , n65210 );
not ( n69541 , n69540 );
and ( n69542 , n69539 , n69541 );
and ( n69543 , n62593 , n64412 );
not ( n69544 , n69543 );
and ( n69545 , n69541 , n69544 );
and ( n69546 , n69539 , n69544 );
or ( n69547 , n69542 , n69545 , n69546 );
and ( n69548 , n59365 , n67411 );
not ( n69549 , n69548 );
and ( n69550 , n69547 , n69549 );
and ( n69551 , n60821 , n66005 );
not ( n69552 , n69551 );
and ( n69553 , n69549 , n69552 );
and ( n69554 , n69547 , n69552 );
or ( n69555 , n69550 , n69553 , n69554 );
xor ( n69556 , n69061 , n69063 );
xor ( n69557 , n69556 , n69066 );
or ( n69558 , n69555 , n69557 );
xor ( n69559 , n68894 , n68896 );
xor ( n69560 , n69559 , n68899 );
xnor ( n69561 , n69131 , n69141 );
and ( n69562 , n69560 , n69561 );
xor ( n69563 , n69159 , n69163 );
and ( n69564 , n69561 , n69563 );
and ( n69565 , n69560 , n69563 );
or ( n69566 , n69562 , n69564 , n69565 );
and ( n69567 , n69558 , n69566 );
and ( n69568 , n58628 , n68752 );
not ( n69569 , n69568 );
and ( n69570 , n63024 , n63766 );
not ( n69571 , n69570 );
and ( n69572 , n69569 , n69571 );
buf ( n69573 , n63492 );
not ( n69574 , n69573 );
and ( n69575 , n69571 , n69574 );
and ( n69576 , n69569 , n69574 );
or ( n69577 , n69572 , n69575 , n69576 );
and ( n69578 , n59615 , n67411 );
not ( n69579 , n69578 );
and ( n69580 , n61008 , n66005 );
not ( n69581 , n69580 );
and ( n69582 , n69579 , n69581 );
and ( n69583 , n61505 , n65586 );
not ( n69584 , n69583 );
and ( n69585 , n69581 , n69584 );
and ( n69586 , n69579 , n69584 );
or ( n69587 , n69582 , n69585 , n69586 );
and ( n69588 , n69577 , n69587 );
and ( n69589 , n69303 , n58444 );
not ( n69590 , n69589 );
and ( n69591 , n69590 , n69478 );
and ( n69592 , n66980 , n59920 );
not ( n69593 , n69592 );
and ( n69594 , n69478 , n69593 );
and ( n69595 , n69590 , n69593 );
or ( n69596 , n69591 , n69594 , n69595 );
and ( n69597 , n69587 , n69596 );
and ( n69598 , n69577 , n69596 );
or ( n69599 , n69588 , n69597 , n69598 );
and ( n69600 , n69059 , n58542 );
not ( n69601 , n69600 );
and ( n69602 , n66720 , n60372 );
not ( n69603 , n69602 );
and ( n69604 , n69601 , n69603 );
and ( n69605 , n65177 , n61914 );
not ( n69606 , n69605 );
and ( n69607 , n69603 , n69606 );
and ( n69608 , n69601 , n69606 );
or ( n69609 , n69604 , n69607 , n69608 );
and ( n69610 , n58292 , n69204 );
not ( n69611 , n69610 );
and ( n69612 , n64221 , n62868 );
not ( n69613 , n69612 );
and ( n69614 , n69611 , n69613 );
and ( n69615 , n63987 , n62998 );
not ( n69616 , n69615 );
and ( n69617 , n69613 , n69616 );
and ( n69618 , n69611 , n69616 );
or ( n69619 , n69614 , n69617 , n69618 );
and ( n69620 , n69609 , n69619 );
and ( n69621 , n64221 , n62151 );
not ( n69622 , n69621 );
and ( n69623 , n69619 , n69622 );
and ( n69624 , n69609 , n69622 );
or ( n69625 , n69620 , n69623 , n69624 );
and ( n69626 , n69599 , n69625 );
and ( n69627 , n49115 , n56503 );
and ( n69628 , n48988 , n56501 );
nor ( n69629 , n69627 , n69628 );
xnor ( n69630 , n69629 , n56178 );
and ( n69631 , n53328 , n51221 );
and ( n69632 , n53041 , n51219 );
nor ( n69633 , n69631 , n69632 );
xnor ( n69634 , n69633 , n51000 );
and ( n69635 , n69630 , n69634 );
xor ( n69636 , n69147 , n69151 );
xor ( n69637 , n69636 , n69156 );
and ( n69638 , n69634 , n69637 );
and ( n69639 , n69630 , n69637 );
or ( n69640 , n69635 , n69638 , n69639 );
and ( n69641 , n69625 , n69640 );
and ( n69642 , n69599 , n69640 );
or ( n69643 , n69626 , n69641 , n69642 );
and ( n69644 , n69566 , n69643 );
and ( n69645 , n69558 , n69643 );
or ( n69646 , n69567 , n69644 , n69645 );
and ( n69647 , n67343 , n59207 );
not ( n69648 , n69647 );
and ( n69649 , n65678 , n60711 );
not ( n69650 , n69649 );
and ( n69651 , n69648 , n69650 );
xor ( n69652 , n69180 , n69182 );
xor ( n69653 , n69652 , n69185 );
and ( n69654 , n69650 , n69653 );
and ( n69655 , n69648 , n69653 );
or ( n69656 , n69651 , n69654 , n69655 );
xor ( n69657 , n69194 , n69196 );
xor ( n69658 , n69657 , n69199 );
xor ( n69659 , n69206 , n69208 );
xor ( n69660 , n69659 , n69211 );
and ( n69661 , n69658 , n69660 );
xor ( n69662 , n69219 , n69223 );
and ( n69663 , n69660 , n69662 );
and ( n69664 , n69658 , n69662 );
or ( n69665 , n69661 , n69663 , n69664 );
and ( n69666 , n69656 , n69665 );
and ( n69667 , n67343 , n59611 );
not ( n69668 , n69667 );
and ( n69669 , n59908 , n67013 );
not ( n69670 , n69669 );
and ( n69671 , n69668 , n69670 );
and ( n69672 , n64548 , n62151 );
not ( n69673 , n69672 );
and ( n69674 , n69670 , n69673 );
and ( n69675 , n69668 , n69673 );
or ( n69676 , n69671 , n69674 , n69675 );
and ( n69677 , n51077 , n53928 );
and ( n69678 , n50726 , n53926 );
nor ( n69679 , n69677 , n69678 );
xnor ( n69680 , n69679 , n53652 );
and ( n69681 , n51510 , n53357 );
and ( n69682 , n51298 , n53355 );
nor ( n69683 , n69681 , n69682 );
xnor ( n69684 , n69683 , n53060 );
or ( n69685 , n69680 , n69684 );
and ( n69686 , n69676 , n69685 );
buf ( n69687 , n10629 );
buf ( n69688 , n69687 );
and ( n69689 , n69688 , n58294 );
not ( n69690 , n69689 );
and ( n69691 , n65678 , n61015 );
not ( n69692 , n69691 );
or ( n69693 , n69690 , n69692 );
and ( n69694 , n69685 , n69693 );
and ( n69695 , n69676 , n69693 );
or ( n69696 , n69686 , n69694 , n69695 );
and ( n69697 , n69665 , n69696 );
and ( n69698 , n69656 , n69696 );
or ( n69699 , n69666 , n69697 , n69698 );
and ( n69700 , n67997 , n59207 );
not ( n69701 , n69700 );
and ( n69702 , n60821 , n66469 );
not ( n69703 , n69702 );
or ( n69704 , n69701 , n69703 );
and ( n69705 , n49781 , n55851 );
and ( n69706 , n49570 , n55849 );
nor ( n69707 , n69705 , n69706 );
xnor ( n69708 , n69707 , n55506 );
and ( n69709 , n50625 , n54535 );
and ( n69710 , n50404 , n54533 );
nor ( n69711 , n69709 , n69710 );
xnor ( n69712 , n69711 , n54237 );
and ( n69713 , n69708 , n69712 );
and ( n69714 , n69704 , n69713 );
and ( n69715 , n48988 , n57187 );
and ( n69716 , n48709 , n57184 );
nor ( n69717 , n69715 , n69716 );
xnor ( n69718 , n69717 , n56175 );
and ( n69719 , n49374 , n56503 );
and ( n69720 , n49115 , n56501 );
nor ( n69721 , n69719 , n69720 );
xnor ( n69722 , n69721 , n56178 );
and ( n69723 , n69718 , n69722 );
and ( n69724 , n50195 , n55159 );
and ( n69725 , n49976 , n55157 );
nor ( n69726 , n69724 , n69725 );
xnor ( n69727 , n69726 , n54864 );
and ( n69728 , n69722 , n69727 );
and ( n69729 , n69718 , n69727 );
or ( n69730 , n69723 , n69728 , n69729 );
and ( n69731 , n69713 , n69730 );
and ( n69732 , n69704 , n69730 );
or ( n69733 , n69714 , n69731 , n69732 );
and ( n69734 , n52082 , n52799 );
and ( n69735 , n51734 , n52797 );
nor ( n69736 , n69734 , n69735 );
xnor ( n69737 , n69736 , n52538 );
and ( n69738 , n52612 , n52269 );
and ( n69739 , n52332 , n52267 );
nor ( n69740 , n69738 , n69739 );
xnor ( n69741 , n69740 , n52008 );
and ( n69742 , n69737 , n69741 );
and ( n69743 , n53041 , n51750 );
and ( n69744 , n52790 , n51748 );
nor ( n69745 , n69743 , n69744 );
xnor ( n69746 , n69745 , n51520 );
and ( n69747 , n69741 , n69746 );
and ( n69748 , n69737 , n69746 );
or ( n69749 , n69742 , n69747 , n69748 );
and ( n69750 , n53639 , n51221 );
and ( n69751 , n53328 , n51219 );
nor ( n69752 , n69750 , n69751 );
xnor ( n69753 , n69752 , n51000 );
and ( n69754 , n54227 , n50783 );
and ( n69755 , n53922 , n50781 );
nor ( n69756 , n69754 , n69755 );
xnor ( n69757 , n69756 , n50557 );
and ( n69758 , n69753 , n69757 );
and ( n69759 , n54942 , n50338 );
and ( n69760 , n54604 , n50336 );
nor ( n69761 , n69759 , n69760 );
xnor ( n69762 , n69761 , n50111 );
and ( n69763 , n69757 , n69762 );
and ( n69764 , n69753 , n69762 );
or ( n69765 , n69758 , n69763 , n69764 );
and ( n69766 , n69749 , n69765 );
and ( n69767 , n55497 , n49896 );
and ( n69768 , n55143 , n49894 );
nor ( n69769 , n69767 , n69768 );
xnor ( n69770 , n69769 , n49711 );
and ( n69771 , n56255 , n49513 );
and ( n69772 , n55756 , n49511 );
nor ( n69773 , n69771 , n69772 );
xnor ( n69774 , n69773 , n49310 );
and ( n69775 , n69770 , n69774 );
and ( n69776 , n56915 , n49121 );
and ( n69777 , n56388 , n49119 );
nor ( n69778 , n69776 , n69777 );
xnor ( n69779 , n69778 , n48932 );
and ( n69780 , n69774 , n69779 );
and ( n69781 , n69770 , n69779 );
or ( n69782 , n69775 , n69780 , n69781 );
and ( n69783 , n69765 , n69782 );
and ( n69784 , n69749 , n69782 );
or ( n69785 , n69766 , n69783 , n69784 );
and ( n69786 , n69733 , n69785 );
xor ( n69787 , n45356 , n45534 );
buf ( n69788 , n69787 );
buf ( n69789 , n69788 );
buf ( n69790 , n69789 );
and ( n69791 , n69291 , n69790 );
and ( n69792 , n68307 , n58911 );
not ( n69793 , n69792 );
and ( n69794 , n69790 , n69793 );
and ( n69795 , n69291 , n69793 );
or ( n69796 , n69791 , n69794 , n69795 );
and ( n69797 , n66415 , n60711 );
not ( n69798 , n69797 );
and ( n69799 , n65606 , n61481 );
not ( n69800 , n69799 );
and ( n69801 , n69798 , n69800 );
buf ( n69802 , n69801 );
and ( n69803 , n69796 , n69802 );
xor ( n69804 , n69238 , n69242 );
xor ( n69805 , n69804 , n69247 );
and ( n69806 , n69802 , n69805 );
and ( n69807 , n69796 , n69805 );
or ( n69808 , n69803 , n69806 , n69807 );
and ( n69809 , n69785 , n69808 );
and ( n69810 , n69733 , n69808 );
or ( n69811 , n69786 , n69809 , n69810 );
and ( n69812 , n69699 , n69811 );
xor ( n69813 , n69254 , n69258 );
xor ( n69814 , n69813 , n69263 );
xor ( n69815 , n69271 , n69275 );
xor ( n69816 , n69815 , n69280 );
and ( n69817 , n69814 , n69816 );
xor ( n69818 , n69290 , n69293 );
xor ( n69819 , n69818 , n69298 );
and ( n69820 , n69816 , n69819 );
and ( n69821 , n69814 , n69819 );
or ( n69822 , n69817 , n69820 , n69821 );
buf ( n69823 , n69170 );
xor ( n69824 , n69823 , n69172 );
and ( n69825 , n69822 , n69824 );
xor ( n69826 , n69176 , n69177 );
xor ( n69827 , n69826 , n69188 );
and ( n69828 , n69824 , n69827 );
and ( n69829 , n69822 , n69827 );
or ( n69830 , n69825 , n69828 , n69829 );
and ( n69831 , n69811 , n69830 );
and ( n69832 , n69699 , n69830 );
or ( n69833 , n69812 , n69831 , n69832 );
and ( n69834 , n69646 , n69833 );
xor ( n69835 , n69202 , n69214 );
xor ( n69836 , n69835 , n69224 );
xor ( n69837 , n69250 , n69266 );
xor ( n69838 , n69837 , n69283 );
and ( n69839 , n69836 , n69838 );
xor ( n69840 , n69301 , n69313 );
xor ( n69841 , n69840 , n69320 );
and ( n69842 , n69838 , n69841 );
and ( n69843 , n69836 , n69841 );
or ( n69844 , n69839 , n69842 , n69843 );
xor ( n69845 , n69111 , n69113 );
xor ( n69846 , n69845 , n69116 );
and ( n69847 , n69844 , n69846 );
xor ( n69848 , n69121 , n69142 );
xor ( n69849 , n69848 , n69164 );
and ( n69850 , n69846 , n69849 );
and ( n69851 , n69844 , n69849 );
or ( n69852 , n69847 , n69850 , n69851 );
and ( n69853 , n69833 , n69852 );
and ( n69854 , n69646 , n69852 );
or ( n69855 , n69834 , n69853 , n69854 );
xor ( n69856 , n69174 , n69191 );
xor ( n69857 , n69856 , n69227 );
xor ( n69858 , n69286 , n69323 );
xor ( n69859 , n69858 , n69334 );
and ( n69860 , n69857 , n69859 );
xor ( n69861 , n69347 , n69349 );
xor ( n69862 , n69861 , n69352 );
and ( n69863 , n69859 , n69862 );
and ( n69864 , n69857 , n69862 );
or ( n69865 , n69860 , n69863 , n69864 );
xor ( n69866 , n69091 , n69092 );
xor ( n69867 , n69866 , n69106 );
and ( n69868 , n69865 , n69867 );
xor ( n69869 , n69119 , n69167 );
xor ( n69870 , n69869 , n69230 );
and ( n69871 , n69867 , n69870 );
and ( n69872 , n69865 , n69870 );
or ( n69873 , n69868 , n69871 , n69872 );
and ( n69874 , n69855 , n69873 );
xor ( n69875 , n69337 , n69355 );
xor ( n69876 , n69875 , n69366 );
xor ( n69877 , n69385 , n69387 );
xor ( n69878 , n69877 , n69390 );
and ( n69879 , n69876 , n69878 );
xor ( n69880 , n69395 , n69397 );
xor ( n69881 , n69880 , n69400 );
and ( n69882 , n69878 , n69881 );
and ( n69883 , n69876 , n69881 );
or ( n69884 , n69879 , n69882 , n69883 );
and ( n69885 , n69873 , n69884 );
and ( n69886 , n69855 , n69884 );
or ( n69887 , n69874 , n69885 , n69886 );
and ( n69888 , n69537 , n69887 );
xor ( n69889 , n69109 , n69233 );
xor ( n69890 , n69889 , n69369 );
xor ( n69891 , n69393 , n69403 );
xor ( n69892 , n69891 , n69406 );
and ( n69893 , n69890 , n69892 );
xor ( n69894 , n69411 , n69413 );
xor ( n69895 , n69894 , n69416 );
and ( n69896 , n69892 , n69895 );
and ( n69897 , n69890 , n69895 );
or ( n69898 , n69893 , n69896 , n69897 );
and ( n69899 , n69887 , n69898 );
and ( n69900 , n69537 , n69898 );
or ( n69901 , n69888 , n69899 , n69900 );
xor ( n69902 , n69057 , n69088 );
xor ( n69903 , n69902 , n69372 );
xor ( n69904 , n69409 , n69419 );
xor ( n69905 , n69904 , n69422 );
and ( n69906 , n69903 , n69905 );
xor ( n69907 , n69428 , n69430 );
xor ( n69908 , n69907 , n69433 );
and ( n69909 , n69905 , n69908 );
and ( n69910 , n69903 , n69908 );
or ( n69911 , n69906 , n69909 , n69910 );
and ( n69912 , n69901 , n69911 );
xor ( n69913 , n69375 , n69425 );
xor ( n69914 , n69913 , n69436 );
and ( n69915 , n69911 , n69914 );
and ( n69916 , n69901 , n69914 );
or ( n69917 , n69912 , n69915 , n69916 );
and ( n69918 , n69466 , n69917 );
and ( n69919 , n69464 , n69917 );
or ( n69920 , n69467 , n69918 , n69919 );
xor ( n69921 , n69053 , n69453 );
xor ( n69922 , n69921 , n69456 );
and ( n69923 , n69920 , n69922 );
xor ( n69924 , n69055 , n69439 );
xor ( n69925 , n69924 , n69450 );
xor ( n69926 , n69442 , n69444 );
xor ( n69927 , n69926 , n69447 );
xor ( n69928 , n69358 , n69360 );
xor ( n69929 , n69928 , n69363 );
xor ( n69930 , n69377 , n69379 );
xor ( n69931 , n69930 , n69382 );
and ( n69932 , n69929 , n69931 );
xor ( n69933 , n69326 , n69328 );
xor ( n69934 , n69933 , n69331 );
xor ( n69935 , n69339 , n69341 );
xor ( n69936 , n69935 , n69344 );
and ( n69937 , n69934 , n69936 );
xor ( n69938 , n69488 , n69498 );
xor ( n69939 , n69938 , n69501 );
and ( n69940 , n69936 , n69939 );
and ( n69941 , n69934 , n69939 );
or ( n69942 , n69937 , n69940 , n69941 );
and ( n69943 , n69931 , n69942 );
and ( n69944 , n69929 , n69942 );
or ( n69945 , n69932 , n69943 , n69944 );
xnor ( n69946 , n69525 , n69527 );
xnor ( n69947 , n69555 , n69557 );
and ( n69948 , n69946 , n69947 );
and ( n69949 , n59615 , n67844 );
not ( n69950 , n69949 );
and ( n69951 , n59908 , n67411 );
not ( n69952 , n69951 );
and ( n69953 , n69950 , n69952 );
and ( n69954 , n62377 , n65210 );
not ( n69955 , n69954 );
and ( n69956 , n69952 , n69955 );
and ( n69957 , n69950 , n69955 );
or ( n69958 , n69953 , n69956 , n69957 );
xor ( n69959 , n69509 , n69511 );
xor ( n69960 , n69959 , n69514 );
and ( n69961 , n69958 , n69960 );
xor ( n69962 , n69539 , n69541 );
xor ( n69963 , n69962 , n69544 );
and ( n69964 , n69960 , n69963 );
and ( n69965 , n69958 , n69963 );
or ( n69966 , n69961 , n69964 , n69965 );
and ( n69967 , n68307 , n59207 );
not ( n69968 , n69967 );
and ( n69969 , n66720 , n60711 );
not ( n69970 , n69969 );
and ( n69971 , n69968 , n69970 );
and ( n69972 , n65678 , n61481 );
not ( n69973 , n69972 );
and ( n69974 , n69970 , n69973 );
and ( n69975 , n69968 , n69973 );
or ( n69976 , n69971 , n69974 , n69975 );
xor ( n69977 , n69579 , n69581 );
xor ( n69978 , n69977 , n69584 );
and ( n69979 , n69976 , n69978 );
xor ( n69980 , n69590 , n69478 );
xor ( n69981 , n69980 , n69593 );
and ( n69982 , n69978 , n69981 );
and ( n69983 , n69976 , n69981 );
or ( n69984 , n69979 , n69982 , n69983 );
and ( n69985 , n69966 , n69984 );
xor ( n69986 , n69517 , n69519 );
xor ( n69987 , n69986 , n69522 );
and ( n69988 , n69984 , n69987 );
and ( n69989 , n69966 , n69987 );
or ( n69990 , n69985 , n69988 , n69989 );
and ( n69991 , n69947 , n69990 );
and ( n69992 , n69946 , n69990 );
or ( n69993 , n69948 , n69991 , n69992 );
xor ( n69994 , n69480 , n69482 );
xor ( n69995 , n69994 , n69485 );
xor ( n69996 , n69490 , n69492 );
xor ( n69997 , n69996 , n69495 );
or ( n69998 , n69995 , n69997 );
xor ( n69999 , n69305 , n69307 );
xor ( n70000 , n69999 , n69310 );
xor ( n70001 , n69316 , n69318 );
buf ( n70002 , n70001 );
and ( n70003 , n70000 , n70002 );
xor ( n70004 , n69577 , n69587 );
xor ( n70005 , n70004 , n69596 );
and ( n70006 , n70002 , n70005 );
and ( n70007 , n70000 , n70005 );
or ( n70008 , n70003 , n70006 , n70007 );
and ( n70009 , n69998 , n70008 );
xor ( n70010 , n69547 , n69549 );
xor ( n70011 , n70010 , n69552 );
xor ( n70012 , n69609 , n69619 );
xor ( n70013 , n70012 , n69622 );
and ( n70014 , n70011 , n70013 );
xor ( n70015 , n69630 , n69634 );
xor ( n70016 , n70015 , n69637 );
and ( n70017 , n70013 , n70016 );
and ( n70018 , n70011 , n70016 );
or ( n70019 , n70014 , n70017 , n70018 );
and ( n70020 , n70008 , n70019 );
and ( n70021 , n69998 , n70019 );
or ( n70022 , n70009 , n70020 , n70021 );
and ( n70023 , n69993 , n70022 );
xor ( n70024 , n69648 , n69650 );
xor ( n70025 , n70024 , n69653 );
and ( n70026 , n69688 , n58444 );
not ( n70027 , n70026 );
and ( n70028 , n62593 , n64811 );
not ( n70029 , n70028 );
and ( n70030 , n70027 , n70029 );
and ( n70031 , n64221 , n62998 );
not ( n70032 , n70031 );
and ( n70033 , n70029 , n70032 );
and ( n70034 , n70027 , n70032 );
or ( n70035 , n70030 , n70033 , n70034 );
xor ( n70036 , n69601 , n69603 );
xor ( n70037 , n70036 , n69606 );
and ( n70038 , n70035 , n70037 );
xor ( n70039 , n69611 , n69613 );
xor ( n70040 , n70039 , n69616 );
and ( n70041 , n70037 , n70040 );
and ( n70042 , n70035 , n70040 );
or ( n70043 , n70038 , n70041 , n70042 );
and ( n70044 , n70025 , n70043 );
and ( n70045 , n58628 , n69204 );
not ( n70046 , n70045 );
and ( n70047 , n61918 , n65586 );
not ( n70048 , n70047 );
and ( n70049 , n70046 , n70048 );
and ( n70050 , n63024 , n64412 );
not ( n70051 , n70050 );
and ( n70052 , n70048 , n70051 );
and ( n70053 , n70046 , n70051 );
or ( n70054 , n70049 , n70052 , n70053 );
xor ( n70055 , n69569 , n69571 );
xor ( n70056 , n70055 , n69574 );
or ( n70057 , n70054 , n70056 );
and ( n70058 , n70043 , n70057 );
and ( n70059 , n70025 , n70057 );
or ( n70060 , n70044 , n70058 , n70059 );
xor ( n70061 , n69668 , n69670 );
xor ( n70062 , n70061 , n69673 );
xnor ( n70063 , n69680 , n69684 );
and ( n70064 , n70062 , n70063 );
xnor ( n70065 , n69690 , n69692 );
and ( n70066 , n70063 , n70065 );
and ( n70067 , n70062 , n70065 );
or ( n70068 , n70064 , n70066 , n70067 );
xnor ( n70069 , n69701 , n69703 );
xor ( n70070 , n69708 , n69712 );
and ( n70071 , n70069 , n70070 );
and ( n70072 , n58292 , n69507 );
not ( n70073 , n70072 );
and ( n70074 , n58915 , n68752 );
not ( n70075 , n70074 );
and ( n70076 , n70073 , n70075 );
and ( n70077 , n63492 , n63766 );
not ( n70078 , n70077 );
and ( n70079 , n70075 , n70078 );
and ( n70080 , n70073 , n70078 );
or ( n70081 , n70076 , n70079 , n70080 );
and ( n70082 , n70070 , n70081 );
and ( n70083 , n70069 , n70081 );
or ( n70084 , n70071 , n70082 , n70083 );
and ( n70085 , n70068 , n70084 );
and ( n70086 , n59365 , n68610 );
not ( n70087 , n70086 );
and ( n70088 , n60821 , n66917 );
not ( n70089 , n70088 );
and ( n70090 , n70087 , n70089 );
and ( n70091 , n61505 , n66005 );
not ( n70092 , n70091 );
and ( n70093 , n70089 , n70092 );
and ( n70094 , n70087 , n70092 );
or ( n70095 , n70090 , n70093 , n70094 );
and ( n70096 , n69303 , n58542 );
not ( n70097 , n70096 );
and ( n70098 , n60376 , n67013 );
not ( n70099 , n70098 );
and ( n70100 , n70097 , n70099 );
and ( n70101 , n65606 , n61914 );
not ( n70102 , n70101 );
and ( n70103 , n70099 , n70102 );
and ( n70104 , n70097 , n70102 );
or ( n70105 , n70100 , n70103 , n70104 );
and ( n70106 , n70095 , n70105 );
buf ( n70107 , n10921 );
buf ( n70108 , n70107 );
and ( n70109 , n57948 , n70108 );
not ( n70110 , n70109 );
and ( n70111 , n67343 , n59920 );
not ( n70112 , n70111 );
and ( n70113 , n70110 , n70112 );
and ( n70114 , n61008 , n66469 );
not ( n70115 , n70114 );
and ( n70116 , n70112 , n70115 );
and ( n70117 , n70110 , n70115 );
or ( n70118 , n70113 , n70116 , n70117 );
and ( n70119 , n70105 , n70118 );
and ( n70120 , n70095 , n70118 );
or ( n70121 , n70106 , n70119 , n70120 );
and ( n70122 , n70084 , n70121 );
and ( n70123 , n70068 , n70121 );
or ( n70124 , n70085 , n70122 , n70123 );
and ( n70125 , n70060 , n70124 );
and ( n70126 , n69059 , n58911 );
not ( n70127 , n70126 );
and ( n70128 , n63987 , n63679 );
not ( n70129 , n70128 );
or ( n70130 , n70127 , n70129 );
and ( n70131 , n67997 , n59611 );
and ( n70132 , n65177 , n62151 );
not ( n70133 , n70132 );
and ( n70134 , n70131 , n70133 );
and ( n70135 , n70130 , n70134 );
not ( n70136 , n70131 );
buf ( n70137 , n70136 );
and ( n70138 , n70134 , n70137 );
and ( n70139 , n70130 , n70137 );
or ( n70140 , n70135 , n70138 , n70139 );
and ( n70141 , n49115 , n57187 );
and ( n70142 , n48988 , n57184 );
nor ( n70143 , n70141 , n70142 );
xnor ( n70144 , n70143 , n56175 );
and ( n70145 , n49570 , n56503 );
and ( n70146 , n49374 , n56501 );
nor ( n70147 , n70145 , n70146 );
xnor ( n70148 , n70147 , n56178 );
and ( n70149 , n70144 , n70148 );
and ( n70150 , n49976 , n55851 );
and ( n70151 , n49781 , n55849 );
nor ( n70152 , n70150 , n70151 );
xnor ( n70153 , n70152 , n55506 );
and ( n70154 , n70148 , n70153 );
and ( n70155 , n70144 , n70153 );
or ( n70156 , n70149 , n70154 , n70155 );
and ( n70157 , n50404 , n55159 );
and ( n70158 , n50195 , n55157 );
nor ( n70159 , n70157 , n70158 );
xnor ( n70160 , n70159 , n54864 );
and ( n70161 , n50726 , n54535 );
and ( n70162 , n50625 , n54533 );
nor ( n70163 , n70161 , n70162 );
xnor ( n70164 , n70163 , n54237 );
and ( n70165 , n70160 , n70164 );
and ( n70166 , n51298 , n53928 );
and ( n70167 , n51077 , n53926 );
nor ( n70168 , n70166 , n70167 );
xnor ( n70169 , n70168 , n53652 );
and ( n70170 , n70164 , n70169 );
and ( n70171 , n70160 , n70169 );
or ( n70172 , n70165 , n70170 , n70171 );
and ( n70173 , n70156 , n70172 );
and ( n70174 , n51734 , n53357 );
and ( n70175 , n51510 , n53355 );
nor ( n70176 , n70174 , n70175 );
xnor ( n70177 , n70176 , n53060 );
and ( n70178 , n52332 , n52799 );
and ( n70179 , n52082 , n52797 );
nor ( n70180 , n70178 , n70179 );
xnor ( n70181 , n70180 , n52538 );
and ( n70182 , n70177 , n70181 );
and ( n70183 , n52790 , n52269 );
and ( n70184 , n52612 , n52267 );
nor ( n70185 , n70183 , n70184 );
xnor ( n70186 , n70185 , n52008 );
and ( n70187 , n70181 , n70186 );
and ( n70188 , n70177 , n70186 );
or ( n70189 , n70182 , n70187 , n70188 );
and ( n70190 , n70172 , n70189 );
and ( n70191 , n70156 , n70189 );
or ( n70192 , n70173 , n70190 , n70191 );
and ( n70193 , n70140 , n70192 );
and ( n70194 , n53328 , n51750 );
and ( n70195 , n53041 , n51748 );
nor ( n70196 , n70194 , n70195 );
xnor ( n70197 , n70196 , n51520 );
and ( n70198 , n53922 , n51221 );
and ( n70199 , n53639 , n51219 );
nor ( n70200 , n70198 , n70199 );
xnor ( n70201 , n70200 , n51000 );
and ( n70202 , n70197 , n70201 );
and ( n70203 , n54604 , n50783 );
and ( n70204 , n54227 , n50781 );
nor ( n70205 , n70203 , n70204 );
xnor ( n70206 , n70205 , n50557 );
and ( n70207 , n70201 , n70206 );
and ( n70208 , n70197 , n70206 );
or ( n70209 , n70202 , n70207 , n70208 );
and ( n70210 , n55143 , n50338 );
and ( n70211 , n54942 , n50336 );
nor ( n70212 , n70210 , n70211 );
xnor ( n70213 , n70212 , n50111 );
and ( n70214 , n55756 , n49896 );
and ( n70215 , n55497 , n49894 );
nor ( n70216 , n70214 , n70215 );
xnor ( n70217 , n70216 , n49711 );
and ( n70218 , n70213 , n70217 );
and ( n70219 , n56388 , n49513 );
and ( n70220 , n56255 , n49511 );
nor ( n70221 , n70219 , n70220 );
xnor ( n70222 , n70221 , n49310 );
and ( n70223 , n70217 , n70222 );
and ( n70224 , n70213 , n70222 );
or ( n70225 , n70218 , n70223 , n70224 );
and ( n70226 , n70209 , n70225 );
and ( n70227 , n57063 , n49121 );
and ( n70228 , n56915 , n49119 );
nor ( n70229 , n70227 , n70228 );
xnor ( n70230 , n70229 , n48932 );
and ( n70231 , n57063 , n49119 );
not ( n70232 , n70231 );
and ( n70233 , n70232 , n48932 );
and ( n70234 , n70230 , n70233 );
xor ( n70235 , n45359 , n45532 );
buf ( n70236 , n70235 );
buf ( n70237 , n70236 );
buf ( n70238 , n70237 );
and ( n70239 , n70233 , n70238 );
and ( n70240 , n70230 , n70238 );
or ( n70241 , n70234 , n70239 , n70240 );
and ( n70242 , n70225 , n70241 );
and ( n70243 , n70209 , n70241 );
or ( n70244 , n70226 , n70242 , n70243 );
and ( n70245 , n70192 , n70244 );
and ( n70246 , n70140 , n70244 );
or ( n70247 , n70193 , n70245 , n70246 );
and ( n70248 , n70124 , n70247 );
and ( n70249 , n70060 , n70247 );
or ( n70250 , n70125 , n70248 , n70249 );
and ( n70251 , n70022 , n70250 );
and ( n70252 , n69993 , n70250 );
or ( n70253 , n70023 , n70251 , n70252 );
and ( n70254 , n69945 , n70253 );
buf ( n70255 , n10921 );
buf ( n70256 , n70255 );
and ( n70257 , n70256 , n58294 );
not ( n70258 , n70257 );
and ( n70259 , n66980 , n60372 );
not ( n70260 , n70259 );
and ( n70261 , n70258 , n70260 );
and ( n70262 , n66415 , n61015 );
not ( n70263 , n70262 );
and ( n70264 , n70260 , n70263 );
and ( n70265 , n70258 , n70263 );
or ( n70266 , n70261 , n70264 , n70265 );
xor ( n70267 , n69718 , n69722 );
xor ( n70268 , n70267 , n69727 );
and ( n70269 , n70266 , n70268 );
xor ( n70270 , n69737 , n69741 );
xor ( n70271 , n70270 , n69746 );
and ( n70272 , n70268 , n70271 );
and ( n70273 , n70266 , n70271 );
or ( n70274 , n70269 , n70272 , n70273 );
xor ( n70275 , n69753 , n69757 );
xor ( n70276 , n70275 , n69762 );
xor ( n70277 , n69770 , n69774 );
xor ( n70278 , n70277 , n69779 );
and ( n70279 , n70276 , n70278 );
xor ( n70280 , n69291 , n69790 );
xor ( n70281 , n70280 , n69793 );
and ( n70282 , n70278 , n70281 );
and ( n70283 , n70276 , n70281 );
or ( n70284 , n70279 , n70282 , n70283 );
and ( n70285 , n70274 , n70284 );
xor ( n70286 , n69658 , n69660 );
xor ( n70287 , n70286 , n69662 );
and ( n70288 , n70284 , n70287 );
and ( n70289 , n70274 , n70287 );
or ( n70290 , n70285 , n70288 , n70289 );
xor ( n70291 , n69676 , n69685 );
xor ( n70292 , n70291 , n69693 );
xor ( n70293 , n69704 , n69713 );
xor ( n70294 , n70293 , n69730 );
and ( n70295 , n70292 , n70294 );
xor ( n70296 , n69749 , n69765 );
xor ( n70297 , n70296 , n69782 );
and ( n70298 , n70294 , n70297 );
and ( n70299 , n70292 , n70297 );
or ( n70300 , n70295 , n70298 , n70299 );
and ( n70301 , n70290 , n70300 );
xor ( n70302 , n69560 , n69561 );
xor ( n70303 , n70302 , n69563 );
and ( n70304 , n70300 , n70303 );
and ( n70305 , n70290 , n70303 );
or ( n70306 , n70301 , n70304 , n70305 );
xor ( n70307 , n69599 , n69625 );
xor ( n70308 , n70307 , n69640 );
xor ( n70309 , n69656 , n69665 );
xor ( n70310 , n70309 , n69696 );
and ( n70311 , n70308 , n70310 );
xor ( n70312 , n69733 , n69785 );
xor ( n70313 , n70312 , n69808 );
and ( n70314 , n70310 , n70313 );
and ( n70315 , n70308 , n70313 );
or ( n70316 , n70311 , n70314 , n70315 );
and ( n70317 , n70306 , n70316 );
xor ( n70318 , n69477 , n69504 );
xor ( n70319 , n70318 , n69528 );
and ( n70320 , n70316 , n70319 );
and ( n70321 , n70306 , n70319 );
or ( n70322 , n70317 , n70320 , n70321 );
and ( n70323 , n70253 , n70322 );
and ( n70324 , n69945 , n70322 );
or ( n70325 , n70254 , n70323 , n70324 );
xor ( n70326 , n69558 , n69566 );
xor ( n70327 , n70326 , n69643 );
xor ( n70328 , n69699 , n69811 );
xor ( n70329 , n70328 , n69830 );
and ( n70330 , n70327 , n70329 );
xor ( n70331 , n69844 , n69846 );
xor ( n70332 , n70331 , n69849 );
and ( n70333 , n70329 , n70332 );
and ( n70334 , n70327 , n70332 );
or ( n70335 , n70330 , n70333 , n70334 );
xor ( n70336 , n69473 , n69475 );
xor ( n70337 , n70336 , n69531 );
and ( n70338 , n70335 , n70337 );
xor ( n70339 , n69646 , n69833 );
xor ( n70340 , n70339 , n69852 );
and ( n70341 , n70337 , n70340 );
and ( n70342 , n70335 , n70340 );
or ( n70343 , n70338 , n70341 , n70342 );
and ( n70344 , n70325 , n70343 );
xor ( n70345 , n69469 , n69470 );
xor ( n70346 , n70345 , n69534 );
and ( n70347 , n70343 , n70346 );
and ( n70348 , n70325 , n70346 );
or ( n70349 , n70344 , n70347 , n70348 );
xor ( n70350 , n69537 , n69887 );
xor ( n70351 , n70350 , n69898 );
and ( n70352 , n70349 , n70351 );
xor ( n70353 , n69903 , n69905 );
xor ( n70354 , n70353 , n69908 );
and ( n70355 , n70351 , n70354 );
and ( n70356 , n70349 , n70354 );
or ( n70357 , n70352 , n70355 , n70356 );
and ( n70358 , n69927 , n70357 );
xor ( n70359 , n69901 , n69911 );
xor ( n70360 , n70359 , n69914 );
and ( n70361 , n70357 , n70360 );
and ( n70362 , n69927 , n70360 );
or ( n70363 , n70358 , n70361 , n70362 );
and ( n70364 , n69925 , n70363 );
xor ( n70365 , n69464 , n69466 );
xor ( n70366 , n70365 , n69917 );
and ( n70367 , n70363 , n70366 );
and ( n70368 , n69925 , n70366 );
or ( n70369 , n70364 , n70367 , n70368 );
and ( n70370 , n69922 , n70369 );
and ( n70371 , n69920 , n70369 );
or ( n70372 , n69923 , n70370 , n70371 );
and ( n70373 , n69461 , n70372 );
and ( n70374 , n69459 , n70372 );
or ( n70375 , n69462 , n70373 , n70374 );
and ( n70376 , n69051 , n70375 );
xor ( n70377 , n69051 , n70375 );
xor ( n70378 , n69459 , n69461 );
xor ( n70379 , n70378 , n70372 );
not ( n70380 , n70379 );
xor ( n70381 , n69920 , n69922 );
xor ( n70382 , n70381 , n70369 );
xor ( n70383 , n69925 , n70363 );
xor ( n70384 , n70383 , n70366 );
xor ( n70385 , n69927 , n70357 );
xor ( n70386 , n70385 , n70360 );
xor ( n70387 , n69855 , n69873 );
xor ( n70388 , n70387 , n69884 );
xor ( n70389 , n69890 , n69892 );
xor ( n70390 , n70389 , n69895 );
and ( n70391 , n70388 , n70390 );
xor ( n70392 , n69865 , n69867 );
xor ( n70393 , n70392 , n69870 );
xor ( n70394 , n69876 , n69878 );
xor ( n70395 , n70394 , n69881 );
and ( n70396 , n70393 , n70395 );
xor ( n70397 , n69857 , n69859 );
xor ( n70398 , n70397 , n69862 );
xor ( n70399 , n69822 , n69824 );
xor ( n70400 , n70399 , n69827 );
xor ( n70401 , n69836 , n69838 );
xor ( n70402 , n70401 , n69841 );
and ( n70403 , n70400 , n70402 );
xor ( n70404 , n69796 , n69802 );
xor ( n70405 , n70404 , n69805 );
xor ( n70406 , n69814 , n69816 );
xor ( n70407 , n70406 , n69819 );
and ( n70408 , n70405 , n70407 );
xor ( n70409 , n69966 , n69984 );
xor ( n70410 , n70409 , n69987 );
and ( n70411 , n70407 , n70410 );
and ( n70412 , n70405 , n70410 );
or ( n70413 , n70408 , n70411 , n70412 );
and ( n70414 , n70402 , n70413 );
and ( n70415 , n70400 , n70413 );
or ( n70416 , n70403 , n70414 , n70415 );
and ( n70417 , n70398 , n70416 );
xnor ( n70418 , n69995 , n69997 );
xor ( n70419 , n69798 , n69800 );
buf ( n70420 , n70419 );
xor ( n70421 , n69958 , n69960 );
xor ( n70422 , n70421 , n69963 );
and ( n70423 , n70420 , n70422 );
xor ( n70424 , n69976 , n69978 );
xor ( n70425 , n70424 , n69981 );
and ( n70426 , n70422 , n70425 );
and ( n70427 , n70420 , n70425 );
or ( n70428 , n70423 , n70426 , n70427 );
and ( n70429 , n70418 , n70428 );
xor ( n70430 , n70035 , n70037 );
xor ( n70431 , n70430 , n70040 );
xnor ( n70432 , n70054 , n70056 );
and ( n70433 , n70431 , n70432 );
and ( n70434 , n58915 , n69204 );
not ( n70435 , n70434 );
and ( n70436 , n60376 , n67411 );
not ( n70437 , n70436 );
and ( n70438 , n70435 , n70437 );
and ( n70439 , n63024 , n64811 );
not ( n70440 , n70439 );
and ( n70441 , n70437 , n70440 );
and ( n70442 , n70435 , n70440 );
or ( n70443 , n70438 , n70441 , n70442 );
and ( n70444 , n58628 , n69507 );
not ( n70445 , n70444 );
and ( n70446 , n61918 , n66005 );
not ( n70447 , n70446 );
and ( n70448 , n70445 , n70447 );
and ( n70449 , n62593 , n65210 );
not ( n70450 , n70449 );
and ( n70451 , n70447 , n70450 );
and ( n70452 , n70445 , n70450 );
or ( n70453 , n70448 , n70451 , n70452 );
and ( n70454 , n70443 , n70453 );
xor ( n70455 , n70073 , n70075 );
xor ( n70456 , n70455 , n70078 );
and ( n70457 , n70453 , n70456 );
and ( n70458 , n70443 , n70456 );
or ( n70459 , n70454 , n70457 , n70458 );
and ( n70460 , n70432 , n70459 );
and ( n70461 , n70431 , n70459 );
or ( n70462 , n70433 , n70460 , n70461 );
and ( n70463 , n70428 , n70462 );
and ( n70464 , n70418 , n70462 );
or ( n70465 , n70429 , n70463 , n70464 );
xor ( n70466 , n69968 , n69970 );
xor ( n70467 , n70466 , n69973 );
xor ( n70468 , n70087 , n70089 );
xor ( n70469 , n70468 , n70092 );
and ( n70470 , n70467 , n70469 );
and ( n70471 , n64548 , n62868 );
not ( n70472 , n70471 );
xor ( n70473 , n70046 , n70048 );
xor ( n70474 , n70473 , n70051 );
and ( n70475 , n70472 , n70474 );
buf ( n70476 , n70475 );
and ( n70477 , n70470 , n70476 );
xor ( n70478 , n69950 , n69952 );
xor ( n70479 , n70478 , n69955 );
xor ( n70480 , n70027 , n70029 );
xor ( n70481 , n70480 , n70032 );
and ( n70482 , n70479 , n70481 );
xor ( n70483 , n70097 , n70099 );
xor ( n70484 , n70483 , n70102 );
and ( n70485 , n70481 , n70484 );
and ( n70486 , n70479 , n70484 );
or ( n70487 , n70482 , n70485 , n70486 );
and ( n70488 , n70476 , n70487 );
and ( n70489 , n70470 , n70487 );
or ( n70490 , n70477 , n70488 , n70489 );
xor ( n70491 , n70110 , n70112 );
xor ( n70492 , n70491 , n70115 );
xnor ( n70493 , n70127 , n70129 );
and ( n70494 , n70492 , n70493 );
xor ( n70495 , n70131 , n70133 );
and ( n70496 , n70493 , n70495 );
and ( n70497 , n70492 , n70495 );
or ( n70498 , n70494 , n70496 , n70497 );
and ( n70499 , n59908 , n67844 );
not ( n70500 , n70499 );
and ( n70501 , n62377 , n65586 );
not ( n70502 , n70501 );
and ( n70503 , n70500 , n70502 );
buf ( n70504 , n63987 );
not ( n70505 , n70504 );
and ( n70506 , n70502 , n70505 );
and ( n70507 , n70500 , n70505 );
or ( n70508 , n70503 , n70506 , n70507 );
and ( n70509 , n59615 , n68610 );
not ( n70510 , n70509 );
and ( n70511 , n61008 , n66917 );
not ( n70512 , n70511 );
and ( n70513 , n70510 , n70512 );
and ( n70514 , n61505 , n66469 );
not ( n70515 , n70514 );
and ( n70516 , n70512 , n70515 );
and ( n70517 , n70510 , n70515 );
or ( n70518 , n70513 , n70516 , n70517 );
and ( n70519 , n70508 , n70518 );
and ( n70520 , n69303 , n58911 );
not ( n70521 , n70520 );
and ( n70522 , n67343 , n60372 );
not ( n70523 , n70522 );
and ( n70524 , n70521 , n70523 );
and ( n70525 , n63492 , n64412 );
not ( n70526 , n70525 );
and ( n70527 , n70523 , n70526 );
and ( n70528 , n70521 , n70526 );
or ( n70529 , n70524 , n70527 , n70528 );
and ( n70530 , n70518 , n70529 );
and ( n70531 , n70508 , n70529 );
or ( n70532 , n70519 , n70530 , n70531 );
and ( n70533 , n70498 , n70532 );
and ( n70534 , n58292 , n70108 );
not ( n70535 , n70534 );
and ( n70536 , n69688 , n58542 );
not ( n70537 , n70536 );
and ( n70538 , n70535 , n70537 );
and ( n70539 , n64548 , n62998 );
not ( n70540 , n70539 );
and ( n70541 , n70537 , n70540 );
and ( n70542 , n70535 , n70540 );
or ( n70543 , n70538 , n70541 , n70542 );
and ( n70544 , n68307 , n59611 );
not ( n70545 , n70544 );
and ( n70546 , n67997 , n59920 );
not ( n70547 , n70546 );
and ( n70548 , n70545 , n70547 );
and ( n70549 , n65606 , n62151 );
not ( n70550 , n70549 );
and ( n70551 , n70547 , n70550 );
and ( n70552 , n70545 , n70550 );
or ( n70553 , n70548 , n70551 , n70552 );
and ( n70554 , n70543 , n70553 );
and ( n70555 , n51077 , n54535 );
and ( n70556 , n50726 , n54533 );
nor ( n70557 , n70555 , n70556 );
xnor ( n70558 , n70557 , n54237 );
and ( n70559 , n53639 , n51750 );
and ( n70560 , n53328 , n51748 );
nor ( n70561 , n70559 , n70560 );
xnor ( n70562 , n70561 , n51520 );
or ( n70563 , n70558 , n70562 );
and ( n70564 , n70553 , n70563 );
and ( n70565 , n70543 , n70563 );
or ( n70566 , n70554 , n70564 , n70565 );
and ( n70567 , n70532 , n70566 );
and ( n70568 , n70498 , n70566 );
or ( n70569 , n70533 , n70567 , n70568 );
and ( n70570 , n70490 , n70569 );
and ( n70571 , n65678 , n61914 );
not ( n70572 , n70571 );
and ( n70573 , n65177 , n62868 );
not ( n70574 , n70573 );
or ( n70575 , n70572 , n70574 );
and ( n70576 , n70256 , n58444 );
not ( n70577 , n70576 );
and ( n70578 , n64221 , n63679 );
not ( n70579 , n70578 );
or ( n70580 , n70577 , n70579 );
and ( n70581 , n70575 , n70580 );
and ( n70582 , n49374 , n57187 );
and ( n70583 , n49115 , n57184 );
nor ( n70584 , n70582 , n70583 );
xnor ( n70585 , n70584 , n56175 );
and ( n70586 , n49781 , n56503 );
and ( n70587 , n49570 , n56501 );
nor ( n70588 , n70586 , n70587 );
xnor ( n70589 , n70588 , n56178 );
and ( n70590 , n70585 , n70589 );
and ( n70591 , n50195 , n55851 );
and ( n70592 , n49976 , n55849 );
nor ( n70593 , n70591 , n70592 );
xnor ( n70594 , n70593 , n55506 );
and ( n70595 , n70589 , n70594 );
and ( n70596 , n70585 , n70594 );
or ( n70597 , n70590 , n70595 , n70596 );
and ( n70598 , n70580 , n70597 );
and ( n70599 , n70575 , n70597 );
or ( n70600 , n70581 , n70598 , n70599 );
and ( n70601 , n50625 , n55159 );
and ( n70602 , n50404 , n55157 );
nor ( n70603 , n70601 , n70602 );
xnor ( n70604 , n70603 , n54864 );
and ( n70605 , n51510 , n53928 );
and ( n70606 , n51298 , n53926 );
nor ( n70607 , n70605 , n70606 );
xnor ( n70608 , n70607 , n53652 );
and ( n70609 , n70604 , n70608 );
and ( n70610 , n52082 , n53357 );
and ( n70611 , n51734 , n53355 );
nor ( n70612 , n70610 , n70611 );
xnor ( n70613 , n70612 , n53060 );
and ( n70614 , n70608 , n70613 );
and ( n70615 , n70604 , n70613 );
or ( n70616 , n70609 , n70614 , n70615 );
and ( n70617 , n52612 , n52799 );
and ( n70618 , n52332 , n52797 );
nor ( n70619 , n70617 , n70618 );
xnor ( n70620 , n70619 , n52538 );
and ( n70621 , n53041 , n52269 );
and ( n70622 , n52790 , n52267 );
nor ( n70623 , n70621 , n70622 );
xnor ( n70624 , n70623 , n52008 );
and ( n70625 , n70620 , n70624 );
and ( n70626 , n54227 , n51221 );
and ( n70627 , n53922 , n51219 );
nor ( n70628 , n70626 , n70627 );
xnor ( n70629 , n70628 , n51000 );
and ( n70630 , n70624 , n70629 );
and ( n70631 , n70620 , n70629 );
or ( n70632 , n70625 , n70630 , n70631 );
and ( n70633 , n70616 , n70632 );
and ( n70634 , n54942 , n50783 );
and ( n70635 , n54604 , n50781 );
nor ( n70636 , n70634 , n70635 );
xnor ( n70637 , n70636 , n50557 );
and ( n70638 , n55497 , n50338 );
and ( n70639 , n55143 , n50336 );
nor ( n70640 , n70638 , n70639 );
xnor ( n70641 , n70640 , n50111 );
and ( n70642 , n70637 , n70641 );
and ( n70643 , n56255 , n49896 );
and ( n70644 , n55756 , n49894 );
nor ( n70645 , n70643 , n70644 );
xnor ( n70646 , n70645 , n49711 );
and ( n70647 , n70641 , n70646 );
and ( n70648 , n70637 , n70646 );
or ( n70649 , n70642 , n70647 , n70648 );
and ( n70650 , n70632 , n70649 );
and ( n70651 , n70616 , n70649 );
or ( n70652 , n70633 , n70650 , n70651 );
and ( n70653 , n70600 , n70652 );
and ( n70654 , n56915 , n49513 );
and ( n70655 , n56388 , n49511 );
nor ( n70656 , n70654 , n70655 );
xnor ( n70657 , n70656 , n49310 );
and ( n70658 , n70657 , n70231 );
xor ( n70659 , n45361 , n45531 );
buf ( n70660 , n70659 );
buf ( n70661 , n70660 );
buf ( n70662 , n70661 );
and ( n70663 , n70231 , n70662 );
and ( n70664 , n70657 , n70662 );
or ( n70665 , n70658 , n70663 , n70664 );
and ( n70666 , n66720 , n61015 );
not ( n70667 , n70666 );
and ( n70668 , n66415 , n61481 );
not ( n70669 , n70668 );
and ( n70670 , n70667 , n70669 );
buf ( n70671 , n70670 );
and ( n70672 , n70665 , n70671 );
xor ( n70673 , n70144 , n70148 );
xor ( n70674 , n70673 , n70153 );
and ( n70675 , n70671 , n70674 );
and ( n70676 , n70665 , n70674 );
or ( n70677 , n70672 , n70675 , n70676 );
and ( n70678 , n70652 , n70677 );
and ( n70679 , n70600 , n70677 );
or ( n70680 , n70653 , n70678 , n70679 );
and ( n70681 , n70569 , n70680 );
and ( n70682 , n70490 , n70680 );
or ( n70683 , n70570 , n70681 , n70682 );
and ( n70684 , n70465 , n70683 );
xor ( n70685 , n70160 , n70164 );
xor ( n70686 , n70685 , n70169 );
xor ( n70687 , n70177 , n70181 );
xor ( n70688 , n70687 , n70186 );
and ( n70689 , n70686 , n70688 );
xor ( n70690 , n70197 , n70201 );
xor ( n70691 , n70690 , n70206 );
and ( n70692 , n70688 , n70691 );
and ( n70693 , n70686 , n70691 );
or ( n70694 , n70689 , n70692 , n70693 );
xor ( n70695 , n70213 , n70217 );
xor ( n70696 , n70695 , n70222 );
xor ( n70697 , n70230 , n70233 );
xor ( n70698 , n70697 , n70238 );
and ( n70699 , n70696 , n70698 );
xor ( n70700 , n70258 , n70260 );
xor ( n70701 , n70700 , n70263 );
and ( n70702 , n70698 , n70701 );
and ( n70703 , n70696 , n70701 );
or ( n70704 , n70699 , n70702 , n70703 );
and ( n70705 , n70694 , n70704 );
xor ( n70706 , n70062 , n70063 );
xor ( n70707 , n70706 , n70065 );
and ( n70708 , n70704 , n70707 );
and ( n70709 , n70694 , n70707 );
or ( n70710 , n70705 , n70708 , n70709 );
xor ( n70711 , n70069 , n70070 );
xor ( n70712 , n70711 , n70081 );
xor ( n70713 , n70095 , n70105 );
xor ( n70714 , n70713 , n70118 );
and ( n70715 , n70712 , n70714 );
xor ( n70716 , n70130 , n70134 );
xor ( n70717 , n70716 , n70137 );
and ( n70718 , n70714 , n70717 );
and ( n70719 , n70712 , n70717 );
or ( n70720 , n70715 , n70718 , n70719 );
and ( n70721 , n70710 , n70720 );
xor ( n70722 , n70156 , n70172 );
xor ( n70723 , n70722 , n70189 );
xor ( n70724 , n70209 , n70225 );
xor ( n70725 , n70724 , n70241 );
and ( n70726 , n70723 , n70725 );
xor ( n70727 , n70266 , n70268 );
xor ( n70728 , n70727 , n70271 );
and ( n70729 , n70725 , n70728 );
and ( n70730 , n70723 , n70728 );
or ( n70731 , n70726 , n70729 , n70730 );
and ( n70732 , n70720 , n70731 );
and ( n70733 , n70710 , n70731 );
or ( n70734 , n70721 , n70732 , n70733 );
and ( n70735 , n70683 , n70734 );
and ( n70736 , n70465 , n70734 );
or ( n70737 , n70684 , n70735 , n70736 );
and ( n70738 , n70416 , n70737 );
and ( n70739 , n70398 , n70737 );
or ( n70740 , n70417 , n70738 , n70739 );
and ( n70741 , n70395 , n70740 );
and ( n70742 , n70393 , n70740 );
or ( n70743 , n70396 , n70741 , n70742 );
and ( n70744 , n70390 , n70743 );
and ( n70745 , n70388 , n70743 );
or ( n70746 , n70391 , n70744 , n70745 );
xor ( n70747 , n70349 , n70351 );
xor ( n70748 , n70747 , n70354 );
and ( n70749 , n70746 , n70748 );
xor ( n70750 , n70000 , n70002 );
xor ( n70751 , n70750 , n70005 );
xor ( n70752 , n70011 , n70013 );
xor ( n70753 , n70752 , n70016 );
and ( n70754 , n70751 , n70753 );
xor ( n70755 , n70025 , n70043 );
xor ( n70756 , n70755 , n70057 );
and ( n70757 , n70753 , n70756 );
and ( n70758 , n70751 , n70756 );
or ( n70759 , n70754 , n70757 , n70758 );
xor ( n70760 , n70068 , n70084 );
xor ( n70761 , n70760 , n70121 );
xor ( n70762 , n70140 , n70192 );
xor ( n70763 , n70762 , n70244 );
and ( n70764 , n70761 , n70763 );
xor ( n70765 , n70274 , n70284 );
xor ( n70766 , n70765 , n70287 );
and ( n70767 , n70763 , n70766 );
and ( n70768 , n70761 , n70766 );
or ( n70769 , n70764 , n70767 , n70768 );
and ( n70770 , n70759 , n70769 );
xor ( n70771 , n69934 , n69936 );
xor ( n70772 , n70771 , n69939 );
and ( n70773 , n70769 , n70772 );
and ( n70774 , n70759 , n70772 );
or ( n70775 , n70770 , n70773 , n70774 );
xor ( n70776 , n69946 , n69947 );
xor ( n70777 , n70776 , n69990 );
xor ( n70778 , n69998 , n70008 );
xor ( n70779 , n70778 , n70019 );
and ( n70780 , n70777 , n70779 );
xor ( n70781 , n70060 , n70124 );
xor ( n70782 , n70781 , n70247 );
and ( n70783 , n70779 , n70782 );
and ( n70784 , n70777 , n70782 );
or ( n70785 , n70780 , n70783 , n70784 );
and ( n70786 , n70775 , n70785 );
xor ( n70787 , n69929 , n69931 );
xor ( n70788 , n70787 , n69942 );
and ( n70789 , n70785 , n70788 );
and ( n70790 , n70775 , n70788 );
or ( n70791 , n70786 , n70789 , n70790 );
xor ( n70792 , n69993 , n70022 );
xor ( n70793 , n70792 , n70250 );
xor ( n70794 , n70306 , n70316 );
xor ( n70795 , n70794 , n70319 );
and ( n70796 , n70793 , n70795 );
xor ( n70797 , n70327 , n70329 );
xor ( n70798 , n70797 , n70332 );
and ( n70799 , n70795 , n70798 );
and ( n70800 , n70793 , n70798 );
or ( n70801 , n70796 , n70799 , n70800 );
and ( n70802 , n70791 , n70801 );
xor ( n70803 , n69945 , n70253 );
xor ( n70804 , n70803 , n70322 );
and ( n70805 , n70801 , n70804 );
and ( n70806 , n70791 , n70804 );
or ( n70807 , n70802 , n70805 , n70806 );
xor ( n70808 , n70325 , n70343 );
xor ( n70809 , n70808 , n70346 );
and ( n70810 , n70807 , n70809 );
xor ( n70811 , n70335 , n70337 );
xor ( n70812 , n70811 , n70340 );
xor ( n70813 , n70290 , n70300 );
xor ( n70814 , n70813 , n70303 );
xor ( n70815 , n70308 , n70310 );
xor ( n70816 , n70815 , n70313 );
and ( n70817 , n70814 , n70816 );
xor ( n70818 , n70292 , n70294 );
xor ( n70819 , n70818 , n70297 );
xor ( n70820 , n70276 , n70278 );
xor ( n70821 , n70820 , n70281 );
and ( n70822 , n58915 , n69507 );
not ( n70823 , n70822 );
and ( n70824 , n63492 , n64811 );
not ( n70825 , n70824 );
and ( n70826 , n70823 , n70825 );
and ( n70827 , n63987 , n64412 );
not ( n70828 , n70827 );
and ( n70829 , n70825 , n70828 );
and ( n70830 , n70823 , n70828 );
or ( n70831 , n70826 , n70829 , n70830 );
and ( n70832 , n69059 , n59207 );
not ( n70833 , n70832 );
and ( n70834 , n70831 , n70833 );
and ( n70835 , n66980 , n60711 );
not ( n70836 , n70835 );
and ( n70837 , n70833 , n70836 );
and ( n70838 , n70831 , n70836 );
or ( n70839 , n70834 , n70837 , n70838 );
and ( n70840 , n69688 , n58911 );
not ( n70841 , n70840 );
and ( n70842 , n64548 , n63679 );
not ( n70843 , n70842 );
and ( n70844 , n70841 , n70843 );
and ( n70845 , n64221 , n63766 );
not ( n70846 , n70845 );
and ( n70847 , n70843 , n70846 );
and ( n70848 , n70841 , n70846 );
or ( n70849 , n70844 , n70847 , n70848 );
and ( n70850 , n59365 , n68752 );
not ( n70851 , n70850 );
and ( n70852 , n70849 , n70851 );
and ( n70853 , n60821 , n67013 );
not ( n70854 , n70853 );
and ( n70855 , n70851 , n70854 );
and ( n70856 , n70849 , n70854 );
or ( n70857 , n70852 , n70855 , n70856 );
and ( n70858 , n70839 , n70857 );
and ( n70859 , n70821 , n70858 );
xor ( n70860 , n70443 , n70453 );
xor ( n70861 , n70860 , n70456 );
xor ( n70862 , n70467 , n70469 );
and ( n70863 , n70861 , n70862 );
and ( n70864 , n58628 , n70108 );
not ( n70865 , n70864 );
and ( n70866 , n67997 , n60372 );
not ( n70867 , n70866 );
and ( n70868 , n70865 , n70867 );
and ( n70869 , n63024 , n65210 );
not ( n70870 , n70869 );
and ( n70871 , n70867 , n70870 );
and ( n70872 , n70865 , n70870 );
or ( n70873 , n70868 , n70871 , n70872 );
xor ( n70874 , n70521 , n70523 );
xor ( n70875 , n70874 , n70526 );
or ( n70876 , n70873 , n70875 );
and ( n70877 , n70862 , n70876 );
and ( n70878 , n70861 , n70876 );
or ( n70879 , n70863 , n70877 , n70878 );
and ( n70880 , n70858 , n70879 );
and ( n70881 , n70821 , n70879 );
or ( n70882 , n70859 , n70880 , n70881 );
and ( n70883 , n70819 , n70882 );
xor ( n70884 , n70435 , n70437 );
xor ( n70885 , n70884 , n70440 );
xor ( n70886 , n70500 , n70502 );
xor ( n70887 , n70886 , n70505 );
and ( n70888 , n70885 , n70887 );
xor ( n70889 , n70510 , n70512 );
xor ( n70890 , n70889 , n70515 );
and ( n70891 , n70887 , n70890 );
and ( n70892 , n70885 , n70890 );
or ( n70893 , n70888 , n70891 , n70892 );
xor ( n70894 , n70535 , n70537 );
xor ( n70895 , n70894 , n70540 );
xor ( n70896 , n70545 , n70547 );
xor ( n70897 , n70896 , n70550 );
and ( n70898 , n70895 , n70897 );
xnor ( n70899 , n70558 , n70562 );
and ( n70900 , n70897 , n70899 );
and ( n70901 , n70895 , n70899 );
or ( n70902 , n70898 , n70900 , n70901 );
and ( n70903 , n70893 , n70902 );
xnor ( n70904 , n70572 , n70574 );
xnor ( n70905 , n70577 , n70579 );
and ( n70906 , n70904 , n70905 );
and ( n70907 , n60376 , n67844 );
not ( n70908 , n70907 );
and ( n70909 , n61918 , n66469 );
not ( n70910 , n70909 );
and ( n70911 , n70908 , n70910 );
and ( n70912 , n62593 , n65586 );
not ( n70913 , n70912 );
and ( n70914 , n70910 , n70913 );
and ( n70915 , n70908 , n70913 );
or ( n70916 , n70911 , n70914 , n70915 );
and ( n70917 , n70905 , n70916 );
and ( n70918 , n70904 , n70916 );
or ( n70919 , n70906 , n70917 , n70918 );
and ( n70920 , n70902 , n70919 );
and ( n70921 , n70893 , n70919 );
or ( n70922 , n70903 , n70920 , n70921 );
and ( n70923 , n68307 , n59920 );
not ( n70924 , n70923 );
and ( n70925 , n61008 , n67013 );
not ( n70926 , n70925 );
and ( n70927 , n70924 , n70926 );
and ( n70928 , n61505 , n66917 );
not ( n70929 , n70928 );
and ( n70930 , n70926 , n70929 );
and ( n70931 , n70924 , n70929 );
or ( n70932 , n70927 , n70930 , n70931 );
and ( n70933 , n70256 , n58542 );
not ( n70934 , n70933 );
and ( n70935 , n65177 , n62998 );
not ( n70936 , n70935 );
or ( n70937 , n70934 , n70936 );
and ( n70938 , n70932 , n70937 );
and ( n70939 , n51298 , n54535 );
and ( n70940 , n51077 , n54533 );
nor ( n70941 , n70939 , n70940 );
xnor ( n70942 , n70941 , n54237 );
and ( n70943 , n53922 , n51750 );
and ( n70944 , n53639 , n51748 );
nor ( n70945 , n70943 , n70944 );
xnor ( n70946 , n70945 , n51520 );
and ( n70947 , n70942 , n70946 );
and ( n70948 , n70937 , n70947 );
and ( n70949 , n70932 , n70947 );
or ( n70950 , n70938 , n70948 , n70949 );
and ( n70951 , n60821 , n67411 );
not ( n70952 , n70951 );
and ( n70953 , n67343 , n60711 );
not ( n70954 , n70953 );
and ( n70955 , n70952 , n70954 );
and ( n70956 , n49570 , n57187 );
and ( n70957 , n49374 , n57184 );
nor ( n70958 , n70956 , n70957 );
xnor ( n70959 , n70958 , n56175 );
and ( n70960 , n49976 , n56503 );
and ( n70961 , n49781 , n56501 );
nor ( n70962 , n70960 , n70961 );
xnor ( n70963 , n70962 , n56178 );
and ( n70964 , n70959 , n70963 );
and ( n70965 , n50404 , n55851 );
and ( n70966 , n50195 , n55849 );
nor ( n70967 , n70965 , n70966 );
xnor ( n70968 , n70967 , n55506 );
and ( n70969 , n70963 , n70968 );
and ( n70970 , n70959 , n70968 );
or ( n70971 , n70964 , n70969 , n70970 );
and ( n70972 , n70955 , n70971 );
and ( n70973 , n50726 , n55159 );
and ( n70974 , n50625 , n55157 );
nor ( n70975 , n70973 , n70974 );
xnor ( n70976 , n70975 , n54864 );
and ( n70977 , n51734 , n53928 );
and ( n70978 , n51510 , n53926 );
nor ( n70979 , n70977 , n70978 );
xnor ( n70980 , n70979 , n53652 );
and ( n70981 , n70976 , n70980 );
and ( n70982 , n52332 , n53357 );
and ( n70983 , n52082 , n53355 );
nor ( n70984 , n70982 , n70983 );
xnor ( n70985 , n70984 , n53060 );
and ( n70986 , n70980 , n70985 );
and ( n70987 , n70976 , n70985 );
or ( n70988 , n70981 , n70986 , n70987 );
and ( n70989 , n70971 , n70988 );
and ( n70990 , n70955 , n70988 );
or ( n70991 , n70972 , n70989 , n70990 );
and ( n70992 , n70950 , n70991 );
and ( n70993 , n52790 , n52799 );
and ( n70994 , n52612 , n52797 );
nor ( n70995 , n70993 , n70994 );
xnor ( n70996 , n70995 , n52538 );
and ( n70997 , n53328 , n52269 );
and ( n70998 , n53041 , n52267 );
nor ( n70999 , n70997 , n70998 );
xnor ( n71000 , n70999 , n52008 );
and ( n71001 , n70996 , n71000 );
and ( n71002 , n54604 , n51221 );
and ( n71003 , n54227 , n51219 );
nor ( n71004 , n71002 , n71003 );
xnor ( n71005 , n71004 , n51000 );
and ( n71006 , n71000 , n71005 );
and ( n71007 , n70996 , n71005 );
or ( n71008 , n71001 , n71006 , n71007 );
and ( n71009 , n55143 , n50783 );
and ( n71010 , n54942 , n50781 );
nor ( n71011 , n71009 , n71010 );
xnor ( n71012 , n71011 , n50557 );
and ( n71013 , n55756 , n50338 );
and ( n71014 , n55497 , n50336 );
nor ( n71015 , n71013 , n71014 );
xnor ( n71016 , n71015 , n50111 );
and ( n71017 , n71012 , n71016 );
and ( n71018 , n56388 , n49896 );
and ( n71019 , n56255 , n49894 );
nor ( n71020 , n71018 , n71019 );
xnor ( n71021 , n71020 , n49711 );
and ( n71022 , n71016 , n71021 );
and ( n71023 , n71012 , n71021 );
or ( n71024 , n71017 , n71022 , n71023 );
and ( n71025 , n71008 , n71024 );
and ( n71026 , n57063 , n49513 );
and ( n71027 , n56915 , n49511 );
nor ( n71028 , n71026 , n71027 );
xnor ( n71029 , n71028 , n49310 );
and ( n71030 , n57063 , n49511 );
not ( n71031 , n71030 );
and ( n71032 , n71031 , n49310 );
and ( n71033 , n71029 , n71032 );
xor ( n71034 , n45364 , n45529 );
buf ( n71035 , n71034 );
buf ( n71036 , n71035 );
buf ( n71037 , n71036 );
and ( n71038 , n71032 , n71037 );
and ( n71039 , n71029 , n71037 );
or ( n71040 , n71033 , n71038 , n71039 );
and ( n71041 , n71024 , n71040 );
and ( n71042 , n71008 , n71040 );
or ( n71043 , n71025 , n71041 , n71042 );
and ( n71044 , n70991 , n71043 );
and ( n71045 , n70950 , n71043 );
or ( n71046 , n70992 , n71044 , n71045 );
and ( n71047 , n70922 , n71046 );
and ( n71048 , n69303 , n59207 );
not ( n71049 , n71048 );
and ( n71050 , n69059 , n59611 );
not ( n71051 , n71050 );
and ( n71052 , n71049 , n71051 );
and ( n71053 , n66980 , n61015 );
not ( n71054 , n71053 );
and ( n71055 , n71051 , n71054 );
and ( n71056 , n71049 , n71054 );
or ( n71057 , n71052 , n71055 , n71056 );
and ( n71058 , n66720 , n61481 );
not ( n71059 , n71058 );
and ( n71060 , n66415 , n61914 );
not ( n71061 , n71060 );
and ( n71062 , n71059 , n71061 );
and ( n71063 , n65678 , n62151 );
not ( n71064 , n71063 );
and ( n71065 , n71061 , n71064 );
and ( n71066 , n71059 , n71064 );
or ( n71067 , n71062 , n71065 , n71066 );
and ( n71068 , n71057 , n71067 );
xor ( n71069 , n70585 , n70589 );
xor ( n71070 , n71069 , n70594 );
and ( n71071 , n71067 , n71070 );
and ( n71072 , n71057 , n71070 );
or ( n71073 , n71068 , n71071 , n71072 );
xor ( n71074 , n70604 , n70608 );
xor ( n71075 , n71074 , n70613 );
xor ( n71076 , n70620 , n70624 );
xor ( n71077 , n71076 , n70629 );
and ( n71078 , n71075 , n71077 );
xor ( n71079 , n70637 , n70641 );
xor ( n71080 , n71079 , n70646 );
and ( n71081 , n71077 , n71080 );
and ( n71082 , n71075 , n71080 );
or ( n71083 , n71078 , n71081 , n71082 );
and ( n71084 , n71073 , n71083 );
buf ( n71085 , n70472 );
xor ( n71086 , n71085 , n70474 );
and ( n71087 , n71083 , n71086 );
and ( n71088 , n71073 , n71086 );
or ( n71089 , n71084 , n71087 , n71088 );
and ( n71090 , n71046 , n71089 );
and ( n71091 , n70922 , n71089 );
or ( n71092 , n71047 , n71090 , n71091 );
and ( n71093 , n70882 , n71092 );
and ( n71094 , n70819 , n71092 );
or ( n71095 , n70883 , n71093 , n71094 );
and ( n71096 , n70816 , n71095 );
and ( n71097 , n70814 , n71095 );
or ( n71098 , n70817 , n71096 , n71097 );
xor ( n71099 , n70479 , n70481 );
xor ( n71100 , n71099 , n70484 );
xor ( n71101 , n70492 , n70493 );
xor ( n71102 , n71101 , n70495 );
and ( n71103 , n71100 , n71102 );
xor ( n71104 , n70508 , n70518 );
xor ( n71105 , n71104 , n70529 );
and ( n71106 , n71102 , n71105 );
and ( n71107 , n71100 , n71105 );
or ( n71108 , n71103 , n71106 , n71107 );
xor ( n71109 , n70543 , n70553 );
xor ( n71110 , n71109 , n70563 );
xor ( n71111 , n70575 , n70580 );
xor ( n71112 , n71111 , n70597 );
and ( n71113 , n71110 , n71112 );
xor ( n71114 , n70616 , n70632 );
xor ( n71115 , n71114 , n70649 );
and ( n71116 , n71112 , n71115 );
and ( n71117 , n71110 , n71115 );
or ( n71118 , n71113 , n71116 , n71117 );
and ( n71119 , n71108 , n71118 );
xor ( n71120 , n70665 , n70671 );
xor ( n71121 , n71120 , n70674 );
xor ( n71122 , n70686 , n70688 );
xor ( n71123 , n71122 , n70691 );
and ( n71124 , n71121 , n71123 );
xor ( n71125 , n70696 , n70698 );
xor ( n71126 , n71125 , n70701 );
and ( n71127 , n71123 , n71126 );
and ( n71128 , n71121 , n71126 );
or ( n71129 , n71124 , n71127 , n71128 );
and ( n71130 , n71118 , n71129 );
and ( n71131 , n71108 , n71129 );
or ( n71132 , n71119 , n71130 , n71131 );
xor ( n71133 , n70420 , n70422 );
xor ( n71134 , n71133 , n70425 );
xor ( n71135 , n70431 , n70432 );
xor ( n71136 , n71135 , n70459 );
and ( n71137 , n71134 , n71136 );
xor ( n71138 , n70470 , n70476 );
xor ( n71139 , n71138 , n70487 );
and ( n71140 , n71136 , n71139 );
and ( n71141 , n71134 , n71139 );
or ( n71142 , n71137 , n71140 , n71141 );
and ( n71143 , n71132 , n71142 );
xor ( n71144 , n70498 , n70532 );
xor ( n71145 , n71144 , n70566 );
xor ( n71146 , n70600 , n70652 );
xor ( n71147 , n71146 , n70677 );
and ( n71148 , n71145 , n71147 );
xor ( n71149 , n70694 , n70704 );
xor ( n71150 , n71149 , n70707 );
and ( n71151 , n71147 , n71150 );
and ( n71152 , n71145 , n71150 );
or ( n71153 , n71148 , n71151 , n71152 );
and ( n71154 , n71142 , n71153 );
and ( n71155 , n71132 , n71153 );
or ( n71156 , n71143 , n71154 , n71155 );
xor ( n71157 , n70405 , n70407 );
xor ( n71158 , n71157 , n70410 );
xor ( n71159 , n70418 , n70428 );
xor ( n71160 , n71159 , n70462 );
and ( n71161 , n71158 , n71160 );
xor ( n71162 , n70490 , n70569 );
xor ( n71163 , n71162 , n70680 );
and ( n71164 , n71160 , n71163 );
and ( n71165 , n71158 , n71163 );
or ( n71166 , n71161 , n71164 , n71165 );
and ( n71167 , n71156 , n71166 );
xor ( n71168 , n70710 , n70720 );
xor ( n71169 , n71168 , n70731 );
xor ( n71170 , n70751 , n70753 );
xor ( n71171 , n71170 , n70756 );
and ( n71172 , n71169 , n71171 );
xor ( n71173 , n70761 , n70763 );
xor ( n71174 , n71173 , n70766 );
and ( n71175 , n71171 , n71174 );
and ( n71176 , n71169 , n71174 );
or ( n71177 , n71172 , n71175 , n71176 );
and ( n71178 , n71166 , n71177 );
and ( n71179 , n71156 , n71177 );
or ( n71180 , n71167 , n71178 , n71179 );
and ( n71181 , n71098 , n71180 );
xor ( n71182 , n70400 , n70402 );
xor ( n71183 , n71182 , n70413 );
xor ( n71184 , n70465 , n70683 );
xor ( n71185 , n71184 , n70734 );
and ( n71186 , n71183 , n71185 );
xor ( n71187 , n70759 , n70769 );
xor ( n71188 , n71187 , n70772 );
and ( n71189 , n71185 , n71188 );
and ( n71190 , n71183 , n71188 );
or ( n71191 , n71186 , n71189 , n71190 );
and ( n71192 , n71180 , n71191 );
and ( n71193 , n71098 , n71191 );
or ( n71194 , n71181 , n71192 , n71193 );
and ( n71195 , n70812 , n71194 );
xor ( n71196 , n70398 , n70416 );
xor ( n71197 , n71196 , n70737 );
xor ( n71198 , n70775 , n70785 );
xor ( n71199 , n71198 , n70788 );
and ( n71200 , n71197 , n71199 );
xor ( n71201 , n70793 , n70795 );
xor ( n71202 , n71201 , n70798 );
and ( n71203 , n71199 , n71202 );
and ( n71204 , n71197 , n71202 );
or ( n71205 , n71200 , n71203 , n71204 );
and ( n71206 , n71194 , n71205 );
and ( n71207 , n70812 , n71205 );
or ( n71208 , n71195 , n71206 , n71207 );
and ( n71209 , n70809 , n71208 );
and ( n71210 , n70807 , n71208 );
or ( n71211 , n70810 , n71209 , n71210 );
and ( n71212 , n70748 , n71211 );
and ( n71213 , n70746 , n71211 );
or ( n71214 , n70749 , n71212 , n71213 );
and ( n71215 , n70386 , n71214 );
xor ( n71216 , n70388 , n70390 );
xor ( n71217 , n71216 , n70743 );
xor ( n71218 , n70393 , n70395 );
xor ( n71219 , n71218 , n70740 );
xor ( n71220 , n70791 , n70801 );
xor ( n71221 , n71220 , n70804 );
and ( n71222 , n71219 , n71221 );
xor ( n71223 , n70777 , n70779 );
xor ( n71224 , n71223 , n70782 );
xor ( n71225 , n70712 , n70714 );
xor ( n71226 , n71225 , n70717 );
xor ( n71227 , n70723 , n70725 );
xor ( n71228 , n71227 , n70728 );
and ( n71229 , n71226 , n71228 );
xor ( n71230 , n70839 , n70857 );
and ( n71231 , n63492 , n65210 );
not ( n71232 , n71231 );
and ( n71233 , n65177 , n63679 );
not ( n71234 , n71233 );
and ( n71235 , n71232 , n71234 );
and ( n71236 , n59908 , n68610 );
not ( n71237 , n71236 );
and ( n71238 , n71235 , n71237 );
and ( n71239 , n62377 , n66005 );
not ( n71240 , n71239 );
and ( n71241 , n71237 , n71240 );
and ( n71242 , n71235 , n71240 );
or ( n71243 , n71238 , n71241 , n71242 );
xor ( n71244 , n70445 , n70447 );
xor ( n71245 , n71244 , n70450 );
or ( n71246 , n71243 , n71245 );
and ( n71247 , n71230 , n71246 );
xor ( n71248 , n70831 , n70833 );
xor ( n71249 , n71248 , n70836 );
xor ( n71250 , n70849 , n70851 );
xor ( n71251 , n71250 , n70854 );
and ( n71252 , n71249 , n71251 );
and ( n71253 , n71246 , n71252 );
and ( n71254 , n71230 , n71252 );
or ( n71255 , n71247 , n71253 , n71254 );
and ( n71256 , n71228 , n71255 );
and ( n71257 , n71226 , n71255 );
or ( n71258 , n71229 , n71256 , n71257 );
xor ( n71259 , n70657 , n70231 );
xor ( n71260 , n71259 , n70662 );
xor ( n71261 , n70667 , n70669 );
buf ( n71262 , n71261 );
and ( n71263 , n71260 , n71262 );
xnor ( n71264 , n70873 , n70875 );
and ( n71265 , n71262 , n71264 );
and ( n71266 , n71260 , n71264 );
or ( n71267 , n71263 , n71265 , n71266 );
and ( n71268 , n68307 , n60372 );
not ( n71269 , n71268 );
and ( n71270 , n61918 , n66917 );
not ( n71271 , n71270 );
and ( n71272 , n71269 , n71271 );
and ( n71273 , n63024 , n65586 );
not ( n71274 , n71273 );
and ( n71275 , n71271 , n71274 );
and ( n71276 , n71269 , n71274 );
or ( n71277 , n71272 , n71275 , n71276 );
and ( n71278 , n59365 , n69204 );
not ( n71279 , n71278 );
and ( n71280 , n71277 , n71279 );
and ( n71281 , n59615 , n68752 );
not ( n71282 , n71281 );
and ( n71283 , n71279 , n71282 );
and ( n71284 , n71277 , n71282 );
or ( n71285 , n71280 , n71283 , n71284 );
and ( n71286 , n59615 , n69204 );
not ( n71287 , n71286 );
and ( n71288 , n59908 , n68752 );
not ( n71289 , n71288 );
and ( n71290 , n71287 , n71289 );
and ( n71291 , n62377 , n66469 );
not ( n71292 , n71291 );
and ( n71293 , n71289 , n71292 );
and ( n71294 , n71287 , n71292 );
or ( n71295 , n71290 , n71293 , n71294 );
xor ( n71296 , n70908 , n70910 );
xor ( n71297 , n71296 , n70913 );
or ( n71298 , n71295 , n71297 );
and ( n71299 , n71285 , n71298 );
and ( n71300 , n70256 , n58911 );
not ( n71301 , n71300 );
and ( n71302 , n64548 , n63766 );
not ( n71303 , n71302 );
or ( n71304 , n71301 , n71303 );
and ( n71305 , n58915 , n70108 );
not ( n71306 , n71305 );
and ( n71307 , n63987 , n64811 );
not ( n71308 , n71307 );
or ( n71309 , n71306 , n71308 );
and ( n71310 , n71304 , n71309 );
and ( n71311 , n71298 , n71310 );
and ( n71312 , n71285 , n71310 );
or ( n71313 , n71299 , n71311 , n71312 );
and ( n71314 , n71267 , n71313 );
xor ( n71315 , n70841 , n70843 );
xor ( n71316 , n71315 , n70846 );
xor ( n71317 , n70823 , n70825 );
xor ( n71318 , n71317 , n70828 );
and ( n71319 , n71316 , n71318 );
and ( n71320 , n65606 , n62868 );
not ( n71321 , n71320 );
xor ( n71322 , n70865 , n70867 );
xor ( n71323 , n71322 , n70870 );
and ( n71324 , n71321 , n71323 );
buf ( n71325 , n71324 );
and ( n71326 , n71319 , n71325 );
xor ( n71327 , n70924 , n70926 );
xor ( n71328 , n71327 , n70929 );
xnor ( n71329 , n70934 , n70936 );
and ( n71330 , n71328 , n71329 );
xor ( n71331 , n70942 , n70946 );
and ( n71332 , n71329 , n71331 );
and ( n71333 , n71328 , n71331 );
or ( n71334 , n71330 , n71332 , n71333 );
and ( n71335 , n71325 , n71334 );
and ( n71336 , n71319 , n71334 );
or ( n71337 , n71326 , n71335 , n71336 );
and ( n71338 , n71313 , n71337 );
and ( n71339 , n71267 , n71337 );
or ( n71340 , n71314 , n71338 , n71339 );
xor ( n71341 , n70952 , n70954 );
and ( n71342 , n60376 , n68610 );
not ( n71343 , n71342 );
and ( n71344 , n62593 , n66005 );
not ( n71345 , n71344 );
and ( n71346 , n71343 , n71345 );
buf ( n71347 , n64221 );
not ( n71348 , n71347 );
and ( n71349 , n71345 , n71348 );
and ( n71350 , n71343 , n71348 );
or ( n71351 , n71346 , n71349 , n71350 );
and ( n71352 , n71341 , n71351 );
and ( n71353 , n69059 , n59920 );
not ( n71354 , n71353 );
and ( n71355 , n61008 , n67411 );
not ( n71356 , n71355 );
and ( n71357 , n71354 , n71356 );
and ( n71358 , n61505 , n67013 );
not ( n71359 , n71358 );
and ( n71360 , n71356 , n71359 );
and ( n71361 , n71354 , n71359 );
or ( n71362 , n71357 , n71360 , n71361 );
and ( n71363 , n71351 , n71362 );
and ( n71364 , n71341 , n71362 );
or ( n71365 , n71352 , n71363 , n71364 );
and ( n71366 , n59365 , n69507 );
not ( n71367 , n71366 );
and ( n71368 , n69688 , n59207 );
not ( n71369 , n71368 );
and ( n71370 , n71367 , n71369 );
and ( n71371 , n60821 , n67844 );
not ( n71372 , n71371 );
and ( n71373 , n67997 , n60711 );
not ( n71374 , n71373 );
and ( n71375 , n71372 , n71374 );
and ( n71376 , n71370 , n71375 );
and ( n71377 , n49781 , n57187 );
and ( n71378 , n49570 , n57184 );
nor ( n71379 , n71377 , n71378 );
xnor ( n71380 , n71379 , n56175 );
and ( n71381 , n50195 , n56503 );
and ( n71382 , n49976 , n56501 );
nor ( n71383 , n71381 , n71382 );
xnor ( n71384 , n71383 , n56178 );
and ( n71385 , n71380 , n71384 );
and ( n71386 , n50625 , n55851 );
and ( n71387 , n50404 , n55849 );
nor ( n71388 , n71386 , n71387 );
xnor ( n71389 , n71388 , n55506 );
and ( n71390 , n71384 , n71389 );
and ( n71391 , n71380 , n71389 );
or ( n71392 , n71385 , n71390 , n71391 );
and ( n71393 , n71375 , n71392 );
and ( n71394 , n71370 , n71392 );
or ( n71395 , n71376 , n71393 , n71394 );
and ( n71396 , n71365 , n71395 );
and ( n71397 , n51077 , n55159 );
and ( n71398 , n50726 , n55157 );
nor ( n71399 , n71397 , n71398 );
xnor ( n71400 , n71399 , n54864 );
and ( n71401 , n51510 , n54535 );
and ( n71402 , n51298 , n54533 );
nor ( n71403 , n71401 , n71402 );
xnor ( n71404 , n71403 , n54237 );
and ( n71405 , n71400 , n71404 );
and ( n71406 , n52082 , n53928 );
and ( n71407 , n51734 , n53926 );
nor ( n71408 , n71406 , n71407 );
xnor ( n71409 , n71408 , n53652 );
and ( n71410 , n71404 , n71409 );
and ( n71411 , n71400 , n71409 );
or ( n71412 , n71405 , n71410 , n71411 );
and ( n71413 , n52612 , n53357 );
and ( n71414 , n52332 , n53355 );
nor ( n71415 , n71413 , n71414 );
xnor ( n71416 , n71415 , n53060 );
and ( n71417 , n53041 , n52799 );
and ( n71418 , n52790 , n52797 );
nor ( n71419 , n71417 , n71418 );
xnor ( n71420 , n71419 , n52538 );
and ( n71421 , n71416 , n71420 );
and ( n71422 , n53639 , n52269 );
and ( n71423 , n53328 , n52267 );
nor ( n71424 , n71422 , n71423 );
xnor ( n71425 , n71424 , n52008 );
and ( n71426 , n71420 , n71425 );
and ( n71427 , n71416 , n71425 );
or ( n71428 , n71421 , n71426 , n71427 );
and ( n71429 , n71412 , n71428 );
and ( n71430 , n54227 , n51750 );
and ( n71431 , n53922 , n51748 );
nor ( n71432 , n71430 , n71431 );
xnor ( n71433 , n71432 , n51520 );
and ( n71434 , n54942 , n51221 );
and ( n71435 , n54604 , n51219 );
nor ( n71436 , n71434 , n71435 );
xnor ( n71437 , n71436 , n51000 );
and ( n71438 , n71433 , n71437 );
and ( n71439 , n55497 , n50783 );
and ( n71440 , n55143 , n50781 );
nor ( n71441 , n71439 , n71440 );
xnor ( n71442 , n71441 , n50557 );
and ( n71443 , n71437 , n71442 );
and ( n71444 , n71433 , n71442 );
or ( n71445 , n71438 , n71443 , n71444 );
and ( n71446 , n71428 , n71445 );
and ( n71447 , n71412 , n71445 );
or ( n71448 , n71429 , n71446 , n71447 );
and ( n71449 , n71395 , n71448 );
and ( n71450 , n71365 , n71448 );
or ( n71451 , n71396 , n71449 , n71450 );
and ( n71452 , n56255 , n50338 );
and ( n71453 , n55756 , n50336 );
nor ( n71454 , n71452 , n71453 );
xnor ( n71455 , n71454 , n50111 );
and ( n71456 , n56915 , n49896 );
and ( n71457 , n56388 , n49894 );
nor ( n71458 , n71456 , n71457 );
xnor ( n71459 , n71458 , n49711 );
and ( n71460 , n71455 , n71459 );
and ( n71461 , n71459 , n71030 );
and ( n71462 , n71455 , n71030 );
or ( n71463 , n71460 , n71461 , n71462 );
xor ( n71464 , n45367 , n45527 );
buf ( n71465 , n71464 );
buf ( n71466 , n71465 );
buf ( n71467 , n71466 );
and ( n71468 , n67343 , n61015 );
not ( n71469 , n71468 );
and ( n71470 , n71467 , n71469 );
and ( n71471 , n66980 , n61481 );
not ( n71472 , n71471 );
and ( n71473 , n71469 , n71472 );
and ( n71474 , n71467 , n71472 );
or ( n71475 , n71470 , n71473 , n71474 );
and ( n71476 , n71463 , n71475 );
and ( n71477 , n66720 , n61914 );
not ( n71478 , n71477 );
and ( n71479 , n65678 , n62868 );
not ( n71480 , n71479 );
and ( n71481 , n71478 , n71480 );
and ( n71482 , n65606 , n62998 );
not ( n71483 , n71482 );
and ( n71484 , n71480 , n71483 );
and ( n71485 , n71478 , n71483 );
or ( n71486 , n71481 , n71484 , n71485 );
and ( n71487 , n71475 , n71486 );
and ( n71488 , n71463 , n71486 );
or ( n71489 , n71476 , n71487 , n71488 );
xor ( n71490 , n70959 , n70963 );
xor ( n71491 , n71490 , n70968 );
xor ( n71492 , n70976 , n70980 );
xor ( n71493 , n71492 , n70985 );
and ( n71494 , n71491 , n71493 );
xor ( n71495 , n70996 , n71000 );
xor ( n71496 , n71495 , n71005 );
and ( n71497 , n71493 , n71496 );
and ( n71498 , n71491 , n71496 );
or ( n71499 , n71494 , n71497 , n71498 );
and ( n71500 , n71489 , n71499 );
xor ( n71501 , n71012 , n71016 );
xor ( n71502 , n71501 , n71021 );
xor ( n71503 , n71029 , n71032 );
xor ( n71504 , n71503 , n71037 );
and ( n71505 , n71502 , n71504 );
xor ( n71506 , n71049 , n71051 );
xor ( n71507 , n71506 , n71054 );
and ( n71508 , n71504 , n71507 );
and ( n71509 , n71502 , n71507 );
or ( n71510 , n71505 , n71508 , n71509 );
and ( n71511 , n71499 , n71510 );
and ( n71512 , n71489 , n71510 );
or ( n71513 , n71500 , n71511 , n71512 );
and ( n71514 , n71451 , n71513 );
xor ( n71515 , n70885 , n70887 );
xor ( n71516 , n71515 , n70890 );
xor ( n71517 , n70895 , n70897 );
xor ( n71518 , n71517 , n70899 );
and ( n71519 , n71516 , n71518 );
xor ( n71520 , n70904 , n70905 );
xor ( n71521 , n71520 , n70916 );
and ( n71522 , n71518 , n71521 );
and ( n71523 , n71516 , n71521 );
or ( n71524 , n71519 , n71522 , n71523 );
and ( n71525 , n71513 , n71524 );
and ( n71526 , n71451 , n71524 );
or ( n71527 , n71514 , n71525 , n71526 );
and ( n71528 , n71340 , n71527 );
xor ( n71529 , n70932 , n70937 );
xor ( n71530 , n71529 , n70947 );
xor ( n71531 , n70955 , n70971 );
xor ( n71532 , n71531 , n70988 );
and ( n71533 , n71530 , n71532 );
xor ( n71534 , n71008 , n71024 );
xor ( n71535 , n71534 , n71040 );
and ( n71536 , n71532 , n71535 );
and ( n71537 , n71530 , n71535 );
or ( n71538 , n71533 , n71536 , n71537 );
xor ( n71539 , n70861 , n70862 );
xor ( n71540 , n71539 , n70876 );
and ( n71541 , n71538 , n71540 );
xor ( n71542 , n70893 , n70902 );
xor ( n71543 , n71542 , n70919 );
and ( n71544 , n71540 , n71543 );
and ( n71545 , n71538 , n71543 );
or ( n71546 , n71541 , n71544 , n71545 );
and ( n71547 , n71527 , n71546 );
and ( n71548 , n71340 , n71546 );
or ( n71549 , n71528 , n71547 , n71548 );
and ( n71550 , n71258 , n71549 );
xor ( n71551 , n70950 , n70991 );
xor ( n71552 , n71551 , n71043 );
xor ( n71553 , n71073 , n71083 );
xor ( n71554 , n71553 , n71086 );
and ( n71555 , n71552 , n71554 );
xor ( n71556 , n71100 , n71102 );
xor ( n71557 , n71556 , n71105 );
and ( n71558 , n71554 , n71557 );
and ( n71559 , n71552 , n71557 );
or ( n71560 , n71555 , n71558 , n71559 );
xor ( n71561 , n70821 , n70858 );
xor ( n71562 , n71561 , n70879 );
and ( n71563 , n71560 , n71562 );
xor ( n71564 , n70922 , n71046 );
xor ( n71565 , n71564 , n71089 );
and ( n71566 , n71562 , n71565 );
and ( n71567 , n71560 , n71565 );
or ( n71568 , n71563 , n71566 , n71567 );
and ( n71569 , n71549 , n71568 );
and ( n71570 , n71258 , n71568 );
or ( n71571 , n71550 , n71569 , n71570 );
and ( n71572 , n71224 , n71571 );
xor ( n71573 , n71108 , n71118 );
xor ( n71574 , n71573 , n71129 );
xor ( n71575 , n71134 , n71136 );
xor ( n71576 , n71575 , n71139 );
and ( n71577 , n71574 , n71576 );
xor ( n71578 , n71145 , n71147 );
xor ( n71579 , n71578 , n71150 );
and ( n71580 , n71576 , n71579 );
and ( n71581 , n71574 , n71579 );
or ( n71582 , n71577 , n71580 , n71581 );
xor ( n71583 , n70819 , n70882 );
xor ( n71584 , n71583 , n71092 );
and ( n71585 , n71582 , n71584 );
xor ( n71586 , n71132 , n71142 );
xor ( n71587 , n71586 , n71153 );
and ( n71588 , n71584 , n71587 );
and ( n71589 , n71582 , n71587 );
or ( n71590 , n71585 , n71588 , n71589 );
and ( n71591 , n71571 , n71590 );
and ( n71592 , n71224 , n71590 );
or ( n71593 , n71572 , n71591 , n71592 );
xor ( n71594 , n70814 , n70816 );
xor ( n71595 , n71594 , n71095 );
xor ( n71596 , n71156 , n71166 );
xor ( n71597 , n71596 , n71177 );
and ( n71598 , n71595 , n71597 );
xor ( n71599 , n71183 , n71185 );
xor ( n71600 , n71599 , n71188 );
and ( n71601 , n71597 , n71600 );
and ( n71602 , n71595 , n71600 );
or ( n71603 , n71598 , n71601 , n71602 );
and ( n71604 , n71593 , n71603 );
xor ( n71605 , n71098 , n71180 );
xor ( n71606 , n71605 , n71191 );
and ( n71607 , n71603 , n71606 );
and ( n71608 , n71593 , n71606 );
or ( n71609 , n71604 , n71607 , n71608 );
and ( n71610 , n71221 , n71609 );
and ( n71611 , n71219 , n71609 );
or ( n71612 , n71222 , n71610 , n71611 );
and ( n71613 , n71217 , n71612 );
xor ( n71614 , n70807 , n70809 );
xor ( n71615 , n71614 , n71208 );
and ( n71616 , n71612 , n71615 );
and ( n71617 , n71217 , n71615 );
or ( n71618 , n71613 , n71616 , n71617 );
xor ( n71619 , n70746 , n70748 );
xor ( n71620 , n71619 , n71211 );
and ( n71621 , n71618 , n71620 );
xor ( n71622 , n70812 , n71194 );
xor ( n71623 , n71622 , n71205 );
xor ( n71624 , n71197 , n71199 );
xor ( n71625 , n71624 , n71202 );
xor ( n71626 , n71158 , n71160 );
xor ( n71627 , n71626 , n71163 );
xor ( n71628 , n71169 , n71171 );
xor ( n71629 , n71628 , n71174 );
and ( n71630 , n71627 , n71629 );
xor ( n71631 , n71110 , n71112 );
xor ( n71632 , n71631 , n71115 );
xor ( n71633 , n71121 , n71123 );
xor ( n71634 , n71633 , n71126 );
and ( n71635 , n71632 , n71634 );
xor ( n71636 , n71057 , n71067 );
xor ( n71637 , n71636 , n71070 );
xor ( n71638 , n71075 , n71077 );
xor ( n71639 , n71638 , n71080 );
and ( n71640 , n71637 , n71639 );
xnor ( n71641 , n71243 , n71245 );
and ( n71642 , n71639 , n71641 );
and ( n71643 , n71637 , n71641 );
or ( n71644 , n71640 , n71642 , n71643 );
and ( n71645 , n71634 , n71644 );
and ( n71646 , n71632 , n71644 );
or ( n71647 , n71635 , n71645 , n71646 );
xor ( n71648 , n71249 , n71251 );
xor ( n71649 , n71059 , n71061 );
xor ( n71650 , n71649 , n71064 );
xor ( n71651 , n71235 , n71237 );
xor ( n71652 , n71651 , n71240 );
and ( n71653 , n71650 , n71652 );
xor ( n71654 , n71277 , n71279 );
xor ( n71655 , n71654 , n71282 );
and ( n71656 , n71652 , n71655 );
and ( n71657 , n71650 , n71655 );
or ( n71658 , n71653 , n71656 , n71657 );
and ( n71659 , n71648 , n71658 );
xnor ( n71660 , n71295 , n71297 );
xor ( n71661 , n71304 , n71309 );
and ( n71662 , n71660 , n71661 );
xor ( n71663 , n71316 , n71318 );
and ( n71664 , n71661 , n71663 );
and ( n71665 , n71660 , n71663 );
or ( n71666 , n71662 , n71664 , n71665 );
and ( n71667 , n71658 , n71666 );
and ( n71668 , n71648 , n71666 );
or ( n71669 , n71659 , n71667 , n71668 );
and ( n71670 , n69059 , n60372 );
not ( n71671 , n71670 );
and ( n71672 , n66415 , n62868 );
not ( n71673 , n71672 );
and ( n71674 , n71671 , n71673 );
and ( n71675 , n63024 , n66005 );
not ( n71676 , n71675 );
and ( n71677 , n71673 , n71676 );
and ( n71678 , n71671 , n71676 );
or ( n71679 , n71674 , n71677 , n71678 );
and ( n71680 , n69303 , n59611 );
not ( n71681 , n71680 );
and ( n71682 , n71679 , n71681 );
and ( n71683 , n66415 , n62151 );
not ( n71684 , n71683 );
and ( n71685 , n71681 , n71684 );
and ( n71686 , n71679 , n71684 );
or ( n71687 , n71682 , n71685 , n71686 );
and ( n71688 , n66980 , n61914 );
not ( n71689 , n71688 );
and ( n71690 , n65177 , n63766 );
not ( n71691 , n71690 );
and ( n71692 , n71689 , n71691 );
and ( n71693 , n61918 , n67013 );
not ( n71694 , n71693 );
and ( n71695 , n63987 , n65210 );
not ( n71696 , n71695 );
and ( n71697 , n71694 , n71696 );
and ( n71698 , n71692 , n71697 );
and ( n71699 , n71687 , n71698 );
xnor ( n71700 , n71301 , n71303 );
xnor ( n71701 , n71306 , n71308 );
and ( n71702 , n71700 , n71701 );
and ( n71703 , n71698 , n71702 );
and ( n71704 , n71687 , n71702 );
or ( n71705 , n71699 , n71703 , n71704 );
xor ( n71706 , n71343 , n71345 );
xor ( n71707 , n71706 , n71348 );
xor ( n71708 , n71287 , n71289 );
xor ( n71709 , n71708 , n71292 );
and ( n71710 , n71707 , n71709 );
buf ( n71711 , n71710 );
xor ( n71712 , n71269 , n71271 );
xor ( n71713 , n71712 , n71274 );
xor ( n71714 , n71354 , n71356 );
xor ( n71715 , n71714 , n71359 );
and ( n71716 , n71713 , n71715 );
xor ( n71717 , n71367 , n71369 );
and ( n71718 , n71715 , n71717 );
and ( n71719 , n71713 , n71717 );
or ( n71720 , n71716 , n71718 , n71719 );
and ( n71721 , n71711 , n71720 );
xor ( n71722 , n71372 , n71374 );
xor ( n71723 , n71232 , n71234 );
and ( n71724 , n71722 , n71723 );
and ( n71725 , n59615 , n69507 );
not ( n71726 , n71725 );
and ( n71727 , n59908 , n69204 );
not ( n71728 , n71727 );
and ( n71729 , n71726 , n71728 );
and ( n71730 , n62377 , n66917 );
not ( n71731 , n71730 );
and ( n71732 , n71728 , n71731 );
and ( n71733 , n71726 , n71731 );
or ( n71734 , n71729 , n71732 , n71733 );
and ( n71735 , n71723 , n71734 );
and ( n71736 , n71722 , n71734 );
or ( n71737 , n71724 , n71735 , n71736 );
and ( n71738 , n71720 , n71737 );
and ( n71739 , n71711 , n71737 );
or ( n71740 , n71721 , n71738 , n71739 );
and ( n71741 , n71705 , n71740 );
and ( n71742 , n60376 , n68752 );
not ( n71743 , n71742 );
and ( n71744 , n61505 , n67411 );
not ( n71745 , n71744 );
and ( n71746 , n71743 , n71745 );
and ( n71747 , n62593 , n66469 );
not ( n71748 , n71747 );
and ( n71749 , n71745 , n71748 );
and ( n71750 , n71743 , n71748 );
or ( n71751 , n71746 , n71749 , n71750 );
and ( n71752 , n67997 , n61015 );
not ( n71753 , n71752 );
and ( n71754 , n67343 , n61481 );
not ( n71755 , n71754 );
or ( n71756 , n71753 , n71755 );
and ( n71757 , n71751 , n71756 );
and ( n71758 , n50726 , n55851 );
and ( n71759 , n50625 , n55849 );
nor ( n71760 , n71758 , n71759 );
xnor ( n71761 , n71760 , n55506 );
and ( n71762 , n51734 , n54535 );
and ( n71763 , n51510 , n54533 );
nor ( n71764 , n71762 , n71763 );
xnor ( n71765 , n71764 , n54237 );
and ( n71766 , n71761 , n71765 );
and ( n71767 , n71756 , n71766 );
and ( n71768 , n71751 , n71766 );
or ( n71769 , n71757 , n71767 , n71768 );
and ( n71770 , n60821 , n68610 );
not ( n71771 , n71770 );
and ( n71772 , n68307 , n60711 );
not ( n71773 , n71772 );
and ( n71774 , n71771 , n71773 );
and ( n71775 , n63492 , n65586 );
not ( n71776 , n71775 );
and ( n71777 , n65606 , n63679 );
not ( n71778 , n71777 );
and ( n71779 , n71776 , n71778 );
and ( n71780 , n71774 , n71779 );
and ( n71781 , n64221 , n64811 );
not ( n71782 , n71781 );
and ( n71783 , n64548 , n64412 );
not ( n71784 , n71783 );
and ( n71785 , n71782 , n71784 );
and ( n71786 , n71779 , n71785 );
and ( n71787 , n71774 , n71785 );
or ( n71788 , n71780 , n71786 , n71787 );
and ( n71789 , n71769 , n71788 );
and ( n71790 , n49976 , n57187 );
and ( n71791 , n49781 , n57184 );
nor ( n71792 , n71790 , n71791 );
xnor ( n71793 , n71792 , n56175 );
and ( n71794 , n50404 , n56503 );
and ( n71795 , n50195 , n56501 );
nor ( n71796 , n71794 , n71795 );
xnor ( n71797 , n71796 , n56178 );
and ( n71798 , n71793 , n71797 );
and ( n71799 , n51298 , n55159 );
and ( n71800 , n51077 , n55157 );
nor ( n71801 , n71799 , n71800 );
xnor ( n71802 , n71801 , n54864 );
and ( n71803 , n71797 , n71802 );
and ( n71804 , n71793 , n71802 );
or ( n71805 , n71798 , n71803 , n71804 );
and ( n71806 , n52790 , n53357 );
and ( n71807 , n52612 , n53355 );
nor ( n71808 , n71806 , n71807 );
xnor ( n71809 , n71808 , n53060 );
and ( n71810 , n53328 , n52799 );
and ( n71811 , n53041 , n52797 );
nor ( n71812 , n71810 , n71811 );
xnor ( n71813 , n71812 , n52538 );
and ( n71814 , n71809 , n71813 );
and ( n71815 , n54604 , n51750 );
and ( n71816 , n54227 , n51748 );
nor ( n71817 , n71815 , n71816 );
xnor ( n71818 , n71817 , n51520 );
and ( n71819 , n71813 , n71818 );
and ( n71820 , n71809 , n71818 );
or ( n71821 , n71814 , n71819 , n71820 );
and ( n71822 , n71805 , n71821 );
and ( n71823 , n55143 , n51221 );
and ( n71824 , n54942 , n51219 );
nor ( n71825 , n71823 , n71824 );
xnor ( n71826 , n71825 , n51000 );
and ( n71827 , n55756 , n50783 );
and ( n71828 , n55497 , n50781 );
nor ( n71829 , n71827 , n71828 );
xnor ( n71830 , n71829 , n50557 );
and ( n71831 , n71826 , n71830 );
and ( n71832 , n56388 , n50338 );
and ( n71833 , n56255 , n50336 );
nor ( n71834 , n71832 , n71833 );
xnor ( n71835 , n71834 , n50111 );
and ( n71836 , n71830 , n71835 );
and ( n71837 , n71826 , n71835 );
or ( n71838 , n71831 , n71836 , n71837 );
and ( n71839 , n71821 , n71838 );
and ( n71840 , n71805 , n71838 );
or ( n71841 , n71822 , n71839 , n71840 );
and ( n71842 , n71788 , n71841 );
and ( n71843 , n71769 , n71841 );
or ( n71844 , n71789 , n71842 , n71843 );
and ( n71845 , n71740 , n71844 );
and ( n71846 , n71705 , n71844 );
or ( n71847 , n71741 , n71845 , n71846 );
and ( n71848 , n71669 , n71847 );
and ( n71849 , n57063 , n49896 );
and ( n71850 , n56915 , n49894 );
nor ( n71851 , n71849 , n71850 );
xnor ( n71852 , n71851 , n49711 );
and ( n71853 , n57063 , n49894 );
not ( n71854 , n71853 );
and ( n71855 , n71854 , n49711 );
and ( n71856 , n71852 , n71855 );
xor ( n71857 , n45370 , n45525 );
buf ( n71858 , n71857 );
buf ( n71859 , n71858 );
buf ( n71860 , n71859 );
and ( n71861 , n71855 , n71860 );
and ( n71862 , n71852 , n71860 );
or ( n71863 , n71856 , n71861 , n71862 );
and ( n71864 , n70256 , n59207 );
not ( n71865 , n71864 );
and ( n71866 , n69688 , n59611 );
not ( n71867 , n71866 );
and ( n71868 , n71865 , n71867 );
and ( n71869 , n66720 , n62151 );
not ( n71870 , n71869 );
and ( n71871 , n71867 , n71870 );
and ( n71872 , n71865 , n71870 );
or ( n71873 , n71868 , n71871 , n71872 );
and ( n71874 , n71863 , n71873 );
xor ( n71875 , n71380 , n71384 );
xor ( n71876 , n71875 , n71389 );
and ( n71877 , n71873 , n71876 );
and ( n71878 , n71863 , n71876 );
or ( n71879 , n71874 , n71877 , n71878 );
xor ( n71880 , n71400 , n71404 );
xor ( n71881 , n71880 , n71409 );
xor ( n71882 , n71416 , n71420 );
xor ( n71883 , n71882 , n71425 );
and ( n71884 , n71881 , n71883 );
xor ( n71885 , n71433 , n71437 );
xor ( n71886 , n71885 , n71442 );
and ( n71887 , n71883 , n71886 );
and ( n71888 , n71881 , n71886 );
or ( n71889 , n71884 , n71887 , n71888 );
and ( n71890 , n71879 , n71889 );
xor ( n71891 , n71455 , n71459 );
xor ( n71892 , n71891 , n71030 );
xor ( n71893 , n71467 , n71469 );
xor ( n71894 , n71893 , n71472 );
and ( n71895 , n71892 , n71894 );
xor ( n71896 , n71478 , n71480 );
xor ( n71897 , n71896 , n71483 );
and ( n71898 , n71894 , n71897 );
and ( n71899 , n71892 , n71897 );
or ( n71900 , n71895 , n71898 , n71899 );
and ( n71901 , n71889 , n71900 );
and ( n71902 , n71879 , n71900 );
or ( n71903 , n71890 , n71901 , n71902 );
buf ( n71904 , n71321 );
xor ( n71905 , n71904 , n71323 );
xor ( n71906 , n71328 , n71329 );
xor ( n71907 , n71906 , n71331 );
and ( n71908 , n71905 , n71907 );
xor ( n71909 , n71341 , n71351 );
xor ( n71910 , n71909 , n71362 );
and ( n71911 , n71907 , n71910 );
and ( n71912 , n71905 , n71910 );
or ( n71913 , n71908 , n71911 , n71912 );
and ( n71914 , n71903 , n71913 );
xor ( n71915 , n71370 , n71375 );
xor ( n71916 , n71915 , n71392 );
xor ( n71917 , n71412 , n71428 );
xor ( n71918 , n71917 , n71445 );
and ( n71919 , n71916 , n71918 );
xor ( n71920 , n71463 , n71475 );
xor ( n71921 , n71920 , n71486 );
and ( n71922 , n71918 , n71921 );
and ( n71923 , n71916 , n71921 );
or ( n71924 , n71919 , n71922 , n71923 );
and ( n71925 , n71913 , n71924 );
and ( n71926 , n71903 , n71924 );
or ( n71927 , n71914 , n71925 , n71926 );
and ( n71928 , n71847 , n71927 );
and ( n71929 , n71669 , n71927 );
or ( n71930 , n71848 , n71928 , n71929 );
and ( n71931 , n71647 , n71930 );
xor ( n71932 , n71260 , n71262 );
xor ( n71933 , n71932 , n71264 );
xor ( n71934 , n71285 , n71298 );
xor ( n71935 , n71934 , n71310 );
and ( n71936 , n71933 , n71935 );
xor ( n71937 , n71319 , n71325 );
xor ( n71938 , n71937 , n71334 );
and ( n71939 , n71935 , n71938 );
and ( n71940 , n71933 , n71938 );
or ( n71941 , n71936 , n71939 , n71940 );
xor ( n71942 , n71365 , n71395 );
xor ( n71943 , n71942 , n71448 );
xor ( n71944 , n71489 , n71499 );
xor ( n71945 , n71944 , n71510 );
and ( n71946 , n71943 , n71945 );
xor ( n71947 , n71516 , n71518 );
xor ( n71948 , n71947 , n71521 );
and ( n71949 , n71945 , n71948 );
and ( n71950 , n71943 , n71948 );
or ( n71951 , n71946 , n71949 , n71950 );
and ( n71952 , n71941 , n71951 );
xor ( n71953 , n71230 , n71246 );
xor ( n71954 , n71953 , n71252 );
and ( n71955 , n71951 , n71954 );
and ( n71956 , n71941 , n71954 );
or ( n71957 , n71952 , n71955 , n71956 );
and ( n71958 , n71930 , n71957 );
and ( n71959 , n71647 , n71957 );
or ( n71960 , n71931 , n71958 , n71959 );
and ( n71961 , n71629 , n71960 );
and ( n71962 , n71627 , n71960 );
or ( n71963 , n71630 , n71961 , n71962 );
xor ( n71964 , n71267 , n71313 );
xor ( n71965 , n71964 , n71337 );
xor ( n71966 , n71451 , n71513 );
xor ( n71967 , n71966 , n71524 );
and ( n71968 , n71965 , n71967 );
xor ( n71969 , n71538 , n71540 );
xor ( n71970 , n71969 , n71543 );
and ( n71971 , n71967 , n71970 );
and ( n71972 , n71965 , n71970 );
or ( n71973 , n71968 , n71971 , n71972 );
xor ( n71974 , n71226 , n71228 );
xor ( n71975 , n71974 , n71255 );
and ( n71976 , n71973 , n71975 );
xor ( n71977 , n71340 , n71527 );
xor ( n71978 , n71977 , n71546 );
and ( n71979 , n71975 , n71978 );
and ( n71980 , n71973 , n71978 );
or ( n71981 , n71976 , n71979 , n71980 );
xor ( n71982 , n71258 , n71549 );
xor ( n71983 , n71982 , n71568 );
and ( n71984 , n71981 , n71983 );
xor ( n71985 , n71582 , n71584 );
xor ( n71986 , n71985 , n71587 );
and ( n71987 , n71983 , n71986 );
and ( n71988 , n71981 , n71986 );
or ( n71989 , n71984 , n71987 , n71988 );
and ( n71990 , n71963 , n71989 );
xor ( n71991 , n71224 , n71571 );
xor ( n71992 , n71991 , n71590 );
and ( n71993 , n71989 , n71992 );
and ( n71994 , n71963 , n71992 );
or ( n71995 , n71990 , n71993 , n71994 );
and ( n71996 , n71625 , n71995 );
xor ( n71997 , n71593 , n71603 );
xor ( n71998 , n71997 , n71606 );
and ( n71999 , n71995 , n71998 );
and ( n72000 , n71625 , n71998 );
or ( n72001 , n71996 , n71999 , n72000 );
and ( n72002 , n71623 , n72001 );
xor ( n72003 , n71219 , n71221 );
xor ( n72004 , n72003 , n71609 );
and ( n72005 , n72001 , n72004 );
and ( n72006 , n71623 , n72004 );
or ( n72007 , n72002 , n72005 , n72006 );
xor ( n72008 , n71217 , n71612 );
xor ( n72009 , n72008 , n71615 );
and ( n72010 , n72007 , n72009 );
xor ( n72011 , n71623 , n72001 );
xor ( n72012 , n72011 , n72004 );
xor ( n72013 , n71595 , n71597 );
xor ( n72014 , n72013 , n71600 );
xor ( n72015 , n71560 , n71562 );
xor ( n72016 , n72015 , n71565 );
xor ( n72017 , n71574 , n71576 );
xor ( n72018 , n72017 , n71579 );
and ( n72019 , n72016 , n72018 );
xor ( n72020 , n71552 , n71554 );
xor ( n72021 , n72020 , n71557 );
xor ( n72022 , n71530 , n71532 );
xor ( n72023 , n72022 , n71535 );
xor ( n72024 , n71491 , n71493 );
xor ( n72025 , n72024 , n71496 );
xor ( n72026 , n71502 , n71504 );
xor ( n72027 , n72026 , n71507 );
and ( n72028 , n72025 , n72027 );
xor ( n72029 , n71679 , n71681 );
xor ( n72030 , n72029 , n71684 );
xor ( n72031 , n71692 , n71697 );
and ( n72032 , n72030 , n72031 );
xor ( n72033 , n71700 , n71701 );
and ( n72034 , n72031 , n72033 );
and ( n72035 , n72030 , n72033 );
or ( n72036 , n72032 , n72034 , n72035 );
and ( n72037 , n72027 , n72036 );
and ( n72038 , n72025 , n72036 );
or ( n72039 , n72028 , n72037 , n72038 );
and ( n72040 , n72023 , n72039 );
and ( n72041 , n69303 , n60372 );
not ( n72042 , n72041 );
and ( n72043 , n66720 , n62868 );
not ( n72044 , n72043 );
and ( n72045 , n72042 , n72044 );
and ( n72046 , n63987 , n65586 );
not ( n72047 , n72046 );
and ( n72048 , n72044 , n72047 );
and ( n72049 , n72042 , n72047 );
or ( n72050 , n72045 , n72048 , n72049 );
and ( n72051 , n59365 , n70108 );
not ( n72052 , n72051 );
and ( n72053 , n72050 , n72052 );
and ( n72054 , n69303 , n59920 );
not ( n72055 , n72054 );
and ( n72056 , n72052 , n72055 );
and ( n72057 , n72050 , n72055 );
or ( n72058 , n72053 , n72056 , n72057 );
and ( n72059 , n64221 , n65210 );
not ( n72060 , n72059 );
buf ( n72061 , n72060 );
and ( n72062 , n61008 , n67844 );
not ( n72063 , n72062 );
or ( n72064 , n72061 , n72063 );
and ( n72065 , n72058 , n72064 );
xor ( n72066 , n71689 , n71691 );
xor ( n72067 , n71694 , n71696 );
and ( n72068 , n72066 , n72067 );
and ( n72069 , n72064 , n72068 );
and ( n72070 , n72058 , n72068 );
or ( n72071 , n72065 , n72069 , n72070 );
and ( n72072 , n65678 , n62998 );
not ( n72073 , n72072 );
xor ( n72074 , n71726 , n71728 );
xor ( n72075 , n72074 , n71731 );
and ( n72076 , n72073 , n72075 );
buf ( n72077 , n72076 );
xor ( n72078 , n71743 , n71745 );
xor ( n72079 , n72078 , n71748 );
xor ( n72080 , n71671 , n71673 );
xor ( n72081 , n72080 , n71676 );
and ( n72082 , n72079 , n72081 );
xnor ( n72083 , n71753 , n71755 );
and ( n72084 , n72081 , n72083 );
and ( n72085 , n72079 , n72083 );
or ( n72086 , n72082 , n72084 , n72085 );
and ( n72087 , n72077 , n72086 );
xor ( n72088 , n71761 , n71765 );
xor ( n72089 , n71771 , n71773 );
and ( n72090 , n72088 , n72089 );
xor ( n72091 , n71776 , n71778 );
and ( n72092 , n72089 , n72091 );
and ( n72093 , n72088 , n72091 );
or ( n72094 , n72090 , n72092 , n72093 );
and ( n72095 , n72086 , n72094 );
and ( n72096 , n72077 , n72094 );
or ( n72097 , n72087 , n72095 , n72096 );
and ( n72098 , n72071 , n72097 );
xor ( n72099 , n71782 , n71784 );
and ( n72100 , n59908 , n69507 );
not ( n72101 , n72100 );
and ( n72102 , n61008 , n68610 );
not ( n72103 , n72102 );
and ( n72104 , n72101 , n72103 );
and ( n72105 , n62377 , n67013 );
not ( n72106 , n72105 );
and ( n72107 , n72103 , n72106 );
and ( n72108 , n72101 , n72106 );
or ( n72109 , n72104 , n72107 , n72108 );
and ( n72110 , n72099 , n72109 );
and ( n72111 , n60376 , n69204 );
not ( n72112 , n72111 );
and ( n72113 , n62593 , n66917 );
not ( n72114 , n72113 );
and ( n72115 , n72112 , n72114 );
buf ( n72116 , n64548 );
not ( n72117 , n72116 );
and ( n72118 , n72114 , n72117 );
and ( n72119 , n72112 , n72117 );
or ( n72120 , n72115 , n72118 , n72119 );
and ( n72121 , n72109 , n72120 );
and ( n72122 , n72099 , n72120 );
or ( n72123 , n72110 , n72121 , n72122 );
and ( n72124 , n69688 , n59920 );
not ( n72125 , n72124 );
and ( n72126 , n68307 , n61015 );
not ( n72127 , n72126 );
and ( n72128 , n72125 , n72127 );
and ( n72129 , n61505 , n67844 );
not ( n72130 , n72129 );
and ( n72131 , n72127 , n72130 );
and ( n72132 , n72125 , n72130 );
or ( n72133 , n72128 , n72131 , n72132 );
and ( n72134 , n59615 , n70108 );
not ( n72135 , n72134 );
and ( n72136 , n60821 , n68752 );
not ( n72137 , n72136 );
and ( n72138 , n72135 , n72137 );
and ( n72139 , n72137 , n72059 );
and ( n72140 , n72135 , n72059 );
or ( n72141 , n72138 , n72139 , n72140 );
and ( n72142 , n72133 , n72141 );
and ( n72143 , n67997 , n61481 );
not ( n72144 , n72143 );
and ( n72145 , n61918 , n67411 );
not ( n72146 , n72145 );
or ( n72147 , n72144 , n72146 );
and ( n72148 , n72141 , n72147 );
and ( n72149 , n72133 , n72147 );
or ( n72150 , n72142 , n72148 , n72149 );
and ( n72151 , n72123 , n72150 );
and ( n72152 , n51077 , n55851 );
and ( n72153 , n50726 , n55849 );
nor ( n72154 , n72152 , n72153 );
xnor ( n72155 , n72154 , n55506 );
and ( n72156 , n54942 , n51750 );
and ( n72157 , n54604 , n51748 );
nor ( n72158 , n72156 , n72157 );
xnor ( n72159 , n72158 , n51520 );
and ( n72160 , n72155 , n72159 );
and ( n72161 , n70256 , n59611 );
not ( n72162 , n72161 );
and ( n72163 , n66980 , n62151 );
not ( n72164 , n72163 );
and ( n72165 , n72162 , n72164 );
and ( n72166 , n72160 , n72165 );
and ( n72167 , n63024 , n66469 );
not ( n72168 , n72167 );
and ( n72169 , n66415 , n62998 );
not ( n72170 , n72169 );
and ( n72171 , n72168 , n72170 );
and ( n72172 , n72165 , n72171 );
and ( n72173 , n72160 , n72171 );
or ( n72174 , n72166 , n72172 , n72173 );
and ( n72175 , n72150 , n72174 );
and ( n72176 , n72123 , n72174 );
or ( n72177 , n72151 , n72175 , n72176 );
and ( n72178 , n72097 , n72177 );
and ( n72179 , n72071 , n72177 );
or ( n72180 , n72098 , n72178 , n72179 );
and ( n72181 , n72039 , n72180 );
and ( n72182 , n72023 , n72180 );
or ( n72183 , n72040 , n72181 , n72182 );
and ( n72184 , n72021 , n72183 );
and ( n72185 , n63492 , n66005 );
not ( n72186 , n72185 );
and ( n72187 , n65678 , n63679 );
not ( n72188 , n72187 );
and ( n72189 , n72186 , n72188 );
and ( n72190 , n50195 , n57187 );
and ( n72191 , n49976 , n57184 );
nor ( n72192 , n72190 , n72191 );
xnor ( n72193 , n72192 , n56175 );
and ( n72194 , n50625 , n56503 );
and ( n72195 , n50404 , n56501 );
nor ( n72196 , n72194 , n72195 );
xnor ( n72197 , n72196 , n56178 );
and ( n72198 , n72193 , n72197 );
and ( n72199 , n52082 , n54535 );
and ( n72200 , n51734 , n54533 );
nor ( n72201 , n72199 , n72200 );
xnor ( n72202 , n72201 , n54237 );
and ( n72203 , n72197 , n72202 );
and ( n72204 , n72193 , n72202 );
or ( n72205 , n72198 , n72203 , n72204 );
and ( n72206 , n72189 , n72205 );
and ( n72207 , n52612 , n53928 );
and ( n72208 , n52332 , n53926 );
nor ( n72209 , n72207 , n72208 );
xnor ( n72210 , n72209 , n53652 );
and ( n72211 , n54227 , n52269 );
and ( n72212 , n53922 , n52267 );
nor ( n72213 , n72211 , n72212 );
xnor ( n72214 , n72213 , n52008 );
and ( n72215 , n72210 , n72214 );
and ( n72216 , n55497 , n51221 );
and ( n72217 , n55143 , n51219 );
nor ( n72218 , n72216 , n72217 );
xnor ( n72219 , n72218 , n51000 );
and ( n72220 , n72214 , n72219 );
and ( n72221 , n72210 , n72219 );
or ( n72222 , n72215 , n72220 , n72221 );
and ( n72223 , n72205 , n72222 );
and ( n72224 , n72189 , n72222 );
or ( n72225 , n72206 , n72223 , n72224 );
and ( n72226 , n56255 , n50783 );
and ( n72227 , n55756 , n50781 );
nor ( n72228 , n72226 , n72227 );
xnor ( n72229 , n72228 , n50557 );
and ( n72230 , n56915 , n50338 );
and ( n72231 , n56388 , n50336 );
nor ( n72232 , n72230 , n72231 );
xnor ( n72233 , n72232 , n50111 );
and ( n72234 , n72229 , n72233 );
and ( n72235 , n72233 , n71853 );
and ( n72236 , n72229 , n71853 );
or ( n72237 , n72234 , n72235 , n72236 );
xor ( n72238 , n45371 , n45524 );
buf ( n72239 , n72238 );
buf ( n72240 , n72239 );
buf ( n72241 , n72240 );
and ( n72242 , n67343 , n61914 );
not ( n72243 , n72242 );
and ( n72244 , n72241 , n72243 );
and ( n72245 , n65606 , n63766 );
not ( n72246 , n72245 );
and ( n72247 , n72243 , n72246 );
and ( n72248 , n72241 , n72246 );
or ( n72249 , n72244 , n72247 , n72248 );
and ( n72250 , n72237 , n72249 );
xor ( n72251 , n71793 , n71797 );
xor ( n72252 , n72251 , n71802 );
and ( n72253 , n72249 , n72252 );
and ( n72254 , n72237 , n72252 );
or ( n72255 , n72250 , n72253 , n72254 );
and ( n72256 , n72225 , n72255 );
xor ( n72257 , n71809 , n71813 );
xor ( n72258 , n72257 , n71818 );
xor ( n72259 , n71826 , n71830 );
xor ( n72260 , n72259 , n71835 );
and ( n72261 , n72258 , n72260 );
xor ( n72262 , n71852 , n71855 );
xor ( n72263 , n72262 , n71860 );
and ( n72264 , n72260 , n72263 );
and ( n72265 , n72258 , n72263 );
or ( n72266 , n72261 , n72264 , n72265 );
and ( n72267 , n72255 , n72266 );
and ( n72268 , n72225 , n72266 );
or ( n72269 , n72256 , n72267 , n72268 );
buf ( n72270 , n71707 );
xor ( n72271 , n72270 , n71709 );
xor ( n72272 , n71713 , n71715 );
xor ( n72273 , n72272 , n71717 );
and ( n72274 , n72271 , n72273 );
xor ( n72275 , n71722 , n71723 );
xor ( n72276 , n72275 , n71734 );
and ( n72277 , n72273 , n72276 );
and ( n72278 , n72271 , n72276 );
or ( n72279 , n72274 , n72277 , n72278 );
and ( n72280 , n72269 , n72279 );
xor ( n72281 , n71751 , n71756 );
xor ( n72282 , n72281 , n71766 );
xor ( n72283 , n71774 , n71779 );
xor ( n72284 , n72283 , n71785 );
and ( n72285 , n72282 , n72284 );
xor ( n72286 , n71805 , n71821 );
xor ( n72287 , n72286 , n71838 );
and ( n72288 , n72284 , n72287 );
and ( n72289 , n72282 , n72287 );
or ( n72290 , n72285 , n72288 , n72289 );
and ( n72291 , n72279 , n72290 );
and ( n72292 , n72269 , n72290 );
or ( n72293 , n72280 , n72291 , n72292 );
xor ( n72294 , n71863 , n71873 );
xor ( n72295 , n72294 , n71876 );
xor ( n72296 , n71881 , n71883 );
xor ( n72297 , n72296 , n71886 );
and ( n72298 , n72295 , n72297 );
xor ( n72299 , n71892 , n71894 );
xor ( n72300 , n72299 , n71897 );
and ( n72301 , n72297 , n72300 );
and ( n72302 , n72295 , n72300 );
or ( n72303 , n72298 , n72301 , n72302 );
xor ( n72304 , n71650 , n71652 );
xor ( n72305 , n72304 , n71655 );
and ( n72306 , n72303 , n72305 );
xor ( n72307 , n71660 , n71661 );
xor ( n72308 , n72307 , n71663 );
and ( n72309 , n72305 , n72308 );
and ( n72310 , n72303 , n72308 );
or ( n72311 , n72306 , n72309 , n72310 );
and ( n72312 , n72293 , n72311 );
xor ( n72313 , n71687 , n71698 );
xor ( n72314 , n72313 , n71702 );
xor ( n72315 , n71711 , n71720 );
xor ( n72316 , n72315 , n71737 );
and ( n72317 , n72314 , n72316 );
xor ( n72318 , n71769 , n71788 );
xor ( n72319 , n72318 , n71841 );
and ( n72320 , n72316 , n72319 );
and ( n72321 , n72314 , n72319 );
or ( n72322 , n72317 , n72320 , n72321 );
and ( n72323 , n72311 , n72322 );
and ( n72324 , n72293 , n72322 );
or ( n72325 , n72312 , n72323 , n72324 );
and ( n72326 , n72183 , n72325 );
and ( n72327 , n72021 , n72325 );
or ( n72328 , n72184 , n72326 , n72327 );
and ( n72329 , n72018 , n72328 );
and ( n72330 , n72016 , n72328 );
or ( n72331 , n72019 , n72329 , n72330 );
xor ( n72332 , n71879 , n71889 );
xor ( n72333 , n72332 , n71900 );
xor ( n72334 , n71905 , n71907 );
xor ( n72335 , n72334 , n71910 );
and ( n72336 , n72333 , n72335 );
xor ( n72337 , n71916 , n71918 );
xor ( n72338 , n72337 , n71921 );
and ( n72339 , n72335 , n72338 );
and ( n72340 , n72333 , n72338 );
or ( n72341 , n72336 , n72339 , n72340 );
xor ( n72342 , n71637 , n71639 );
xor ( n72343 , n72342 , n71641 );
and ( n72344 , n72341 , n72343 );
xor ( n72345 , n71648 , n71658 );
xor ( n72346 , n72345 , n71666 );
and ( n72347 , n72343 , n72346 );
and ( n72348 , n72341 , n72346 );
or ( n72349 , n72344 , n72347 , n72348 );
xor ( n72350 , n71705 , n71740 );
xor ( n72351 , n72350 , n71844 );
xor ( n72352 , n71903 , n71913 );
xor ( n72353 , n72352 , n71924 );
and ( n72354 , n72351 , n72353 );
xor ( n72355 , n71933 , n71935 );
xor ( n72356 , n72355 , n71938 );
and ( n72357 , n72353 , n72356 );
and ( n72358 , n72351 , n72356 );
or ( n72359 , n72354 , n72357 , n72358 );
and ( n72360 , n72349 , n72359 );
xor ( n72361 , n71632 , n71634 );
xor ( n72362 , n72361 , n71644 );
and ( n72363 , n72359 , n72362 );
and ( n72364 , n72349 , n72362 );
or ( n72365 , n72360 , n72363 , n72364 );
xor ( n72366 , n71669 , n71847 );
xor ( n72367 , n72366 , n71927 );
xor ( n72368 , n71941 , n71951 );
xor ( n72369 , n72368 , n71954 );
and ( n72370 , n72367 , n72369 );
xor ( n72371 , n71965 , n71967 );
xor ( n72372 , n72371 , n71970 );
and ( n72373 , n72369 , n72372 );
and ( n72374 , n72367 , n72372 );
or ( n72375 , n72370 , n72373 , n72374 );
and ( n72376 , n72365 , n72375 );
xor ( n72377 , n71647 , n71930 );
xor ( n72378 , n72377 , n71957 );
and ( n72379 , n72375 , n72378 );
and ( n72380 , n72365 , n72378 );
or ( n72381 , n72376 , n72379 , n72380 );
and ( n72382 , n72331 , n72381 );
xor ( n72383 , n71627 , n71629 );
xor ( n72384 , n72383 , n71960 );
and ( n72385 , n72381 , n72384 );
and ( n72386 , n72331 , n72384 );
or ( n72387 , n72382 , n72385 , n72386 );
and ( n72388 , n72014 , n72387 );
xor ( n72389 , n71963 , n71989 );
xor ( n72390 , n72389 , n71992 );
and ( n72391 , n72387 , n72390 );
and ( n72392 , n72014 , n72390 );
or ( n72393 , n72388 , n72391 , n72392 );
xor ( n72394 , n71625 , n71995 );
xor ( n72395 , n72394 , n71998 );
and ( n72396 , n72393 , n72395 );
xor ( n72397 , n71981 , n71983 );
xor ( n72398 , n72397 , n71986 );
xor ( n72399 , n71973 , n71975 );
xor ( n72400 , n72399 , n71978 );
xor ( n72401 , n71943 , n71945 );
xor ( n72402 , n72401 , n71948 );
xor ( n72403 , n71865 , n71867 );
xor ( n72404 , n72403 , n71870 );
xor ( n72405 , n72050 , n72052 );
xor ( n72406 , n72405 , n72055 );
and ( n72407 , n72404 , n72406 );
xnor ( n72408 , n72061 , n72063 );
and ( n72409 , n72406 , n72408 );
and ( n72410 , n72404 , n72408 );
or ( n72411 , n72407 , n72409 , n72410 );
xor ( n72412 , n72066 , n72067 );
and ( n72413 , n59908 , n70108 );
not ( n72414 , n72413 );
and ( n72415 , n70256 , n59920 );
not ( n72416 , n72415 );
and ( n72417 , n72414 , n72416 );
and ( n72418 , n62377 , n67411 );
not ( n72419 , n72418 );
and ( n72420 , n67343 , n62151 );
not ( n72421 , n72420 );
and ( n72422 , n72419 , n72421 );
and ( n72423 , n72417 , n72422 );
and ( n72424 , n53041 , n53357 );
and ( n72425 , n52790 , n53355 );
nor ( n72426 , n72424 , n72425 );
xnor ( n72427 , n72426 , n53060 );
and ( n72428 , n72422 , n72427 );
and ( n72429 , n72417 , n72427 );
or ( n72430 , n72423 , n72428 , n72429 );
and ( n72431 , n72412 , n72430 );
and ( n72432 , n69688 , n60372 );
not ( n72433 , n72432 );
and ( n72434 , n66980 , n62868 );
not ( n72435 , n72434 );
and ( n72436 , n72433 , n72435 );
and ( n72437 , n65606 , n64412 );
not ( n72438 , n72437 );
and ( n72439 , n72435 , n72438 );
and ( n72440 , n72433 , n72438 );
or ( n72441 , n72436 , n72439 , n72440 );
and ( n72442 , n69059 , n60711 );
not ( n72443 , n72442 );
and ( n72444 , n72441 , n72443 );
xor ( n72445 , n72042 , n72044 );
xor ( n72446 , n72445 , n72047 );
and ( n72447 , n72443 , n72446 );
and ( n72448 , n72441 , n72446 );
or ( n72449 , n72444 , n72447 , n72448 );
and ( n72450 , n72430 , n72449 );
and ( n72451 , n72412 , n72449 );
or ( n72452 , n72431 , n72450 , n72451 );
and ( n72453 , n72411 , n72452 );
and ( n72454 , n65177 , n64412 );
not ( n72455 , n72454 );
xor ( n72456 , n72101 , n72103 );
xor ( n72457 , n72456 , n72106 );
and ( n72458 , n72455 , n72457 );
buf ( n72459 , n72458 );
xor ( n72460 , n72112 , n72114 );
xor ( n72461 , n72460 , n72117 );
xor ( n72462 , n72125 , n72127 );
xor ( n72463 , n72462 , n72130 );
and ( n72464 , n72461 , n72463 );
xor ( n72465 , n72135 , n72137 );
xor ( n72466 , n72465 , n72059 );
and ( n72467 , n72463 , n72466 );
and ( n72468 , n72461 , n72466 );
or ( n72469 , n72464 , n72467 , n72468 );
and ( n72470 , n72459 , n72469 );
xnor ( n72471 , n72144 , n72146 );
xor ( n72472 , n72155 , n72159 );
and ( n72473 , n72471 , n72472 );
xor ( n72474 , n72162 , n72164 );
and ( n72475 , n72472 , n72474 );
and ( n72476 , n72471 , n72474 );
or ( n72477 , n72473 , n72475 , n72476 );
and ( n72478 , n72469 , n72477 );
and ( n72479 , n72459 , n72477 );
or ( n72480 , n72470 , n72478 , n72479 );
and ( n72481 , n72452 , n72480 );
and ( n72482 , n72411 , n72480 );
or ( n72483 , n72453 , n72481 , n72482 );
xor ( n72484 , n72168 , n72170 );
xor ( n72485 , n72186 , n72188 );
and ( n72486 , n72484 , n72485 );
and ( n72487 , n51734 , n55159 );
and ( n72488 , n51510 , n55157 );
nor ( n72489 , n72487 , n72488 );
xnor ( n72490 , n72489 , n54864 );
and ( n72491 , n52332 , n54535 );
and ( n72492 , n52082 , n54533 );
nor ( n72493 , n72491 , n72492 );
xnor ( n72494 , n72493 , n54237 );
and ( n72495 , n72490 , n72494 );
and ( n72496 , n54604 , n52269 );
and ( n72497 , n54227 , n52267 );
nor ( n72498 , n72496 , n72497 );
xnor ( n72499 , n72498 , n52008 );
and ( n72500 , n72494 , n72499 );
and ( n72501 , n72490 , n72499 );
or ( n72502 , n72495 , n72500 , n72501 );
and ( n72503 , n72485 , n72502 );
and ( n72504 , n72484 , n72502 );
or ( n72505 , n72486 , n72503 , n72504 );
and ( n72506 , n60376 , n69507 );
not ( n72507 , n72506 );
and ( n72508 , n62593 , n67013 );
not ( n72509 , n72508 );
and ( n72510 , n72507 , n72509 );
and ( n72511 , n63024 , n66917 );
not ( n72512 , n72511 );
and ( n72513 , n72509 , n72512 );
and ( n72514 , n72507 , n72512 );
or ( n72515 , n72510 , n72513 , n72514 );
and ( n72516 , n61918 , n67844 );
not ( n72517 , n72516 );
and ( n72518 , n63987 , n66005 );
not ( n72519 , n72518 );
and ( n72520 , n72517 , n72519 );
and ( n72521 , n64221 , n65586 );
not ( n72522 , n72521 );
and ( n72523 , n72519 , n72522 );
and ( n72524 , n72517 , n72522 );
or ( n72525 , n72520 , n72523 , n72524 );
and ( n72526 , n72515 , n72525 );
and ( n72527 , n67997 , n61914 );
not ( n72528 , n72527 );
and ( n72529 , n66720 , n62998 );
not ( n72530 , n72529 );
and ( n72531 , n72528 , n72530 );
and ( n72532 , n65678 , n63766 );
not ( n72533 , n72532 );
and ( n72534 , n72530 , n72533 );
and ( n72535 , n72528 , n72533 );
or ( n72536 , n72531 , n72534 , n72535 );
and ( n72537 , n72525 , n72536 );
and ( n72538 , n72515 , n72536 );
or ( n72539 , n72526 , n72537 , n72538 );
and ( n72540 , n72505 , n72539 );
and ( n72541 , n56388 , n50783 );
and ( n72542 , n56255 , n50781 );
nor ( n72543 , n72541 , n72542 );
xnor ( n72544 , n72543 , n50557 );
and ( n72545 , n57063 , n50336 );
not ( n72546 , n72545 );
and ( n72547 , n72546 , n50111 );
or ( n72548 , n72544 , n72547 );
and ( n72549 , n51298 , n55851 );
and ( n72550 , n51077 , n55849 );
nor ( n72551 , n72549 , n72550 );
xnor ( n72552 , n72551 , n55506 );
and ( n72553 , n55143 , n51750 );
and ( n72554 , n54942 , n51748 );
nor ( n72555 , n72553 , n72554 );
xnor ( n72556 , n72555 , n51520 );
and ( n72557 , n72552 , n72556 );
and ( n72558 , n72548 , n72557 );
and ( n72559 , n61008 , n68752 );
not ( n72560 , n72559 );
and ( n72561 , n69059 , n61015 );
not ( n72562 , n72561 );
and ( n72563 , n72560 , n72562 );
and ( n72564 , n72557 , n72563 );
and ( n72565 , n72548 , n72563 );
or ( n72566 , n72558 , n72564 , n72565 );
and ( n72567 , n72539 , n72566 );
and ( n72568 , n72505 , n72566 );
or ( n72569 , n72540 , n72567 , n72568 );
and ( n72570 , n63492 , n66469 );
not ( n72571 , n72570 );
and ( n72572 , n66415 , n63679 );
not ( n72573 , n72572 );
and ( n72574 , n72571 , n72573 );
and ( n72575 , n64548 , n65210 );
not ( n72576 , n72575 );
and ( n72577 , n65177 , n64811 );
not ( n72578 , n72577 );
and ( n72579 , n72576 , n72578 );
and ( n72580 , n72574 , n72579 );
and ( n72581 , n50404 , n57187 );
and ( n72582 , n50195 , n57184 );
nor ( n72583 , n72581 , n72582 );
xnor ( n72584 , n72583 , n56175 );
and ( n72585 , n50726 , n56503 );
and ( n72586 , n50625 , n56501 );
nor ( n72587 , n72585 , n72586 );
xnor ( n72588 , n72587 , n56178 );
and ( n72589 , n72584 , n72588 );
and ( n72590 , n53922 , n52799 );
and ( n72591 , n53639 , n52797 );
nor ( n72592 , n72590 , n72591 );
xnor ( n72593 , n72592 , n52538 );
and ( n72594 , n72588 , n72593 );
and ( n72595 , n72584 , n72593 );
or ( n72596 , n72589 , n72594 , n72595 );
and ( n72597 , n72579 , n72596 );
and ( n72598 , n72574 , n72596 );
or ( n72599 , n72580 , n72597 , n72598 );
and ( n72600 , n55756 , n51221 );
and ( n72601 , n55497 , n51219 );
nor ( n72602 , n72600 , n72601 );
xnor ( n72603 , n72602 , n51000 );
and ( n72604 , n57063 , n50338 );
and ( n72605 , n56915 , n50336 );
nor ( n72606 , n72604 , n72605 );
xnor ( n72607 , n72606 , n50111 );
and ( n72608 , n72603 , n72607 );
xor ( n72609 , n45374 , n45522 );
buf ( n72610 , n72609 );
buf ( n72611 , n72610 );
buf ( n72612 , n72611 );
and ( n72613 , n72607 , n72612 );
and ( n72614 , n72603 , n72612 );
or ( n72615 , n72608 , n72613 , n72614 );
xor ( n72616 , n72193 , n72197 );
xor ( n72617 , n72616 , n72202 );
and ( n72618 , n72615 , n72617 );
xor ( n72619 , n72210 , n72214 );
xor ( n72620 , n72619 , n72219 );
and ( n72621 , n72617 , n72620 );
and ( n72622 , n72615 , n72620 );
or ( n72623 , n72618 , n72621 , n72622 );
and ( n72624 , n72599 , n72623 );
buf ( n72625 , n72073 );
xor ( n72626 , n72625 , n72075 );
and ( n72627 , n72623 , n72626 );
and ( n72628 , n72599 , n72626 );
or ( n72629 , n72624 , n72627 , n72628 );
and ( n72630 , n72569 , n72629 );
xor ( n72631 , n72079 , n72081 );
xor ( n72632 , n72631 , n72083 );
xor ( n72633 , n72088 , n72089 );
xor ( n72634 , n72633 , n72091 );
and ( n72635 , n72632 , n72634 );
xor ( n72636 , n72099 , n72109 );
xor ( n72637 , n72636 , n72120 );
and ( n72638 , n72634 , n72637 );
and ( n72639 , n72632 , n72637 );
or ( n72640 , n72635 , n72638 , n72639 );
and ( n72641 , n72629 , n72640 );
and ( n72642 , n72569 , n72640 );
or ( n72643 , n72630 , n72641 , n72642 );
and ( n72644 , n72483 , n72643 );
xor ( n72645 , n72133 , n72141 );
xor ( n72646 , n72645 , n72147 );
xor ( n72647 , n72160 , n72165 );
xor ( n72648 , n72647 , n72171 );
and ( n72649 , n72646 , n72648 );
xor ( n72650 , n72189 , n72205 );
xor ( n72651 , n72650 , n72222 );
and ( n72652 , n72648 , n72651 );
and ( n72653 , n72646 , n72651 );
or ( n72654 , n72649 , n72652 , n72653 );
xor ( n72655 , n72030 , n72031 );
xor ( n72656 , n72655 , n72033 );
and ( n72657 , n72654 , n72656 );
xor ( n72658 , n72058 , n72064 );
xor ( n72659 , n72658 , n72068 );
and ( n72660 , n72656 , n72659 );
and ( n72661 , n72654 , n72659 );
or ( n72662 , n72657 , n72660 , n72661 );
and ( n72663 , n72643 , n72662 );
and ( n72664 , n72483 , n72662 );
or ( n72665 , n72644 , n72663 , n72664 );
and ( n72666 , n72402 , n72665 );
xor ( n72667 , n72077 , n72086 );
xor ( n72668 , n72667 , n72094 );
xor ( n72669 , n72123 , n72150 );
xor ( n72670 , n72669 , n72174 );
and ( n72671 , n72668 , n72670 );
xor ( n72672 , n72225 , n72255 );
xor ( n72673 , n72672 , n72266 );
and ( n72674 , n72670 , n72673 );
and ( n72675 , n72668 , n72673 );
or ( n72676 , n72671 , n72674 , n72675 );
xor ( n72677 , n72271 , n72273 );
xor ( n72678 , n72677 , n72276 );
xor ( n72679 , n72282 , n72284 );
xor ( n72680 , n72679 , n72287 );
and ( n72681 , n72678 , n72680 );
xor ( n72682 , n72295 , n72297 );
xor ( n72683 , n72682 , n72300 );
and ( n72684 , n72680 , n72683 );
and ( n72685 , n72678 , n72683 );
or ( n72686 , n72681 , n72684 , n72685 );
and ( n72687 , n72676 , n72686 );
xor ( n72688 , n72025 , n72027 );
xor ( n72689 , n72688 , n72036 );
and ( n72690 , n72686 , n72689 );
and ( n72691 , n72676 , n72689 );
or ( n72692 , n72687 , n72690 , n72691 );
and ( n72693 , n72665 , n72692 );
and ( n72694 , n72402 , n72692 );
or ( n72695 , n72666 , n72693 , n72694 );
xor ( n72696 , n72071 , n72097 );
xor ( n72697 , n72696 , n72177 );
xor ( n72698 , n72269 , n72279 );
xor ( n72699 , n72698 , n72290 );
and ( n72700 , n72697 , n72699 );
xor ( n72701 , n72303 , n72305 );
xor ( n72702 , n72701 , n72308 );
and ( n72703 , n72699 , n72702 );
and ( n72704 , n72697 , n72702 );
or ( n72705 , n72700 , n72703 , n72704 );
xor ( n72706 , n72023 , n72039 );
xor ( n72707 , n72706 , n72180 );
and ( n72708 , n72705 , n72707 );
xor ( n72709 , n72293 , n72311 );
xor ( n72710 , n72709 , n72322 );
and ( n72711 , n72707 , n72710 );
and ( n72712 , n72705 , n72710 );
or ( n72713 , n72708 , n72711 , n72712 );
and ( n72714 , n72695 , n72713 );
xor ( n72715 , n72021 , n72183 );
xor ( n72716 , n72715 , n72325 );
and ( n72717 , n72713 , n72716 );
and ( n72718 , n72695 , n72716 );
or ( n72719 , n72714 , n72717 , n72718 );
and ( n72720 , n72400 , n72719 );
xor ( n72721 , n72016 , n72018 );
xor ( n72722 , n72721 , n72328 );
and ( n72723 , n72719 , n72722 );
and ( n72724 , n72400 , n72722 );
or ( n72725 , n72720 , n72723 , n72724 );
and ( n72726 , n72398 , n72725 );
xor ( n72727 , n72331 , n72381 );
xor ( n72728 , n72727 , n72384 );
and ( n72729 , n72725 , n72728 );
and ( n72730 , n72398 , n72728 );
or ( n72731 , n72726 , n72729 , n72730 );
xor ( n72732 , n72014 , n72387 );
xor ( n72733 , n72732 , n72390 );
and ( n72734 , n72731 , n72733 );
xor ( n72735 , n72365 , n72375 );
xor ( n72736 , n72735 , n72378 );
xor ( n72737 , n72349 , n72359 );
xor ( n72738 , n72737 , n72362 );
xor ( n72739 , n72367 , n72369 );
xor ( n72740 , n72739 , n72372 );
and ( n72741 , n72738 , n72740 );
xor ( n72742 , n72341 , n72343 );
xor ( n72743 , n72742 , n72346 );
xor ( n72744 , n72351 , n72353 );
xor ( n72745 , n72744 , n72356 );
and ( n72746 , n72743 , n72745 );
xor ( n72747 , n72314 , n72316 );
xor ( n72748 , n72747 , n72319 );
xor ( n72749 , n72333 , n72335 );
xor ( n72750 , n72749 , n72338 );
and ( n72751 , n72748 , n72750 );
and ( n72752 , n68307 , n61914 );
not ( n72753 , n72752 );
and ( n72754 , n66415 , n63766 );
not ( n72755 , n72754 );
and ( n72756 , n72753 , n72755 );
and ( n72757 , n65606 , n64811 );
not ( n72758 , n72757 );
and ( n72759 , n72755 , n72758 );
and ( n72760 , n72753 , n72758 );
or ( n72761 , n72756 , n72759 , n72760 );
and ( n72762 , n61918 , n68610 );
not ( n72763 , n72762 );
and ( n72764 , n63987 , n66469 );
not ( n72765 , n72764 );
and ( n72766 , n72763 , n72765 );
and ( n72767 , n64548 , n65586 );
not ( n72768 , n72767 );
and ( n72769 , n72765 , n72768 );
and ( n72770 , n72763 , n72768 );
or ( n72771 , n72766 , n72769 , n72770 );
and ( n72772 , n72761 , n72771 );
and ( n72773 , n61505 , n68610 );
not ( n72774 , n72773 );
and ( n72775 , n68307 , n61481 );
not ( n72776 , n72775 );
and ( n72777 , n72774 , n72776 );
and ( n72778 , n72772 , n72777 );
and ( n72779 , n53639 , n52799 );
and ( n72780 , n53328 , n52797 );
nor ( n72781 , n72779 , n72780 );
xnor ( n72782 , n72781 , n52538 );
and ( n72783 , n72777 , n72782 );
and ( n72784 , n72772 , n72782 );
or ( n72785 , n72778 , n72783 , n72784 );
and ( n72786 , n52332 , n53928 );
and ( n72787 , n52082 , n53926 );
nor ( n72788 , n72786 , n72787 );
xnor ( n72789 , n72788 , n53652 );
and ( n72790 , n72785 , n72789 );
and ( n72791 , n53922 , n52269 );
and ( n72792 , n53639 , n52267 );
nor ( n72793 , n72791 , n72792 );
xnor ( n72794 , n72793 , n52008 );
and ( n72795 , n72789 , n72794 );
and ( n72796 , n72785 , n72794 );
or ( n72797 , n72790 , n72795 , n72796 );
xor ( n72798 , n72237 , n72249 );
xor ( n72799 , n72798 , n72252 );
xor ( n72800 , n72258 , n72260 );
xor ( n72801 , n72800 , n72263 );
and ( n72802 , n72799 , n72801 );
xor ( n72803 , n72229 , n72233 );
xor ( n72804 , n72803 , n71853 );
xor ( n72805 , n72241 , n72243 );
xor ( n72806 , n72805 , n72246 );
and ( n72807 , n72804 , n72806 );
xor ( n72808 , n72441 , n72443 );
xor ( n72809 , n72808 , n72446 );
and ( n72810 , n72806 , n72809 );
and ( n72811 , n72804 , n72809 );
or ( n72812 , n72807 , n72810 , n72811 );
and ( n72813 , n72801 , n72812 );
and ( n72814 , n72799 , n72812 );
or ( n72815 , n72802 , n72813 , n72814 );
and ( n72816 , n72797 , n72815 );
and ( n72817 , n60376 , n70108 );
not ( n72818 , n72817 );
and ( n72819 , n61505 , n68752 );
not ( n72820 , n72819 );
and ( n72821 , n72818 , n72820 );
and ( n72822 , n62593 , n67411 );
not ( n72823 , n72822 );
and ( n72824 , n72820 , n72823 );
and ( n72825 , n72818 , n72823 );
or ( n72826 , n72821 , n72824 , n72825 );
xor ( n72827 , n72507 , n72509 );
xor ( n72828 , n72827 , n72512 );
and ( n72829 , n72826 , n72828 );
xor ( n72830 , n72517 , n72519 );
xor ( n72831 , n72830 , n72522 );
and ( n72832 , n72828 , n72831 );
and ( n72833 , n72826 , n72831 );
or ( n72834 , n72829 , n72832 , n72833 );
and ( n72835 , n70256 , n60372 );
not ( n72836 , n72835 );
and ( n72837 , n67343 , n62868 );
not ( n72838 , n72837 );
and ( n72839 , n72836 , n72838 );
and ( n72840 , n63024 , n67013 );
not ( n72841 , n72840 );
and ( n72842 , n72838 , n72841 );
and ( n72843 , n72836 , n72841 );
or ( n72844 , n72839 , n72842 , n72843 );
and ( n72845 , n60821 , n69204 );
not ( n72846 , n72845 );
and ( n72847 , n72844 , n72846 );
xor ( n72848 , n72528 , n72530 );
xor ( n72849 , n72848 , n72533 );
and ( n72850 , n72846 , n72849 );
and ( n72851 , n72844 , n72849 );
or ( n72852 , n72847 , n72850 , n72851 );
and ( n72853 , n72834 , n72852 );
and ( n72854 , n61008 , n69204 );
not ( n72855 , n72854 );
and ( n72856 , n69303 , n61015 );
not ( n72857 , n72856 );
and ( n72858 , n72855 , n72857 );
and ( n72859 , n53328 , n53357 );
and ( n72860 , n53041 , n53355 );
nor ( n72861 , n72859 , n72860 );
xnor ( n72862 , n72861 , n53060 );
and ( n72863 , n72858 , n72862 );
and ( n72864 , n72852 , n72863 );
and ( n72865 , n72834 , n72863 );
or ( n72866 , n72853 , n72864 , n72865 );
and ( n72867 , n69303 , n60711 );
not ( n72868 , n72867 );
xor ( n72869 , n72490 , n72494 );
xor ( n72870 , n72869 , n72499 );
and ( n72871 , n72868 , n72870 );
buf ( n72872 , n72871 );
xor ( n72873 , n72433 , n72435 );
xor ( n72874 , n72873 , n72438 );
xnor ( n72875 , n72544 , n72547 );
and ( n72876 , n72874 , n72875 );
xor ( n72877 , n72552 , n72556 );
and ( n72878 , n72875 , n72877 );
and ( n72879 , n72874 , n72877 );
or ( n72880 , n72876 , n72878 , n72879 );
and ( n72881 , n72872 , n72880 );
xor ( n72882 , n72414 , n72416 );
xor ( n72883 , n72560 , n72562 );
and ( n72884 , n72882 , n72883 );
xor ( n72885 , n72774 , n72776 );
and ( n72886 , n72883 , n72885 );
and ( n72887 , n72882 , n72885 );
or ( n72888 , n72884 , n72886 , n72887 );
and ( n72889 , n72880 , n72888 );
and ( n72890 , n72872 , n72888 );
or ( n72891 , n72881 , n72889 , n72890 );
and ( n72892 , n72866 , n72891 );
xor ( n72893 , n72419 , n72421 );
xor ( n72894 , n72571 , n72573 );
and ( n72895 , n72893 , n72894 );
xor ( n72896 , n72576 , n72578 );
and ( n72897 , n72894 , n72896 );
and ( n72898 , n72893 , n72896 );
or ( n72899 , n72895 , n72897 , n72898 );
and ( n72900 , n63492 , n66917 );
not ( n72901 , n72900 );
and ( n72902 , n64221 , n66005 );
not ( n72903 , n72902 );
and ( n72904 , n72901 , n72903 );
buf ( n72905 , n65177 );
not ( n72906 , n72905 );
and ( n72907 , n72903 , n72906 );
and ( n72908 , n72901 , n72906 );
or ( n72909 , n72904 , n72907 , n72908 );
and ( n72910 , n56915 , n50783 );
and ( n72911 , n56388 , n50781 );
nor ( n72912 , n72910 , n72911 );
xnor ( n72913 , n72912 , n50557 );
or ( n72914 , n72913 , n72545 );
and ( n72915 , n72909 , n72914 );
and ( n72916 , n51077 , n56503 );
and ( n72917 , n50726 , n56501 );
nor ( n72918 , n72916 , n72917 );
xnor ( n72919 , n72918 , n56178 );
and ( n72920 , n51510 , n55851 );
and ( n72921 , n51298 , n55849 );
nor ( n72922 , n72920 , n72921 );
xnor ( n72923 , n72922 , n55506 );
and ( n72924 , n72919 , n72923 );
and ( n72925 , n72914 , n72924 );
and ( n72926 , n72909 , n72924 );
or ( n72927 , n72915 , n72925 , n72926 );
and ( n72928 , n72899 , n72927 );
and ( n72929 , n62377 , n67844 );
not ( n72930 , n72929 );
and ( n72931 , n67997 , n62151 );
not ( n72932 , n72931 );
and ( n72933 , n72930 , n72932 );
and ( n72934 , n50625 , n57187 );
and ( n72935 , n50404 , n57184 );
nor ( n72936 , n72934 , n72935 );
xnor ( n72937 , n72936 , n56175 );
and ( n72938 , n52612 , n54535 );
and ( n72939 , n52332 , n54533 );
nor ( n72940 , n72938 , n72939 );
xnor ( n72941 , n72940 , n54237 );
and ( n72942 , n72937 , n72941 );
and ( n72943 , n53639 , n53357 );
and ( n72944 , n53328 , n53355 );
nor ( n72945 , n72943 , n72944 );
xnor ( n72946 , n72945 , n53060 );
and ( n72947 , n72941 , n72946 );
and ( n72948 , n72937 , n72946 );
or ( n72949 , n72942 , n72947 , n72948 );
and ( n72950 , n72933 , n72949 );
and ( n72951 , n54227 , n52799 );
and ( n72952 , n53922 , n52797 );
nor ( n72953 , n72951 , n72952 );
xnor ( n72954 , n72953 , n52538 );
and ( n72955 , n55497 , n51750 );
and ( n72956 , n55143 , n51748 );
nor ( n72957 , n72955 , n72956 );
xnor ( n72958 , n72957 , n51520 );
and ( n72959 , n72954 , n72958 );
and ( n72960 , n56255 , n51221 );
and ( n72961 , n55756 , n51219 );
nor ( n72962 , n72960 , n72961 );
xnor ( n72963 , n72962 , n51000 );
and ( n72964 , n72958 , n72963 );
and ( n72965 , n72954 , n72963 );
or ( n72966 , n72959 , n72964 , n72965 );
and ( n72967 , n72949 , n72966 );
and ( n72968 , n72933 , n72966 );
or ( n72969 , n72950 , n72967 , n72968 );
and ( n72970 , n72927 , n72969 );
and ( n72971 , n72899 , n72969 );
or ( n72972 , n72928 , n72970 , n72971 );
and ( n72973 , n72891 , n72972 );
and ( n72974 , n72866 , n72972 );
or ( n72975 , n72892 , n72973 , n72974 );
and ( n72976 , n72815 , n72975 );
and ( n72977 , n72797 , n72975 );
or ( n72978 , n72816 , n72976 , n72977 );
and ( n72979 , n72750 , n72978 );
and ( n72980 , n72748 , n72978 );
or ( n72981 , n72751 , n72979 , n72980 );
and ( n72982 , n72745 , n72981 );
and ( n72983 , n72743 , n72981 );
or ( n72984 , n72746 , n72982 , n72983 );
and ( n72985 , n72740 , n72984 );
and ( n72986 , n72738 , n72984 );
or ( n72987 , n72741 , n72985 , n72986 );
and ( n72988 , n72736 , n72987 );
xor ( n72989 , n72400 , n72719 );
xor ( n72990 , n72989 , n72722 );
and ( n72991 , n72987 , n72990 );
and ( n72992 , n72736 , n72990 );
or ( n72993 , n72988 , n72991 , n72992 );
xor ( n72994 , n72398 , n72725 );
xor ( n72995 , n72994 , n72728 );
and ( n72996 , n72993 , n72995 );
xor ( n72997 , n45377 , n45520 );
buf ( n72998 , n72997 );
buf ( n72999 , n72998 );
buf ( n73000 , n72999 );
and ( n73001 , n69059 , n61481 );
not ( n73002 , n73001 );
and ( n73003 , n73000 , n73002 );
and ( n73004 , n66980 , n62998 );
not ( n73005 , n73004 );
and ( n73006 , n73002 , n73005 );
and ( n73007 , n73000 , n73005 );
or ( n73008 , n73003 , n73006 , n73007 );
and ( n73009 , n66720 , n63679 );
not ( n73010 , n73009 );
and ( n73011 , n65678 , n64412 );
not ( n73012 , n73011 );
and ( n73013 , n73010 , n73012 );
buf ( n73014 , n73013 );
and ( n73015 , n73008 , n73014 );
xor ( n73016 , n72584 , n72588 );
xor ( n73017 , n73016 , n72593 );
and ( n73018 , n73014 , n73017 );
and ( n73019 , n73008 , n73017 );
or ( n73020 , n73015 , n73018 , n73019 );
buf ( n73021 , n72455 );
xor ( n73022 , n73021 , n72457 );
and ( n73023 , n73020 , n73022 );
xor ( n73024 , n72461 , n72463 );
xor ( n73025 , n73024 , n72466 );
and ( n73026 , n73022 , n73025 );
and ( n73027 , n73020 , n73025 );
or ( n73028 , n73023 , n73026 , n73027 );
xor ( n73029 , n72471 , n72472 );
xor ( n73030 , n73029 , n72474 );
xor ( n73031 , n72484 , n72485 );
xor ( n73032 , n73031 , n72502 );
and ( n73033 , n73030 , n73032 );
xor ( n73034 , n72515 , n72525 );
xor ( n73035 , n73034 , n72536 );
and ( n73036 , n73032 , n73035 );
and ( n73037 , n73030 , n73035 );
or ( n73038 , n73033 , n73036 , n73037 );
and ( n73039 , n73028 , n73038 );
xor ( n73040 , n72548 , n72557 );
xor ( n73041 , n73040 , n72563 );
xor ( n73042 , n72574 , n72579 );
xor ( n73043 , n73042 , n72596 );
and ( n73044 , n73041 , n73043 );
xor ( n73045 , n72615 , n72617 );
xor ( n73046 , n73045 , n72620 );
and ( n73047 , n73043 , n73046 );
and ( n73048 , n73041 , n73046 );
or ( n73049 , n73044 , n73047 , n73048 );
and ( n73050 , n73038 , n73049 );
and ( n73051 , n73028 , n73049 );
or ( n73052 , n73039 , n73050 , n73051 );
xor ( n73053 , n72404 , n72406 );
xor ( n73054 , n73053 , n72408 );
xor ( n73055 , n72412 , n72430 );
xor ( n73056 , n73055 , n72449 );
and ( n73057 , n73054 , n73056 );
xor ( n73058 , n72459 , n72469 );
xor ( n73059 , n73058 , n72477 );
and ( n73060 , n73056 , n73059 );
and ( n73061 , n73054 , n73059 );
or ( n73062 , n73057 , n73060 , n73061 );
and ( n73063 , n73052 , n73062 );
xor ( n73064 , n72505 , n72539 );
xor ( n73065 , n73064 , n72566 );
xor ( n73066 , n72599 , n72623 );
xor ( n73067 , n73066 , n72626 );
and ( n73068 , n73065 , n73067 );
xor ( n73069 , n72632 , n72634 );
xor ( n73070 , n73069 , n72637 );
and ( n73071 , n73067 , n73070 );
and ( n73072 , n73065 , n73070 );
or ( n73073 , n73068 , n73071 , n73072 );
and ( n73074 , n73062 , n73073 );
and ( n73075 , n73052 , n73073 );
or ( n73076 , n73063 , n73074 , n73075 );
xor ( n73077 , n72411 , n72452 );
xor ( n73078 , n73077 , n72480 );
xor ( n73079 , n72569 , n72629 );
xor ( n73080 , n73079 , n72640 );
and ( n73081 , n73078 , n73080 );
xor ( n73082 , n72654 , n72656 );
xor ( n73083 , n73082 , n72659 );
and ( n73084 , n73080 , n73083 );
and ( n73085 , n73078 , n73083 );
or ( n73086 , n73081 , n73084 , n73085 );
and ( n73087 , n73076 , n73086 );
xor ( n73088 , n72483 , n72643 );
xor ( n73089 , n73088 , n72662 );
and ( n73090 , n73086 , n73089 );
and ( n73091 , n73076 , n73089 );
or ( n73092 , n73087 , n73090 , n73091 );
xor ( n73093 , n72402 , n72665 );
xor ( n73094 , n73093 , n72692 );
and ( n73095 , n73092 , n73094 );
xor ( n73096 , n72705 , n72707 );
xor ( n73097 , n73096 , n72710 );
and ( n73098 , n73094 , n73097 );
and ( n73099 , n73092 , n73097 );
or ( n73100 , n73095 , n73098 , n73099 );
xor ( n73101 , n72695 , n72713 );
xor ( n73102 , n73101 , n72716 );
and ( n73103 , n73100 , n73102 );
xor ( n73104 , n72676 , n72686 );
xor ( n73105 , n73104 , n72689 );
xor ( n73106 , n72697 , n72699 );
xor ( n73107 , n73106 , n72702 );
and ( n73108 , n73105 , n73107 );
xor ( n73109 , n72668 , n72670 );
xor ( n73110 , n73109 , n72673 );
xor ( n73111 , n72678 , n72680 );
xor ( n73112 , n73111 , n72683 );
and ( n73113 , n73110 , n73112 );
and ( n73114 , n61918 , n68752 );
not ( n73115 , n73114 );
and ( n73116 , n62593 , n67844 );
not ( n73117 , n73116 );
and ( n73118 , n73115 , n73117 );
and ( n73119 , n63987 , n66917 );
not ( n73120 , n73119 );
and ( n73121 , n73117 , n73120 );
and ( n73122 , n73115 , n73120 );
or ( n73123 , n73118 , n73121 , n73122 );
and ( n73124 , n69688 , n60711 );
not ( n73125 , n73124 );
and ( n73126 , n73123 , n73125 );
xor ( n73127 , n72753 , n72755 );
xor ( n73128 , n73127 , n72758 );
and ( n73129 , n73125 , n73128 );
and ( n73130 , n73123 , n73128 );
or ( n73131 , n73126 , n73129 , n73130 );
and ( n73132 , n69059 , n61914 );
not ( n73133 , n73132 );
and ( n73134 , n67997 , n62868 );
not ( n73135 , n73134 );
and ( n73136 , n73133 , n73135 );
and ( n73137 , n66720 , n63766 );
not ( n73138 , n73137 );
and ( n73139 , n73135 , n73138 );
and ( n73140 , n73133 , n73138 );
or ( n73141 , n73136 , n73139 , n73140 );
and ( n73142 , n60821 , n69507 );
not ( n73143 , n73142 );
and ( n73144 , n73141 , n73143 );
xor ( n73145 , n72763 , n72765 );
xor ( n73146 , n73145 , n72768 );
and ( n73147 , n73143 , n73146 );
and ( n73148 , n73141 , n73146 );
or ( n73149 , n73144 , n73147 , n73148 );
and ( n73150 , n73131 , n73149 );
and ( n73151 , n51510 , n55159 );
and ( n73152 , n51298 , n55157 );
nor ( n73153 , n73151 , n73152 );
xnor ( n73154 , n73153 , n54864 );
and ( n73155 , n73150 , n73154 );
xor ( n73156 , n72417 , n72422 );
xor ( n73157 , n73156 , n72427 );
and ( n73158 , n73154 , n73157 );
and ( n73159 , n73150 , n73157 );
or ( n73160 , n73155 , n73158 , n73159 );
xor ( n73161 , n72785 , n72789 );
xor ( n73162 , n73161 , n72794 );
and ( n73163 , n73160 , n73162 );
and ( n73164 , n73112 , n73163 );
and ( n73165 , n73110 , n73163 );
or ( n73166 , n73113 , n73164 , n73165 );
and ( n73167 , n73107 , n73166 );
and ( n73168 , n73105 , n73166 );
or ( n73169 , n73108 , n73167 , n73168 );
xor ( n73170 , n72646 , n72648 );
xor ( n73171 , n73170 , n72651 );
xor ( n73172 , n72772 , n72777 );
xor ( n73173 , n73172 , n72782 );
and ( n73174 , n67343 , n62998 );
not ( n73175 , n73174 );
and ( n73176 , n66415 , n64412 );
not ( n73177 , n73176 );
and ( n73178 , n73175 , n73177 );
and ( n73179 , n65678 , n64811 );
not ( n73180 , n73179 );
and ( n73181 , n73177 , n73180 );
and ( n73182 , n73175 , n73180 );
or ( n73183 , n73178 , n73181 , n73182 );
and ( n73184 , n63024 , n67411 );
not ( n73185 , n73184 );
and ( n73186 , n64221 , n66469 );
not ( n73187 , n73186 );
and ( n73188 , n73185 , n73187 );
and ( n73189 , n64548 , n66005 );
not ( n73190 , n73189 );
and ( n73191 , n73187 , n73190 );
and ( n73192 , n73185 , n73190 );
or ( n73193 , n73188 , n73191 , n73192 );
and ( n73194 , n73183 , n73193 );
and ( n73195 , n52790 , n53928 );
and ( n73196 , n52612 , n53926 );
nor ( n73197 , n73195 , n73196 );
xnor ( n73198 , n73197 , n53652 );
and ( n73199 , n73194 , n73198 );
and ( n73200 , n73173 , n73199 );
xor ( n73201 , n72603 , n72607 );
xor ( n73202 , n73201 , n72612 );
xor ( n73203 , n72826 , n72828 );
xor ( n73204 , n73203 , n72831 );
and ( n73205 , n73202 , n73204 );
xor ( n73206 , n72844 , n72846 );
xor ( n73207 , n73206 , n72849 );
and ( n73208 , n73204 , n73207 );
and ( n73209 , n73202 , n73207 );
or ( n73210 , n73205 , n73208 , n73209 );
and ( n73211 , n73199 , n73210 );
and ( n73212 , n73173 , n73210 );
or ( n73213 , n73200 , n73211 , n73212 );
and ( n73214 , n73171 , n73213 );
xor ( n73215 , n72858 , n72862 );
xor ( n73216 , n72761 , n72771 );
and ( n73217 , n73215 , n73216 );
and ( n73218 , n61008 , n69507 );
not ( n73219 , n73218 );
and ( n73220 , n69688 , n61015 );
not ( n73221 , n73220 );
and ( n73222 , n73219 , n73221 );
and ( n73223 , n62377 , n68610 );
not ( n73224 , n73223 );
and ( n73225 , n68307 , n62151 );
not ( n73226 , n73225 );
and ( n73227 , n73224 , n73226 );
and ( n73228 , n73222 , n73227 );
and ( n73229 , n53041 , n53928 );
and ( n73230 , n52790 , n53926 );
nor ( n73231 , n73229 , n73230 );
xnor ( n73232 , n73231 , n53652 );
and ( n73233 , n73227 , n73232 );
and ( n73234 , n73222 , n73232 );
or ( n73235 , n73228 , n73233 , n73234 );
and ( n73236 , n73216 , n73235 );
and ( n73237 , n73215 , n73235 );
or ( n73238 , n73217 , n73236 , n73237 );
xor ( n73239 , n72818 , n72820 );
xor ( n73240 , n73239 , n72823 );
xor ( n73241 , n72901 , n72903 );
xor ( n73242 , n73241 , n72906 );
and ( n73243 , n73240 , n73242 );
xor ( n73244 , n72836 , n72838 );
xor ( n73245 , n73244 , n72841 );
and ( n73246 , n73242 , n73245 );
and ( n73247 , n73240 , n73245 );
or ( n73248 , n73243 , n73246 , n73247 );
xnor ( n73249 , n72913 , n72545 );
xor ( n73250 , n72919 , n72923 );
and ( n73251 , n73249 , n73250 );
xor ( n73252 , n72855 , n72857 );
and ( n73253 , n73250 , n73252 );
and ( n73254 , n73249 , n73252 );
or ( n73255 , n73251 , n73253 , n73254 );
and ( n73256 , n73248 , n73255 );
xor ( n73257 , n72930 , n72932 );
and ( n73258 , n50726 , n57187 );
and ( n73259 , n50625 , n57184 );
nor ( n73260 , n73258 , n73259 );
xnor ( n73261 , n73260 , n56175 );
and ( n73262 , n51298 , n56503 );
and ( n73263 , n51077 , n56501 );
nor ( n73264 , n73262 , n73263 );
xnor ( n73265 , n73264 , n56178 );
and ( n73266 , n73261 , n73265 );
and ( n73267 , n55756 , n51750 );
and ( n73268 , n55497 , n51748 );
nor ( n73269 , n73267 , n73268 );
xnor ( n73270 , n73269 , n51520 );
and ( n73271 , n73265 , n73270 );
and ( n73272 , n73261 , n73270 );
or ( n73273 , n73266 , n73271 , n73272 );
and ( n73274 , n73257 , n73273 );
and ( n73275 , n61505 , n69204 );
not ( n73276 , n73275 );
and ( n73277 , n69303 , n61481 );
not ( n73278 , n73277 );
and ( n73279 , n73276 , n73278 );
and ( n73280 , n73273 , n73279 );
and ( n73281 , n73257 , n73279 );
or ( n73282 , n73274 , n73280 , n73281 );
and ( n73283 , n73255 , n73282 );
and ( n73284 , n73248 , n73282 );
or ( n73285 , n73256 , n73283 , n73284 );
and ( n73286 , n73238 , n73285 );
and ( n73287 , n63492 , n67013 );
not ( n73288 , n73287 );
and ( n73289 , n66980 , n63679 );
not ( n73290 , n73289 );
and ( n73291 , n73288 , n73290 );
and ( n73292 , n65177 , n65586 );
not ( n73293 , n73292 );
and ( n73294 , n65606 , n65210 );
not ( n73295 , n73294 );
and ( n73296 , n73293 , n73295 );
and ( n73297 , n73291 , n73296 );
and ( n73298 , n51734 , n55851 );
and ( n73299 , n51510 , n55849 );
nor ( n73300 , n73298 , n73299 );
xnor ( n73301 , n73300 , n55506 );
and ( n73302 , n52332 , n55159 );
and ( n73303 , n52082 , n55157 );
nor ( n73304 , n73302 , n73303 );
xnor ( n73305 , n73304 , n54864 );
and ( n73306 , n73301 , n73305 );
and ( n73307 , n53328 , n53928 );
and ( n73308 , n53041 , n53926 );
nor ( n73309 , n73307 , n73308 );
xnor ( n73310 , n73309 , n53652 );
and ( n73311 , n73305 , n73310 );
and ( n73312 , n73301 , n73310 );
or ( n73313 , n73306 , n73311 , n73312 );
and ( n73314 , n73296 , n73313 );
and ( n73315 , n73291 , n73313 );
or ( n73316 , n73297 , n73314 , n73315 );
and ( n73317 , n54604 , n52799 );
and ( n73318 , n54227 , n52797 );
nor ( n73319 , n73317 , n73318 );
xnor ( n73320 , n73319 , n52538 );
and ( n73321 , n55143 , n52269 );
and ( n73322 , n54942 , n52267 );
nor ( n73323 , n73321 , n73322 );
xnor ( n73324 , n73323 , n52008 );
and ( n73325 , n73320 , n73324 );
and ( n73326 , n56388 , n51221 );
and ( n73327 , n56255 , n51219 );
nor ( n73328 , n73326 , n73327 );
xnor ( n73329 , n73328 , n51000 );
and ( n73330 , n73324 , n73329 );
and ( n73331 , n73320 , n73329 );
or ( n73332 , n73325 , n73330 , n73331 );
and ( n73333 , n57063 , n50783 );
and ( n73334 , n56915 , n50781 );
nor ( n73335 , n73333 , n73334 );
xnor ( n73336 , n73335 , n50557 );
and ( n73337 , n57063 , n50781 );
not ( n73338 , n73337 );
and ( n73339 , n73338 , n50557 );
and ( n73340 , n73336 , n73339 );
xor ( n73341 , n45378 , n45519 );
buf ( n73342 , n73341 );
buf ( n73343 , n73342 );
buf ( n73344 , n73343 );
and ( n73345 , n73339 , n73344 );
and ( n73346 , n73336 , n73344 );
or ( n73347 , n73340 , n73345 , n73346 );
and ( n73348 , n73332 , n73347 );
xor ( n73349 , n72937 , n72941 );
xor ( n73350 , n73349 , n72946 );
and ( n73351 , n73347 , n73350 );
and ( n73352 , n73332 , n73350 );
or ( n73353 , n73348 , n73351 , n73352 );
and ( n73354 , n73316 , n73353 );
xor ( n73355 , n72954 , n72958 );
xor ( n73356 , n73355 , n72963 );
xor ( n73357 , n73000 , n73002 );
xor ( n73358 , n73357 , n73005 );
and ( n73359 , n73356 , n73358 );
xor ( n73360 , n73010 , n73012 );
buf ( n73361 , n73360 );
and ( n73362 , n73358 , n73361 );
and ( n73363 , n73356 , n73361 );
or ( n73364 , n73359 , n73362 , n73363 );
and ( n73365 , n73353 , n73364 );
and ( n73366 , n73316 , n73364 );
or ( n73367 , n73354 , n73365 , n73366 );
and ( n73368 , n73285 , n73367 );
and ( n73369 , n73238 , n73367 );
or ( n73370 , n73286 , n73368 , n73369 );
and ( n73371 , n73213 , n73370 );
and ( n73372 , n73171 , n73370 );
or ( n73373 , n73214 , n73371 , n73372 );
buf ( n73374 , n72868 );
xor ( n73375 , n73374 , n72870 );
xor ( n73376 , n72874 , n72875 );
xor ( n73377 , n73376 , n72877 );
and ( n73378 , n73375 , n73377 );
xor ( n73379 , n72882 , n72883 );
xor ( n73380 , n73379 , n72885 );
and ( n73381 , n73377 , n73380 );
and ( n73382 , n73375 , n73380 );
or ( n73383 , n73378 , n73381 , n73382 );
xor ( n73384 , n72893 , n72894 );
xor ( n73385 , n73384 , n72896 );
xor ( n73386 , n72909 , n72914 );
xor ( n73387 , n73386 , n72924 );
and ( n73388 , n73385 , n73387 );
xor ( n73389 , n72933 , n72949 );
xor ( n73390 , n73389 , n72966 );
and ( n73391 , n73387 , n73390 );
and ( n73392 , n73385 , n73390 );
or ( n73393 , n73388 , n73391 , n73392 );
and ( n73394 , n73383 , n73393 );
xor ( n73395 , n72804 , n72806 );
xor ( n73396 , n73395 , n72809 );
and ( n73397 , n73393 , n73396 );
and ( n73398 , n73383 , n73396 );
or ( n73399 , n73394 , n73397 , n73398 );
xor ( n73400 , n72834 , n72852 );
xor ( n73401 , n73400 , n72863 );
xor ( n73402 , n72872 , n72880 );
xor ( n73403 , n73402 , n72888 );
and ( n73404 , n73401 , n73403 );
xor ( n73405 , n72899 , n72927 );
xor ( n73406 , n73405 , n72969 );
and ( n73407 , n73403 , n73406 );
and ( n73408 , n73401 , n73406 );
or ( n73409 , n73404 , n73407 , n73408 );
and ( n73410 , n73399 , n73409 );
xor ( n73411 , n73020 , n73022 );
xor ( n73412 , n73411 , n73025 );
xor ( n73413 , n73030 , n73032 );
xor ( n73414 , n73413 , n73035 );
and ( n73415 , n73412 , n73414 );
xor ( n73416 , n73041 , n73043 );
xor ( n73417 , n73416 , n73046 );
and ( n73418 , n73414 , n73417 );
and ( n73419 , n73412 , n73417 );
or ( n73420 , n73415 , n73418 , n73419 );
and ( n73421 , n73409 , n73420 );
and ( n73422 , n73399 , n73420 );
or ( n73423 , n73410 , n73421 , n73422 );
and ( n73424 , n73373 , n73423 );
xor ( n73425 , n72799 , n72801 );
xor ( n73426 , n73425 , n72812 );
xor ( n73427 , n72866 , n72891 );
xor ( n73428 , n73427 , n72972 );
and ( n73429 , n73426 , n73428 );
xor ( n73430 , n73028 , n73038 );
xor ( n73431 , n73430 , n73049 );
and ( n73432 , n73428 , n73431 );
and ( n73433 , n73426 , n73431 );
or ( n73434 , n73429 , n73432 , n73433 );
and ( n73435 , n73423 , n73434 );
and ( n73436 , n73373 , n73434 );
or ( n73437 , n73424 , n73435 , n73436 );
xor ( n73438 , n72797 , n72815 );
xor ( n73439 , n73438 , n72975 );
xor ( n73440 , n73052 , n73062 );
xor ( n73441 , n73440 , n73073 );
and ( n73442 , n73439 , n73441 );
xor ( n73443 , n73078 , n73080 );
xor ( n73444 , n73443 , n73083 );
and ( n73445 , n73441 , n73444 );
and ( n73446 , n73439 , n73444 );
or ( n73447 , n73442 , n73445 , n73446 );
and ( n73448 , n73437 , n73447 );
xor ( n73449 , n72748 , n72750 );
xor ( n73450 , n73449 , n72978 );
and ( n73451 , n73447 , n73450 );
and ( n73452 , n73437 , n73450 );
or ( n73453 , n73448 , n73451 , n73452 );
and ( n73454 , n73169 , n73453 );
xor ( n73455 , n72743 , n72745 );
xor ( n73456 , n73455 , n72981 );
and ( n73457 , n73453 , n73456 );
and ( n73458 , n73169 , n73456 );
or ( n73459 , n73454 , n73457 , n73458 );
and ( n73460 , n73102 , n73459 );
and ( n73461 , n73100 , n73459 );
or ( n73462 , n73103 , n73460 , n73461 );
xor ( n73463 , n72736 , n72987 );
xor ( n73464 , n73463 , n72990 );
and ( n73465 , n73462 , n73464 );
xor ( n73466 , n72738 , n72740 );
xor ( n73467 , n73466 , n72984 );
xor ( n73468 , n73092 , n73094 );
xor ( n73469 , n73468 , n73097 );
xor ( n73470 , n73076 , n73086 );
xor ( n73471 , n73470 , n73089 );
xor ( n73472 , n73054 , n73056 );
xor ( n73473 , n73472 , n73059 );
xor ( n73474 , n73065 , n73067 );
xor ( n73475 , n73474 , n73070 );
and ( n73476 , n73473 , n73475 );
xor ( n73477 , n73160 , n73162 );
and ( n73478 , n73475 , n73477 );
and ( n73479 , n73473 , n73477 );
or ( n73480 , n73476 , n73478 , n73479 );
xor ( n73481 , n73150 , n73154 );
xor ( n73482 , n73481 , n73157 );
xor ( n73483 , n73008 , n73014 );
xor ( n73484 , n73483 , n73017 );
xor ( n73485 , n73194 , n73198 );
and ( n73486 , n73484 , n73485 );
xor ( n73487 , n73131 , n73149 );
and ( n73488 , n73485 , n73487 );
and ( n73489 , n73484 , n73487 );
or ( n73490 , n73486 , n73488 , n73489 );
and ( n73491 , n73482 , n73490 );
and ( n73492 , n52082 , n55159 );
and ( n73493 , n51734 , n55157 );
nor ( n73494 , n73492 , n73493 );
xnor ( n73495 , n73494 , n54864 );
and ( n73496 , n54942 , n52269 );
and ( n73497 , n54604 , n52267 );
nor ( n73498 , n73496 , n73497 );
xnor ( n73499 , n73498 , n52008 );
and ( n73500 , n73495 , n73499 );
xor ( n73501 , n73222 , n73227 );
xor ( n73502 , n73501 , n73232 );
and ( n73503 , n73499 , n73502 );
and ( n73504 , n73495 , n73502 );
or ( n73505 , n73500 , n73503 , n73504 );
and ( n73506 , n70256 , n60711 );
not ( n73507 , n73506 );
xor ( n73508 , n73115 , n73117 );
xor ( n73509 , n73508 , n73120 );
and ( n73510 , n73507 , n73509 );
and ( n73511 , n60821 , n70108 );
not ( n73512 , n73511 );
xor ( n73513 , n73133 , n73135 );
xor ( n73514 , n73513 , n73138 );
and ( n73515 , n73512 , n73514 );
and ( n73516 , n73510 , n73515 );
and ( n73517 , n73505 , n73516 );
xor ( n73518 , n73123 , n73125 );
xor ( n73519 , n73518 , n73128 );
xor ( n73520 , n73141 , n73143 );
xor ( n73521 , n73520 , n73146 );
and ( n73522 , n73519 , n73521 );
and ( n73523 , n73516 , n73522 );
and ( n73524 , n73505 , n73522 );
or ( n73525 , n73517 , n73523 , n73524 );
and ( n73526 , n73490 , n73525 );
and ( n73527 , n73482 , n73525 );
or ( n73528 , n73491 , n73526 , n73527 );
xor ( n73529 , n73183 , n73193 );
and ( n73530 , n63492 , n67411 );
not ( n73531 , n73530 );
and ( n73532 , n67343 , n63679 );
not ( n73533 , n73532 );
and ( n73534 , n73531 , n73533 );
and ( n73535 , n64548 , n66469 );
not ( n73536 , n73535 );
and ( n73537 , n66415 , n64811 );
not ( n73538 , n73537 );
and ( n73539 , n73536 , n73538 );
and ( n73540 , n73534 , n73539 );
and ( n73541 , n53922 , n53357 );
and ( n73542 , n53639 , n53355 );
nor ( n73543 , n73541 , n73542 );
xnor ( n73544 , n73543 , n53060 );
and ( n73545 , n73539 , n73544 );
and ( n73546 , n73534 , n73544 );
or ( n73547 , n73540 , n73545 , n73546 );
and ( n73548 , n73529 , n73547 );
and ( n73549 , n69688 , n61481 );
not ( n73550 , n73549 );
and ( n73551 , n69059 , n62151 );
not ( n73552 , n73551 );
and ( n73553 , n73550 , n73552 );
and ( n73554 , n68307 , n62868 );
not ( n73555 , n73554 );
and ( n73556 , n73552 , n73555 );
and ( n73557 , n73550 , n73555 );
or ( n73558 , n73553 , n73556 , n73557 );
and ( n73559 , n61505 , n69507 );
not ( n73560 , n73559 );
and ( n73561 , n62377 , n68752 );
not ( n73562 , n73561 );
and ( n73563 , n73560 , n73562 );
and ( n73564 , n62593 , n68610 );
not ( n73565 , n73564 );
and ( n73566 , n73562 , n73565 );
and ( n73567 , n73560 , n73565 );
or ( n73568 , n73563 , n73566 , n73567 );
and ( n73569 , n73558 , n73568 );
and ( n73570 , n73547 , n73569 );
and ( n73571 , n73529 , n73569 );
or ( n73572 , n73548 , n73570 , n73571 );
xor ( n73573 , n73175 , n73177 );
xor ( n73574 , n73573 , n73180 );
xor ( n73575 , n73185 , n73187 );
xor ( n73576 , n73575 , n73190 );
and ( n73577 , n73574 , n73576 );
xor ( n73578 , n73261 , n73265 );
xor ( n73579 , n73578 , n73270 );
xor ( n73580 , n73219 , n73221 );
and ( n73581 , n73579 , n73580 );
buf ( n73582 , n73581 );
and ( n73583 , n73577 , n73582 );
xor ( n73584 , n73276 , n73278 );
xor ( n73585 , n73224 , n73226 );
and ( n73586 , n73584 , n73585 );
xor ( n73587 , n73288 , n73290 );
and ( n73588 , n73585 , n73587 );
and ( n73589 , n73584 , n73587 );
or ( n73590 , n73586 , n73588 , n73589 );
and ( n73591 , n73582 , n73590 );
and ( n73592 , n73577 , n73590 );
or ( n73593 , n73583 , n73591 , n73592 );
and ( n73594 , n73572 , n73593 );
xor ( n73595 , n73293 , n73295 );
and ( n73596 , n51510 , n56503 );
and ( n73597 , n51298 , n56501 );
nor ( n73598 , n73596 , n73597 );
xnor ( n73599 , n73598 , n56178 );
and ( n73600 , n52082 , n55851 );
and ( n73601 , n51734 , n55849 );
nor ( n73602 , n73600 , n73601 );
xnor ( n73603 , n73602 , n55506 );
and ( n73604 , n73599 , n73603 );
and ( n73605 , n55497 , n52269 );
and ( n73606 , n55143 , n52267 );
nor ( n73607 , n73605 , n73606 );
xnor ( n73608 , n73607 , n52008 );
and ( n73609 , n73603 , n73608 );
and ( n73610 , n73599 , n73608 );
or ( n73611 , n73604 , n73609 , n73610 );
and ( n73612 , n73595 , n73611 );
and ( n73613 , n61918 , n69204 );
not ( n73614 , n73613 );
and ( n73615 , n63987 , n67013 );
not ( n73616 , n73615 );
and ( n73617 , n73614 , n73616 );
and ( n73618 , n64221 , n66917 );
not ( n73619 , n73618 );
and ( n73620 , n73616 , n73619 );
and ( n73621 , n73614 , n73619 );
or ( n73622 , n73617 , n73620 , n73621 );
and ( n73623 , n73611 , n73622 );
and ( n73624 , n73595 , n73622 );
or ( n73625 , n73612 , n73623 , n73624 );
and ( n73626 , n66720 , n64412 );
not ( n73627 , n73626 );
and ( n73628 , n65177 , n66005 );
not ( n73629 , n73628 );
and ( n73630 , n73627 , n73629 );
buf ( n73631 , n65606 );
not ( n73632 , n73631 );
and ( n73633 , n73629 , n73632 );
and ( n73634 , n73627 , n73632 );
or ( n73635 , n73630 , n73633 , n73634 );
and ( n73636 , n63024 , n67844 );
not ( n73637 , n73636 );
and ( n73638 , n66980 , n63766 );
not ( n73639 , n73638 );
and ( n73640 , n73637 , n73639 );
and ( n73641 , n73635 , n73640 );
and ( n73642 , n61008 , n70108 );
not ( n73643 , n73642 );
and ( n73644 , n70256 , n61015 );
not ( n73645 , n73644 );
and ( n73646 , n73643 , n73645 );
and ( n73647 , n73640 , n73646 );
and ( n73648 , n73635 , n73646 );
or ( n73649 , n73641 , n73647 , n73648 );
and ( n73650 , n73625 , n73649 );
and ( n73651 , n51077 , n57187 );
and ( n73652 , n50726 , n57184 );
nor ( n73653 , n73651 , n73652 );
xnor ( n73654 , n73653 , n56175 );
and ( n73655 , n52612 , n55159 );
and ( n73656 , n52332 , n55157 );
nor ( n73657 , n73655 , n73656 );
xnor ( n73658 , n73657 , n54864 );
and ( n73659 , n73654 , n73658 );
and ( n73660 , n53639 , n53928 );
and ( n73661 , n53328 , n53926 );
nor ( n73662 , n73660 , n73661 );
xnor ( n73663 , n73662 , n53652 );
and ( n73664 , n73658 , n73663 );
and ( n73665 , n73654 , n73663 );
or ( n73666 , n73659 , n73664 , n73665 );
and ( n73667 , n54227 , n53357 );
and ( n73668 , n53922 , n53355 );
nor ( n73669 , n73667 , n73668 );
xnor ( n73670 , n73669 , n53060 );
and ( n73671 , n54942 , n52799 );
and ( n73672 , n54604 , n52797 );
nor ( n73673 , n73671 , n73672 );
xnor ( n73674 , n73673 , n52538 );
and ( n73675 , n73670 , n73674 );
and ( n73676 , n56255 , n51750 );
and ( n73677 , n55756 , n51748 );
nor ( n73678 , n73676 , n73677 );
xnor ( n73679 , n73678 , n51520 );
and ( n73680 , n73674 , n73679 );
and ( n73681 , n73670 , n73679 );
or ( n73682 , n73675 , n73680 , n73681 );
and ( n73683 , n73666 , n73682 );
and ( n73684 , n56915 , n51221 );
and ( n73685 , n56388 , n51219 );
nor ( n73686 , n73684 , n73685 );
xnor ( n73687 , n73686 , n51000 );
and ( n73688 , n73687 , n73337 );
xor ( n73689 , n45381 , n45517 );
buf ( n73690 , n73689 );
buf ( n73691 , n73690 );
buf ( n73692 , n73691 );
and ( n73693 , n73337 , n73692 );
and ( n73694 , n73687 , n73692 );
or ( n73695 , n73688 , n73693 , n73694 );
and ( n73696 , n73682 , n73695 );
and ( n73697 , n73666 , n73695 );
or ( n73698 , n73683 , n73696 , n73697 );
and ( n73699 , n73649 , n73698 );
and ( n73700 , n73625 , n73698 );
or ( n73701 , n73650 , n73699 , n73700 );
and ( n73702 , n73593 , n73701 );
and ( n73703 , n73572 , n73701 );
or ( n73704 , n73594 , n73702 , n73703 );
and ( n73705 , n69303 , n61914 );
not ( n73706 , n73705 );
and ( n73707 , n67997 , n62998 );
not ( n73708 , n73707 );
and ( n73709 , n73706 , n73708 );
and ( n73710 , n65678 , n65210 );
not ( n73711 , n73710 );
and ( n73712 , n73708 , n73711 );
and ( n73713 , n73706 , n73711 );
or ( n73714 , n73709 , n73712 , n73713 );
xor ( n73715 , n73301 , n73305 );
xor ( n73716 , n73715 , n73310 );
and ( n73717 , n73714 , n73716 );
xor ( n73718 , n73320 , n73324 );
xor ( n73719 , n73718 , n73329 );
and ( n73720 , n73716 , n73719 );
and ( n73721 , n73714 , n73719 );
or ( n73722 , n73717 , n73720 , n73721 );
xor ( n73723 , n73240 , n73242 );
xor ( n73724 , n73723 , n73245 );
and ( n73725 , n73722 , n73724 );
xor ( n73726 , n73249 , n73250 );
xor ( n73727 , n73726 , n73252 );
and ( n73728 , n73724 , n73727 );
and ( n73729 , n73722 , n73727 );
or ( n73730 , n73725 , n73728 , n73729 );
xor ( n73731 , n73257 , n73273 );
xor ( n73732 , n73731 , n73279 );
xor ( n73733 , n73291 , n73296 );
xor ( n73734 , n73733 , n73313 );
and ( n73735 , n73732 , n73734 );
xor ( n73736 , n73332 , n73347 );
xor ( n73737 , n73736 , n73350 );
and ( n73738 , n73734 , n73737 );
and ( n73739 , n73732 , n73737 );
or ( n73740 , n73735 , n73738 , n73739 );
and ( n73741 , n73730 , n73740 );
xor ( n73742 , n73202 , n73204 );
xor ( n73743 , n73742 , n73207 );
and ( n73744 , n73740 , n73743 );
and ( n73745 , n73730 , n73743 );
or ( n73746 , n73741 , n73744 , n73745 );
and ( n73747 , n73704 , n73746 );
xor ( n73748 , n73215 , n73216 );
xor ( n73749 , n73748 , n73235 );
xor ( n73750 , n73248 , n73255 );
xor ( n73751 , n73750 , n73282 );
and ( n73752 , n73749 , n73751 );
xor ( n73753 , n73316 , n73353 );
xor ( n73754 , n73753 , n73364 );
and ( n73755 , n73751 , n73754 );
and ( n73756 , n73749 , n73754 );
or ( n73757 , n73752 , n73755 , n73756 );
and ( n73758 , n73746 , n73757 );
and ( n73759 , n73704 , n73757 );
or ( n73760 , n73747 , n73758 , n73759 );
and ( n73761 , n73528 , n73760 );
xor ( n73762 , n73173 , n73199 );
xor ( n73763 , n73762 , n73210 );
xor ( n73764 , n73238 , n73285 );
xor ( n73765 , n73764 , n73367 );
and ( n73766 , n73763 , n73765 );
xor ( n73767 , n73383 , n73393 );
xor ( n73768 , n73767 , n73396 );
and ( n73769 , n73765 , n73768 );
and ( n73770 , n73763 , n73768 );
or ( n73771 , n73766 , n73769 , n73770 );
and ( n73772 , n73760 , n73771 );
and ( n73773 , n73528 , n73771 );
or ( n73774 , n73761 , n73772 , n73773 );
and ( n73775 , n73480 , n73774 );
xor ( n73776 , n73171 , n73213 );
xor ( n73777 , n73776 , n73370 );
xor ( n73778 , n73399 , n73409 );
xor ( n73779 , n73778 , n73420 );
and ( n73780 , n73777 , n73779 );
xor ( n73781 , n73426 , n73428 );
xor ( n73782 , n73781 , n73431 );
and ( n73783 , n73779 , n73782 );
and ( n73784 , n73777 , n73782 );
or ( n73785 , n73780 , n73783 , n73784 );
and ( n73786 , n73774 , n73785 );
and ( n73787 , n73480 , n73785 );
or ( n73788 , n73775 , n73786 , n73787 );
and ( n73789 , n73471 , n73788 );
xor ( n73790 , n73110 , n73112 );
xor ( n73791 , n73790 , n73163 );
xor ( n73792 , n73373 , n73423 );
xor ( n73793 , n73792 , n73434 );
and ( n73794 , n73791 , n73793 );
xor ( n73795 , n73439 , n73441 );
xor ( n73796 , n73795 , n73444 );
and ( n73797 , n73793 , n73796 );
and ( n73798 , n73791 , n73796 );
or ( n73799 , n73794 , n73797 , n73798 );
and ( n73800 , n73788 , n73799 );
and ( n73801 , n73471 , n73799 );
or ( n73802 , n73789 , n73800 , n73801 );
and ( n73803 , n73469 , n73802 );
xor ( n73804 , n73169 , n73453 );
xor ( n73805 , n73804 , n73456 );
and ( n73806 , n73802 , n73805 );
and ( n73807 , n73469 , n73805 );
or ( n73808 , n73803 , n73806 , n73807 );
and ( n73809 , n73467 , n73808 );
xor ( n73810 , n73100 , n73102 );
xor ( n73811 , n73810 , n73459 );
and ( n73812 , n73808 , n73811 );
and ( n73813 , n73467 , n73811 );
or ( n73814 , n73809 , n73812 , n73813 );
and ( n73815 , n73464 , n73814 );
and ( n73816 , n73462 , n73814 );
or ( n73817 , n73465 , n73815 , n73816 );
and ( n73818 , n72995 , n73817 );
and ( n73819 , n72993 , n73817 );
or ( n73820 , n72996 , n73818 , n73819 );
and ( n73821 , n72733 , n73820 );
and ( n73822 , n72731 , n73820 );
or ( n73823 , n72734 , n73821 , n73822 );
and ( n73824 , n72395 , n73823 );
and ( n73825 , n72393 , n73823 );
or ( n73826 , n72396 , n73824 , n73825 );
or ( n73827 , n72012 , n73826 );
and ( n73828 , n72009 , n73827 );
and ( n73829 , n72007 , n73827 );
or ( n73830 , n72010 , n73828 , n73829 );
and ( n73831 , n71620 , n73830 );
and ( n73832 , n71618 , n73830 );
or ( n73833 , n71621 , n73831 , n73832 );
and ( n73834 , n71214 , n73833 );
and ( n73835 , n70386 , n73833 );
or ( n73836 , n71215 , n73834 , n73835 );
and ( n73837 , n70384 , n73836 );
xor ( n73838 , n70384 , n73836 );
xor ( n73839 , n70386 , n71214 );
xor ( n73840 , n73839 , n73833 );
xor ( n73841 , n71618 , n71620 );
xor ( n73842 , n73841 , n73830 );
xor ( n73843 , n72007 , n72009 );
xor ( n73844 , n73843 , n73827 );
xnor ( n73845 , n72012 , n73826 );
xor ( n73846 , n72393 , n72395 );
xor ( n73847 , n73846 , n73823 );
xor ( n73848 , n72731 , n72733 );
xor ( n73849 , n73848 , n73820 );
not ( n73850 , n73849 );
xor ( n73851 , n72993 , n72995 );
xor ( n73852 , n73851 , n73817 );
xor ( n73853 , n73462 , n73464 );
xor ( n73854 , n73853 , n73814 );
xor ( n73855 , n73467 , n73808 );
xor ( n73856 , n73855 , n73811 );
xor ( n73857 , n73105 , n73107 );
xor ( n73858 , n73857 , n73166 );
xor ( n73859 , n73437 , n73447 );
xor ( n73860 , n73859 , n73450 );
and ( n73861 , n73858 , n73860 );
xor ( n73862 , n73401 , n73403 );
xor ( n73863 , n73862 , n73406 );
xor ( n73864 , n73412 , n73414 );
xor ( n73865 , n73864 , n73417 );
and ( n73866 , n73863 , n73865 );
xor ( n73867 , n73375 , n73377 );
xor ( n73868 , n73867 , n73380 );
xor ( n73869 , n73385 , n73387 );
xor ( n73870 , n73869 , n73390 );
and ( n73871 , n73868 , n73870 );
xor ( n73872 , n73356 , n73358 );
xor ( n73873 , n73872 , n73361 );
xor ( n73874 , n73495 , n73499 );
xor ( n73875 , n73874 , n73502 );
and ( n73876 , n73873 , n73875 );
xor ( n73877 , n73510 , n73515 );
and ( n73878 , n73875 , n73877 );
and ( n73879 , n73873 , n73877 );
or ( n73880 , n73876 , n73878 , n73879 );
and ( n73881 , n73870 , n73880 );
and ( n73882 , n73868 , n73880 );
or ( n73883 , n73871 , n73881 , n73882 );
and ( n73884 , n73865 , n73883 );
and ( n73885 , n73863 , n73883 );
or ( n73886 , n73866 , n73884 , n73885 );
xor ( n73887 , n73519 , n73521 );
and ( n73888 , n69059 , n62868 );
not ( n73889 , n73888 );
and ( n73890 , n68307 , n62998 );
not ( n73891 , n73890 );
and ( n73892 , n73889 , n73891 );
and ( n73893 , n66720 , n64811 );
not ( n73894 , n73893 );
and ( n73895 , n73891 , n73894 );
and ( n73896 , n73889 , n73894 );
or ( n73897 , n73892 , n73895 , n73896 );
and ( n73898 , n62593 , n68752 );
not ( n73899 , n73898 );
and ( n73900 , n63024 , n68610 );
not ( n73901 , n73900 );
and ( n73902 , n73899 , n73901 );
and ( n73903 , n64548 , n66917 );
not ( n73904 , n73903 );
and ( n73905 , n73901 , n73904 );
and ( n73906 , n73899 , n73904 );
or ( n73907 , n73902 , n73905 , n73906 );
and ( n73908 , n73897 , n73907 );
and ( n73909 , n52790 , n54535 );
and ( n73910 , n52612 , n54533 );
nor ( n73911 , n73909 , n73910 );
xnor ( n73912 , n73911 , n54237 );
and ( n73913 , n73908 , n73912 );
and ( n73914 , n73887 , n73913 );
xor ( n73915 , n73507 , n73509 );
xor ( n73916 , n73512 , n73514 );
and ( n73917 , n73915 , n73916 );
and ( n73918 , n73913 , n73917 );
and ( n73919 , n73887 , n73917 );
or ( n73920 , n73914 , n73918 , n73919 );
xor ( n73921 , n73336 , n73339 );
xor ( n73922 , n73921 , n73344 );
xor ( n73923 , n73534 , n73539 );
xor ( n73924 , n73923 , n73544 );
and ( n73925 , n73922 , n73924 );
xor ( n73926 , n73558 , n73568 );
and ( n73927 , n73924 , n73926 );
and ( n73928 , n73922 , n73926 );
or ( n73929 , n73925 , n73927 , n73928 );
xor ( n73930 , n73574 , n73576 );
and ( n73931 , n67997 , n63679 );
not ( n73932 , n73931 );
and ( n73933 , n66980 , n64412 );
not ( n73934 , n73933 );
and ( n73935 , n73932 , n73934 );
and ( n73936 , n65678 , n65586 );
not ( n73937 , n73936 );
and ( n73938 , n73934 , n73937 );
and ( n73939 , n73932 , n73937 );
or ( n73940 , n73935 , n73938 , n73939 );
and ( n73941 , n63492 , n67844 );
not ( n73942 , n73941 );
and ( n73943 , n64221 , n67013 );
not ( n73944 , n73943 );
and ( n73945 , n73942 , n73944 );
and ( n73946 , n65606 , n66005 );
not ( n73947 , n73946 );
and ( n73948 , n73944 , n73947 );
and ( n73949 , n73942 , n73947 );
or ( n73950 , n73945 , n73948 , n73949 );
and ( n73951 , n73940 , n73950 );
and ( n73952 , n73930 , n73951 );
and ( n73953 , n70256 , n61481 );
not ( n73954 , n73953 );
and ( n73955 , n69303 , n62151 );
not ( n73956 , n73955 );
or ( n73957 , n73954 , n73956 );
and ( n73958 , n61505 , n70108 );
not ( n73959 , n73958 );
and ( n73960 , n62377 , n69204 );
not ( n73961 , n73960 );
or ( n73962 , n73959 , n73961 );
and ( n73963 , n73957 , n73962 );
and ( n73964 , n73951 , n73963 );
and ( n73965 , n73930 , n73963 );
or ( n73966 , n73952 , n73964 , n73965 );
and ( n73967 , n73929 , n73966 );
and ( n73968 , n69688 , n61914 );
not ( n73969 , n73968 );
and ( n73970 , n67343 , n63766 );
not ( n73971 , n73970 );
and ( n73972 , n73969 , n73971 );
and ( n73973 , n61918 , n69507 );
not ( n73974 , n73973 );
and ( n73975 , n63987 , n67411 );
not ( n73976 , n73975 );
and ( n73977 , n73974 , n73976 );
and ( n73978 , n73972 , n73977 );
xor ( n73979 , n73550 , n73552 );
xor ( n73980 , n73979 , n73555 );
xor ( n73981 , n73560 , n73562 );
xor ( n73982 , n73981 , n73565 );
and ( n73983 , n73980 , n73982 );
and ( n73984 , n73978 , n73983 );
xor ( n73985 , n73599 , n73603 );
xor ( n73986 , n73985 , n73608 );
xor ( n73987 , n73614 , n73616 );
xor ( n73988 , n73987 , n73619 );
and ( n73989 , n73986 , n73988 );
buf ( n73990 , n73989 );
and ( n73991 , n73983 , n73990 );
and ( n73992 , n73978 , n73990 );
or ( n73993 , n73984 , n73991 , n73992 );
and ( n73994 , n73966 , n73993 );
and ( n73995 , n73929 , n73993 );
or ( n73996 , n73967 , n73994 , n73995 );
and ( n73997 , n73920 , n73996 );
xor ( n73998 , n73627 , n73629 );
xor ( n73999 , n73998 , n73632 );
xor ( n74000 , n73637 , n73639 );
and ( n74001 , n73999 , n74000 );
xor ( n74002 , n73643 , n73645 );
and ( n74003 , n74000 , n74002 );
and ( n74004 , n73999 , n74002 );
or ( n74005 , n74001 , n74003 , n74004 );
xor ( n74006 , n73531 , n73533 );
xor ( n74007 , n73536 , n73538 );
and ( n74008 , n74006 , n74007 );
and ( n74009 , n65177 , n66469 );
not ( n74010 , n74009 );
and ( n74011 , n66415 , n65210 );
not ( n74012 , n74011 );
and ( n74013 , n74010 , n74012 );
and ( n74014 , n74007 , n74013 );
and ( n74015 , n74006 , n74013 );
or ( n74016 , n74008 , n74014 , n74015 );
and ( n74017 , n74005 , n74016 );
and ( n74018 , n51298 , n57187 );
and ( n74019 , n51077 , n57184 );
nor ( n74020 , n74018 , n74019 );
xnor ( n74021 , n74020 , n56175 );
and ( n74022 , n51734 , n56503 );
and ( n74023 , n51510 , n56501 );
nor ( n74024 , n74022 , n74023 );
xnor ( n74025 , n74024 , n56178 );
and ( n74026 , n74021 , n74025 );
and ( n74027 , n52332 , n55851 );
and ( n74028 , n52082 , n55849 );
nor ( n74029 , n74027 , n74028 );
xnor ( n74030 , n74029 , n55506 );
and ( n74031 , n74025 , n74030 );
and ( n74032 , n74021 , n74030 );
or ( n74033 , n74026 , n74031 , n74032 );
and ( n74034 , n52790 , n55159 );
and ( n74035 , n52612 , n55157 );
nor ( n74036 , n74034 , n74035 );
xnor ( n74037 , n74036 , n54864 );
and ( n74038 , n53922 , n53928 );
and ( n74039 , n53639 , n53926 );
nor ( n74040 , n74038 , n74039 );
xnor ( n74041 , n74040 , n53652 );
and ( n74042 , n74037 , n74041 );
and ( n74043 , n54604 , n53357 );
and ( n74044 , n54227 , n53355 );
nor ( n74045 , n74043 , n74044 );
xnor ( n74046 , n74045 , n53060 );
and ( n74047 , n74041 , n74046 );
and ( n74048 , n74037 , n74046 );
or ( n74049 , n74042 , n74047 , n74048 );
and ( n74050 , n74033 , n74049 );
and ( n74051 , n55143 , n52799 );
and ( n74052 , n54942 , n52797 );
nor ( n74053 , n74051 , n74052 );
xnor ( n74054 , n74053 , n52538 );
and ( n74055 , n55756 , n52269 );
and ( n74056 , n55497 , n52267 );
nor ( n74057 , n74055 , n74056 );
xnor ( n74058 , n74057 , n52008 );
and ( n74059 , n74054 , n74058 );
and ( n74060 , n56388 , n51750 );
and ( n74061 , n56255 , n51748 );
nor ( n74062 , n74060 , n74061 );
xnor ( n74063 , n74062 , n51520 );
and ( n74064 , n74058 , n74063 );
and ( n74065 , n74054 , n74063 );
or ( n74066 , n74059 , n74064 , n74065 );
and ( n74067 , n74049 , n74066 );
and ( n74068 , n74033 , n74066 );
or ( n74069 , n74050 , n74067 , n74068 );
and ( n74070 , n74016 , n74069 );
and ( n74071 , n74005 , n74069 );
or ( n74072 , n74017 , n74070 , n74071 );
and ( n74073 , n57063 , n51221 );
and ( n74074 , n56915 , n51219 );
nor ( n74075 , n74073 , n74074 );
xnor ( n74076 , n74075 , n51000 );
and ( n74077 , n57063 , n51219 );
not ( n74078 , n74077 );
and ( n74079 , n74078 , n51000 );
and ( n74080 , n74076 , n74079 );
xor ( n74081 , n45384 , n45515 );
buf ( n74082 , n74081 );
buf ( n74083 , n74082 );
buf ( n74084 , n74083 );
and ( n74085 , n74079 , n74084 );
and ( n74086 , n74076 , n74084 );
or ( n74087 , n74080 , n74085 , n74086 );
xor ( n74088 , n73654 , n73658 );
xor ( n74089 , n74088 , n73663 );
and ( n74090 , n74087 , n74089 );
xor ( n74091 , n73670 , n73674 );
xor ( n74092 , n74091 , n73679 );
and ( n74093 , n74089 , n74092 );
and ( n74094 , n74087 , n74092 );
or ( n74095 , n74090 , n74093 , n74094 );
buf ( n74096 , n73579 );
xor ( n74097 , n74096 , n73580 );
and ( n74098 , n74095 , n74097 );
xor ( n74099 , n73584 , n73585 );
xor ( n74100 , n74099 , n73587 );
and ( n74101 , n74097 , n74100 );
and ( n74102 , n74095 , n74100 );
or ( n74103 , n74098 , n74101 , n74102 );
and ( n74104 , n74072 , n74103 );
xor ( n74105 , n73595 , n73611 );
xor ( n74106 , n74105 , n73622 );
xor ( n74107 , n73635 , n73640 );
xor ( n74108 , n74107 , n73646 );
and ( n74109 , n74106 , n74108 );
xor ( n74110 , n73666 , n73682 );
xor ( n74111 , n74110 , n73695 );
and ( n74112 , n74108 , n74111 );
and ( n74113 , n74106 , n74111 );
or ( n74114 , n74109 , n74112 , n74113 );
and ( n74115 , n74103 , n74114 );
and ( n74116 , n74072 , n74114 );
or ( n74117 , n74104 , n74115 , n74116 );
and ( n74118 , n73996 , n74117 );
and ( n74119 , n73920 , n74117 );
or ( n74120 , n73997 , n74118 , n74119 );
xor ( n74121 , n73529 , n73547 );
xor ( n74122 , n74121 , n73569 );
xor ( n74123 , n73577 , n73582 );
xor ( n74124 , n74123 , n73590 );
and ( n74125 , n74122 , n74124 );
xor ( n74126 , n73625 , n73649 );
xor ( n74127 , n74126 , n73698 );
and ( n74128 , n74124 , n74127 );
and ( n74129 , n74122 , n74127 );
or ( n74130 , n74125 , n74128 , n74129 );
xor ( n74131 , n73484 , n73485 );
xor ( n74132 , n74131 , n73487 );
and ( n74133 , n74130 , n74132 );
xor ( n74134 , n73505 , n73516 );
xor ( n74135 , n74134 , n73522 );
and ( n74136 , n74132 , n74135 );
and ( n74137 , n74130 , n74135 );
or ( n74138 , n74133 , n74136 , n74137 );
and ( n74139 , n74120 , n74138 );
xor ( n74140 , n73572 , n73593 );
xor ( n74141 , n74140 , n73701 );
xor ( n74142 , n73730 , n73740 );
xor ( n74143 , n74142 , n73743 );
and ( n74144 , n74141 , n74143 );
xor ( n74145 , n73749 , n73751 );
xor ( n74146 , n74145 , n73754 );
and ( n74147 , n74143 , n74146 );
and ( n74148 , n74141 , n74146 );
or ( n74149 , n74144 , n74147 , n74148 );
and ( n74150 , n74138 , n74149 );
and ( n74151 , n74120 , n74149 );
or ( n74152 , n74139 , n74150 , n74151 );
and ( n74153 , n73886 , n74152 );
xor ( n74154 , n73482 , n73490 );
xor ( n74155 , n74154 , n73525 );
xor ( n74156 , n73704 , n73746 );
xor ( n74157 , n74156 , n73757 );
and ( n74158 , n74155 , n74157 );
xor ( n74159 , n73763 , n73765 );
xor ( n74160 , n74159 , n73768 );
and ( n74161 , n74157 , n74160 );
and ( n74162 , n74155 , n74160 );
or ( n74163 , n74158 , n74161 , n74162 );
and ( n74164 , n74152 , n74163 );
and ( n74165 , n73886 , n74163 );
or ( n74166 , n74153 , n74164 , n74165 );
xor ( n74167 , n73473 , n73475 );
xor ( n74168 , n74167 , n73477 );
xor ( n74169 , n73528 , n73760 );
xor ( n74170 , n74169 , n73771 );
and ( n74171 , n74168 , n74170 );
xor ( n74172 , n73777 , n73779 );
xor ( n74173 , n74172 , n73782 );
and ( n74174 , n74170 , n74173 );
and ( n74175 , n74168 , n74173 );
or ( n74176 , n74171 , n74174 , n74175 );
and ( n74177 , n74166 , n74176 );
xor ( n74178 , n73480 , n73774 );
xor ( n74179 , n74178 , n73785 );
and ( n74180 , n74176 , n74179 );
and ( n74181 , n74166 , n74179 );
or ( n74182 , n74177 , n74180 , n74181 );
and ( n74183 , n73860 , n74182 );
and ( n74184 , n73858 , n74182 );
or ( n74185 , n73861 , n74183 , n74184 );
xor ( n74186 , n73469 , n73802 );
xor ( n74187 , n74186 , n73805 );
and ( n74188 , n74185 , n74187 );
xor ( n74189 , n73471 , n73788 );
xor ( n74190 , n74189 , n73799 );
xor ( n74191 , n73791 , n73793 );
xor ( n74192 , n74191 , n73796 );
xor ( n74193 , n73722 , n73724 );
xor ( n74194 , n74193 , n73727 );
xor ( n74195 , n73732 , n73734 );
xor ( n74196 , n74195 , n73737 );
and ( n74197 , n74194 , n74196 );
xor ( n74198 , n73714 , n73716 );
xor ( n74199 , n74198 , n73719 );
xor ( n74200 , n73908 , n73912 );
and ( n74201 , n74199 , n74200 );
xor ( n74202 , n73915 , n73916 );
and ( n74203 , n74200 , n74202 );
and ( n74204 , n74199 , n74202 );
or ( n74205 , n74201 , n74203 , n74204 );
and ( n74206 , n74196 , n74205 );
and ( n74207 , n74194 , n74205 );
or ( n74208 , n74197 , n74206 , n74207 );
and ( n74209 , n70256 , n61914 );
not ( n74210 , n74209 );
and ( n74211 , n69303 , n62868 );
not ( n74212 , n74211 );
and ( n74213 , n74210 , n74212 );
and ( n74214 , n67997 , n63766 );
not ( n74215 , n74214 );
and ( n74216 , n74212 , n74215 );
and ( n74217 , n74210 , n74215 );
or ( n74218 , n74213 , n74216 , n74217 );
and ( n74219 , n61918 , n70108 );
not ( n74220 , n74219 );
and ( n74221 , n62593 , n69204 );
not ( n74222 , n74221 );
and ( n74223 , n74220 , n74222 );
and ( n74224 , n63987 , n67844 );
not ( n74225 , n74224 );
and ( n74226 , n74222 , n74225 );
and ( n74227 , n74220 , n74225 );
or ( n74228 , n74223 , n74226 , n74227 );
and ( n74229 , n74218 , n74228 );
and ( n74230 , n53041 , n54535 );
and ( n74231 , n52790 , n54533 );
nor ( n74232 , n74230 , n74231 );
xnor ( n74233 , n74232 , n54237 );
and ( n74234 , n74229 , n74233 );
xor ( n74235 , n73687 , n73337 );
xor ( n74236 , n74235 , n73692 );
xor ( n74237 , n73706 , n73708 );
xor ( n74238 , n74237 , n73711 );
and ( n74239 , n74236 , n74238 );
xor ( n74240 , n73940 , n73950 );
and ( n74241 , n74238 , n74240 );
and ( n74242 , n74236 , n74240 );
or ( n74243 , n74239 , n74241 , n74242 );
and ( n74244 , n74234 , n74243 );
xor ( n74245 , n73897 , n73907 );
xor ( n74246 , n73957 , n73962 );
and ( n74247 , n74245 , n74246 );
xor ( n74248 , n73972 , n73977 );
and ( n74249 , n74246 , n74248 );
and ( n74250 , n74245 , n74248 );
or ( n74251 , n74247 , n74249 , n74250 );
and ( n74252 , n74243 , n74251 );
and ( n74253 , n74234 , n74251 );
or ( n74254 , n74244 , n74252 , n74253 );
xor ( n74255 , n73980 , n73982 );
and ( n74256 , n62377 , n69507 );
not ( n74257 , n74256 );
and ( n74258 , n69688 , n62151 );
not ( n74259 , n74258 );
and ( n74260 , n74257 , n74259 );
and ( n74261 , n53328 , n54535 );
and ( n74262 , n53041 , n54533 );
nor ( n74263 , n74261 , n74262 );
xnor ( n74264 , n74263 , n54237 );
and ( n74265 , n74260 , n74264 );
and ( n74266 , n74255 , n74265 );
xor ( n74267 , n73932 , n73934 );
xor ( n74268 , n74267 , n73937 );
xor ( n74269 , n73942 , n73944 );
xor ( n74270 , n74269 , n73947 );
and ( n74271 , n74268 , n74270 );
and ( n74272 , n74265 , n74271 );
and ( n74273 , n74255 , n74271 );
or ( n74274 , n74266 , n74272 , n74273 );
xor ( n74275 , n73889 , n73891 );
xor ( n74276 , n74275 , n73894 );
xor ( n74277 , n73899 , n73901 );
xor ( n74278 , n74277 , n73904 );
and ( n74279 , n74276 , n74278 );
xnor ( n74280 , n73954 , n73956 );
xnor ( n74281 , n73959 , n73961 );
and ( n74282 , n74280 , n74281 );
and ( n74283 , n74279 , n74282 );
xor ( n74284 , n73969 , n73971 );
xor ( n74285 , n73974 , n73976 );
and ( n74286 , n74284 , n74285 );
and ( n74287 , n74282 , n74286 );
and ( n74288 , n74279 , n74286 );
or ( n74289 , n74283 , n74287 , n74288 );
and ( n74290 , n74274 , n74289 );
xor ( n74291 , n74010 , n74012 );
and ( n74292 , n53041 , n55159 );
and ( n74293 , n52790 , n55157 );
nor ( n74294 , n74292 , n74293 );
xnor ( n74295 , n74294 , n54864 );
and ( n74296 , n53639 , n54535 );
and ( n74297 , n53328 , n54533 );
nor ( n74298 , n74296 , n74297 );
xnor ( n74299 , n74298 , n54237 );
and ( n74300 , n74295 , n74299 );
and ( n74301 , n55497 , n52799 );
and ( n74302 , n55143 , n52797 );
nor ( n74303 , n74301 , n74302 );
xnor ( n74304 , n74303 , n52538 );
and ( n74305 , n74299 , n74304 );
and ( n74306 , n74295 , n74304 );
or ( n74307 , n74300 , n74305 , n74306 );
and ( n74308 , n74291 , n74307 );
buf ( n74309 , n74308 );
and ( n74310 , n63492 , n68610 );
not ( n74311 , n74310 );
and ( n74312 , n64548 , n67013 );
not ( n74313 , n74312 );
and ( n74314 , n74311 , n74313 );
buf ( n74315 , n65678 );
not ( n74316 , n74315 );
and ( n74317 , n74313 , n74316 );
and ( n74318 , n74311 , n74316 );
or ( n74319 , n74314 , n74317 , n74318 );
and ( n74320 , n68307 , n63679 );
not ( n74321 , n74320 );
and ( n74322 , n64221 , n67411 );
not ( n74323 , n74322 );
and ( n74324 , n74321 , n74323 );
and ( n74325 , n65606 , n66469 );
not ( n74326 , n74325 );
and ( n74327 , n74323 , n74326 );
and ( n74328 , n74321 , n74326 );
or ( n74329 , n74324 , n74327 , n74328 );
and ( n74330 , n74319 , n74329 );
and ( n74331 , n67343 , n64412 );
and ( n74332 , n66415 , n65586 );
not ( n74333 , n74332 );
and ( n74334 , n74331 , n74333 );
and ( n74335 , n74329 , n74334 );
and ( n74336 , n74319 , n74334 );
or ( n74337 , n74330 , n74335 , n74336 );
and ( n74338 , n74309 , n74337 );
not ( n74339 , n74331 );
buf ( n74340 , n74339 );
and ( n74341 , n63024 , n68752 );
not ( n74342 , n74341 );
and ( n74343 , n69059 , n62998 );
not ( n74344 , n74343 );
and ( n74345 , n74342 , n74344 );
and ( n74346 , n74340 , n74345 );
and ( n74347 , n65177 , n66917 );
not ( n74348 , n74347 );
and ( n74349 , n66720 , n65210 );
not ( n74350 , n74349 );
and ( n74351 , n74348 , n74350 );
and ( n74352 , n74345 , n74351 );
and ( n74353 , n74340 , n74351 );
or ( n74354 , n74346 , n74352 , n74353 );
and ( n74355 , n74337 , n74354 );
and ( n74356 , n74309 , n74354 );
or ( n74357 , n74338 , n74355 , n74356 );
and ( n74358 , n74289 , n74357 );
and ( n74359 , n74274 , n74357 );
or ( n74360 , n74290 , n74358 , n74359 );
and ( n74361 , n74254 , n74360 );
and ( n74362 , n51510 , n57187 );
and ( n74363 , n51298 , n57184 );
nor ( n74364 , n74362 , n74363 );
xnor ( n74365 , n74364 , n56175 );
and ( n74366 , n52082 , n56503 );
and ( n74367 , n51734 , n56501 );
nor ( n74368 , n74366 , n74367 );
xnor ( n74369 , n74368 , n56178 );
and ( n74370 , n74365 , n74369 );
and ( n74371 , n54227 , n53928 );
and ( n74372 , n53922 , n53926 );
nor ( n74373 , n74371 , n74372 );
xnor ( n74374 , n74373 , n53652 );
and ( n74375 , n74369 , n74374 );
and ( n74376 , n74365 , n74374 );
or ( n74377 , n74370 , n74375 , n74376 );
and ( n74378 , n54942 , n53357 );
and ( n74379 , n54604 , n53355 );
nor ( n74380 , n74378 , n74379 );
xnor ( n74381 , n74380 , n53060 );
and ( n74382 , n56255 , n52269 );
and ( n74383 , n55756 , n52267 );
nor ( n74384 , n74382 , n74383 );
xnor ( n74385 , n74384 , n52008 );
and ( n74386 , n74381 , n74385 );
and ( n74387 , n56915 , n51750 );
and ( n74388 , n56388 , n51748 );
nor ( n74389 , n74387 , n74388 );
xnor ( n74390 , n74389 , n51520 );
and ( n74391 , n74385 , n74390 );
and ( n74392 , n74381 , n74390 );
or ( n74393 , n74386 , n74391 , n74392 );
and ( n74394 , n74377 , n74393 );
xor ( n74395 , n45385 , n45514 );
buf ( n74396 , n74395 );
buf ( n74397 , n74396 );
buf ( n74398 , n74397 );
and ( n74399 , n74077 , n74398 );
and ( n74400 , n66980 , n64811 );
not ( n74401 , n74400 );
and ( n74402 , n74398 , n74401 );
and ( n74403 , n74077 , n74401 );
or ( n74404 , n74399 , n74402 , n74403 );
and ( n74405 , n74393 , n74404 );
and ( n74406 , n74377 , n74404 );
or ( n74407 , n74394 , n74405 , n74406 );
xor ( n74408 , n74021 , n74025 );
xor ( n74409 , n74408 , n74030 );
xor ( n74410 , n74037 , n74041 );
xor ( n74411 , n74410 , n74046 );
and ( n74412 , n74409 , n74411 );
xor ( n74413 , n74054 , n74058 );
xor ( n74414 , n74413 , n74063 );
and ( n74415 , n74411 , n74414 );
and ( n74416 , n74409 , n74414 );
or ( n74417 , n74412 , n74415 , n74416 );
and ( n74418 , n74407 , n74417 );
buf ( n74419 , n73986 );
xor ( n74420 , n74419 , n73988 );
and ( n74421 , n74417 , n74420 );
and ( n74422 , n74407 , n74420 );
or ( n74423 , n74418 , n74421 , n74422 );
xor ( n74424 , n73999 , n74000 );
xor ( n74425 , n74424 , n74002 );
xor ( n74426 , n74006 , n74007 );
xor ( n74427 , n74426 , n74013 );
and ( n74428 , n74425 , n74427 );
xor ( n74429 , n74033 , n74049 );
xor ( n74430 , n74429 , n74066 );
and ( n74431 , n74427 , n74430 );
and ( n74432 , n74425 , n74430 );
or ( n74433 , n74428 , n74431 , n74432 );
and ( n74434 , n74423 , n74433 );
xor ( n74435 , n73922 , n73924 );
xor ( n74436 , n74435 , n73926 );
and ( n74437 , n74433 , n74436 );
and ( n74438 , n74423 , n74436 );
or ( n74439 , n74434 , n74437 , n74438 );
and ( n74440 , n74360 , n74439 );
and ( n74441 , n74254 , n74439 );
or ( n74442 , n74361 , n74440 , n74441 );
and ( n74443 , n74208 , n74442 );
xor ( n74444 , n73930 , n73951 );
xor ( n74445 , n74444 , n73963 );
xor ( n74446 , n73978 , n73983 );
xor ( n74447 , n74446 , n73990 );
and ( n74448 , n74445 , n74447 );
xor ( n74449 , n74005 , n74016 );
xor ( n74450 , n74449 , n74069 );
and ( n74451 , n74447 , n74450 );
and ( n74452 , n74445 , n74450 );
or ( n74453 , n74448 , n74451 , n74452 );
xor ( n74454 , n73873 , n73875 );
xor ( n74455 , n74454 , n73877 );
and ( n74456 , n74453 , n74455 );
xor ( n74457 , n73887 , n73913 );
xor ( n74458 , n74457 , n73917 );
and ( n74459 , n74455 , n74458 );
and ( n74460 , n74453 , n74458 );
or ( n74461 , n74456 , n74459 , n74460 );
and ( n74462 , n74442 , n74461 );
and ( n74463 , n74208 , n74461 );
or ( n74464 , n74443 , n74462 , n74463 );
xor ( n74465 , n73929 , n73966 );
xor ( n74466 , n74465 , n73993 );
xor ( n74467 , n74072 , n74103 );
xor ( n74468 , n74467 , n74114 );
and ( n74469 , n74466 , n74468 );
xor ( n74470 , n74122 , n74124 );
xor ( n74471 , n74470 , n74127 );
and ( n74472 , n74468 , n74471 );
and ( n74473 , n74466 , n74471 );
or ( n74474 , n74469 , n74472 , n74473 );
xor ( n74475 , n73868 , n73870 );
xor ( n74476 , n74475 , n73880 );
and ( n74477 , n74474 , n74476 );
xor ( n74478 , n73920 , n73996 );
xor ( n74479 , n74478 , n74117 );
and ( n74480 , n74476 , n74479 );
and ( n74481 , n74474 , n74479 );
or ( n74482 , n74477 , n74480 , n74481 );
and ( n74483 , n74464 , n74482 );
xor ( n74484 , n73863 , n73865 );
xor ( n74485 , n74484 , n73883 );
and ( n74486 , n74482 , n74485 );
and ( n74487 , n74464 , n74485 );
or ( n74488 , n74483 , n74486 , n74487 );
xor ( n74489 , n73886 , n74152 );
xor ( n74490 , n74489 , n74163 );
and ( n74491 , n74488 , n74490 );
xor ( n74492 , n74168 , n74170 );
xor ( n74493 , n74492 , n74173 );
and ( n74494 , n74490 , n74493 );
and ( n74495 , n74488 , n74493 );
or ( n74496 , n74491 , n74494 , n74495 );
and ( n74497 , n74192 , n74496 );
xor ( n74498 , n74166 , n74176 );
xor ( n74499 , n74498 , n74179 );
and ( n74500 , n74496 , n74499 );
and ( n74501 , n74192 , n74499 );
or ( n74502 , n74497 , n74500 , n74501 );
and ( n74503 , n74190 , n74502 );
xor ( n74504 , n73858 , n73860 );
xor ( n74505 , n74504 , n74182 );
and ( n74506 , n74502 , n74505 );
and ( n74507 , n74190 , n74505 );
or ( n74508 , n74503 , n74506 , n74507 );
and ( n74509 , n74187 , n74508 );
and ( n74510 , n74185 , n74508 );
or ( n74511 , n74188 , n74509 , n74510 );
and ( n74512 , n73856 , n74511 );
xor ( n74513 , n73856 , n74511 );
xor ( n74514 , n74185 , n74187 );
xor ( n74515 , n74514 , n74508 );
not ( n74516 , n74515 );
xor ( n74517 , n74190 , n74502 );
xor ( n74518 , n74517 , n74505 );
xor ( n74519 , n74192 , n74496 );
xor ( n74520 , n74519 , n74499 );
xor ( n74521 , n74120 , n74138 );
xor ( n74522 , n74521 , n74149 );
xor ( n74523 , n74155 , n74157 );
xor ( n74524 , n74523 , n74160 );
and ( n74525 , n74522 , n74524 );
xor ( n74526 , n74130 , n74132 );
xor ( n74527 , n74526 , n74135 );
xor ( n74528 , n74141 , n74143 );
xor ( n74529 , n74528 , n74146 );
and ( n74530 , n74527 , n74529 );
xor ( n74531 , n74095 , n74097 );
xor ( n74532 , n74531 , n74100 );
xor ( n74533 , n74106 , n74108 );
xor ( n74534 , n74533 , n74111 );
and ( n74535 , n74532 , n74534 );
xor ( n74536 , n74087 , n74089 );
xor ( n74537 , n74536 , n74092 );
xor ( n74538 , n74229 , n74233 );
and ( n74539 , n74537 , n74538 );
xor ( n74540 , n74076 , n74079 );
xor ( n74541 , n74540 , n74084 );
xor ( n74542 , n74260 , n74264 );
and ( n74543 , n74541 , n74542 );
xor ( n74544 , n74218 , n74228 );
and ( n74545 , n74542 , n74544 );
and ( n74546 , n74541 , n74544 );
or ( n74547 , n74543 , n74545 , n74546 );
and ( n74548 , n74538 , n74547 );
and ( n74549 , n74537 , n74547 );
or ( n74550 , n74539 , n74548 , n74549 );
and ( n74551 , n74534 , n74550 );
and ( n74552 , n74532 , n74550 );
or ( n74553 , n74535 , n74551 , n74552 );
xor ( n74554 , n74268 , n74270 );
xor ( n74555 , n74276 , n74278 );
and ( n74556 , n74554 , n74555 );
xor ( n74557 , n74280 , n74281 );
and ( n74558 , n74555 , n74557 );
and ( n74559 , n74554 , n74557 );
or ( n74560 , n74556 , n74558 , n74559 );
xor ( n74561 , n74284 , n74285 );
and ( n74562 , n52612 , n55851 );
and ( n74563 , n52332 , n55849 );
nor ( n74564 , n74562 , n74563 );
xnor ( n74565 , n74564 , n55506 );
xor ( n74566 , n74295 , n74299 );
xor ( n74567 , n74566 , n74304 );
and ( n74568 , n74565 , n74567 );
and ( n74569 , n74561 , n74568 );
and ( n74570 , n69059 , n63679 );
not ( n74571 , n74570 );
and ( n74572 , n66980 , n65210 );
not ( n74573 , n74572 );
and ( n74574 , n74571 , n74573 );
and ( n74575 , n66415 , n66005 );
not ( n74576 , n74575 );
and ( n74577 , n74573 , n74576 );
and ( n74578 , n74571 , n74576 );
or ( n74579 , n74574 , n74577 , n74578 );
and ( n74580 , n63492 , n68752 );
not ( n74581 , n74580 );
and ( n74582 , n65177 , n67013 );
not ( n74583 , n74582 );
and ( n74584 , n74581 , n74583 );
and ( n74585 , n65678 , n66469 );
not ( n74586 , n74585 );
and ( n74587 , n74583 , n74586 );
and ( n74588 , n74581 , n74586 );
or ( n74589 , n74584 , n74587 , n74588 );
and ( n74590 , n74579 , n74589 );
and ( n74591 , n74568 , n74590 );
and ( n74592 , n74561 , n74590 );
or ( n74593 , n74569 , n74591 , n74592 );
and ( n74594 , n74560 , n74593 );
and ( n74595 , n68307 , n63766 );
not ( n74596 , n74595 );
and ( n74597 , n67997 , n64412 );
not ( n74598 , n74597 );
and ( n74599 , n74596 , n74598 );
and ( n74600 , n67343 , n64811 );
not ( n74601 , n74600 );
and ( n74602 , n74598 , n74601 );
and ( n74603 , n74596 , n74601 );
or ( n74604 , n74599 , n74602 , n74603 );
and ( n74605 , n63987 , n68610 );
not ( n74606 , n74605 );
and ( n74607 , n64221 , n67844 );
not ( n74608 , n74607 );
and ( n74609 , n74606 , n74608 );
and ( n74610 , n64548 , n67411 );
not ( n74611 , n74610 );
and ( n74612 , n74608 , n74611 );
and ( n74613 , n74606 , n74611 );
or ( n74614 , n74609 , n74612 , n74613 );
and ( n74615 , n74604 , n74614 );
xor ( n74616 , n74210 , n74212 );
xor ( n74617 , n74616 , n74215 );
xor ( n74618 , n74220 , n74222 );
xor ( n74619 , n74618 , n74225 );
and ( n74620 , n74617 , n74619 );
and ( n74621 , n74615 , n74620 );
xor ( n74622 , n74311 , n74313 );
xor ( n74623 , n74622 , n74316 );
xor ( n74624 , n74321 , n74323 );
xor ( n74625 , n74624 , n74326 );
and ( n74626 , n74623 , n74625 );
buf ( n74627 , n74626 );
and ( n74628 , n74620 , n74627 );
and ( n74629 , n74615 , n74627 );
or ( n74630 , n74621 , n74628 , n74629 );
and ( n74631 , n74593 , n74630 );
and ( n74632 , n74560 , n74630 );
or ( n74633 , n74594 , n74631 , n74632 );
xor ( n74634 , n74331 , n74333 );
xor ( n74635 , n74257 , n74259 );
and ( n74636 , n74634 , n74635 );
xor ( n74637 , n74342 , n74344 );
and ( n74638 , n74635 , n74637 );
and ( n74639 , n74634 , n74637 );
or ( n74640 , n74636 , n74638 , n74639 );
xor ( n74641 , n74348 , n74350 );
and ( n74642 , n65606 , n66917 );
not ( n74643 , n74642 );
and ( n74644 , n66720 , n65586 );
not ( n74645 , n74644 );
and ( n74646 , n74643 , n74645 );
and ( n74647 , n74641 , n74646 );
and ( n74648 , n51734 , n57187 );
and ( n74649 , n51510 , n57184 );
nor ( n74650 , n74648 , n74649 );
xnor ( n74651 , n74650 , n56175 );
and ( n74652 , n52332 , n56503 );
and ( n74653 , n52082 , n56501 );
nor ( n74654 , n74652 , n74653 );
xnor ( n74655 , n74654 , n56178 );
and ( n74656 , n74651 , n74655 );
and ( n74657 , n52790 , n55851 );
and ( n74658 , n52612 , n55849 );
nor ( n74659 , n74657 , n74658 );
xnor ( n74660 , n74659 , n55506 );
and ( n74661 , n74655 , n74660 );
and ( n74662 , n74651 , n74660 );
or ( n74663 , n74656 , n74661 , n74662 );
and ( n74664 , n74646 , n74663 );
and ( n74665 , n74641 , n74663 );
or ( n74666 , n74647 , n74664 , n74665 );
and ( n74667 , n74640 , n74666 );
and ( n74668 , n53328 , n55159 );
and ( n74669 , n53041 , n55157 );
nor ( n74670 , n74668 , n74669 );
xnor ( n74671 , n74670 , n54864 );
and ( n74672 , n53922 , n54535 );
and ( n74673 , n53639 , n54533 );
nor ( n74674 , n74672 , n74673 );
xnor ( n74675 , n74674 , n54237 );
and ( n74676 , n74671 , n74675 );
and ( n74677 , n54604 , n53928 );
and ( n74678 , n54227 , n53926 );
nor ( n74679 , n74677 , n74678 );
xnor ( n74680 , n74679 , n53652 );
and ( n74681 , n74675 , n74680 );
and ( n74682 , n74671 , n74680 );
or ( n74683 , n74676 , n74681 , n74682 );
and ( n74684 , n55756 , n52799 );
and ( n74685 , n55497 , n52797 );
nor ( n74686 , n74684 , n74685 );
xnor ( n74687 , n74686 , n52538 );
and ( n74688 , n56388 , n52269 );
and ( n74689 , n56255 , n52267 );
nor ( n74690 , n74688 , n74689 );
xnor ( n74691 , n74690 , n52008 );
and ( n74692 , n74687 , n74691 );
and ( n74693 , n57063 , n51750 );
and ( n74694 , n56915 , n51748 );
nor ( n74695 , n74693 , n74694 );
xnor ( n74696 , n74695 , n51520 );
and ( n74697 , n74691 , n74696 );
and ( n74698 , n74687 , n74696 );
or ( n74699 , n74692 , n74697 , n74698 );
and ( n74700 , n74683 , n74699 );
and ( n74701 , n57063 , n51748 );
not ( n74702 , n74701 );
and ( n74703 , n74702 , n51520 );
xor ( n74704 , n45387 , n45513 );
buf ( n74705 , n74704 );
buf ( n74706 , n74705 );
buf ( n74707 , n74706 );
and ( n74708 , n74703 , n74707 );
and ( n74709 , n70256 , n62151 );
not ( n74710 , n74709 );
and ( n74711 , n74707 , n74710 );
and ( n74712 , n74703 , n74710 );
or ( n74713 , n74708 , n74711 , n74712 );
and ( n74714 , n74699 , n74713 );
and ( n74715 , n74683 , n74713 );
or ( n74716 , n74700 , n74714 , n74715 );
and ( n74717 , n74666 , n74716 );
and ( n74718 , n74640 , n74716 );
or ( n74719 , n74667 , n74717 , n74718 );
xor ( n74720 , n74365 , n74369 );
xor ( n74721 , n74720 , n74374 );
xor ( n74722 , n74381 , n74385 );
xor ( n74723 , n74722 , n74390 );
and ( n74724 , n74721 , n74723 );
xor ( n74725 , n74077 , n74398 );
xor ( n74726 , n74725 , n74401 );
and ( n74727 , n74723 , n74726 );
and ( n74728 , n74721 , n74726 );
or ( n74729 , n74724 , n74727 , n74728 );
buf ( n74730 , n74291 );
xor ( n74731 , n74730 , n74307 );
and ( n74732 , n74729 , n74731 );
xor ( n74733 , n74319 , n74329 );
xor ( n74734 , n74733 , n74334 );
and ( n74735 , n74731 , n74734 );
and ( n74736 , n74729 , n74734 );
or ( n74737 , n74732 , n74735 , n74736 );
and ( n74738 , n74719 , n74737 );
xor ( n74739 , n74340 , n74345 );
xor ( n74740 , n74739 , n74351 );
xor ( n74741 , n74377 , n74393 );
xor ( n74742 , n74741 , n74404 );
and ( n74743 , n74740 , n74742 );
xor ( n74744 , n74409 , n74411 );
xor ( n74745 , n74744 , n74414 );
and ( n74746 , n74742 , n74745 );
and ( n74747 , n74740 , n74745 );
or ( n74748 , n74743 , n74746 , n74747 );
and ( n74749 , n74737 , n74748 );
and ( n74750 , n74719 , n74748 );
or ( n74751 , n74738 , n74749 , n74750 );
and ( n74752 , n74633 , n74751 );
xor ( n74753 , n74236 , n74238 );
xor ( n74754 , n74753 , n74240 );
xor ( n74755 , n74245 , n74246 );
xor ( n74756 , n74755 , n74248 );
and ( n74757 , n74754 , n74756 );
xor ( n74758 , n74255 , n74265 );
xor ( n74759 , n74758 , n74271 );
and ( n74760 , n74756 , n74759 );
and ( n74761 , n74754 , n74759 );
or ( n74762 , n74757 , n74760 , n74761 );
and ( n74763 , n74751 , n74762 );
and ( n74764 , n74633 , n74762 );
or ( n74765 , n74752 , n74763 , n74764 );
and ( n74766 , n74553 , n74765 );
xor ( n74767 , n74279 , n74282 );
xor ( n74768 , n74767 , n74286 );
xor ( n74769 , n74309 , n74337 );
xor ( n74770 , n74769 , n74354 );
and ( n74771 , n74768 , n74770 );
xor ( n74772 , n74407 , n74417 );
xor ( n74773 , n74772 , n74420 );
and ( n74774 , n74770 , n74773 );
and ( n74775 , n74768 , n74773 );
or ( n74776 , n74771 , n74774 , n74775 );
xor ( n74777 , n74199 , n74200 );
xor ( n74778 , n74777 , n74202 );
and ( n74779 , n74776 , n74778 );
xor ( n74780 , n74234 , n74243 );
xor ( n74781 , n74780 , n74251 );
and ( n74782 , n74778 , n74781 );
and ( n74783 , n74776 , n74781 );
or ( n74784 , n74779 , n74782 , n74783 );
and ( n74785 , n74765 , n74784 );
and ( n74786 , n74553 , n74784 );
or ( n74787 , n74766 , n74785 , n74786 );
and ( n74788 , n74529 , n74787 );
and ( n74789 , n74527 , n74787 );
or ( n74790 , n74530 , n74788 , n74789 );
and ( n74791 , n74524 , n74790 );
and ( n74792 , n74522 , n74790 );
or ( n74793 , n74525 , n74791 , n74792 );
xor ( n74794 , n74488 , n74490 );
xor ( n74795 , n74794 , n74493 );
and ( n74796 , n74793 , n74795 );
xor ( n74797 , n74274 , n74289 );
xor ( n74798 , n74797 , n74357 );
xor ( n74799 , n74423 , n74433 );
xor ( n74800 , n74799 , n74436 );
and ( n74801 , n74798 , n74800 );
xor ( n74802 , n74445 , n74447 );
xor ( n74803 , n74802 , n74450 );
and ( n74804 , n74800 , n74803 );
and ( n74805 , n74798 , n74803 );
or ( n74806 , n74801 , n74804 , n74805 );
xor ( n74807 , n74194 , n74196 );
xor ( n74808 , n74807 , n74205 );
and ( n74809 , n74806 , n74808 );
xor ( n74810 , n74254 , n74360 );
xor ( n74811 , n74810 , n74439 );
and ( n74812 , n74808 , n74811 );
and ( n74813 , n74806 , n74811 );
or ( n74814 , n74809 , n74812 , n74813 );
xor ( n74815 , n74208 , n74442 );
xor ( n74816 , n74815 , n74461 );
and ( n74817 , n74814 , n74816 );
xor ( n74818 , n74474 , n74476 );
xor ( n74819 , n74818 , n74479 );
and ( n74820 , n74816 , n74819 );
and ( n74821 , n74814 , n74819 );
or ( n74822 , n74817 , n74820 , n74821 );
xor ( n74823 , n74464 , n74482 );
xor ( n74824 , n74823 , n74485 );
and ( n74825 , n74822 , n74824 );
xor ( n74826 , n74453 , n74455 );
xor ( n74827 , n74826 , n74458 );
xor ( n74828 , n74466 , n74468 );
xor ( n74829 , n74828 , n74471 );
and ( n74830 , n74827 , n74829 );
xor ( n74831 , n74425 , n74427 );
xor ( n74832 , n74831 , n74430 );
and ( n74833 , n65678 , n66917 );
not ( n74834 , n74833 );
buf ( n74835 , n74834 );
and ( n74836 , n55143 , n53357 );
and ( n74837 , n54942 , n53355 );
nor ( n74838 , n74836 , n74837 );
xnor ( n74839 , n74838 , n53060 );
and ( n74840 , n74835 , n74839 );
buf ( n74841 , n20817 );
and ( n74842 , n74839 , n74841 );
and ( n74843 , n74835 , n74841 );
or ( n74844 , n74840 , n74842 , n74843 );
and ( n74845 , n62593 , n69507 );
not ( n74846 , n74845 );
and ( n74847 , n69688 , n62868 );
not ( n74848 , n74847 );
and ( n74849 , n74846 , n74848 );
and ( n74850 , n74844 , n74849 );
and ( n74851 , n63024 , n69204 );
not ( n74852 , n74851 );
and ( n74853 , n69303 , n62998 );
not ( n74854 , n74853 );
and ( n74855 , n74852 , n74854 );
and ( n74856 , n74849 , n74855 );
and ( n74857 , n74844 , n74855 );
or ( n74858 , n74850 , n74856 , n74857 );
xor ( n74859 , n74565 , n74567 );
xor ( n74860 , n74579 , n74589 );
and ( n74861 , n74859 , n74860 );
xor ( n74862 , n74604 , n74614 );
and ( n74863 , n74860 , n74862 );
and ( n74864 , n74859 , n74862 );
or ( n74865 , n74861 , n74863 , n74864 );
and ( n74866 , n74858 , n74865 );
xor ( n74867 , n74617 , n74619 );
and ( n74868 , n63492 , n69204 );
not ( n74869 , n74868 );
and ( n74870 , n68307 , n64412 );
not ( n74871 , n74870 );
and ( n74872 , n74869 , n74871 );
and ( n74873 , n66980 , n65586 );
not ( n74874 , n74873 );
and ( n74875 , n74871 , n74874 );
and ( n74876 , n74869 , n74874 );
or ( n74877 , n74872 , n74875 , n74876 );
and ( n74878 , n62377 , n70108 );
not ( n74879 , n74878 );
and ( n74880 , n74877 , n74879 );
and ( n74881 , n74867 , n74880 );
and ( n74882 , n70256 , n62868 );
not ( n74883 , n74882 );
and ( n74884 , n69059 , n63766 );
not ( n74885 , n74884 );
and ( n74886 , n74883 , n74885 );
and ( n74887 , n62593 , n70108 );
not ( n74888 , n74887 );
and ( n74889 , n63987 , n68752 );
not ( n74890 , n74889 );
and ( n74891 , n74888 , n74890 );
and ( n74892 , n74886 , n74891 );
and ( n74893 , n74880 , n74892 );
and ( n74894 , n74867 , n74892 );
or ( n74895 , n74881 , n74893 , n74894 );
and ( n74896 , n74865 , n74895 );
and ( n74897 , n74858 , n74895 );
or ( n74898 , n74866 , n74896 , n74897 );
and ( n74899 , n74832 , n74898 );
xor ( n74900 , n74571 , n74573 );
xor ( n74901 , n74900 , n74576 );
xor ( n74902 , n74581 , n74583 );
xor ( n74903 , n74902 , n74586 );
and ( n74904 , n74901 , n74903 );
xor ( n74905 , n74596 , n74598 );
xor ( n74906 , n74905 , n74601 );
xor ( n74907 , n74606 , n74608 );
xor ( n74908 , n74907 , n74611 );
and ( n74909 , n74906 , n74908 );
and ( n74910 , n74904 , n74909 );
xor ( n74911 , n74846 , n74848 );
xor ( n74912 , n74852 , n74854 );
and ( n74913 , n74911 , n74912 );
xor ( n74914 , n74643 , n74645 );
and ( n74915 , n74912 , n74914 );
and ( n74916 , n74911 , n74914 );
or ( n74917 , n74913 , n74915 , n74916 );
and ( n74918 , n74909 , n74917 );
and ( n74919 , n74904 , n74917 );
or ( n74920 , n74910 , n74918 , n74919 );
and ( n74921 , n64221 , n68610 );
not ( n74922 , n74921 );
and ( n74923 , n65606 , n67013 );
not ( n74924 , n74923 );
and ( n74925 , n74922 , n74924 );
buf ( n74926 , n66415 );
not ( n74927 , n74926 );
and ( n74928 , n74924 , n74927 );
and ( n74929 , n74922 , n74927 );
or ( n74930 , n74925 , n74928 , n74929 );
and ( n74931 , n63024 , n69507 );
not ( n74932 , n74931 );
and ( n74933 , n69303 , n63679 );
not ( n74934 , n74933 );
and ( n74935 , n74932 , n74934 );
and ( n74936 , n74934 , n74833 );
and ( n74937 , n74932 , n74833 );
or ( n74938 , n74935 , n74936 , n74937 );
and ( n74939 , n74930 , n74938 );
and ( n74940 , n54942 , n53928 );
and ( n74941 , n54604 , n53926 );
nor ( n74942 , n74940 , n74941 );
xnor ( n74943 , n74942 , n53652 );
and ( n74944 , n55497 , n53357 );
and ( n74945 , n55143 , n53355 );
nor ( n74946 , n74944 , n74945 );
xnor ( n74947 , n74946 , n53060 );
and ( n74948 , n74943 , n74947 );
and ( n74949 , n74938 , n74948 );
and ( n74950 , n74930 , n74948 );
or ( n74951 , n74939 , n74949 , n74950 );
and ( n74952 , n53041 , n55851 );
and ( n74953 , n52790 , n55849 );
nor ( n74954 , n74952 , n74953 );
xnor ( n74955 , n74954 , n55506 );
and ( n74956 , n53639 , n55159 );
and ( n74957 , n53328 , n55157 );
nor ( n74958 , n74956 , n74957 );
xnor ( n74959 , n74958 , n54864 );
and ( n74960 , n74955 , n74959 );
and ( n74961 , n64548 , n67844 );
not ( n74962 , n74961 );
and ( n74963 , n67997 , n64811 );
not ( n74964 , n74963 );
and ( n74965 , n74962 , n74964 );
and ( n74966 , n74960 , n74965 );
and ( n74967 , n65177 , n67411 );
not ( n74968 , n74967 );
and ( n74969 , n67343 , n65210 );
not ( n74970 , n74969 );
and ( n74971 , n74968 , n74970 );
and ( n74972 , n74965 , n74971 );
and ( n74973 , n74960 , n74971 );
or ( n74974 , n74966 , n74972 , n74973 );
and ( n74975 , n74951 , n74974 );
and ( n74976 , n52082 , n57187 );
and ( n74977 , n51734 , n57184 );
nor ( n74978 , n74976 , n74977 );
xnor ( n74979 , n74978 , n56175 );
and ( n74980 , n52612 , n56503 );
and ( n74981 , n52332 , n56501 );
nor ( n74982 , n74980 , n74981 );
xnor ( n74983 , n74982 , n56178 );
and ( n74984 , n74979 , n74983 );
and ( n74985 , n54227 , n54535 );
and ( n74986 , n53922 , n54533 );
nor ( n74987 , n74985 , n74986 );
xnor ( n74988 , n74987 , n54237 );
and ( n74989 , n74983 , n74988 );
and ( n74990 , n74979 , n74988 );
or ( n74991 , n74984 , n74989 , n74990 );
and ( n74992 , n56915 , n52269 );
and ( n74993 , n56388 , n52267 );
nor ( n74994 , n74992 , n74993 );
xnor ( n74995 , n74994 , n52008 );
and ( n74996 , n74995 , n74701 );
xor ( n74997 , n45388 , n45512 );
buf ( n74998 , n74997 );
buf ( n74999 , n74998 );
buf ( n75000 , n74999 );
and ( n75001 , n74701 , n75000 );
and ( n75002 , n74995 , n75000 );
or ( n75003 , n74996 , n75001 , n75002 );
and ( n75004 , n74991 , n75003 );
and ( n75005 , n69688 , n62998 );
not ( n75006 , n75005 );
and ( n75007 , n66720 , n66005 );
not ( n75008 , n75007 );
and ( n75009 , n75006 , n75008 );
buf ( n75010 , n20818 );
and ( n75011 , n75008 , n75010 );
and ( n75012 , n75006 , n75010 );
or ( n75013 , n75009 , n75011 , n75012 );
and ( n75014 , n75003 , n75013 );
and ( n75015 , n74991 , n75013 );
or ( n75016 , n75004 , n75014 , n75015 );
and ( n75017 , n74974 , n75016 );
and ( n75018 , n74951 , n75016 );
or ( n75019 , n74975 , n75017 , n75018 );
and ( n75020 , n74920 , n75019 );
xor ( n75021 , n74651 , n74655 );
xor ( n75022 , n75021 , n74660 );
xor ( n75023 , n74671 , n74675 );
xor ( n75024 , n75023 , n74680 );
and ( n75025 , n75022 , n75024 );
xor ( n75026 , n74687 , n74691 );
xor ( n75027 , n75026 , n74696 );
and ( n75028 , n75024 , n75027 );
and ( n75029 , n75022 , n75027 );
or ( n75030 , n75025 , n75028 , n75029 );
buf ( n75031 , n74623 );
xor ( n75032 , n75031 , n74625 );
and ( n75033 , n75030 , n75032 );
xor ( n75034 , n74634 , n74635 );
xor ( n75035 , n75034 , n74637 );
and ( n75036 , n75032 , n75035 );
and ( n75037 , n75030 , n75035 );
or ( n75038 , n75033 , n75036 , n75037 );
and ( n75039 , n75019 , n75038 );
and ( n75040 , n74920 , n75038 );
or ( n75041 , n75020 , n75039 , n75040 );
and ( n75042 , n74898 , n75041 );
and ( n75043 , n74832 , n75041 );
or ( n75044 , n74899 , n75042 , n75043 );
xor ( n75045 , n74641 , n74646 );
xor ( n75046 , n75045 , n74663 );
xor ( n75047 , n74683 , n74699 );
xor ( n75048 , n75047 , n74713 );
and ( n75049 , n75046 , n75048 );
xor ( n75050 , n74721 , n74723 );
xor ( n75051 , n75050 , n74726 );
and ( n75052 , n75048 , n75051 );
and ( n75053 , n75046 , n75051 );
or ( n75054 , n75049 , n75052 , n75053 );
xor ( n75055 , n74541 , n74542 );
xor ( n75056 , n75055 , n74544 );
and ( n75057 , n75054 , n75056 );
xor ( n75058 , n74554 , n74555 );
xor ( n75059 , n75058 , n74557 );
and ( n75060 , n75056 , n75059 );
and ( n75061 , n75054 , n75059 );
or ( n75062 , n75057 , n75060 , n75061 );
xor ( n75063 , n74561 , n74568 );
xor ( n75064 , n75063 , n74590 );
xor ( n75065 , n74615 , n74620 );
xor ( n75066 , n75065 , n74627 );
and ( n75067 , n75064 , n75066 );
xor ( n75068 , n74640 , n74666 );
xor ( n75069 , n75068 , n74716 );
and ( n75070 , n75066 , n75069 );
and ( n75071 , n75064 , n75069 );
or ( n75072 , n75067 , n75070 , n75071 );
and ( n75073 , n75062 , n75072 );
xor ( n75074 , n74537 , n74538 );
xor ( n75075 , n75074 , n74547 );
and ( n75076 , n75072 , n75075 );
and ( n75077 , n75062 , n75075 );
or ( n75078 , n75073 , n75076 , n75077 );
and ( n75079 , n75044 , n75078 );
xor ( n75080 , n74560 , n74593 );
xor ( n75081 , n75080 , n74630 );
xor ( n75082 , n74719 , n74737 );
xor ( n75083 , n75082 , n74748 );
and ( n75084 , n75081 , n75083 );
xor ( n75085 , n74754 , n74756 );
xor ( n75086 , n75085 , n74759 );
and ( n75087 , n75083 , n75086 );
and ( n75088 , n75081 , n75086 );
or ( n75089 , n75084 , n75087 , n75088 );
and ( n75090 , n75078 , n75089 );
and ( n75091 , n75044 , n75089 );
or ( n75092 , n75079 , n75090 , n75091 );
and ( n75093 , n74829 , n75092 );
and ( n75094 , n74827 , n75092 );
or ( n75095 , n74830 , n75093 , n75094 );
xor ( n75096 , n74532 , n74534 );
xor ( n75097 , n75096 , n74550 );
xor ( n75098 , n74633 , n74751 );
xor ( n75099 , n75098 , n74762 );
and ( n75100 , n75097 , n75099 );
xor ( n75101 , n74776 , n74778 );
xor ( n75102 , n75101 , n74781 );
and ( n75103 , n75099 , n75102 );
and ( n75104 , n75097 , n75102 );
or ( n75105 , n75100 , n75103 , n75104 );
xor ( n75106 , n74553 , n74765 );
xor ( n75107 , n75106 , n74784 );
and ( n75108 , n75105 , n75107 );
xor ( n75109 , n74806 , n74808 );
xor ( n75110 , n75109 , n74811 );
and ( n75111 , n75107 , n75110 );
and ( n75112 , n75105 , n75110 );
or ( n75113 , n75108 , n75111 , n75112 );
and ( n75114 , n75095 , n75113 );
xor ( n75115 , n74527 , n74529 );
xor ( n75116 , n75115 , n74787 );
and ( n75117 , n75113 , n75116 );
and ( n75118 , n75095 , n75116 );
or ( n75119 , n75114 , n75117 , n75118 );
and ( n75120 , n74824 , n75119 );
and ( n75121 , n74822 , n75119 );
or ( n75122 , n74825 , n75120 , n75121 );
and ( n75123 , n74795 , n75122 );
and ( n75124 , n74793 , n75122 );
or ( n75125 , n74796 , n75123 , n75124 );
and ( n75126 , n74520 , n75125 );
xor ( n75127 , n74520 , n75125 );
xor ( n75128 , n74522 , n74524 );
xor ( n75129 , n75128 , n74790 );
xor ( n75130 , n74814 , n74816 );
xor ( n75131 , n75130 , n74819 );
xor ( n75132 , n74798 , n74800 );
xor ( n75133 , n75132 , n74803 );
xor ( n75134 , n74768 , n74770 );
xor ( n75135 , n75134 , n74773 );
xor ( n75136 , n74729 , n74731 );
xor ( n75137 , n75136 , n74734 );
xor ( n75138 , n74740 , n74742 );
xor ( n75139 , n75138 , n74745 );
and ( n75140 , n75137 , n75139 );
xor ( n75141 , n74844 , n74849 );
xor ( n75142 , n75141 , n74855 );
xor ( n75143 , n74703 , n74707 );
xor ( n75144 , n75143 , n74710 );
xor ( n75145 , n74835 , n74839 );
xor ( n75146 , n75145 , n74841 );
and ( n75147 , n75144 , n75146 );
xor ( n75148 , n74877 , n74879 );
and ( n75149 , n75146 , n75148 );
and ( n75150 , n75144 , n75148 );
or ( n75151 , n75147 , n75149 , n75150 );
and ( n75152 , n75142 , n75151 );
xor ( n75153 , n74886 , n74891 );
xor ( n75154 , n74901 , n74903 );
and ( n75155 , n75153 , n75154 );
xor ( n75156 , n74906 , n74908 );
and ( n75157 , n75154 , n75156 );
and ( n75158 , n75153 , n75156 );
or ( n75159 , n75155 , n75157 , n75158 );
and ( n75160 , n75151 , n75159 );
and ( n75161 , n75142 , n75159 );
or ( n75162 , n75152 , n75160 , n75161 );
and ( n75163 , n75139 , n75162 );
and ( n75164 , n75137 , n75162 );
or ( n75165 , n75140 , n75163 , n75164 );
and ( n75166 , n75135 , n75165 );
and ( n75167 , n67997 , n65210 );
not ( n75168 , n75167 );
and ( n75169 , n66980 , n66005 );
not ( n75170 , n75169 );
and ( n75171 , n75168 , n75170 );
and ( n75172 , n66720 , n66469 );
not ( n75173 , n75172 );
and ( n75174 , n75170 , n75173 );
and ( n75175 , n75168 , n75173 );
or ( n75176 , n75171 , n75174 , n75175 );
and ( n75177 , n65177 , n67844 );
not ( n75178 , n75177 );
and ( n75179 , n65678 , n67013 );
not ( n75180 , n75179 );
and ( n75181 , n75178 , n75180 );
and ( n75182 , n66415 , n66917 );
not ( n75183 , n75182 );
and ( n75184 , n75180 , n75183 );
and ( n75185 , n75178 , n75183 );
or ( n75186 , n75181 , n75184 , n75185 );
and ( n75187 , n75176 , n75186 );
and ( n75188 , n69688 , n63679 );
not ( n75189 , n75188 );
and ( n75190 , n69059 , n64412 );
not ( n75191 , n75190 );
and ( n75192 , n75189 , n75191 );
and ( n75193 , n68307 , n64811 );
not ( n75194 , n75193 );
and ( n75195 , n75191 , n75194 );
and ( n75196 , n75189 , n75194 );
or ( n75197 , n75192 , n75195 , n75196 );
and ( n75198 , n63492 , n69507 );
not ( n75199 , n75198 );
and ( n75200 , n64221 , n68752 );
not ( n75201 , n75200 );
and ( n75202 , n75199 , n75201 );
and ( n75203 , n64548 , n68610 );
not ( n75204 , n75203 );
and ( n75205 , n75201 , n75204 );
and ( n75206 , n75199 , n75204 );
or ( n75207 , n75202 , n75205 , n75206 );
and ( n75208 , n75197 , n75207 );
and ( n75209 , n75187 , n75208 );
xor ( n75210 , n74883 , n74885 );
xor ( n75211 , n74888 , n74890 );
and ( n75212 , n75210 , n75211 );
and ( n75213 , n75208 , n75212 );
and ( n75214 , n75187 , n75212 );
or ( n75215 , n75209 , n75213 , n75214 );
xor ( n75216 , n74922 , n74924 );
xor ( n75217 , n75216 , n74927 );
xor ( n75218 , n74869 , n74871 );
xor ( n75219 , n75218 , n74874 );
and ( n75220 , n75217 , n75219 );
xor ( n75221 , n74932 , n74934 );
xor ( n75222 , n75221 , n74833 );
and ( n75223 , n75219 , n75222 );
and ( n75224 , n75217 , n75222 );
or ( n75225 , n75220 , n75223 , n75224 );
xor ( n75226 , n74943 , n74947 );
xor ( n75227 , n74955 , n74959 );
and ( n75228 , n75226 , n75227 );
xor ( n75229 , n74962 , n74964 );
and ( n75230 , n75227 , n75229 );
and ( n75231 , n75226 , n75229 );
or ( n75232 , n75228 , n75230 , n75231 );
and ( n75233 , n75225 , n75232 );
xor ( n75234 , n74968 , n74970 );
and ( n75235 , n63987 , n69204 );
not ( n75236 , n75235 );
and ( n75237 , n69303 , n63766 );
not ( n75238 , n75237 );
and ( n75239 , n75236 , n75238 );
and ( n75240 , n75234 , n75239 );
and ( n75241 , n65606 , n67411 );
not ( n75242 , n75241 );
and ( n75243 , n67343 , n65586 );
not ( n75244 , n75243 );
and ( n75245 , n75242 , n75244 );
and ( n75246 , n75239 , n75245 );
and ( n75247 , n75234 , n75245 );
or ( n75248 , n75240 , n75246 , n75247 );
and ( n75249 , n75232 , n75248 );
and ( n75250 , n75225 , n75248 );
or ( n75251 , n75233 , n75249 , n75250 );
and ( n75252 , n75215 , n75251 );
and ( n75253 , n52332 , n57187 );
and ( n75254 , n52082 , n57184 );
nor ( n75255 , n75253 , n75254 );
xnor ( n75256 , n75255 , n56175 );
and ( n75257 , n52790 , n56503 );
and ( n75258 , n52612 , n56501 );
nor ( n75259 , n75257 , n75258 );
xnor ( n75260 , n75259 , n56178 );
and ( n75261 , n75256 , n75260 );
and ( n75262 , n53328 , n55851 );
and ( n75263 , n53041 , n55849 );
nor ( n75264 , n75262 , n75263 );
xnor ( n75265 , n75264 , n55506 );
and ( n75266 , n75260 , n75265 );
and ( n75267 , n75256 , n75265 );
or ( n75268 , n75261 , n75266 , n75267 );
and ( n75269 , n53922 , n55159 );
and ( n75270 , n53639 , n55157 );
nor ( n75271 , n75269 , n75270 );
xnor ( n75272 , n75271 , n54864 );
and ( n75273 , n55756 , n53357 );
and ( n75274 , n55497 , n53355 );
nor ( n75275 , n75273 , n75274 );
xnor ( n75276 , n75275 , n53060 );
and ( n75277 , n75272 , n75276 );
and ( n75278 , n56388 , n52799 );
and ( n75279 , n56255 , n52797 );
nor ( n75280 , n75278 , n75279 );
xnor ( n75281 , n75280 , n52538 );
and ( n75282 , n75276 , n75281 );
and ( n75283 , n75272 , n75281 );
or ( n75284 , n75277 , n75282 , n75283 );
and ( n75285 , n75268 , n75284 );
and ( n75286 , n57063 , n52269 );
and ( n75287 , n56915 , n52267 );
nor ( n75288 , n75286 , n75287 );
xnor ( n75289 , n75288 , n52008 );
and ( n75290 , n57063 , n52267 );
not ( n75291 , n75290 );
and ( n75292 , n75291 , n52008 );
and ( n75293 , n75289 , n75292 );
xor ( n75294 , n45389 , n45511 );
buf ( n75295 , n75294 );
buf ( n75296 , n75295 );
buf ( n75297 , n75296 );
and ( n75298 , n75292 , n75297 );
and ( n75299 , n75289 , n75297 );
or ( n75300 , n75293 , n75298 , n75299 );
and ( n75301 , n75284 , n75300 );
and ( n75302 , n75268 , n75300 );
or ( n75303 , n75285 , n75301 , n75302 );
xor ( n75304 , n74979 , n74983 );
xor ( n75305 , n75304 , n74988 );
xor ( n75306 , n74995 , n74701 );
xor ( n75307 , n75306 , n75000 );
and ( n75308 , n75305 , n75307 );
xor ( n75309 , n75006 , n75008 );
xor ( n75310 , n75309 , n75010 );
and ( n75311 , n75307 , n75310 );
and ( n75312 , n75305 , n75310 );
or ( n75313 , n75308 , n75311 , n75312 );
and ( n75314 , n75303 , n75313 );
xor ( n75315 , n74911 , n74912 );
xor ( n75316 , n75315 , n74914 );
and ( n75317 , n75313 , n75316 );
and ( n75318 , n75303 , n75316 );
or ( n75319 , n75314 , n75317 , n75318 );
and ( n75320 , n75251 , n75319 );
and ( n75321 , n75215 , n75319 );
or ( n75322 , n75252 , n75320 , n75321 );
xor ( n75323 , n74930 , n74938 );
xor ( n75324 , n75323 , n74948 );
xor ( n75325 , n74960 , n74965 );
xor ( n75326 , n75325 , n74971 );
and ( n75327 , n75324 , n75326 );
xor ( n75328 , n74991 , n75003 );
xor ( n75329 , n75328 , n75013 );
and ( n75330 , n75326 , n75329 );
and ( n75331 , n75324 , n75329 );
or ( n75332 , n75327 , n75330 , n75331 );
xor ( n75333 , n74859 , n74860 );
xor ( n75334 , n75333 , n74862 );
and ( n75335 , n75332 , n75334 );
xor ( n75336 , n74867 , n74880 );
xor ( n75337 , n75336 , n74892 );
and ( n75338 , n75334 , n75337 );
and ( n75339 , n75332 , n75337 );
or ( n75340 , n75335 , n75338 , n75339 );
and ( n75341 , n75322 , n75340 );
xor ( n75342 , n74904 , n74909 );
xor ( n75343 , n75342 , n74917 );
xor ( n75344 , n74951 , n74974 );
xor ( n75345 , n75344 , n75016 );
and ( n75346 , n75343 , n75345 );
xor ( n75347 , n75030 , n75032 );
xor ( n75348 , n75347 , n75035 );
and ( n75349 , n75345 , n75348 );
and ( n75350 , n75343 , n75348 );
or ( n75351 , n75346 , n75349 , n75350 );
and ( n75352 , n75340 , n75351 );
and ( n75353 , n75322 , n75351 );
or ( n75354 , n75341 , n75352 , n75353 );
and ( n75355 , n75165 , n75354 );
and ( n75356 , n75135 , n75354 );
or ( n75357 , n75166 , n75355 , n75356 );
and ( n75358 , n75133 , n75357 );
xor ( n75359 , n74858 , n74865 );
xor ( n75360 , n75359 , n74895 );
xor ( n75361 , n74920 , n75019 );
xor ( n75362 , n75361 , n75038 );
and ( n75363 , n75360 , n75362 );
xor ( n75364 , n75054 , n75056 );
xor ( n75365 , n75364 , n75059 );
and ( n75366 , n75362 , n75365 );
and ( n75367 , n75360 , n75365 );
or ( n75368 , n75363 , n75366 , n75367 );
xor ( n75369 , n74832 , n74898 );
xor ( n75370 , n75369 , n75041 );
and ( n75371 , n75368 , n75370 );
xor ( n75372 , n75062 , n75072 );
xor ( n75373 , n75372 , n75075 );
and ( n75374 , n75370 , n75373 );
and ( n75375 , n75368 , n75373 );
or ( n75376 , n75371 , n75374 , n75375 );
and ( n75377 , n75357 , n75376 );
and ( n75378 , n75133 , n75376 );
or ( n75379 , n75358 , n75377 , n75378 );
xor ( n75380 , n74827 , n74829 );
xor ( n75381 , n75380 , n75092 );
and ( n75382 , n75379 , n75381 );
xor ( n75383 , n75105 , n75107 );
xor ( n75384 , n75383 , n75110 );
and ( n75385 , n75381 , n75384 );
and ( n75386 , n75379 , n75384 );
or ( n75387 , n75382 , n75385 , n75386 );
and ( n75388 , n75131 , n75387 );
xor ( n75389 , n75095 , n75113 );
xor ( n75390 , n75389 , n75116 );
and ( n75391 , n75387 , n75390 );
and ( n75392 , n75131 , n75390 );
or ( n75393 , n75388 , n75391 , n75392 );
or ( n75394 , n75129 , n75393 );
xor ( n75395 , n74793 , n74795 );
xor ( n75396 , n75395 , n75122 );
and ( n75397 , n75394 , n75396 );
xor ( n75398 , n75394 , n75396 );
xor ( n75399 , n74822 , n74824 );
xor ( n75400 , n75399 , n75119 );
xnor ( n75401 , n75129 , n75393 );
and ( n75402 , n75400 , n75401 );
xor ( n75403 , n75400 , n75401 );
xor ( n75404 , n75131 , n75387 );
xor ( n75405 , n75404 , n75390 );
xor ( n75406 , n75044 , n75078 );
xor ( n75407 , n75406 , n75089 );
xor ( n75408 , n75097 , n75099 );
xor ( n75409 , n75408 , n75102 );
and ( n75410 , n75407 , n75409 );
xor ( n75411 , n75081 , n75083 );
xor ( n75412 , n75411 , n75086 );
xor ( n75413 , n75064 , n75066 );
xor ( n75414 , n75413 , n75069 );
xor ( n75415 , n75046 , n75048 );
xor ( n75416 , n75415 , n75051 );
xor ( n75417 , n75022 , n75024 );
xor ( n75418 , n75417 , n75027 );
and ( n75419 , n68307 , n65210 );
not ( n75420 , n75419 );
and ( n75421 , n67343 , n66005 );
not ( n75422 , n75421 );
and ( n75423 , n75420 , n75422 );
and ( n75424 , n66980 , n66469 );
not ( n75425 , n75424 );
and ( n75426 , n75422 , n75425 );
and ( n75427 , n75420 , n75425 );
or ( n75428 , n75423 , n75426 , n75427 );
and ( n75429 , n65177 , n68610 );
not ( n75430 , n75429 );
and ( n75431 , n65678 , n67411 );
not ( n75432 , n75431 );
and ( n75433 , n75430 , n75432 );
and ( n75434 , n66415 , n67013 );
not ( n75435 , n75434 );
and ( n75436 , n75432 , n75435 );
and ( n75437 , n75430 , n75435 );
or ( n75438 , n75433 , n75436 , n75437 );
and ( n75439 , n75428 , n75438 );
and ( n75440 , n63024 , n70108 );
not ( n75441 , n75440 );
and ( n75442 , n70256 , n62998 );
not ( n75443 , n75442 );
and ( n75444 , n75441 , n75443 );
and ( n75445 , n75439 , n75444 );
and ( n75446 , n56255 , n52799 );
and ( n75447 , n55756 , n52797 );
nor ( n75448 , n75446 , n75447 );
xnor ( n75449 , n75448 , n52538 );
and ( n75450 , n75444 , n75449 );
and ( n75451 , n75439 , n75449 );
or ( n75452 , n75445 , n75450 , n75451 );
and ( n75453 , n75418 , n75452 );
xor ( n75454 , n75176 , n75186 );
xor ( n75455 , n75197 , n75207 );
and ( n75456 , n75454 , n75455 );
xor ( n75457 , n75210 , n75211 );
and ( n75458 , n75455 , n75457 );
and ( n75459 , n75454 , n75457 );
or ( n75460 , n75456 , n75458 , n75459 );
and ( n75461 , n75452 , n75460 );
and ( n75462 , n75418 , n75460 );
or ( n75463 , n75453 , n75461 , n75462 );
and ( n75464 , n75416 , n75463 );
buf ( n75465 , n66720 );
not ( n75466 , n75465 );
buf ( n75467 , n75466 );
and ( n75468 , n55143 , n53928 );
and ( n75469 , n54942 , n53926 );
nor ( n75470 , n75468 , n75469 );
xnor ( n75471 , n75470 , n53652 );
and ( n75472 , n75467 , n75471 );
buf ( n75473 , n20819 );
and ( n75474 , n75471 , n75473 );
and ( n75475 , n75467 , n75473 );
or ( n75476 , n75472 , n75474 , n75475 );
and ( n75477 , n70256 , n63679 );
and ( n75478 , n69059 , n64811 );
not ( n75479 , n75478 );
and ( n75480 , n75477 , n75479 );
and ( n75481 , n63492 , n70108 );
and ( n75482 , n64548 , n68752 );
not ( n75483 , n75482 );
and ( n75484 , n75481 , n75483 );
and ( n75485 , n75480 , n75484 );
and ( n75486 , n75476 , n75485 );
not ( n75487 , n75477 );
buf ( n75488 , n75487 );
not ( n75489 , n75481 );
buf ( n75490 , n75489 );
and ( n75491 , n75488 , n75490 );
and ( n75492 , n75485 , n75491 );
and ( n75493 , n75476 , n75491 );
or ( n75494 , n75486 , n75492 , n75493 );
xor ( n75495 , n75168 , n75170 );
xor ( n75496 , n75495 , n75173 );
xor ( n75497 , n75178 , n75180 );
xor ( n75498 , n75497 , n75183 );
and ( n75499 , n75496 , n75498 );
xor ( n75500 , n75189 , n75191 );
xor ( n75501 , n75500 , n75194 );
xor ( n75502 , n75199 , n75201 );
xor ( n75503 , n75502 , n75204 );
and ( n75504 , n75501 , n75503 );
and ( n75505 , n75499 , n75504 );
xor ( n75506 , n75441 , n75443 );
xor ( n75507 , n75236 , n75238 );
and ( n75508 , n75506 , n75507 );
xor ( n75509 , n75242 , n75244 );
and ( n75510 , n75507 , n75509 );
and ( n75511 , n75506 , n75509 );
or ( n75512 , n75508 , n75510 , n75511 );
and ( n75513 , n75504 , n75512 );
and ( n75514 , n75499 , n75512 );
or ( n75515 , n75505 , n75513 , n75514 );
and ( n75516 , n75494 , n75515 );
and ( n75517 , n64221 , n69204 );
not ( n75518 , n75517 );
and ( n75519 , n65606 , n67844 );
not ( n75520 , n75519 );
and ( n75521 , n75518 , n75520 );
and ( n75522 , n75520 , n75465 );
and ( n75523 , n75518 , n75465 );
or ( n75524 , n75521 , n75522 , n75523 );
and ( n75525 , n55497 , n53928 );
and ( n75526 , n55143 , n53926 );
nor ( n75527 , n75525 , n75526 );
xnor ( n75528 , n75527 , n53652 );
buf ( n75529 , n20820 );
and ( n75530 , n75528 , n75529 );
and ( n75531 , n75524 , n75530 );
and ( n75532 , n63987 , n69507 );
not ( n75533 , n75532 );
and ( n75534 , n69688 , n63766 );
not ( n75535 , n75534 );
and ( n75536 , n75533 , n75535 );
and ( n75537 , n75530 , n75536 );
and ( n75538 , n75524 , n75536 );
or ( n75539 , n75531 , n75537 , n75538 );
and ( n75540 , n52612 , n57187 );
and ( n75541 , n52332 , n57184 );
nor ( n75542 , n75540 , n75541 );
xnor ( n75543 , n75542 , n56175 );
and ( n75544 , n53041 , n56503 );
and ( n75545 , n52790 , n56501 );
nor ( n75546 , n75544 , n75545 );
xnor ( n75547 , n75546 , n56178 );
and ( n75548 , n75543 , n75547 );
and ( n75549 , n53639 , n55851 );
and ( n75550 , n53328 , n55849 );
nor ( n75551 , n75549 , n75550 );
xnor ( n75552 , n75551 , n55506 );
and ( n75553 , n75547 , n75552 );
and ( n75554 , n75543 , n75552 );
or ( n75555 , n75548 , n75553 , n75554 );
and ( n75556 , n54227 , n55159 );
and ( n75557 , n53922 , n55157 );
nor ( n75558 , n75556 , n75557 );
xnor ( n75559 , n75558 , n54864 );
and ( n75560 , n56915 , n52799 );
and ( n75561 , n56388 , n52797 );
nor ( n75562 , n75560 , n75561 );
xnor ( n75563 , n75562 , n52538 );
and ( n75564 , n75559 , n75563 );
and ( n75565 , n75563 , n75290 );
and ( n75566 , n75559 , n75290 );
or ( n75567 , n75564 , n75565 , n75566 );
and ( n75568 , n75555 , n75567 );
xor ( n75569 , n45390 , n45510 );
buf ( n75570 , n75569 );
buf ( n75571 , n75570 );
buf ( n75572 , n75571 );
and ( n75573 , n69303 , n64412 );
not ( n75574 , n75573 );
and ( n75575 , n75572 , n75574 );
and ( n75576 , n67997 , n65586 );
not ( n75577 , n75576 );
and ( n75578 , n75574 , n75577 );
and ( n75579 , n75572 , n75577 );
or ( n75580 , n75575 , n75578 , n75579 );
and ( n75581 , n75567 , n75580 );
and ( n75582 , n75555 , n75580 );
or ( n75583 , n75568 , n75581 , n75582 );
and ( n75584 , n75539 , n75583 );
xor ( n75585 , n75256 , n75260 );
xor ( n75586 , n75585 , n75265 );
xor ( n75587 , n75272 , n75276 );
xor ( n75588 , n75587 , n75281 );
and ( n75589 , n75586 , n75588 );
xor ( n75590 , n75289 , n75292 );
xor ( n75591 , n75590 , n75297 );
and ( n75592 , n75588 , n75591 );
and ( n75593 , n75586 , n75591 );
or ( n75594 , n75589 , n75592 , n75593 );
and ( n75595 , n75583 , n75594 );
and ( n75596 , n75539 , n75594 );
or ( n75597 , n75584 , n75595 , n75596 );
and ( n75598 , n75515 , n75597 );
and ( n75599 , n75494 , n75597 );
or ( n75600 , n75516 , n75598 , n75599 );
and ( n75601 , n75463 , n75600 );
and ( n75602 , n75416 , n75600 );
or ( n75603 , n75464 , n75601 , n75602 );
and ( n75604 , n75414 , n75603 );
xor ( n75605 , n75217 , n75219 );
xor ( n75606 , n75605 , n75222 );
xor ( n75607 , n75226 , n75227 );
xor ( n75608 , n75607 , n75229 );
and ( n75609 , n75606 , n75608 );
xor ( n75610 , n75234 , n75239 );
xor ( n75611 , n75610 , n75245 );
and ( n75612 , n75608 , n75611 );
and ( n75613 , n75606 , n75611 );
or ( n75614 , n75609 , n75612 , n75613 );
xor ( n75615 , n75144 , n75146 );
xor ( n75616 , n75615 , n75148 );
and ( n75617 , n75614 , n75616 );
xor ( n75618 , n75153 , n75154 );
xor ( n75619 , n75618 , n75156 );
and ( n75620 , n75616 , n75619 );
and ( n75621 , n75614 , n75619 );
or ( n75622 , n75617 , n75620 , n75621 );
xor ( n75623 , n75187 , n75208 );
xor ( n75624 , n75623 , n75212 );
xor ( n75625 , n75225 , n75232 );
xor ( n75626 , n75625 , n75248 );
and ( n75627 , n75624 , n75626 );
xor ( n75628 , n75303 , n75313 );
xor ( n75629 , n75628 , n75316 );
and ( n75630 , n75626 , n75629 );
and ( n75631 , n75624 , n75629 );
or ( n75632 , n75627 , n75630 , n75631 );
and ( n75633 , n75622 , n75632 );
xor ( n75634 , n75142 , n75151 );
xor ( n75635 , n75634 , n75159 );
and ( n75636 , n75632 , n75635 );
and ( n75637 , n75622 , n75635 );
or ( n75638 , n75633 , n75636 , n75637 );
and ( n75639 , n75603 , n75638 );
and ( n75640 , n75414 , n75638 );
or ( n75641 , n75604 , n75639 , n75640 );
and ( n75642 , n75412 , n75641 );
xor ( n75643 , n75215 , n75251 );
xor ( n75644 , n75643 , n75319 );
xor ( n75645 , n75332 , n75334 );
xor ( n75646 , n75645 , n75337 );
and ( n75647 , n75644 , n75646 );
xor ( n75648 , n75343 , n75345 );
xor ( n75649 , n75648 , n75348 );
and ( n75650 , n75646 , n75649 );
and ( n75651 , n75644 , n75649 );
or ( n75652 , n75647 , n75650 , n75651 );
xor ( n75653 , n75137 , n75139 );
xor ( n75654 , n75653 , n75162 );
and ( n75655 , n75652 , n75654 );
xor ( n75656 , n75322 , n75340 );
xor ( n75657 , n75656 , n75351 );
and ( n75658 , n75654 , n75657 );
and ( n75659 , n75652 , n75657 );
or ( n75660 , n75655 , n75658 , n75659 );
and ( n75661 , n75641 , n75660 );
and ( n75662 , n75412 , n75660 );
or ( n75663 , n75642 , n75661 , n75662 );
and ( n75664 , n75409 , n75663 );
and ( n75665 , n75407 , n75663 );
or ( n75666 , n75410 , n75664 , n75665 );
xor ( n75667 , n75379 , n75381 );
xor ( n75668 , n75667 , n75384 );
and ( n75669 , n75666 , n75668 );
xor ( n75670 , n75133 , n75357 );
xor ( n75671 , n75670 , n75376 );
xor ( n75672 , n75135 , n75165 );
xor ( n75673 , n75672 , n75354 );
xor ( n75674 , n75368 , n75370 );
xor ( n75675 , n75674 , n75373 );
and ( n75676 , n75673 , n75675 );
xor ( n75677 , n75360 , n75362 );
xor ( n75678 , n75677 , n75365 );
xor ( n75679 , n75324 , n75326 );
xor ( n75680 , n75679 , n75329 );
xor ( n75681 , n75268 , n75284 );
xor ( n75682 , n75681 , n75300 );
xor ( n75683 , n75305 , n75307 );
xor ( n75684 , n75683 , n75310 );
and ( n75685 , n75682 , n75684 );
xor ( n75686 , n75439 , n75444 );
xor ( n75687 , n75686 , n75449 );
and ( n75688 , n75684 , n75687 );
and ( n75689 , n75682 , n75687 );
or ( n75690 , n75685 , n75688 , n75689 );
and ( n75691 , n75680 , n75690 );
and ( n75692 , n54604 , n54535 );
and ( n75693 , n54227 , n54533 );
nor ( n75694 , n75692 , n75693 );
xnor ( n75695 , n75694 , n54237 );
xor ( n75696 , n75467 , n75471 );
xor ( n75697 , n75696 , n75473 );
and ( n75698 , n75695 , n75697 );
and ( n75699 , n64221 , n69507 );
not ( n75700 , n75699 );
and ( n75701 , n65177 , n68752 );
not ( n75702 , n75701 );
and ( n75703 , n75700 , n75702 );
and ( n75704 , n66415 , n67411 );
not ( n75705 , n75704 );
and ( n75706 , n75702 , n75705 );
and ( n75707 , n75700 , n75705 );
or ( n75708 , n75703 , n75706 , n75707 );
xor ( n75709 , n75430 , n75432 );
xor ( n75710 , n75709 , n75435 );
or ( n75711 , n75708 , n75710 );
and ( n75712 , n69688 , n64412 );
not ( n75713 , n75712 );
and ( n75714 , n69059 , n65210 );
not ( n75715 , n75714 );
and ( n75716 , n75713 , n75715 );
and ( n75717 , n67343 , n66469 );
not ( n75718 , n75717 );
and ( n75719 , n75715 , n75718 );
and ( n75720 , n75713 , n75718 );
or ( n75721 , n75716 , n75719 , n75720 );
xor ( n75722 , n75420 , n75422 );
xor ( n75723 , n75722 , n75425 );
or ( n75724 , n75721 , n75723 );
and ( n75725 , n75711 , n75724 );
and ( n75726 , n75698 , n75725 );
xor ( n75727 , n75428 , n75438 );
xor ( n75728 , n75480 , n75484 );
and ( n75729 , n75727 , n75728 );
xor ( n75730 , n75488 , n75490 );
and ( n75731 , n75728 , n75730 );
and ( n75732 , n75727 , n75730 );
or ( n75733 , n75729 , n75731 , n75732 );
and ( n75734 , n75725 , n75733 );
and ( n75735 , n75698 , n75733 );
or ( n75736 , n75726 , n75734 , n75735 );
and ( n75737 , n75690 , n75736 );
and ( n75738 , n75680 , n75736 );
or ( n75739 , n75691 , n75737 , n75738 );
xor ( n75740 , n75496 , n75498 );
xor ( n75741 , n75501 , n75503 );
and ( n75742 , n75740 , n75741 );
and ( n75743 , n65678 , n67844 );
not ( n75744 , n75743 );
and ( n75745 , n67997 , n66005 );
not ( n75746 , n75745 );
and ( n75747 , n75744 , n75746 );
and ( n75748 , n54942 , n54535 );
and ( n75749 , n54604 , n54533 );
nor ( n75750 , n75748 , n75749 );
xnor ( n75751 , n75750 , n54237 );
and ( n75752 , n75747 , n75751 );
and ( n75753 , n56255 , n53357 );
and ( n75754 , n55756 , n53355 );
nor ( n75755 , n75753 , n75754 );
xnor ( n75756 , n75755 , n53060 );
and ( n75757 , n75751 , n75756 );
and ( n75758 , n75747 , n75756 );
or ( n75759 , n75752 , n75757 , n75758 );
and ( n75760 , n75741 , n75759 );
and ( n75761 , n75740 , n75759 );
or ( n75762 , n75742 , n75760 , n75761 );
xor ( n75763 , n75477 , n75479 );
xor ( n75764 , n75481 , n75483 );
and ( n75765 , n75763 , n75764 );
xor ( n75766 , n75518 , n75520 );
xor ( n75767 , n75766 , n75465 );
xor ( n75768 , n75528 , n75529 );
and ( n75769 , n75767 , n75768 );
xor ( n75770 , n75533 , n75535 );
and ( n75771 , n75768 , n75770 );
and ( n75772 , n75767 , n75770 );
or ( n75773 , n75769 , n75771 , n75772 );
and ( n75774 , n75765 , n75773 );
and ( n75775 , n56388 , n53357 );
and ( n75776 , n56255 , n53355 );
nor ( n75777 , n75775 , n75776 );
xnor ( n75778 , n75777 , n53060 );
and ( n75779 , n57063 , n52797 );
not ( n75780 , n75779 );
and ( n75781 , n75780 , n52538 );
and ( n75782 , n75778 , n75781 );
and ( n75783 , n65606 , n68610 );
not ( n75784 , n75783 );
and ( n75785 , n68307 , n65586 );
not ( n75786 , n75785 );
and ( n75787 , n75784 , n75786 );
and ( n75788 , n75782 , n75787 );
and ( n75789 , n66720 , n67013 );
not ( n75790 , n75789 );
and ( n75791 , n66980 , n66917 );
not ( n75792 , n75791 );
and ( n75793 , n75790 , n75792 );
and ( n75794 , n75787 , n75793 );
and ( n75795 , n75782 , n75793 );
or ( n75796 , n75788 , n75794 , n75795 );
and ( n75797 , n75773 , n75796 );
and ( n75798 , n75765 , n75796 );
or ( n75799 , n75774 , n75797 , n75798 );
and ( n75800 , n75762 , n75799 );
and ( n75801 , n52790 , n57187 );
and ( n75802 , n52612 , n57184 );
nor ( n75803 , n75801 , n75802 );
xnor ( n75804 , n75803 , n56175 );
and ( n75805 , n53328 , n56503 );
and ( n75806 , n53041 , n56501 );
nor ( n75807 , n75805 , n75806 );
xnor ( n75808 , n75807 , n56178 );
and ( n75809 , n75804 , n75808 );
and ( n75810 , n53922 , n55851 );
and ( n75811 , n53639 , n55849 );
nor ( n75812 , n75810 , n75811 );
xnor ( n75813 , n75812 , n55506 );
and ( n75814 , n75808 , n75813 );
and ( n75815 , n75804 , n75813 );
or ( n75816 , n75809 , n75814 , n75815 );
and ( n75817 , n54604 , n55159 );
and ( n75818 , n54227 , n55157 );
nor ( n75819 , n75817 , n75818 );
xnor ( n75820 , n75819 , n54864 );
and ( n75821 , n55143 , n54535 );
and ( n75822 , n54942 , n54533 );
nor ( n75823 , n75821 , n75822 );
xnor ( n75824 , n75823 , n54237 );
and ( n75825 , n75820 , n75824 );
and ( n75826 , n55756 , n53928 );
and ( n75827 , n55497 , n53926 );
nor ( n75828 , n75826 , n75827 );
xnor ( n75829 , n75828 , n53652 );
and ( n75830 , n75824 , n75829 );
and ( n75831 , n75820 , n75829 );
or ( n75832 , n75825 , n75830 , n75831 );
and ( n75833 , n75816 , n75832 );
and ( n75834 , n57063 , n52799 );
and ( n75835 , n56915 , n52797 );
nor ( n75836 , n75834 , n75835 );
xnor ( n75837 , n75836 , n52538 );
xor ( n75838 , n45391 , n45509 );
buf ( n75839 , n75838 );
buf ( n75840 , n75839 );
buf ( n75841 , n75840 );
and ( n75842 , n75837 , n75841 );
and ( n75843 , n70256 , n63766 );
not ( n75844 , n75843 );
and ( n75845 , n75841 , n75844 );
and ( n75846 , n75837 , n75844 );
or ( n75847 , n75842 , n75845 , n75846 );
and ( n75848 , n75832 , n75847 );
and ( n75849 , n75816 , n75847 );
or ( n75850 , n75833 , n75848 , n75849 );
xor ( n75851 , n75543 , n75547 );
xor ( n75852 , n75851 , n75552 );
xor ( n75853 , n75559 , n75563 );
xor ( n75854 , n75853 , n75290 );
and ( n75855 , n75852 , n75854 );
xor ( n75856 , n75572 , n75574 );
xor ( n75857 , n75856 , n75577 );
and ( n75858 , n75854 , n75857 );
and ( n75859 , n75852 , n75857 );
or ( n75860 , n75855 , n75858 , n75859 );
and ( n75861 , n75850 , n75860 );
xor ( n75862 , n75506 , n75507 );
xor ( n75863 , n75862 , n75509 );
and ( n75864 , n75860 , n75863 );
and ( n75865 , n75850 , n75863 );
or ( n75866 , n75861 , n75864 , n75865 );
and ( n75867 , n75799 , n75866 );
and ( n75868 , n75762 , n75866 );
or ( n75869 , n75800 , n75867 , n75868 );
xor ( n75870 , n75524 , n75530 );
xor ( n75871 , n75870 , n75536 );
xor ( n75872 , n75555 , n75567 );
xor ( n75873 , n75872 , n75580 );
and ( n75874 , n75871 , n75873 );
xor ( n75875 , n75586 , n75588 );
xor ( n75876 , n75875 , n75591 );
and ( n75877 , n75873 , n75876 );
and ( n75878 , n75871 , n75876 );
or ( n75879 , n75874 , n75877 , n75878 );
xor ( n75880 , n75454 , n75455 );
xor ( n75881 , n75880 , n75457 );
and ( n75882 , n75879 , n75881 );
xor ( n75883 , n75476 , n75485 );
xor ( n75884 , n75883 , n75491 );
and ( n75885 , n75881 , n75884 );
and ( n75886 , n75879 , n75884 );
or ( n75887 , n75882 , n75885 , n75886 );
and ( n75888 , n75869 , n75887 );
xor ( n75889 , n75499 , n75504 );
xor ( n75890 , n75889 , n75512 );
xor ( n75891 , n75539 , n75583 );
xor ( n75892 , n75891 , n75594 );
and ( n75893 , n75890 , n75892 );
xor ( n75894 , n75606 , n75608 );
xor ( n75895 , n75894 , n75611 );
and ( n75896 , n75892 , n75895 );
and ( n75897 , n75890 , n75895 );
or ( n75898 , n75893 , n75896 , n75897 );
and ( n75899 , n75887 , n75898 );
and ( n75900 , n75869 , n75898 );
or ( n75901 , n75888 , n75899 , n75900 );
and ( n75902 , n75739 , n75901 );
xor ( n75903 , n75418 , n75452 );
xor ( n75904 , n75903 , n75460 );
xor ( n75905 , n75494 , n75515 );
xor ( n75906 , n75905 , n75597 );
and ( n75907 , n75904 , n75906 );
xor ( n75908 , n75614 , n75616 );
xor ( n75909 , n75908 , n75619 );
and ( n75910 , n75906 , n75909 );
and ( n75911 , n75904 , n75909 );
or ( n75912 , n75907 , n75910 , n75911 );
and ( n75913 , n75901 , n75912 );
and ( n75914 , n75739 , n75912 );
or ( n75915 , n75902 , n75913 , n75914 );
and ( n75916 , n75678 , n75915 );
xor ( n75917 , n75416 , n75463 );
xor ( n75918 , n75917 , n75600 );
xor ( n75919 , n75622 , n75632 );
xor ( n75920 , n75919 , n75635 );
and ( n75921 , n75918 , n75920 );
xor ( n75922 , n75644 , n75646 );
xor ( n75923 , n75922 , n75649 );
and ( n75924 , n75920 , n75923 );
and ( n75925 , n75918 , n75923 );
or ( n75926 , n75921 , n75924 , n75925 );
and ( n75927 , n75915 , n75926 );
and ( n75928 , n75678 , n75926 );
or ( n75929 , n75916 , n75927 , n75928 );
and ( n75930 , n75675 , n75929 );
and ( n75931 , n75673 , n75929 );
or ( n75932 , n75676 , n75930 , n75931 );
and ( n75933 , n75671 , n75932 );
xor ( n75934 , n75407 , n75409 );
xor ( n75935 , n75934 , n75663 );
and ( n75936 , n75932 , n75935 );
and ( n75937 , n75671 , n75935 );
or ( n75938 , n75933 , n75936 , n75937 );
and ( n75939 , n75668 , n75938 );
and ( n75940 , n75666 , n75938 );
or ( n75941 , n75669 , n75939 , n75940 );
and ( n75942 , n75405 , n75941 );
xor ( n75943 , n75405 , n75941 );
xor ( n75944 , n75666 , n75668 );
xor ( n75945 , n75944 , n75938 );
xor ( n75946 , n75412 , n75641 );
xor ( n75947 , n75946 , n75660 );
xor ( n75948 , n75414 , n75603 );
xor ( n75949 , n75948 , n75638 );
xor ( n75950 , n75652 , n75654 );
xor ( n75951 , n75950 , n75657 );
and ( n75952 , n75949 , n75951 );
xor ( n75953 , n75624 , n75626 );
xor ( n75954 , n75953 , n75629 );
xor ( n75955 , n75695 , n75697 );
xor ( n75956 , n75711 , n75724 );
and ( n75957 , n75955 , n75956 );
xnor ( n75958 , n75708 , n75710 );
xnor ( n75959 , n75721 , n75723 );
and ( n75960 , n75958 , n75959 );
and ( n75961 , n75956 , n75960 );
and ( n75962 , n75955 , n75960 );
or ( n75963 , n75957 , n75961 , n75962 );
xor ( n75964 , n75747 , n75751 );
xor ( n75965 , n75964 , n75756 );
xor ( n75966 , n75763 , n75764 );
and ( n75967 , n75965 , n75966 );
and ( n75968 , n66720 , n67411 );
not ( n75969 , n75968 );
buf ( n75970 , n75969 );
and ( n75971 , n63987 , n70108 );
not ( n75972 , n75971 );
and ( n75973 , n75970 , n75972 );
and ( n75974 , n64548 , n69204 );
not ( n75975 , n75974 );
and ( n75976 , n75972 , n75975 );
and ( n75977 , n75970 , n75975 );
or ( n75978 , n75973 , n75976 , n75977 );
and ( n75979 , n75966 , n75978 );
and ( n75980 , n75965 , n75978 );
or ( n75981 , n75967 , n75979 , n75980 );
and ( n75982 , n69303 , n65210 );
not ( n75983 , n75982 );
and ( n75984 , n68307 , n66005 );
not ( n75985 , n75984 );
and ( n75986 , n75983 , n75985 );
and ( n75987 , n67997 , n66469 );
not ( n75988 , n75987 );
and ( n75989 , n75985 , n75988 );
and ( n75990 , n75983 , n75988 );
or ( n75991 , n75986 , n75989 , n75990 );
and ( n75992 , n65177 , n69204 );
not ( n75993 , n75992 );
and ( n75994 , n65678 , n68610 );
not ( n75995 , n75994 );
and ( n75996 , n75993 , n75995 );
and ( n75997 , n66415 , n67844 );
not ( n75998 , n75997 );
and ( n75999 , n75995 , n75998 );
and ( n76000 , n75993 , n75998 );
or ( n76001 , n75996 , n75999 , n76000 );
and ( n76002 , n75991 , n76001 );
xor ( n76003 , n75713 , n75715 );
xor ( n76004 , n76003 , n75718 );
xor ( n76005 , n75700 , n75702 );
xor ( n76006 , n76005 , n75705 );
and ( n76007 , n76004 , n76006 );
and ( n76008 , n76002 , n76007 );
and ( n76009 , n69303 , n64811 );
not ( n76010 , n76009 );
buf ( n76011 , n20821 );
and ( n76012 , n76010 , n76011 );
xor ( n76013 , n75778 , n75781 );
and ( n76014 , n76011 , n76013 );
and ( n76015 , n76010 , n76013 );
or ( n76016 , n76012 , n76014 , n76015 );
and ( n76017 , n76007 , n76016 );
and ( n76018 , n76002 , n76016 );
or ( n76019 , n76008 , n76017 , n76018 );
and ( n76020 , n75981 , n76019 );
xor ( n76021 , n75784 , n75786 );
xor ( n76022 , n75744 , n75746 );
and ( n76023 , n76021 , n76022 );
xor ( n76024 , n75790 , n75792 );
and ( n76025 , n76022 , n76024 );
and ( n76026 , n76021 , n76024 );
or ( n76027 , n76023 , n76025 , n76026 );
and ( n76028 , n64221 , n70108 );
not ( n76029 , n76028 );
and ( n76030 , n69688 , n64811 );
not ( n76031 , n76030 );
or ( n76032 , n76029 , n76031 );
and ( n76033 , n53041 , n57187 );
and ( n76034 , n52790 , n57184 );
nor ( n76035 , n76033 , n76034 );
xnor ( n76036 , n76035 , n56175 );
and ( n76037 , n53639 , n56503 );
and ( n76038 , n53328 , n56501 );
nor ( n76039 , n76037 , n76038 );
xnor ( n76040 , n76039 , n56178 );
and ( n76041 , n76036 , n76040 );
and ( n76042 , n76032 , n76041 );
and ( n76043 , n65606 , n68752 );
not ( n76044 , n76043 );
and ( n76045 , n69059 , n65586 );
not ( n76046 , n76045 );
and ( n76047 , n76044 , n76046 );
and ( n76048 , n76041 , n76047 );
and ( n76049 , n76032 , n76047 );
or ( n76050 , n76042 , n76048 , n76049 );
and ( n76051 , n76027 , n76050 );
and ( n76052 , n54227 , n55851 );
and ( n76053 , n53922 , n55849 );
nor ( n76054 , n76052 , n76053 );
xnor ( n76055 , n76054 , n55506 );
and ( n76056 , n54942 , n55159 );
and ( n76057 , n54604 , n55157 );
nor ( n76058 , n76056 , n76057 );
xnor ( n76059 , n76058 , n54864 );
and ( n76060 , n76055 , n76059 );
and ( n76061 , n55497 , n54535 );
and ( n76062 , n55143 , n54533 );
nor ( n76063 , n76061 , n76062 );
xnor ( n76064 , n76063 , n54237 );
and ( n76065 , n76059 , n76064 );
and ( n76066 , n76055 , n76064 );
or ( n76067 , n76060 , n76065 , n76066 );
and ( n76068 , n56255 , n53928 );
and ( n76069 , n55756 , n53926 );
nor ( n76070 , n76068 , n76069 );
xnor ( n76071 , n76070 , n53652 );
and ( n76072 , n56915 , n53357 );
and ( n76073 , n56388 , n53355 );
nor ( n76074 , n76072 , n76073 );
xnor ( n76075 , n76074 , n53060 );
and ( n76076 , n76071 , n76075 );
and ( n76077 , n76075 , n75779 );
and ( n76078 , n76071 , n75779 );
or ( n76079 , n76076 , n76077 , n76078 );
and ( n76080 , n76067 , n76079 );
xor ( n76081 , n45394 , n45507 );
buf ( n76082 , n76081 );
buf ( n76083 , n76082 );
buf ( n76084 , n76083 );
and ( n76085 , n70256 , n64412 );
not ( n76086 , n76085 );
and ( n76087 , n76084 , n76086 );
and ( n76088 , n67343 , n66917 );
not ( n76089 , n76088 );
and ( n76090 , n76086 , n76089 );
and ( n76091 , n76084 , n76089 );
or ( n76092 , n76087 , n76090 , n76091 );
and ( n76093 , n76079 , n76092 );
and ( n76094 , n76067 , n76092 );
or ( n76095 , n76080 , n76093 , n76094 );
and ( n76096 , n76050 , n76095 );
and ( n76097 , n76027 , n76095 );
or ( n76098 , n76051 , n76096 , n76097 );
and ( n76099 , n76019 , n76098 );
and ( n76100 , n75981 , n76098 );
or ( n76101 , n76020 , n76099 , n76100 );
and ( n76102 , n75963 , n76101 );
xor ( n76103 , n75804 , n75808 );
xor ( n76104 , n76103 , n75813 );
xor ( n76105 , n75820 , n75824 );
xor ( n76106 , n76105 , n75829 );
and ( n76107 , n76104 , n76106 );
xor ( n76108 , n75837 , n75841 );
xor ( n76109 , n76108 , n75844 );
and ( n76110 , n76106 , n76109 );
and ( n76111 , n76104 , n76109 );
or ( n76112 , n76107 , n76110 , n76111 );
xor ( n76113 , n75767 , n75768 );
xor ( n76114 , n76113 , n75770 );
and ( n76115 , n76112 , n76114 );
xor ( n76116 , n75782 , n75787 );
xor ( n76117 , n76116 , n75793 );
and ( n76118 , n76114 , n76117 );
and ( n76119 , n76112 , n76117 );
or ( n76120 , n76115 , n76118 , n76119 );
xor ( n76121 , n75727 , n75728 );
xor ( n76122 , n76121 , n75730 );
and ( n76123 , n76120 , n76122 );
xor ( n76124 , n75740 , n75741 );
xor ( n76125 , n76124 , n75759 );
and ( n76126 , n76122 , n76125 );
and ( n76127 , n76120 , n76125 );
or ( n76128 , n76123 , n76126 , n76127 );
and ( n76129 , n76101 , n76128 );
and ( n76130 , n75963 , n76128 );
or ( n76131 , n76102 , n76129 , n76130 );
and ( n76132 , n75954 , n76131 );
xor ( n76133 , n75765 , n75773 );
xor ( n76134 , n76133 , n75796 );
xor ( n76135 , n75850 , n75860 );
xor ( n76136 , n76135 , n75863 );
and ( n76137 , n76134 , n76136 );
xor ( n76138 , n75871 , n75873 );
xor ( n76139 , n76138 , n75876 );
and ( n76140 , n76136 , n76139 );
and ( n76141 , n76134 , n76139 );
or ( n76142 , n76137 , n76140 , n76141 );
xor ( n76143 , n75682 , n75684 );
xor ( n76144 , n76143 , n75687 );
and ( n76145 , n76142 , n76144 );
xor ( n76146 , n75698 , n75725 );
xor ( n76147 , n76146 , n75733 );
and ( n76148 , n76144 , n76147 );
and ( n76149 , n76142 , n76147 );
or ( n76150 , n76145 , n76148 , n76149 );
and ( n76151 , n76131 , n76150 );
and ( n76152 , n75954 , n76150 );
or ( n76153 , n76132 , n76151 , n76152 );
xor ( n76154 , n75762 , n75799 );
xor ( n76155 , n76154 , n75866 );
xor ( n76156 , n75879 , n75881 );
xor ( n76157 , n76156 , n75884 );
and ( n76158 , n76155 , n76157 );
xor ( n76159 , n75890 , n75892 );
xor ( n76160 , n76159 , n75895 );
and ( n76161 , n76157 , n76160 );
and ( n76162 , n76155 , n76160 );
or ( n76163 , n76158 , n76161 , n76162 );
xor ( n76164 , n75680 , n75690 );
xor ( n76165 , n76164 , n75736 );
and ( n76166 , n76163 , n76165 );
xor ( n76167 , n75869 , n75887 );
xor ( n76168 , n76167 , n75898 );
and ( n76169 , n76165 , n76168 );
and ( n76170 , n76163 , n76168 );
or ( n76171 , n76166 , n76169 , n76170 );
and ( n76172 , n76153 , n76171 );
xor ( n76173 , n75739 , n75901 );
xor ( n76174 , n76173 , n75912 );
and ( n76175 , n76171 , n76174 );
and ( n76176 , n76153 , n76174 );
or ( n76177 , n76172 , n76175 , n76176 );
and ( n76178 , n75951 , n76177 );
and ( n76179 , n75949 , n76177 );
or ( n76180 , n75952 , n76178 , n76179 );
and ( n76181 , n75947 , n76180 );
xor ( n76182 , n75673 , n75675 );
xor ( n76183 , n76182 , n75929 );
and ( n76184 , n76180 , n76183 );
and ( n76185 , n75947 , n76183 );
or ( n76186 , n76181 , n76184 , n76185 );
xor ( n76187 , n75671 , n75932 );
xor ( n76188 , n76187 , n75935 );
and ( n76189 , n76186 , n76188 );
xor ( n76190 , n75678 , n75915 );
xor ( n76191 , n76190 , n75926 );
xor ( n76192 , n75918 , n75920 );
xor ( n76193 , n76192 , n75923 );
xor ( n76194 , n75904 , n75906 );
xor ( n76195 , n76194 , n75909 );
xor ( n76196 , n75816 , n75832 );
xor ( n76197 , n76196 , n75847 );
xor ( n76198 , n75852 , n75854 );
xor ( n76199 , n76198 , n75857 );
and ( n76200 , n76197 , n76199 );
xor ( n76201 , n75958 , n75959 );
and ( n76202 , n76199 , n76201 );
and ( n76203 , n76197 , n76201 );
or ( n76204 , n76200 , n76202 , n76203 );
and ( n76205 , n64548 , n69507 );
not ( n76206 , n76205 );
and ( n76207 , n76206 , n75968 );
buf ( n76208 , n66980 );
not ( n76209 , n76208 );
and ( n76210 , n75968 , n76209 );
and ( n76211 , n76206 , n76209 );
or ( n76212 , n76207 , n76210 , n76211 );
xor ( n76213 , n75970 , n75972 );
xor ( n76214 , n76213 , n75975 );
or ( n76215 , n76212 , n76214 );
xor ( n76216 , n75991 , n76001 );
xor ( n76217 , n76004 , n76006 );
and ( n76218 , n76216 , n76217 );
xor ( n76219 , n75983 , n75985 );
xor ( n76220 , n76219 , n75988 );
xor ( n76221 , n75993 , n75995 );
xor ( n76222 , n76221 , n75998 );
and ( n76223 , n76220 , n76222 );
and ( n76224 , n76217 , n76223 );
and ( n76225 , n76216 , n76223 );
or ( n76226 , n76218 , n76224 , n76225 );
and ( n76227 , n76215 , n76226 );
buf ( n76228 , n20822 );
xor ( n76229 , n76206 , n75968 );
xor ( n76230 , n76229 , n76209 );
and ( n76231 , n76228 , n76230 );
xnor ( n76232 , n76029 , n76031 );
and ( n76233 , n76230 , n76232 );
and ( n76234 , n76228 , n76232 );
or ( n76235 , n76231 , n76233 , n76234 );
xor ( n76236 , n76036 , n76040 );
xor ( n76237 , n76044 , n76046 );
and ( n76238 , n76236 , n76237 );
and ( n76239 , n66415 , n68610 );
not ( n76240 , n76239 );
and ( n76241 , n66720 , n67844 );
not ( n76242 , n76241 );
and ( n76243 , n76240 , n76242 );
and ( n76244 , n66980 , n67411 );
not ( n76245 , n76244 );
and ( n76246 , n76242 , n76245 );
and ( n76247 , n76240 , n76245 );
or ( n76248 , n76243 , n76246 , n76247 );
and ( n76249 , n76237 , n76248 );
and ( n76250 , n76236 , n76248 );
or ( n76251 , n76238 , n76249 , n76250 );
and ( n76252 , n76235 , n76251 );
and ( n76253 , n64548 , n70108 );
not ( n76254 , n76253 );
and ( n76255 , n70256 , n64811 );
not ( n76256 , n76255 );
and ( n76257 , n76254 , n76256 );
and ( n76258 , n65606 , n69204 );
not ( n76259 , n76258 );
and ( n76260 , n69303 , n65586 );
not ( n76261 , n76260 );
and ( n76262 , n76259 , n76261 );
and ( n76263 , n76257 , n76262 );
and ( n76264 , n53328 , n57187 );
and ( n76265 , n53041 , n57184 );
nor ( n76266 , n76264 , n76265 );
xnor ( n76267 , n76266 , n56175 );
and ( n76268 , n53922 , n56503 );
and ( n76269 , n53639 , n56501 );
nor ( n76270 , n76268 , n76269 );
xnor ( n76271 , n76270 , n56178 );
and ( n76272 , n76267 , n76271 );
and ( n76273 , n55143 , n55159 );
and ( n76274 , n54942 , n55157 );
nor ( n76275 , n76273 , n76274 );
xnor ( n76276 , n76275 , n54864 );
and ( n76277 , n76271 , n76276 );
and ( n76278 , n76267 , n76276 );
or ( n76279 , n76272 , n76277 , n76278 );
and ( n76280 , n76262 , n76279 );
and ( n76281 , n76257 , n76279 );
or ( n76282 , n76263 , n76280 , n76281 );
and ( n76283 , n76251 , n76282 );
and ( n76284 , n76235 , n76282 );
or ( n76285 , n76252 , n76283 , n76284 );
and ( n76286 , n76226 , n76285 );
and ( n76287 , n76215 , n76285 );
or ( n76288 , n76227 , n76286 , n76287 );
and ( n76289 , n76204 , n76288 );
and ( n76290 , n55756 , n54535 );
and ( n76291 , n55497 , n54533 );
nor ( n76292 , n76290 , n76291 );
xnor ( n76293 , n76292 , n54237 );
and ( n76294 , n56388 , n53928 );
and ( n76295 , n56255 , n53926 );
nor ( n76296 , n76294 , n76295 );
xnor ( n76297 , n76296 , n53652 );
and ( n76298 , n76293 , n76297 );
and ( n76299 , n57063 , n53357 );
and ( n76300 , n56915 , n53355 );
nor ( n76301 , n76299 , n76300 );
xnor ( n76302 , n76301 , n53060 );
and ( n76303 , n76297 , n76302 );
and ( n76304 , n76293 , n76302 );
or ( n76305 , n76298 , n76303 , n76304 );
and ( n76306 , n57063 , n53355 );
not ( n76307 , n76306 );
and ( n76308 , n76307 , n53060 );
xor ( n76309 , n45395 , n45506 );
buf ( n76310 , n76309 );
buf ( n76311 , n76310 );
buf ( n76312 , n76311 );
and ( n76313 , n76308 , n76312 );
and ( n76314 , n69688 , n65210 );
not ( n76315 , n76314 );
and ( n76316 , n76312 , n76315 );
and ( n76317 , n76308 , n76315 );
or ( n76318 , n76313 , n76316 , n76317 );
and ( n76319 , n76305 , n76318 );
xor ( n76320 , n76055 , n76059 );
xor ( n76321 , n76320 , n76064 );
and ( n76322 , n76318 , n76321 );
and ( n76323 , n76305 , n76321 );
or ( n76324 , n76319 , n76322 , n76323 );
xor ( n76325 , n76010 , n76011 );
xor ( n76326 , n76325 , n76013 );
and ( n76327 , n76324 , n76326 );
xor ( n76328 , n76021 , n76022 );
xor ( n76329 , n76328 , n76024 );
and ( n76330 , n76326 , n76329 );
and ( n76331 , n76324 , n76329 );
or ( n76332 , n76327 , n76330 , n76331 );
xor ( n76333 , n76032 , n76041 );
xor ( n76334 , n76333 , n76047 );
xor ( n76335 , n76067 , n76079 );
xor ( n76336 , n76335 , n76092 );
and ( n76337 , n76334 , n76336 );
xor ( n76338 , n76104 , n76106 );
xor ( n76339 , n76338 , n76109 );
and ( n76340 , n76336 , n76339 );
and ( n76341 , n76334 , n76339 );
or ( n76342 , n76337 , n76340 , n76341 );
and ( n76343 , n76332 , n76342 );
xor ( n76344 , n75965 , n75966 );
xor ( n76345 , n76344 , n75978 );
and ( n76346 , n76342 , n76345 );
and ( n76347 , n76332 , n76345 );
or ( n76348 , n76343 , n76346 , n76347 );
and ( n76349 , n76288 , n76348 );
and ( n76350 , n76204 , n76348 );
or ( n76351 , n76289 , n76349 , n76350 );
xor ( n76352 , n76002 , n76007 );
xor ( n76353 , n76352 , n76016 );
xor ( n76354 , n76027 , n76050 );
xor ( n76355 , n76354 , n76095 );
and ( n76356 , n76353 , n76355 );
xor ( n76357 , n76112 , n76114 );
xor ( n76358 , n76357 , n76117 );
and ( n76359 , n76355 , n76358 );
and ( n76360 , n76353 , n76358 );
or ( n76361 , n76356 , n76359 , n76360 );
xor ( n76362 , n75955 , n75956 );
xor ( n76363 , n76362 , n75960 );
and ( n76364 , n76361 , n76363 );
xor ( n76365 , n75981 , n76019 );
xor ( n76366 , n76365 , n76098 );
and ( n76367 , n76363 , n76366 );
and ( n76368 , n76361 , n76366 );
or ( n76369 , n76364 , n76367 , n76368 );
and ( n76370 , n76351 , n76369 );
xor ( n76371 , n75963 , n76101 );
xor ( n76372 , n76371 , n76128 );
and ( n76373 , n76369 , n76372 );
and ( n76374 , n76351 , n76372 );
or ( n76375 , n76370 , n76373 , n76374 );
and ( n76376 , n76195 , n76375 );
xor ( n76377 , n75954 , n76131 );
xor ( n76378 , n76377 , n76150 );
and ( n76379 , n76375 , n76378 );
and ( n76380 , n76195 , n76378 );
or ( n76381 , n76376 , n76379 , n76380 );
and ( n76382 , n76193 , n76381 );
xor ( n76383 , n76153 , n76171 );
xor ( n76384 , n76383 , n76174 );
and ( n76385 , n76381 , n76384 );
and ( n76386 , n76193 , n76384 );
or ( n76387 , n76382 , n76385 , n76386 );
and ( n76388 , n76191 , n76387 );
xor ( n76389 , n75949 , n75951 );
xor ( n76390 , n76389 , n76177 );
and ( n76391 , n76387 , n76390 );
and ( n76392 , n76191 , n76390 );
or ( n76393 , n76388 , n76391 , n76392 );
xor ( n76394 , n75947 , n76180 );
xor ( n76395 , n76394 , n76183 );
and ( n76396 , n76393 , n76395 );
xor ( n76397 , n76191 , n76387 );
xor ( n76398 , n76397 , n76390 );
xor ( n76399 , n76163 , n76165 );
xor ( n76400 , n76399 , n76168 );
xor ( n76401 , n76142 , n76144 );
xor ( n76402 , n76401 , n76147 );
xor ( n76403 , n76155 , n76157 );
xor ( n76404 , n76403 , n76160 );
and ( n76405 , n76402 , n76404 );
xor ( n76406 , n76120 , n76122 );
xor ( n76407 , n76406 , n76125 );
xor ( n76408 , n76134 , n76136 );
xor ( n76409 , n76408 , n76139 );
and ( n76410 , n76407 , n76409 );
xnor ( n76411 , n76212 , n76214 );
and ( n76412 , n66720 , n68610 );
not ( n76413 , n76412 );
and ( n76414 , n68307 , n66917 );
not ( n76415 , n76414 );
and ( n76416 , n76413 , n76415 );
and ( n76417 , n65177 , n69507 );
not ( n76418 , n76417 );
and ( n76419 , n76416 , n76418 );
and ( n76420 , n65678 , n68752 );
not ( n76421 , n76420 );
and ( n76422 , n76418 , n76421 );
and ( n76423 , n76416 , n76421 );
or ( n76424 , n76419 , n76422 , n76423 );
not ( n76425 , n76424 );
and ( n76426 , n68307 , n66469 );
not ( n76427 , n76426 );
and ( n76428 , n67997 , n66917 );
not ( n76429 , n76428 );
and ( n76430 , n76427 , n76429 );
and ( n76431 , n67343 , n67013 );
not ( n76432 , n76431 );
and ( n76433 , n76429 , n76432 );
and ( n76434 , n76427 , n76432 );
or ( n76435 , n76430 , n76433 , n76434 );
and ( n76436 , n76425 , n76435 );
and ( n76437 , n76411 , n76436 );
buf ( n76438 , n76424 );
and ( n76439 , n76436 , n76438 );
and ( n76440 , n76411 , n76438 );
or ( n76441 , n76437 , n76439 , n76440 );
xor ( n76442 , n76071 , n76075 );
xor ( n76443 , n76442 , n75779 );
xor ( n76444 , n76084 , n76086 );
xor ( n76445 , n76444 , n76089 );
and ( n76446 , n76443 , n76445 );
xor ( n76447 , n76220 , n76222 );
and ( n76448 , n76445 , n76447 );
and ( n76449 , n76443 , n76447 );
or ( n76450 , n76446 , n76448 , n76449 );
and ( n76451 , n65177 , n70108 );
not ( n76452 , n76451 );
and ( n76453 , n70256 , n65210 );
not ( n76454 , n76453 );
and ( n76455 , n76452 , n76454 );
and ( n76456 , n54604 , n55851 );
and ( n76457 , n54227 , n55849 );
nor ( n76458 , n76456 , n76457 );
xnor ( n76459 , n76458 , n55506 );
and ( n76460 , n76455 , n76459 );
and ( n76461 , n69303 , n66005 );
not ( n76462 , n76461 );
and ( n76463 , n69059 , n66469 );
not ( n76464 , n76463 );
and ( n76465 , n76462 , n76464 );
and ( n76466 , n67997 , n67013 );
not ( n76467 , n76466 );
and ( n76468 , n76464 , n76467 );
and ( n76469 , n76462 , n76467 );
or ( n76470 , n76465 , n76468 , n76469 );
and ( n76471 , n65678 , n69204 );
not ( n76472 , n76471 );
and ( n76473 , n66415 , n68752 );
not ( n76474 , n76473 );
and ( n76475 , n76472 , n76474 );
and ( n76476 , n66980 , n67844 );
not ( n76477 , n76476 );
and ( n76478 , n76474 , n76477 );
and ( n76479 , n76472 , n76477 );
or ( n76480 , n76475 , n76478 , n76479 );
and ( n76481 , n76470 , n76480 );
and ( n76482 , n76460 , n76481 );
xor ( n76483 , n76427 , n76429 );
xor ( n76484 , n76483 , n76432 );
xor ( n76485 , n76240 , n76242 );
xor ( n76486 , n76485 , n76245 );
and ( n76487 , n76484 , n76486 );
and ( n76488 , n76481 , n76487 );
and ( n76489 , n76460 , n76487 );
or ( n76490 , n76482 , n76488 , n76489 );
and ( n76491 , n76450 , n76490 );
and ( n76492 , n69059 , n66005 );
not ( n76493 , n76492 );
buf ( n76494 , n20823 );
and ( n76495 , n76493 , n76494 );
xor ( n76496 , n76254 , n76256 );
and ( n76497 , n76494 , n76496 );
and ( n76498 , n76493 , n76496 );
or ( n76499 , n76495 , n76497 , n76498 );
xor ( n76500 , n76259 , n76261 );
and ( n76501 , n65606 , n69507 );
not ( n76502 , n76501 );
and ( n76503 , n69688 , n65586 );
not ( n76504 , n76503 );
and ( n76505 , n76502 , n76504 );
and ( n76506 , n76500 , n76505 );
and ( n76507 , n53639 , n57187 );
and ( n76508 , n53328 , n57184 );
nor ( n76509 , n76507 , n76508 );
xnor ( n76510 , n76509 , n56175 );
and ( n76511 , n54942 , n55851 );
and ( n76512 , n54604 , n55849 );
nor ( n76513 , n76511 , n76512 );
xnor ( n76514 , n76513 , n55506 );
and ( n76515 , n76510 , n76514 );
and ( n76516 , n55497 , n55159 );
and ( n76517 , n55143 , n55157 );
nor ( n76518 , n76516 , n76517 );
xnor ( n76519 , n76518 , n54864 );
and ( n76520 , n76514 , n76519 );
and ( n76521 , n76510 , n76519 );
or ( n76522 , n76515 , n76520 , n76521 );
and ( n76523 , n76505 , n76522 );
and ( n76524 , n76500 , n76522 );
or ( n76525 , n76506 , n76523 , n76524 );
and ( n76526 , n76499 , n76525 );
and ( n76527 , n56255 , n54535 );
and ( n76528 , n55756 , n54533 );
nor ( n76529 , n76527 , n76528 );
xnor ( n76530 , n76529 , n54237 );
and ( n76531 , n56915 , n53928 );
and ( n76532 , n56388 , n53926 );
nor ( n76533 , n76531 , n76532 );
xnor ( n76534 , n76533 , n53652 );
and ( n76535 , n76530 , n76534 );
and ( n76536 , n76534 , n76306 );
and ( n76537 , n76530 , n76306 );
or ( n76538 , n76535 , n76536 , n76537 );
xor ( n76539 , n76267 , n76271 );
xor ( n76540 , n76539 , n76276 );
and ( n76541 , n76538 , n76540 );
xor ( n76542 , n76293 , n76297 );
xor ( n76543 , n76542 , n76302 );
and ( n76544 , n76540 , n76543 );
and ( n76545 , n76538 , n76543 );
or ( n76546 , n76541 , n76544 , n76545 );
and ( n76547 , n76525 , n76546 );
and ( n76548 , n76499 , n76546 );
or ( n76549 , n76526 , n76547 , n76548 );
and ( n76550 , n76490 , n76549 );
and ( n76551 , n76450 , n76549 );
or ( n76552 , n76491 , n76550 , n76551 );
and ( n76553 , n76441 , n76552 );
xor ( n76554 , n76228 , n76230 );
xor ( n76555 , n76554 , n76232 );
xor ( n76556 , n76236 , n76237 );
xor ( n76557 , n76556 , n76248 );
and ( n76558 , n76555 , n76557 );
xor ( n76559 , n76257 , n76262 );
xor ( n76560 , n76559 , n76279 );
and ( n76561 , n76557 , n76560 );
and ( n76562 , n76555 , n76560 );
or ( n76563 , n76558 , n76561 , n76562 );
xor ( n76564 , n76216 , n76217 );
xor ( n76565 , n76564 , n76223 );
and ( n76566 , n76563 , n76565 );
xor ( n76567 , n76235 , n76251 );
xor ( n76568 , n76567 , n76282 );
and ( n76569 , n76565 , n76568 );
and ( n76570 , n76563 , n76568 );
or ( n76571 , n76566 , n76569 , n76570 );
and ( n76572 , n76552 , n76571 );
and ( n76573 , n76441 , n76571 );
or ( n76574 , n76553 , n76572 , n76573 );
and ( n76575 , n76409 , n76574 );
and ( n76576 , n76407 , n76574 );
or ( n76577 , n76410 , n76575 , n76576 );
and ( n76578 , n76404 , n76577 );
and ( n76579 , n76402 , n76577 );
or ( n76580 , n76405 , n76578 , n76579 );
and ( n76581 , n76400 , n76580 );
xor ( n76582 , n76195 , n76375 );
xor ( n76583 , n76582 , n76378 );
and ( n76584 , n76580 , n76583 );
and ( n76585 , n76400 , n76583 );
or ( n76586 , n76581 , n76584 , n76585 );
xor ( n76587 , n76193 , n76381 );
xor ( n76588 , n76587 , n76384 );
and ( n76589 , n76586 , n76588 );
xor ( n76590 , n76197 , n76199 );
xor ( n76591 , n76590 , n76201 );
xor ( n76592 , n76215 , n76226 );
xor ( n76593 , n76592 , n76285 );
and ( n76594 , n76591 , n76593 );
xor ( n76595 , n76332 , n76342 );
xor ( n76596 , n76595 , n76345 );
and ( n76597 , n76593 , n76596 );
and ( n76598 , n76591 , n76596 );
or ( n76599 , n76594 , n76597 , n76598 );
xor ( n76600 , n76204 , n76288 );
xor ( n76601 , n76600 , n76348 );
and ( n76602 , n76599 , n76601 );
xor ( n76603 , n76361 , n76363 );
xor ( n76604 , n76603 , n76366 );
and ( n76605 , n76601 , n76604 );
and ( n76606 , n76599 , n76604 );
or ( n76607 , n76602 , n76605 , n76606 );
xor ( n76608 , n76351 , n76369 );
xor ( n76609 , n76608 , n76372 );
and ( n76610 , n76607 , n76609 );
xor ( n76611 , n76353 , n76355 );
xor ( n76612 , n76611 , n76358 );
xor ( n76613 , n76324 , n76326 );
xor ( n76614 , n76613 , n76329 );
xor ( n76615 , n76334 , n76336 );
xor ( n76616 , n76615 , n76339 );
and ( n76617 , n76614 , n76616 );
xor ( n76618 , n76305 , n76318 );
xor ( n76619 , n76618 , n76321 );
xor ( n76620 , n76425 , n76435 );
and ( n76621 , n76619 , n76620 );
xor ( n76622 , n76308 , n76312 );
xor ( n76623 , n76622 , n76315 );
xor ( n76624 , n76416 , n76418 );
xor ( n76625 , n76624 , n76421 );
and ( n76626 , n76623 , n76625 );
xor ( n76627 , n76455 , n76459 );
and ( n76628 , n76625 , n76627 );
and ( n76629 , n76623 , n76627 );
or ( n76630 , n76626 , n76628 , n76629 );
and ( n76631 , n76620 , n76630 );
and ( n76632 , n76619 , n76630 );
or ( n76633 , n76621 , n76631 , n76632 );
and ( n76634 , n76616 , n76633 );
and ( n76635 , n76614 , n76633 );
or ( n76636 , n76617 , n76634 , n76635 );
and ( n76637 , n76612 , n76636 );
xor ( n76638 , n76470 , n76480 );
xor ( n76639 , n76484 , n76486 );
and ( n76640 , n76638 , n76639 );
and ( n76641 , n65606 , n70108 );
not ( n76642 , n76641 );
and ( n76643 , n70256 , n65586 );
not ( n76644 , n76643 );
and ( n76645 , n76642 , n76644 );
and ( n76646 , n66980 , n68610 );
not ( n76647 , n76646 );
and ( n76648 , n68307 , n67013 );
not ( n76649 , n76648 );
and ( n76650 , n76647 , n76649 );
and ( n76651 , n76645 , n76650 );
and ( n76652 , n54227 , n56503 );
and ( n76653 , n53922 , n56501 );
nor ( n76654 , n76652 , n76653 );
xnor ( n76655 , n76654 , n56178 );
and ( n76656 , n76650 , n76655 );
and ( n76657 , n76645 , n76655 );
or ( n76658 , n76651 , n76656 , n76657 );
and ( n76659 , n76639 , n76658 );
and ( n76660 , n76638 , n76658 );
or ( n76661 , n76640 , n76659 , n76660 );
and ( n76662 , n69059 , n66917 );
not ( n76663 , n76662 );
and ( n76664 , n67997 , n67411 );
not ( n76665 , n76664 );
or ( n76666 , n76663 , n76665 );
and ( n76667 , n66720 , n68752 );
not ( n76668 , n76667 );
and ( n76669 , n67343 , n67844 );
not ( n76670 , n76669 );
or ( n76671 , n76668 , n76670 );
and ( n76672 , n76666 , n76671 );
and ( n76673 , n69688 , n66005 );
and ( n76674 , n69303 , n66469 );
not ( n76675 , n76674 );
and ( n76676 , n76673 , n76675 );
and ( n76677 , n65678 , n69507 );
and ( n76678 , n66415 , n69204 );
not ( n76679 , n76678 );
and ( n76680 , n76677 , n76679 );
and ( n76681 , n76676 , n76680 );
and ( n76682 , n76672 , n76681 );
not ( n76683 , n76673 );
buf ( n76684 , n76683 );
not ( n76685 , n76677 );
buf ( n76686 , n76685 );
and ( n76687 , n76684 , n76686 );
and ( n76688 , n76681 , n76687 );
and ( n76689 , n76672 , n76687 );
or ( n76690 , n76682 , n76688 , n76689 );
and ( n76691 , n76661 , n76690 );
xor ( n76692 , n76462 , n76464 );
xor ( n76693 , n76692 , n76467 );
xor ( n76694 , n76472 , n76474 );
xor ( n76695 , n76694 , n76477 );
and ( n76696 , n76693 , n76695 );
xor ( n76697 , n45396 , n45505 );
buf ( n76698 , n76697 );
buf ( n76699 , n76698 );
buf ( n76700 , n76699 );
buf ( n76701 , n20824 );
and ( n76702 , n76700 , n76701 );
xor ( n76703 , n76452 , n76454 );
and ( n76704 , n76701 , n76703 );
and ( n76705 , n76700 , n76703 );
or ( n76706 , n76702 , n76704 , n76705 );
and ( n76707 , n76696 , n76706 );
xor ( n76708 , n76502 , n76504 );
xor ( n76709 , n76413 , n76415 );
and ( n76710 , n76708 , n76709 );
and ( n76711 , n55756 , n55159 );
and ( n76712 , n55497 , n55157 );
nor ( n76713 , n76711 , n76712 );
xnor ( n76714 , n76713 , n54864 );
and ( n76715 , n57063 , n53928 );
and ( n76716 , n56915 , n53926 );
nor ( n76717 , n76715 , n76716 );
xnor ( n76718 , n76717 , n53652 );
and ( n76719 , n76714 , n76718 );
and ( n76720 , n76709 , n76719 );
and ( n76721 , n76708 , n76719 );
or ( n76722 , n76710 , n76720 , n76721 );
and ( n76723 , n76706 , n76722 );
and ( n76724 , n76696 , n76722 );
or ( n76725 , n76707 , n76723 , n76724 );
and ( n76726 , n76690 , n76725 );
and ( n76727 , n76661 , n76725 );
or ( n76728 , n76691 , n76726 , n76727 );
and ( n76729 , n53922 , n57187 );
and ( n76730 , n53639 , n57184 );
nor ( n76731 , n76729 , n76730 );
xnor ( n76732 , n76731 , n56175 );
and ( n76733 , n54604 , n56503 );
and ( n76734 , n54227 , n56501 );
nor ( n76735 , n76733 , n76734 );
xnor ( n76736 , n76735 , n56178 );
and ( n76737 , n76732 , n76736 );
and ( n76738 , n55143 , n55851 );
and ( n76739 , n54942 , n55849 );
nor ( n76740 , n76738 , n76739 );
xnor ( n76741 , n76740 , n55506 );
and ( n76742 , n76736 , n76741 );
and ( n76743 , n76732 , n76741 );
or ( n76744 , n76737 , n76742 , n76743 );
and ( n76745 , n56388 , n54535 );
and ( n76746 , n56255 , n54533 );
nor ( n76747 , n76745 , n76746 );
xnor ( n76748 , n76747 , n54237 );
and ( n76749 , n57063 , n53926 );
not ( n76750 , n76749 );
and ( n76751 , n76750 , n53652 );
and ( n76752 , n76748 , n76751 );
xor ( n76753 , n45398 , n45504 );
buf ( n76754 , n76753 );
buf ( n76755 , n76754 );
buf ( n76756 , n76755 );
and ( n76757 , n76751 , n76756 );
and ( n76758 , n76748 , n76756 );
or ( n76759 , n76752 , n76757 , n76758 );
and ( n76760 , n76744 , n76759 );
xor ( n76761 , n76510 , n76514 );
xor ( n76762 , n76761 , n76519 );
and ( n76763 , n76759 , n76762 );
and ( n76764 , n76744 , n76762 );
or ( n76765 , n76760 , n76763 , n76764 );
xor ( n76766 , n76493 , n76494 );
xor ( n76767 , n76766 , n76496 );
and ( n76768 , n76765 , n76767 );
xor ( n76769 , n76500 , n76505 );
xor ( n76770 , n76769 , n76522 );
and ( n76771 , n76767 , n76770 );
and ( n76772 , n76765 , n76770 );
or ( n76773 , n76768 , n76771 , n76772 );
xor ( n76774 , n76443 , n76445 );
xor ( n76775 , n76774 , n76447 );
and ( n76776 , n76773 , n76775 );
xor ( n76777 , n76460 , n76481 );
xor ( n76778 , n76777 , n76487 );
and ( n76779 , n76775 , n76778 );
and ( n76780 , n76773 , n76778 );
or ( n76781 , n76776 , n76779 , n76780 );
and ( n76782 , n76728 , n76781 );
xor ( n76783 , n76411 , n76436 );
xor ( n76784 , n76783 , n76438 );
and ( n76785 , n76781 , n76784 );
and ( n76786 , n76728 , n76784 );
or ( n76787 , n76782 , n76785 , n76786 );
and ( n76788 , n76636 , n76787 );
and ( n76789 , n76612 , n76787 );
or ( n76790 , n76637 , n76788 , n76789 );
xor ( n76791 , n76407 , n76409 );
xor ( n76792 , n76791 , n76574 );
and ( n76793 , n76790 , n76792 );
xor ( n76794 , n76599 , n76601 );
xor ( n76795 , n76794 , n76604 );
and ( n76796 , n76792 , n76795 );
and ( n76797 , n76790 , n76795 );
or ( n76798 , n76793 , n76796 , n76797 );
and ( n76799 , n76609 , n76798 );
and ( n76800 , n76607 , n76798 );
or ( n76801 , n76610 , n76799 , n76800 );
xor ( n76802 , n76400 , n76580 );
xor ( n76803 , n76802 , n76583 );
and ( n76804 , n76801 , n76803 );
xor ( n76805 , n76402 , n76404 );
xor ( n76806 , n76805 , n76577 );
xor ( n76807 , n76607 , n76609 );
xor ( n76808 , n76807 , n76798 );
and ( n76809 , n76806 , n76808 );
xor ( n76810 , n76441 , n76552 );
xor ( n76811 , n76810 , n76571 );
xor ( n76812 , n76591 , n76593 );
xor ( n76813 , n76812 , n76596 );
and ( n76814 , n76811 , n76813 );
xor ( n76815 , n76450 , n76490 );
xor ( n76816 , n76815 , n76549 );
xor ( n76817 , n76563 , n76565 );
xor ( n76818 , n76817 , n76568 );
and ( n76819 , n76816 , n76818 );
xor ( n76820 , n76499 , n76525 );
xor ( n76821 , n76820 , n76546 );
xor ( n76822 , n76555 , n76557 );
xor ( n76823 , n76822 , n76560 );
and ( n76824 , n76821 , n76823 );
xor ( n76825 , n76538 , n76540 );
xor ( n76826 , n76825 , n76543 );
xor ( n76827 , n76673 , n76675 );
xor ( n76828 , n76677 , n76679 );
and ( n76829 , n76827 , n76828 );
buf ( n76830 , n67343 );
not ( n76831 , n76830 );
or ( n76832 , n76829 , n76831 );
and ( n76833 , n76826 , n76832 );
xor ( n76834 , n76530 , n76534 );
xor ( n76835 , n76834 , n76306 );
xor ( n76836 , n76645 , n76650 );
xor ( n76837 , n76836 , n76655 );
and ( n76838 , n76835 , n76837 );
xor ( n76839 , n76666 , n76671 );
and ( n76840 , n76837 , n76839 );
and ( n76841 , n76835 , n76839 );
or ( n76842 , n76838 , n76840 , n76841 );
and ( n76843 , n76832 , n76842 );
and ( n76844 , n76826 , n76842 );
or ( n76845 , n76833 , n76843 , n76844 );
and ( n76846 , n76823 , n76845 );
and ( n76847 , n76821 , n76845 );
or ( n76848 , n76824 , n76846 , n76847 );
and ( n76849 , n76818 , n76848 );
and ( n76850 , n76816 , n76848 );
or ( n76851 , n76819 , n76849 , n76850 );
and ( n76852 , n76813 , n76851 );
and ( n76853 , n76811 , n76851 );
or ( n76854 , n76814 , n76852 , n76853 );
xor ( n76855 , n76790 , n76792 );
xor ( n76856 , n76855 , n76795 );
and ( n76857 , n76854 , n76856 );
xor ( n76858 , n76676 , n76680 );
xor ( n76859 , n76684 , n76686 );
and ( n76860 , n76858 , n76859 );
xor ( n76861 , n76693 , n76695 );
and ( n76862 , n76859 , n76861 );
and ( n76863 , n76858 , n76861 );
or ( n76864 , n76860 , n76862 , n76863 );
xnor ( n76865 , n76663 , n76665 );
xnor ( n76866 , n76668 , n76670 );
and ( n76867 , n76865 , n76866 );
buf ( n76868 , n20825 );
xor ( n76869 , n76714 , n76718 );
and ( n76870 , n76868 , n76869 );
xor ( n76871 , n76642 , n76644 );
and ( n76872 , n76869 , n76871 );
and ( n76873 , n76868 , n76871 );
or ( n76874 , n76870 , n76872 , n76873 );
and ( n76875 , n76867 , n76874 );
xor ( n76876 , n76647 , n76649 );
and ( n76877 , n66415 , n69507 );
not ( n76878 , n76877 );
and ( n76879 , n66980 , n68752 );
not ( n76880 , n76879 );
and ( n76881 , n76878 , n76880 );
and ( n76882 , n67343 , n68610 );
not ( n76883 , n76882 );
and ( n76884 , n76880 , n76883 );
and ( n76885 , n76878 , n76883 );
or ( n76886 , n76881 , n76884 , n76885 );
and ( n76887 , n76876 , n76886 );
and ( n76888 , n65678 , n70108 );
not ( n76889 , n76888 );
and ( n76890 , n69688 , n66469 );
not ( n76891 , n76890 );
and ( n76892 , n76889 , n76891 );
and ( n76893 , n68307 , n67411 );
not ( n76894 , n76893 );
and ( n76895 , n76891 , n76894 );
and ( n76896 , n76889 , n76894 );
or ( n76897 , n76892 , n76895 , n76896 );
and ( n76898 , n76886 , n76897 );
and ( n76899 , n76876 , n76897 );
or ( n76900 , n76887 , n76898 , n76899 );
and ( n76901 , n76874 , n76900 );
and ( n76902 , n76867 , n76900 );
or ( n76903 , n76875 , n76901 , n76902 );
and ( n76904 , n76864 , n76903 );
and ( n76905 , n70256 , n66005 );
and ( n76906 , n66720 , n69204 );
not ( n76907 , n76906 );
and ( n76908 , n76905 , n76907 );
not ( n76909 , n76905 );
buf ( n76910 , n76909 );
and ( n76911 , n76908 , n76910 );
and ( n76912 , n54227 , n57187 );
and ( n76913 , n53922 , n57184 );
nor ( n76914 , n76912 , n76913 );
xnor ( n76915 , n76914 , n56175 );
and ( n76916 , n55497 , n55851 );
and ( n76917 , n55143 , n55849 );
nor ( n76918 , n76916 , n76917 );
xnor ( n76919 , n76918 , n55506 );
and ( n76920 , n76915 , n76919 );
and ( n76921 , n56255 , n55159 );
and ( n76922 , n55756 , n55157 );
nor ( n76923 , n76921 , n76922 );
xnor ( n76924 , n76923 , n54864 );
and ( n76925 , n76919 , n76924 );
and ( n76926 , n76915 , n76924 );
or ( n76927 , n76920 , n76925 , n76926 );
and ( n76928 , n76910 , n76927 );
and ( n76929 , n76908 , n76927 );
or ( n76930 , n76911 , n76928 , n76929 );
and ( n76931 , n56915 , n54535 );
and ( n76932 , n56388 , n54533 );
nor ( n76933 , n76931 , n76932 );
xnor ( n76934 , n76933 , n54237 );
and ( n76935 , n76934 , n76749 );
xor ( n76936 , n45401 , n45502 );
buf ( n76937 , n76936 );
buf ( n76938 , n76937 );
buf ( n76939 , n76938 );
and ( n76940 , n76749 , n76939 );
and ( n76941 , n76934 , n76939 );
or ( n76942 , n76935 , n76940 , n76941 );
and ( n76943 , n69303 , n66917 );
not ( n76944 , n76943 );
and ( n76945 , n69059 , n67013 );
not ( n76946 , n76945 );
and ( n76947 , n76944 , n76946 );
buf ( n76948 , n67997 );
not ( n76949 , n76948 );
and ( n76950 , n76946 , n76949 );
and ( n76951 , n76944 , n76949 );
or ( n76952 , n76947 , n76950 , n76951 );
and ( n76953 , n76942 , n76952 );
xor ( n76954 , n76732 , n76736 );
xor ( n76955 , n76954 , n76741 );
and ( n76956 , n76952 , n76955 );
and ( n76957 , n76942 , n76955 );
or ( n76958 , n76953 , n76956 , n76957 );
and ( n76959 , n76930 , n76958 );
xor ( n76960 , n76700 , n76701 );
xor ( n76961 , n76960 , n76703 );
and ( n76962 , n76958 , n76961 );
and ( n76963 , n76930 , n76961 );
or ( n76964 , n76959 , n76962 , n76963 );
and ( n76965 , n76903 , n76964 );
and ( n76966 , n76864 , n76964 );
or ( n76967 , n76904 , n76965 , n76966 );
xor ( n76968 , n76623 , n76625 );
xor ( n76969 , n76968 , n76627 );
xor ( n76970 , n76638 , n76639 );
xor ( n76971 , n76970 , n76658 );
and ( n76972 , n76969 , n76971 );
xor ( n76973 , n76672 , n76681 );
xor ( n76974 , n76973 , n76687 );
and ( n76975 , n76971 , n76974 );
and ( n76976 , n76969 , n76974 );
or ( n76977 , n76972 , n76975 , n76976 );
and ( n76978 , n76967 , n76977 );
xor ( n76979 , n76619 , n76620 );
xor ( n76980 , n76979 , n76630 );
and ( n76981 , n76977 , n76980 );
and ( n76982 , n76967 , n76980 );
or ( n76983 , n76978 , n76981 , n76982 );
xor ( n76984 , n76614 , n76616 );
xor ( n76985 , n76984 , n76633 );
and ( n76986 , n76983 , n76985 );
xor ( n76987 , n76728 , n76781 );
xor ( n76988 , n76987 , n76784 );
and ( n76989 , n76985 , n76988 );
and ( n76990 , n76983 , n76988 );
or ( n76991 , n76986 , n76989 , n76990 );
xor ( n76992 , n76612 , n76636 );
xor ( n76993 , n76992 , n76787 );
and ( n76994 , n76991 , n76993 );
xor ( n76995 , n76661 , n76690 );
xor ( n76996 , n76995 , n76725 );
xor ( n76997 , n76773 , n76775 );
xor ( n76998 , n76997 , n76778 );
and ( n76999 , n76996 , n76998 );
xor ( n77000 , n76696 , n76706 );
xor ( n77001 , n77000 , n76722 );
xor ( n77002 , n76765 , n76767 );
xor ( n77003 , n77002 , n76770 );
and ( n77004 , n77001 , n77003 );
xor ( n77005 , n76708 , n76709 );
xor ( n77006 , n77005 , n76719 );
xor ( n77007 , n76744 , n76759 );
xor ( n77008 , n77007 , n76762 );
and ( n77009 , n77006 , n77008 );
xnor ( n77010 , n76829 , n76831 );
and ( n77011 , n77008 , n77010 );
and ( n77012 , n77006 , n77010 );
or ( n77013 , n77009 , n77011 , n77012 );
and ( n77014 , n77003 , n77013 );
and ( n77015 , n77001 , n77013 );
or ( n77016 , n77004 , n77014 , n77015 );
and ( n77017 , n76998 , n77016 );
and ( n77018 , n76996 , n77016 );
or ( n77019 , n76999 , n77017 , n77018 );
xor ( n77020 , n76748 , n76751 );
xor ( n77021 , n77020 , n76756 );
xor ( n77022 , n76865 , n76866 );
and ( n77023 , n77021 , n77022 );
xor ( n77024 , n76827 , n76828 );
and ( n77025 , n77022 , n77024 );
and ( n77026 , n77021 , n77024 );
or ( n77027 , n77023 , n77025 , n77026 );
and ( n77028 , n66415 , n70108 );
not ( n77029 , n77028 );
and ( n77030 , n70256 , n66469 );
not ( n77031 , n77030 );
and ( n77032 , n77029 , n77031 );
and ( n77033 , n67343 , n68752 );
not ( n77034 , n77033 );
and ( n77035 , n69059 , n67411 );
not ( n77036 , n77035 );
and ( n77037 , n77034 , n77036 );
and ( n77038 , n77032 , n77037 );
and ( n77039 , n54942 , n56503 );
and ( n77040 , n54604 , n56501 );
nor ( n77041 , n77039 , n77040 );
xnor ( n77042 , n77041 , n56178 );
and ( n77043 , n77037 , n77042 );
and ( n77044 , n77032 , n77042 );
or ( n77045 , n77038 , n77043 , n77044 );
buf ( n77046 , n20826 );
xor ( n77047 , n76878 , n76880 );
xor ( n77048 , n77047 , n76883 );
and ( n77049 , n77046 , n77048 );
xor ( n77050 , n76889 , n76891 );
xor ( n77051 , n77050 , n76894 );
and ( n77052 , n77048 , n77051 );
and ( n77053 , n77046 , n77051 );
or ( n77054 , n77049 , n77052 , n77053 );
and ( n77055 , n77045 , n77054 );
xor ( n77056 , n76905 , n76907 );
and ( n77057 , n66720 , n69507 );
not ( n77058 , n77057 );
and ( n77059 , n69688 , n66917 );
not ( n77060 , n77059 );
and ( n77061 , n77058 , n77060 );
and ( n77062 , n77056 , n77061 );
and ( n77063 , n66980 , n69204 );
not ( n77064 , n77063 );
and ( n77065 , n69303 , n67013 );
not ( n77066 , n77065 );
and ( n77067 , n77064 , n77066 );
and ( n77068 , n77061 , n77067 );
and ( n77069 , n77056 , n77067 );
or ( n77070 , n77062 , n77068 , n77069 );
and ( n77071 , n77054 , n77070 );
and ( n77072 , n77045 , n77070 );
or ( n77073 , n77055 , n77071 , n77072 );
and ( n77074 , n77027 , n77073 );
and ( n77075 , n54604 , n57187 );
and ( n77076 , n54227 , n57184 );
nor ( n77077 , n77075 , n77076 );
xnor ( n77078 , n77077 , n56175 );
and ( n77079 , n55143 , n56503 );
and ( n77080 , n54942 , n56501 );
nor ( n77081 , n77079 , n77080 );
xnor ( n77082 , n77081 , n56178 );
and ( n77083 , n77078 , n77082 );
and ( n77084 , n55756 , n55851 );
and ( n77085 , n55497 , n55849 );
nor ( n77086 , n77084 , n77085 );
xnor ( n77087 , n77086 , n55506 );
and ( n77088 , n77082 , n77087 );
and ( n77089 , n77078 , n77087 );
or ( n77090 , n77083 , n77088 , n77089 );
and ( n77091 , n56388 , n55159 );
and ( n77092 , n56255 , n55157 );
nor ( n77093 , n77091 , n77092 );
xnor ( n77094 , n77093 , n54864 );
and ( n77095 , n57063 , n54535 );
and ( n77096 , n56915 , n54533 );
nor ( n77097 , n77095 , n77096 );
xnor ( n77098 , n77097 , n54237 );
and ( n77099 , n77094 , n77098 );
and ( n77100 , n57063 , n54533 );
not ( n77101 , n77100 );
and ( n77102 , n77101 , n54237 );
and ( n77103 , n77098 , n77102 );
and ( n77104 , n77094 , n77102 );
or ( n77105 , n77099 , n77103 , n77104 );
and ( n77106 , n77090 , n77105 );
xor ( n77107 , n45402 , n45501 );
buf ( n77108 , n77107 );
buf ( n77109 , n77108 );
buf ( n77110 , n77109 );
and ( n77111 , n68307 , n67844 );
not ( n77112 , n77111 );
and ( n77113 , n77110 , n77112 );
and ( n77114 , n67997 , n68610 );
not ( n77115 , n77114 );
and ( n77116 , n77112 , n77115 );
and ( n77117 , n77110 , n77115 );
or ( n77118 , n77113 , n77116 , n77117 );
and ( n77119 , n77105 , n77118 );
and ( n77120 , n77090 , n77118 );
or ( n77121 , n77106 , n77119 , n77120 );
xor ( n77122 , n76915 , n76919 );
xor ( n77123 , n77122 , n76924 );
xor ( n77124 , n76934 , n76749 );
xor ( n77125 , n77124 , n76939 );
and ( n77126 , n77123 , n77125 );
xor ( n77127 , n76944 , n76946 );
xor ( n77128 , n77127 , n76949 );
and ( n77129 , n77125 , n77128 );
and ( n77130 , n77123 , n77128 );
or ( n77131 , n77126 , n77129 , n77130 );
and ( n77132 , n77121 , n77131 );
xor ( n77133 , n76868 , n76869 );
xor ( n77134 , n77133 , n76871 );
and ( n77135 , n77131 , n77134 );
and ( n77136 , n77121 , n77134 );
or ( n77137 , n77132 , n77135 , n77136 );
and ( n77138 , n77073 , n77137 );
and ( n77139 , n77027 , n77137 );
or ( n77140 , n77074 , n77138 , n77139 );
xor ( n77141 , n76876 , n76886 );
xor ( n77142 , n77141 , n76897 );
xor ( n77143 , n76908 , n76910 );
xor ( n77144 , n77143 , n76927 );
and ( n77145 , n77142 , n77144 );
xor ( n77146 , n76942 , n76952 );
xor ( n77147 , n77146 , n76955 );
and ( n77148 , n77144 , n77147 );
and ( n77149 , n77142 , n77147 );
or ( n77150 , n77145 , n77148 , n77149 );
xor ( n77151 , n76835 , n76837 );
xor ( n77152 , n77151 , n76839 );
and ( n77153 , n77150 , n77152 );
xor ( n77154 , n76858 , n76859 );
xor ( n77155 , n77154 , n76861 );
and ( n77156 , n77152 , n77155 );
and ( n77157 , n77150 , n77155 );
or ( n77158 , n77153 , n77156 , n77157 );
and ( n77159 , n77140 , n77158 );
xor ( n77160 , n76826 , n76832 );
xor ( n77161 , n77160 , n76842 );
and ( n77162 , n77158 , n77161 );
and ( n77163 , n77140 , n77161 );
or ( n77164 , n77159 , n77162 , n77163 );
xor ( n77165 , n76821 , n76823 );
xor ( n77166 , n77165 , n76845 );
and ( n77167 , n77164 , n77166 );
xor ( n77168 , n76967 , n76977 );
xor ( n77169 , n77168 , n76980 );
and ( n77170 , n77166 , n77169 );
and ( n77171 , n77164 , n77169 );
or ( n77172 , n77167 , n77170 , n77171 );
and ( n77173 , n77019 , n77172 );
xor ( n77174 , n76816 , n76818 );
xor ( n77175 , n77174 , n76848 );
and ( n77176 , n77172 , n77175 );
and ( n77177 , n77019 , n77175 );
or ( n77178 , n77173 , n77176 , n77177 );
and ( n77179 , n76993 , n77178 );
and ( n77180 , n76991 , n77178 );
or ( n77181 , n76994 , n77179 , n77180 );
and ( n77182 , n76856 , n77181 );
and ( n77183 , n76854 , n77181 );
or ( n77184 , n76857 , n77182 , n77183 );
and ( n77185 , n76808 , n77184 );
and ( n77186 , n76806 , n77184 );
or ( n77187 , n76809 , n77185 , n77186 );
and ( n77188 , n76803 , n77187 );
and ( n77189 , n76801 , n77187 );
or ( n77190 , n76804 , n77188 , n77189 );
and ( n77191 , n76588 , n77190 );
and ( n77192 , n76586 , n77190 );
or ( n77193 , n76589 , n77191 , n77192 );
or ( n77194 , n76398 , n77193 );
and ( n77195 , n76395 , n77194 );
and ( n77196 , n76393 , n77194 );
or ( n77197 , n76396 , n77195 , n77196 );
and ( n77198 , n76188 , n77197 );
and ( n77199 , n76186 , n77197 );
or ( n77200 , n76189 , n77198 , n77199 );
and ( n77201 , n75945 , n77200 );
xor ( n77202 , n75945 , n77200 );
xor ( n77203 , n76186 , n76188 );
xor ( n77204 , n77203 , n77197 );
not ( n77205 , n77204 );
xor ( n77206 , n76393 , n76395 );
xor ( n77207 , n77206 , n77194 );
xnor ( n77208 , n76398 , n77193 );
xor ( n77209 , n76586 , n76588 );
xor ( n77210 , n77209 , n77190 );
xor ( n77211 , n76801 , n76803 );
xor ( n77212 , n77211 , n77187 );
xor ( n77213 , n76806 , n76808 );
xor ( n77214 , n77213 , n77184 );
xor ( n77215 , n76811 , n76813 );
xor ( n77216 , n77215 , n76851 );
xor ( n77217 , n76983 , n76985 );
xor ( n77218 , n77217 , n76988 );
xor ( n77219 , n76864 , n76903 );
xor ( n77220 , n77219 , n76964 );
xor ( n77221 , n76969 , n76971 );
xor ( n77222 , n77221 , n76974 );
and ( n77223 , n77220 , n77222 );
xor ( n77224 , n76867 , n76874 );
xor ( n77225 , n77224 , n76900 );
xor ( n77226 , n76930 , n76958 );
xor ( n77227 , n77226 , n76961 );
and ( n77228 , n77225 , n77227 );
xor ( n77229 , n77032 , n77037 );
xor ( n77230 , n77229 , n77042 );
buf ( n77231 , n20827 );
xor ( n77232 , n77029 , n77031 );
and ( n77233 , n77231 , n77232 );
xor ( n77234 , n77058 , n77060 );
and ( n77235 , n77232 , n77234 );
and ( n77236 , n77231 , n77234 );
or ( n77237 , n77233 , n77235 , n77236 );
and ( n77238 , n77230 , n77237 );
xor ( n77239 , n77064 , n77066 );
xor ( n77240 , n77034 , n77036 );
and ( n77241 , n77239 , n77240 );
and ( n77242 , n67343 , n69204 );
not ( n77243 , n77242 );
and ( n77244 , n67997 , n68752 );
not ( n77245 , n77244 );
and ( n77246 , n77243 , n77245 );
buf ( n77247 , n68307 );
not ( n77248 , n77247 );
and ( n77249 , n77245 , n77248 );
and ( n77250 , n77243 , n77248 );
or ( n77251 , n77246 , n77249 , n77250 );
and ( n77252 , n77240 , n77251 );
and ( n77253 , n77239 , n77251 );
or ( n77254 , n77241 , n77252 , n77253 );
and ( n77255 , n77237 , n77254 );
and ( n77256 , n77230 , n77254 );
or ( n77257 , n77238 , n77255 , n77256 );
and ( n77258 , n66720 , n70108 );
not ( n77259 , n77258 );
and ( n77260 , n69303 , n67411 );
not ( n77261 , n77260 );
and ( n77262 , n77259 , n77261 );
and ( n77263 , n69059 , n67844 );
not ( n77264 , n77263 );
and ( n77265 , n77261 , n77264 );
and ( n77266 , n77259 , n77264 );
or ( n77267 , n77262 , n77265 , n77266 );
and ( n77268 , n70256 , n66917 );
not ( n77269 , n77268 );
and ( n77270 , n66980 , n69507 );
and ( n77271 , n77269 , n77270 );
and ( n77272 , n77267 , n77271 );
not ( n77273 , n77270 );
buf ( n77274 , n77273 );
and ( n77275 , n77271 , n77274 );
and ( n77276 , n77267 , n77274 );
or ( n77277 , n77272 , n77275 , n77276 );
and ( n77278 , n54942 , n57187 );
and ( n77279 , n54604 , n57184 );
nor ( n77280 , n77278 , n77279 );
xnor ( n77281 , n77280 , n56175 );
and ( n77282 , n55497 , n56503 );
and ( n77283 , n55143 , n56501 );
nor ( n77284 , n77282 , n77283 );
xnor ( n77285 , n77284 , n56178 );
and ( n77286 , n77281 , n77285 );
and ( n77287 , n56255 , n55851 );
and ( n77288 , n55756 , n55849 );
nor ( n77289 , n77287 , n77288 );
xnor ( n77290 , n77289 , n55506 );
and ( n77291 , n77285 , n77290 );
and ( n77292 , n77281 , n77290 );
or ( n77293 , n77286 , n77291 , n77292 );
and ( n77294 , n56915 , n55159 );
and ( n77295 , n56388 , n55157 );
nor ( n77296 , n77294 , n77295 );
xnor ( n77297 , n77296 , n54864 );
and ( n77298 , n77297 , n77100 );
xor ( n77299 , n45404 , n45500 );
buf ( n77300 , n77299 );
buf ( n77301 , n77300 );
buf ( n77302 , n77301 );
and ( n77303 , n77100 , n77302 );
and ( n77304 , n77297 , n77302 );
or ( n77305 , n77298 , n77303 , n77304 );
and ( n77306 , n77293 , n77305 );
xor ( n77307 , n77078 , n77082 );
xor ( n77308 , n77307 , n77087 );
and ( n77309 , n77305 , n77308 );
and ( n77310 , n77293 , n77308 );
or ( n77311 , n77306 , n77309 , n77310 );
and ( n77312 , n77277 , n77311 );
xor ( n77313 , n77046 , n77048 );
xor ( n77314 , n77313 , n77051 );
and ( n77315 , n77311 , n77314 );
and ( n77316 , n77277 , n77314 );
or ( n77317 , n77312 , n77315 , n77316 );
and ( n77318 , n77257 , n77317 );
xor ( n77319 , n77056 , n77061 );
xor ( n77320 , n77319 , n77067 );
xor ( n77321 , n77090 , n77105 );
xor ( n77322 , n77321 , n77118 );
and ( n77323 , n77320 , n77322 );
xor ( n77324 , n77123 , n77125 );
xor ( n77325 , n77324 , n77128 );
and ( n77326 , n77322 , n77325 );
and ( n77327 , n77320 , n77325 );
or ( n77328 , n77323 , n77326 , n77327 );
and ( n77329 , n77317 , n77328 );
and ( n77330 , n77257 , n77328 );
or ( n77331 , n77318 , n77329 , n77330 );
and ( n77332 , n77227 , n77331 );
and ( n77333 , n77225 , n77331 );
or ( n77334 , n77228 , n77332 , n77333 );
and ( n77335 , n77222 , n77334 );
and ( n77336 , n77220 , n77334 );
or ( n77337 , n77223 , n77335 , n77336 );
xor ( n77338 , n77021 , n77022 );
xor ( n77339 , n77338 , n77024 );
xor ( n77340 , n77045 , n77054 );
xor ( n77341 , n77340 , n77070 );
and ( n77342 , n77339 , n77341 );
xor ( n77343 , n77121 , n77131 );
xor ( n77344 , n77343 , n77134 );
and ( n77345 , n77341 , n77344 );
and ( n77346 , n77339 , n77344 );
or ( n77347 , n77342 , n77345 , n77346 );
xor ( n77348 , n77006 , n77008 );
xor ( n77349 , n77348 , n77010 );
and ( n77350 , n77347 , n77349 );
xor ( n77351 , n77027 , n77073 );
xor ( n77352 , n77351 , n77137 );
and ( n77353 , n77349 , n77352 );
and ( n77354 , n77347 , n77352 );
or ( n77355 , n77350 , n77353 , n77354 );
xor ( n77356 , n77001 , n77003 );
xor ( n77357 , n77356 , n77013 );
and ( n77358 , n77355 , n77357 );
xor ( n77359 , n77140 , n77158 );
xor ( n77360 , n77359 , n77161 );
and ( n77361 , n77357 , n77360 );
and ( n77362 , n77355 , n77360 );
or ( n77363 , n77358 , n77361 , n77362 );
and ( n77364 , n77337 , n77363 );
xor ( n77365 , n76996 , n76998 );
xor ( n77366 , n77365 , n77016 );
and ( n77367 , n77363 , n77366 );
and ( n77368 , n77337 , n77366 );
or ( n77369 , n77364 , n77367 , n77368 );
and ( n77370 , n77218 , n77369 );
xor ( n77371 , n77019 , n77172 );
xor ( n77372 , n77371 , n77175 );
and ( n77373 , n77369 , n77372 );
and ( n77374 , n77218 , n77372 );
or ( n77375 , n77370 , n77373 , n77374 );
and ( n77376 , n77216 , n77375 );
xor ( n77377 , n76991 , n76993 );
xor ( n77378 , n77377 , n77178 );
and ( n77379 , n77375 , n77378 );
and ( n77380 , n77216 , n77378 );
or ( n77381 , n77376 , n77379 , n77380 );
xor ( n77382 , n76854 , n76856 );
xor ( n77383 , n77382 , n77181 );
and ( n77384 , n77381 , n77383 );
xor ( n77385 , n77164 , n77166 );
xor ( n77386 , n77385 , n77169 );
xor ( n77387 , n77150 , n77152 );
xor ( n77388 , n77387 , n77155 );
xor ( n77389 , n77142 , n77144 );
xor ( n77390 , n77389 , n77147 );
xor ( n77391 , n77094 , n77098 );
xor ( n77392 , n77391 , n77102 );
xor ( n77393 , n77110 , n77112 );
xor ( n77394 , n77393 , n77115 );
and ( n77395 , n77392 , n77394 );
and ( n77396 , n69688 , n67411 );
not ( n77397 , n77396 );
and ( n77398 , n69303 , n67844 );
not ( n77399 , n77398 );
or ( n77400 , n77397 , n77399 );
and ( n77401 , n67343 , n69507 );
not ( n77402 , n77401 );
and ( n77403 , n67997 , n69204 );
not ( n77404 , n77403 );
or ( n77405 , n77402 , n77404 );
and ( n77406 , n77400 , n77405 );
and ( n77407 , n77394 , n77406 );
and ( n77408 , n77392 , n77406 );
or ( n77409 , n77395 , n77407 , n77408 );
and ( n77410 , n69688 , n67013 );
not ( n77411 , n77410 );
buf ( n77412 , n20828 );
and ( n77413 , n77411 , n77412 );
xor ( n77414 , n77243 , n77245 );
xor ( n77415 , n77414 , n77248 );
and ( n77416 , n77412 , n77415 );
and ( n77417 , n77411 , n77415 );
or ( n77418 , n77413 , n77416 , n77417 );
xor ( n77419 , n77259 , n77261 );
xor ( n77420 , n77419 , n77264 );
xor ( n77421 , n77269 , n77270 );
and ( n77422 , n77420 , n77421 );
and ( n77423 , n66980 , n70108 );
not ( n77424 , n77423 );
and ( n77425 , n70256 , n67013 );
not ( n77426 , n77425 );
and ( n77427 , n77424 , n77426 );
and ( n77428 , n77421 , n77427 );
and ( n77429 , n77420 , n77427 );
or ( n77430 , n77422 , n77428 , n77429 );
and ( n77431 , n77418 , n77430 );
and ( n77432 , n68307 , n68752 );
not ( n77433 , n77432 );
and ( n77434 , n69059 , n68610 );
not ( n77435 , n77434 );
and ( n77436 , n77433 , n77435 );
and ( n77437 , n55143 , n57187 );
and ( n77438 , n54942 , n57184 );
nor ( n77439 , n77437 , n77438 );
xnor ( n77440 , n77439 , n56175 );
and ( n77441 , n55756 , n56503 );
and ( n77442 , n55497 , n56501 );
nor ( n77443 , n77441 , n77442 );
xnor ( n77444 , n77443 , n56178 );
and ( n77445 , n77440 , n77444 );
and ( n77446 , n56388 , n55851 );
and ( n77447 , n56255 , n55849 );
nor ( n77448 , n77446 , n77447 );
xnor ( n77449 , n77448 , n55506 );
and ( n77450 , n77444 , n77449 );
and ( n77451 , n77440 , n77449 );
or ( n77452 , n77445 , n77450 , n77451 );
and ( n77453 , n77436 , n77452 );
and ( n77454 , n57063 , n55159 );
and ( n77455 , n56915 , n55157 );
nor ( n77456 , n77454 , n77455 );
xnor ( n77457 , n77456 , n54864 );
and ( n77458 , n57063 , n55157 );
not ( n77459 , n77458 );
and ( n77460 , n77459 , n54864 );
and ( n77461 , n77457 , n77460 );
xor ( n77462 , n45406 , n45499 );
buf ( n77463 , n77462 );
buf ( n77464 , n77463 );
buf ( n77465 , n77464 );
and ( n77466 , n77460 , n77465 );
and ( n77467 , n77457 , n77465 );
or ( n77468 , n77461 , n77466 , n77467 );
and ( n77469 , n77452 , n77468 );
and ( n77470 , n77436 , n77468 );
or ( n77471 , n77453 , n77469 , n77470 );
and ( n77472 , n77430 , n77471 );
and ( n77473 , n77418 , n77471 );
or ( n77474 , n77431 , n77472 , n77473 );
and ( n77475 , n77409 , n77474 );
xor ( n77476 , n77231 , n77232 );
xor ( n77477 , n77476 , n77234 );
xor ( n77478 , n77239 , n77240 );
xor ( n77479 , n77478 , n77251 );
and ( n77480 , n77477 , n77479 );
xor ( n77481 , n77267 , n77271 );
xor ( n77482 , n77481 , n77274 );
and ( n77483 , n77479 , n77482 );
and ( n77484 , n77477 , n77482 );
or ( n77485 , n77480 , n77483 , n77484 );
and ( n77486 , n77474 , n77485 );
and ( n77487 , n77409 , n77485 );
or ( n77488 , n77475 , n77486 , n77487 );
and ( n77489 , n77390 , n77488 );
xor ( n77490 , n77230 , n77237 );
xor ( n77491 , n77490 , n77254 );
xor ( n77492 , n77277 , n77311 );
xor ( n77493 , n77492 , n77314 );
and ( n77494 , n77491 , n77493 );
xor ( n77495 , n77320 , n77322 );
xor ( n77496 , n77495 , n77325 );
and ( n77497 , n77493 , n77496 );
and ( n77498 , n77491 , n77496 );
or ( n77499 , n77494 , n77497 , n77498 );
and ( n77500 , n77488 , n77499 );
and ( n77501 , n77390 , n77499 );
or ( n77502 , n77489 , n77500 , n77501 );
and ( n77503 , n77388 , n77502 );
xor ( n77504 , n77225 , n77227 );
xor ( n77505 , n77504 , n77331 );
and ( n77506 , n77502 , n77505 );
and ( n77507 , n77388 , n77505 );
or ( n77508 , n77503 , n77506 , n77507 );
xor ( n77509 , n77220 , n77222 );
xor ( n77510 , n77509 , n77334 );
and ( n77511 , n77508 , n77510 );
xor ( n77512 , n77355 , n77357 );
xor ( n77513 , n77512 , n77360 );
and ( n77514 , n77510 , n77513 );
and ( n77515 , n77508 , n77513 );
or ( n77516 , n77511 , n77514 , n77515 );
and ( n77517 , n77386 , n77516 );
xor ( n77518 , n77337 , n77363 );
xor ( n77519 , n77518 , n77366 );
and ( n77520 , n77516 , n77519 );
and ( n77521 , n77386 , n77519 );
or ( n77522 , n77517 , n77520 , n77521 );
xor ( n77523 , n77218 , n77369 );
xor ( n77524 , n77523 , n77372 );
or ( n77525 , n77522 , n77524 );
xor ( n77526 , n77216 , n77375 );
xor ( n77527 , n77526 , n77378 );
or ( n77528 , n77525 , n77527 );
and ( n77529 , n77383 , n77528 );
and ( n77530 , n77381 , n77528 );
or ( n77531 , n77384 , n77529 , n77530 );
or ( n77532 , n77214 , n77531 );
and ( n77533 , n77212 , n77532 );
xor ( n77534 , n77212 , n77532 );
xnor ( n77535 , n77214 , n77531 );
xor ( n77536 , n77381 , n77383 );
xor ( n77537 , n77536 , n77528 );
xnor ( n77538 , n77525 , n77527 );
xnor ( n77539 , n77522 , n77524 );
xor ( n77540 , n77386 , n77516 );
xor ( n77541 , n77540 , n77519 );
xor ( n77542 , n77347 , n77349 );
xor ( n77543 , n77542 , n77352 );
xor ( n77544 , n77257 , n77317 );
xor ( n77545 , n77544 , n77328 );
xor ( n77546 , n77339 , n77341 );
xor ( n77547 , n77546 , n77344 );
and ( n77548 , n77545 , n77547 );
xor ( n77549 , n77293 , n77305 );
xor ( n77550 , n77549 , n77308 );
xor ( n77551 , n77281 , n77285 );
xor ( n77552 , n77551 , n77290 );
xor ( n77553 , n77297 , n77100 );
xor ( n77554 , n77553 , n77302 );
and ( n77555 , n77552 , n77554 );
xor ( n77556 , n77400 , n77405 );
and ( n77557 , n77554 , n77556 );
and ( n77558 , n77552 , n77556 );
or ( n77559 , n77555 , n77557 , n77558 );
and ( n77560 , n77550 , n77559 );
and ( n77561 , n70256 , n67411 );
not ( n77562 , n77561 );
and ( n77563 , n69688 , n67844 );
not ( n77564 , n77563 );
and ( n77565 , n77562 , n77564 );
and ( n77566 , n69303 , n68610 );
not ( n77567 , n77566 );
and ( n77568 , n77564 , n77567 );
and ( n77569 , n77562 , n77567 );
or ( n77570 , n77565 , n77568 , n77569 );
and ( n77571 , n67343 , n70108 );
not ( n77572 , n77571 );
and ( n77573 , n67997 , n69507 );
not ( n77574 , n77573 );
and ( n77575 , n77572 , n77574 );
and ( n77576 , n68307 , n69204 );
not ( n77577 , n77576 );
and ( n77578 , n77574 , n77577 );
and ( n77579 , n77572 , n77577 );
or ( n77580 , n77575 , n77578 , n77579 );
and ( n77581 , n77570 , n77580 );
xnor ( n77582 , n77397 , n77399 );
xnor ( n77583 , n77402 , n77404 );
and ( n77584 , n77582 , n77583 );
and ( n77585 , n77581 , n77584 );
buf ( n77586 , n20829 );
xor ( n77587 , n77424 , n77426 );
and ( n77588 , n77586 , n77587 );
xor ( n77589 , n77433 , n77435 );
and ( n77590 , n77587 , n77589 );
and ( n77591 , n77586 , n77589 );
or ( n77592 , n77588 , n77590 , n77591 );
and ( n77593 , n77584 , n77592 );
and ( n77594 , n77581 , n77592 );
or ( n77595 , n77585 , n77593 , n77594 );
and ( n77596 , n77559 , n77595 );
and ( n77597 , n77550 , n77595 );
or ( n77598 , n77560 , n77596 , n77597 );
and ( n77599 , n55497 , n57187 );
and ( n77600 , n55143 , n57184 );
nor ( n77601 , n77599 , n77600 );
xnor ( n77602 , n77601 , n56175 );
and ( n77603 , n56255 , n56503 );
and ( n77604 , n55756 , n56501 );
nor ( n77605 , n77603 , n77604 );
xnor ( n77606 , n77605 , n56178 );
and ( n77607 , n77602 , n77606 );
and ( n77608 , n56915 , n55851 );
and ( n77609 , n56388 , n55849 );
nor ( n77610 , n77608 , n77609 );
xnor ( n77611 , n77610 , n55506 );
and ( n77612 , n77606 , n77611 );
and ( n77613 , n77602 , n77611 );
or ( n77614 , n77607 , n77612 , n77613 );
xor ( n77615 , n45457 , n45497 );
buf ( n77616 , n77615 );
buf ( n77617 , n77616 );
buf ( n77618 , n77617 );
and ( n77619 , n77458 , n77618 );
buf ( n77620 , n69059 );
not ( n77621 , n77620 );
and ( n77622 , n77618 , n77621 );
and ( n77623 , n77458 , n77621 );
or ( n77624 , n77619 , n77622 , n77623 );
and ( n77625 , n77614 , n77624 );
xor ( n77626 , n77440 , n77444 );
xor ( n77627 , n77626 , n77449 );
and ( n77628 , n77624 , n77627 );
and ( n77629 , n77614 , n77627 );
or ( n77630 , n77625 , n77628 , n77629 );
xor ( n77631 , n77411 , n77412 );
xor ( n77632 , n77631 , n77415 );
and ( n77633 , n77630 , n77632 );
xor ( n77634 , n77420 , n77421 );
xor ( n77635 , n77634 , n77427 );
and ( n77636 , n77632 , n77635 );
and ( n77637 , n77630 , n77635 );
or ( n77638 , n77633 , n77636 , n77637 );
xor ( n77639 , n77392 , n77394 );
xor ( n77640 , n77639 , n77406 );
and ( n77641 , n77638 , n77640 );
xor ( n77642 , n77418 , n77430 );
xor ( n77643 , n77642 , n77471 );
and ( n77644 , n77640 , n77643 );
and ( n77645 , n77638 , n77643 );
or ( n77646 , n77641 , n77644 , n77645 );
and ( n77647 , n77598 , n77646 );
xor ( n77648 , n77409 , n77474 );
xor ( n77649 , n77648 , n77485 );
and ( n77650 , n77646 , n77649 );
and ( n77651 , n77598 , n77649 );
or ( n77652 , n77647 , n77650 , n77651 );
and ( n77653 , n77547 , n77652 );
and ( n77654 , n77545 , n77652 );
or ( n77655 , n77548 , n77653 , n77654 );
and ( n77656 , n77543 , n77655 );
xor ( n77657 , n77388 , n77502 );
xor ( n77658 , n77657 , n77505 );
and ( n77659 , n77655 , n77658 );
and ( n77660 , n77543 , n77658 );
or ( n77661 , n77656 , n77659 , n77660 );
xor ( n77662 , n77508 , n77510 );
xor ( n77663 , n77662 , n77513 );
and ( n77664 , n77661 , n77663 );
xor ( n77665 , n77390 , n77488 );
xor ( n77666 , n77665 , n77499 );
xor ( n77667 , n77491 , n77493 );
xor ( n77668 , n77667 , n77496 );
xor ( n77669 , n77477 , n77479 );
xor ( n77670 , n77669 , n77482 );
xor ( n77671 , n77436 , n77452 );
xor ( n77672 , n77671 , n77468 );
xor ( n77673 , n77457 , n77460 );
xor ( n77674 , n77673 , n77465 );
xor ( n77675 , n77570 , n77580 );
and ( n77676 , n77674 , n77675 );
xor ( n77677 , n77582 , n77583 );
and ( n77678 , n77675 , n77677 );
and ( n77679 , n77674 , n77677 );
or ( n77680 , n77676 , n77678 , n77679 );
and ( n77681 , n77672 , n77680 );
and ( n77682 , n70256 , n67844 );
not ( n77683 , n77682 );
and ( n77684 , n69688 , n68610 );
not ( n77685 , n77684 );
and ( n77686 , n77683 , n77685 );
and ( n77687 , n67997 , n70108 );
not ( n77688 , n77687 );
and ( n77689 , n68307 , n69507 );
not ( n77690 , n77689 );
and ( n77691 , n77688 , n77690 );
and ( n77692 , n77686 , n77691 );
xor ( n77693 , n77562 , n77564 );
xor ( n77694 , n77693 , n77567 );
xor ( n77695 , n77572 , n77574 );
xor ( n77696 , n77695 , n77577 );
and ( n77697 , n77694 , n77696 );
and ( n77698 , n77692 , n77697 );
buf ( n77699 , n20830 );
and ( n77700 , n69059 , n69204 );
not ( n77701 , n77700 );
and ( n77702 , n69303 , n68752 );
not ( n77703 , n77702 );
and ( n77704 , n77701 , n77703 );
and ( n77705 , n77699 , n77704 );
and ( n77706 , n55756 , n57187 );
and ( n77707 , n55497 , n57184 );
nor ( n77708 , n77706 , n77707 );
xnor ( n77709 , n77708 , n56175 );
and ( n77710 , n56388 , n56503 );
and ( n77711 , n56255 , n56501 );
nor ( n77712 , n77710 , n77711 );
xnor ( n77713 , n77712 , n56178 );
and ( n77714 , n77709 , n77713 );
and ( n77715 , n57063 , n55851 );
and ( n77716 , n56915 , n55849 );
nor ( n77717 , n77715 , n77716 );
xnor ( n77718 , n77717 , n55506 );
and ( n77719 , n77713 , n77718 );
and ( n77720 , n77709 , n77718 );
or ( n77721 , n77714 , n77719 , n77720 );
and ( n77722 , n77704 , n77721 );
and ( n77723 , n77699 , n77721 );
or ( n77724 , n77705 , n77722 , n77723 );
and ( n77725 , n77697 , n77724 );
and ( n77726 , n77692 , n77724 );
or ( n77727 , n77698 , n77725 , n77726 );
and ( n77728 , n77680 , n77727 );
and ( n77729 , n77672 , n77727 );
or ( n77730 , n77681 , n77728 , n77729 );
and ( n77731 , n77670 , n77730 );
and ( n77732 , n57063 , n55849 );
not ( n77733 , n77732 );
and ( n77734 , n77733 , n55506 );
xor ( n77735 , n45459 , n45496 );
buf ( n77736 , n77735 );
buf ( n77737 , n77736 );
buf ( n77738 , n77737 );
and ( n77739 , n77734 , n77738 );
buf ( n77740 , n20831 );
and ( n77741 , n77738 , n77740 );
and ( n77742 , n77734 , n77740 );
or ( n77743 , n77739 , n77741 , n77742 );
xor ( n77744 , n77602 , n77606 );
xor ( n77745 , n77744 , n77611 );
and ( n77746 , n77743 , n77745 );
xor ( n77747 , n77458 , n77618 );
xor ( n77748 , n77747 , n77621 );
and ( n77749 , n77745 , n77748 );
and ( n77750 , n77743 , n77748 );
or ( n77751 , n77746 , n77749 , n77750 );
xor ( n77752 , n77586 , n77587 );
xor ( n77753 , n77752 , n77589 );
and ( n77754 , n77751 , n77753 );
xor ( n77755 , n77614 , n77624 );
xor ( n77756 , n77755 , n77627 );
and ( n77757 , n77753 , n77756 );
and ( n77758 , n77751 , n77756 );
or ( n77759 , n77754 , n77757 , n77758 );
xor ( n77760 , n77552 , n77554 );
xor ( n77761 , n77760 , n77556 );
and ( n77762 , n77759 , n77761 );
xor ( n77763 , n77581 , n77584 );
xor ( n77764 , n77763 , n77592 );
and ( n77765 , n77761 , n77764 );
and ( n77766 , n77759 , n77764 );
or ( n77767 , n77762 , n77765 , n77766 );
and ( n77768 , n77730 , n77767 );
and ( n77769 , n77670 , n77767 );
or ( n77770 , n77731 , n77768 , n77769 );
and ( n77771 , n77668 , n77770 );
xor ( n77772 , n77598 , n77646 );
xor ( n77773 , n77772 , n77649 );
and ( n77774 , n77770 , n77773 );
and ( n77775 , n77668 , n77773 );
or ( n77776 , n77771 , n77774 , n77775 );
and ( n77777 , n77666 , n77776 );
xor ( n77778 , n77545 , n77547 );
xor ( n77779 , n77778 , n77652 );
and ( n77780 , n77776 , n77779 );
and ( n77781 , n77666 , n77779 );
or ( n77782 , n77777 , n77780 , n77781 );
xor ( n77783 , n77543 , n77655 );
xor ( n77784 , n77783 , n77658 );
and ( n77785 , n77782 , n77784 );
xor ( n77786 , n77666 , n77776 );
xor ( n77787 , n77786 , n77779 );
xor ( n77788 , n77550 , n77559 );
xor ( n77789 , n77788 , n77595 );
xor ( n77790 , n77638 , n77640 );
xor ( n77791 , n77790 , n77643 );
and ( n77792 , n77789 , n77791 );
xor ( n77793 , n77630 , n77632 );
xor ( n77794 , n77793 , n77635 );
xor ( n77795 , n77686 , n77691 );
xor ( n77796 , n77694 , n77696 );
and ( n77797 , n77795 , n77796 );
xor ( n77798 , n77683 , n77685 );
xor ( n77799 , n77688 , n77690 );
and ( n77800 , n77798 , n77799 );
and ( n77801 , n77796 , n77800 );
and ( n77802 , n77795 , n77800 );
or ( n77803 , n77797 , n77801 , n77802 );
xor ( n77804 , n77701 , n77703 );
and ( n77805 , n68307 , n70108 );
not ( n77806 , n77805 );
and ( n77807 , n70256 , n68610 );
not ( n77808 , n77807 );
and ( n77809 , n77806 , n77808 );
and ( n77810 , n77804 , n77809 );
and ( n77811 , n69059 , n69507 );
not ( n77812 , n77811 );
and ( n77813 , n69688 , n68752 );
not ( n77814 , n77813 );
and ( n77815 , n77812 , n77814 );
and ( n77816 , n77809 , n77815 );
and ( n77817 , n77804 , n77815 );
or ( n77818 , n77810 , n77816 , n77817 );
and ( n77819 , n56255 , n57187 );
and ( n77820 , n55756 , n57184 );
nor ( n77821 , n77819 , n77820 );
xnor ( n77822 , n77821 , n56175 );
and ( n77823 , n56915 , n56503 );
and ( n77824 , n56388 , n56501 );
nor ( n77825 , n77823 , n77824 );
xnor ( n77826 , n77825 , n56178 );
and ( n77827 , n77822 , n77826 );
and ( n77828 , n77826 , n77732 );
and ( n77829 , n77822 , n77732 );
or ( n77830 , n77827 , n77828 , n77829 );
xor ( n77831 , n45461 , n45495 );
buf ( n77832 , n77831 );
buf ( n77833 , n77832 );
buf ( n77834 , n77833 );
buf ( n77835 , n69303 );
not ( n77836 , n77835 );
and ( n77837 , n77834 , n77836 );
buf ( n77838 , n20832 );
and ( n77839 , n77836 , n77838 );
and ( n77840 , n77834 , n77838 );
or ( n77841 , n77837 , n77839 , n77840 );
and ( n77842 , n77830 , n77841 );
xor ( n77843 , n77709 , n77713 );
xor ( n77844 , n77843 , n77718 );
and ( n77845 , n77841 , n77844 );
and ( n77846 , n77830 , n77844 );
or ( n77847 , n77842 , n77845 , n77846 );
and ( n77848 , n77818 , n77847 );
xor ( n77849 , n77699 , n77704 );
xor ( n77850 , n77849 , n77721 );
and ( n77851 , n77847 , n77850 );
and ( n77852 , n77818 , n77850 );
or ( n77853 , n77848 , n77851 , n77852 );
and ( n77854 , n77803 , n77853 );
xor ( n77855 , n77674 , n77675 );
xor ( n77856 , n77855 , n77677 );
and ( n77857 , n77853 , n77856 );
and ( n77858 , n77803 , n77856 );
or ( n77859 , n77854 , n77857 , n77858 );
and ( n77860 , n77794 , n77859 );
xor ( n77861 , n77672 , n77680 );
xor ( n77862 , n77861 , n77727 );
and ( n77863 , n77859 , n77862 );
and ( n77864 , n77794 , n77862 );
or ( n77865 , n77860 , n77863 , n77864 );
and ( n77866 , n77791 , n77865 );
and ( n77867 , n77789 , n77865 );
or ( n77868 , n77792 , n77866 , n77867 );
xor ( n77869 , n77668 , n77770 );
xor ( n77870 , n77869 , n77773 );
and ( n77871 , n77868 , n77870 );
xor ( n77872 , n77670 , n77730 );
xor ( n77873 , n77872 , n77767 );
xor ( n77874 , n77759 , n77761 );
xor ( n77875 , n77874 , n77764 );
xor ( n77876 , n77692 , n77697 );
xor ( n77877 , n77876 , n77724 );
xor ( n77878 , n77751 , n77753 );
xor ( n77879 , n77878 , n77756 );
and ( n77880 , n77877 , n77879 );
xor ( n77881 , n77743 , n77745 );
xor ( n77882 , n77881 , n77748 );
xor ( n77883 , n77734 , n77738 );
xor ( n77884 , n77883 , n77740 );
xor ( n77885 , n77798 , n77799 );
and ( n77886 , n77884 , n77885 );
xor ( n77887 , n77806 , n77808 );
xor ( n77888 , n77812 , n77814 );
and ( n77889 , n77887 , n77888 );
and ( n77890 , n69059 , n70108 );
not ( n77891 , n77890 );
and ( n77892 , n70256 , n68752 );
not ( n77893 , n77892 );
and ( n77894 , n77891 , n77893 );
and ( n77895 , n77888 , n77894 );
and ( n77896 , n77887 , n77894 );
or ( n77897 , n77889 , n77895 , n77896 );
and ( n77898 , n77885 , n77897 );
and ( n77899 , n77884 , n77897 );
or ( n77900 , n77886 , n77898 , n77899 );
and ( n77901 , n77882 , n77900 );
and ( n77902 , n69303 , n69507 );
not ( n77903 , n77902 );
and ( n77904 , n69688 , n69204 );
not ( n77905 , n77904 );
and ( n77906 , n77903 , n77905 );
and ( n77907 , n56388 , n57187 );
and ( n77908 , n56255 , n57184 );
nor ( n77909 , n77907 , n77908 );
xnor ( n77910 , n77909 , n56175 );
and ( n77911 , n57063 , n56503 );
and ( n77912 , n56915 , n56501 );
nor ( n77913 , n77911 , n77912 );
xnor ( n77914 , n77913 , n56178 );
and ( n77915 , n77910 , n77914 );
and ( n77916 , n57063 , n56501 );
not ( n77917 , n77916 );
and ( n77918 , n77917 , n56178 );
and ( n77919 , n77914 , n77918 );
and ( n77920 , n77910 , n77918 );
or ( n77921 , n77915 , n77919 , n77920 );
and ( n77922 , n77906 , n77921 );
xor ( n77923 , n77822 , n77826 );
xor ( n77924 , n77923 , n77732 );
and ( n77925 , n77921 , n77924 );
and ( n77926 , n77906 , n77924 );
or ( n77927 , n77922 , n77925 , n77926 );
xor ( n77928 , n77804 , n77809 );
xor ( n77929 , n77928 , n77815 );
and ( n77930 , n77927 , n77929 );
xor ( n77931 , n77830 , n77841 );
xor ( n77932 , n77931 , n77844 );
and ( n77933 , n77929 , n77932 );
and ( n77934 , n77927 , n77932 );
or ( n77935 , n77930 , n77933 , n77934 );
and ( n77936 , n77900 , n77935 );
and ( n77937 , n77882 , n77935 );
or ( n77938 , n77901 , n77936 , n77937 );
and ( n77939 , n77879 , n77938 );
and ( n77940 , n77877 , n77938 );
or ( n77941 , n77880 , n77939 , n77940 );
and ( n77942 , n77875 , n77941 );
xor ( n77943 , n77794 , n77859 );
xor ( n77944 , n77943 , n77862 );
and ( n77945 , n77941 , n77944 );
and ( n77946 , n77875 , n77944 );
or ( n77947 , n77942 , n77945 , n77946 );
and ( n77948 , n77873 , n77947 );
xor ( n77949 , n77789 , n77791 );
xor ( n77950 , n77949 , n77865 );
and ( n77951 , n77947 , n77950 );
and ( n77952 , n77873 , n77950 );
or ( n77953 , n77948 , n77951 , n77952 );
and ( n77954 , n77870 , n77953 );
and ( n77955 , n77868 , n77953 );
or ( n77956 , n77871 , n77954 , n77955 );
or ( n77957 , n77787 , n77956 );
and ( n77958 , n77784 , n77957 );
and ( n77959 , n77782 , n77957 );
or ( n77960 , n77785 , n77958 , n77959 );
and ( n77961 , n77663 , n77960 );
and ( n77962 , n77661 , n77960 );
or ( n77963 , n77664 , n77961 , n77962 );
and ( n77964 , n77541 , n77963 );
xor ( n77965 , n77541 , n77963 );
xor ( n77966 , n77661 , n77663 );
xor ( n77967 , n77966 , n77960 );
xor ( n77968 , n77782 , n77784 );
xor ( n77969 , n77968 , n77957 );
xnor ( n77970 , n77787 , n77956 );
xor ( n77971 , n77868 , n77870 );
xor ( n77972 , n77971 , n77953 );
xor ( n77973 , n77873 , n77947 );
xor ( n77974 , n77973 , n77950 );
xor ( n77975 , n77803 , n77853 );
xor ( n77976 , n77975 , n77856 );
xor ( n77977 , n77795 , n77796 );
xor ( n77978 , n77977 , n77800 );
xor ( n77979 , n77818 , n77847 );
xor ( n77980 , n77979 , n77850 );
and ( n77981 , n77978 , n77980 );
xor ( n77982 , n77834 , n77836 );
xor ( n77983 , n77982 , n77838 );
xor ( n77984 , n45477 , n45493 );
buf ( n77985 , n77984 );
buf ( n77986 , n77985 );
buf ( n77987 , n77986 );
buf ( n77988 , n77987 );
xor ( n77989 , n77891 , n77893 );
buf ( n77990 , n77989 );
and ( n77991 , n77987 , n77989 );
or ( n77992 , n77988 , n77990 , n77991 );
and ( n77993 , n77983 , n77992 );
xor ( n77994 , n77903 , n77905 );
and ( n77995 , n69303 , n70108 );
not ( n77996 , n77995 );
and ( n77997 , n70256 , n69204 );
not ( n77998 , n77997 );
and ( n77999 , n77996 , n77998 );
and ( n78000 , n77994 , n77999 );
and ( n78001 , n56915 , n57187 );
and ( n78002 , n56388 , n57184 );
nor ( n78003 , n78001 , n78002 );
xnor ( n78004 , n78003 , n56175 );
and ( n78005 , n78004 , n77916 );
xor ( n78006 , n45479 , n45492 );
buf ( n78007 , n78006 );
buf ( n78008 , n78007 );
buf ( n78009 , n78008 );
and ( n78010 , n77916 , n78009 );
and ( n78011 , n78004 , n78009 );
or ( n78012 , n78005 , n78010 , n78011 );
and ( n78013 , n77999 , n78012 );
and ( n78014 , n77994 , n78012 );
or ( n78015 , n78000 , n78013 , n78014 );
and ( n78016 , n77992 , n78015 );
and ( n78017 , n77983 , n78015 );
or ( n78018 , n77993 , n78016 , n78017 );
xor ( n78019 , n77884 , n77885 );
xor ( n78020 , n78019 , n77897 );
and ( n78021 , n78018 , n78020 );
xor ( n78022 , n77927 , n77929 );
xor ( n78023 , n78022 , n77932 );
and ( n78024 , n78020 , n78023 );
and ( n78025 , n78018 , n78023 );
or ( n78026 , n78021 , n78024 , n78025 );
and ( n78027 , n77980 , n78026 );
and ( n78028 , n77978 , n78026 );
or ( n78029 , n77981 , n78027 , n78028 );
and ( n78030 , n77976 , n78029 );
xor ( n78031 , n77877 , n77879 );
xor ( n78032 , n78031 , n77938 );
and ( n78033 , n78029 , n78032 );
and ( n78034 , n77976 , n78032 );
or ( n78035 , n78030 , n78033 , n78034 );
xor ( n78036 , n77875 , n77941 );
xor ( n78037 , n78036 , n77944 );
and ( n78038 , n78035 , n78037 );
xor ( n78039 , n77976 , n78029 );
xor ( n78040 , n78039 , n78032 );
xor ( n78041 , n77882 , n77900 );
xor ( n78042 , n78041 , n77935 );
xor ( n78043 , n77978 , n77980 );
xor ( n78044 , n78043 , n78026 );
and ( n78045 , n78042 , n78044 );
xor ( n78046 , n77887 , n77888 );
xor ( n78047 , n78046 , n77894 );
xor ( n78048 , n77906 , n77921 );
xor ( n78049 , n78048 , n77924 );
and ( n78050 , n78047 , n78049 );
xor ( n78051 , n77910 , n77914 );
xor ( n78052 , n78051 , n77918 );
buf ( n78053 , n69688 );
not ( n78054 , n78053 );
xor ( n78055 , n77996 , n77998 );
and ( n78056 , n78054 , n78055 );
buf ( n78057 , n78056 );
and ( n78058 , n78052 , n78057 );
and ( n78059 , n69688 , n70108 );
not ( n78060 , n78059 );
and ( n78061 , n70256 , n69507 );
not ( n78062 , n78061 );
and ( n78063 , n78060 , n78062 );
and ( n78064 , n57063 , n57187 );
and ( n78065 , n56915 , n57184 );
nor ( n78066 , n78064 , n78065 );
xnor ( n78067 , n78066 , n56175 );
and ( n78068 , n57063 , n57184 );
not ( n78069 , n78068 );
and ( n78070 , n78069 , n56175 );
and ( n78071 , n78067 , n78070 );
xor ( n78072 , n45488 , n45490 );
buf ( n78073 , n78072 );
buf ( n78074 , n78073 );
buf ( n78075 , n78074 );
and ( n78076 , n78070 , n78075 );
and ( n78077 , n78067 , n78075 );
or ( n78078 , n78071 , n78076 , n78077 );
and ( n78079 , n78063 , n78078 );
xor ( n78080 , n78004 , n77916 );
xor ( n78081 , n78080 , n78009 );
and ( n78082 , n78078 , n78081 );
and ( n78083 , n78063 , n78081 );
or ( n78084 , n78079 , n78082 , n78083 );
and ( n78085 , n78057 , n78084 );
and ( n78086 , n78052 , n78084 );
or ( n78087 , n78058 , n78085 , n78086 );
and ( n78088 , n78049 , n78087 );
and ( n78089 , n78047 , n78087 );
or ( n78090 , n78050 , n78088 , n78089 );
xor ( n78091 , n78018 , n78020 );
xor ( n78092 , n78091 , n78023 );
and ( n78093 , n78090 , n78092 );
xor ( n78094 , n77983 , n77992 );
xor ( n78095 , n78094 , n78015 );
not ( n78096 , n77987 );
xor ( n78097 , n78096 , n77989 );
xor ( n78098 , n77994 , n77999 );
xor ( n78099 , n78098 , n78012 );
and ( n78100 , n78097 , n78099 );
xor ( n78101 , n78060 , n78062 );
xor ( n78102 , n45489 , n45484 );
buf ( n78103 , n78102 );
buf ( n78104 , n78103 );
buf ( n78105 , n78104 );
and ( n78106 , n78068 , n78105 );
buf ( n78107 , n70256 );
not ( n78108 , n78107 );
and ( n78109 , n78105 , n78108 );
and ( n78110 , n78068 , n78108 );
or ( n78111 , n78106 , n78109 , n78110 );
and ( n78112 , n78101 , n78111 );
buf ( n78113 , n78112 );
buf ( n78114 , n78054 );
xor ( n78115 , n78114 , n78055 );
and ( n78116 , n78113 , n78115 );
xor ( n78117 , n78063 , n78078 );
xor ( n78118 , n78117 , n78081 );
and ( n78119 , n78115 , n78118 );
and ( n78120 , n78113 , n78118 );
or ( n78121 , n78116 , n78119 , n78120 );
and ( n78122 , n78099 , n78121 );
and ( n78123 , n78097 , n78121 );
or ( n78124 , n78100 , n78122 , n78123 );
and ( n78125 , n78095 , n78124 );
xor ( n78126 , n78047 , n78049 );
xor ( n78127 , n78126 , n78087 );
and ( n78128 , n78124 , n78127 );
and ( n78129 , n78095 , n78127 );
or ( n78130 , n78125 , n78128 , n78129 );
and ( n78131 , n78092 , n78130 );
and ( n78132 , n78090 , n78130 );
or ( n78133 , n78093 , n78131 , n78132 );
and ( n78134 , n78044 , n78133 );
and ( n78135 , n78042 , n78133 );
or ( n78136 , n78045 , n78134 , n78135 );
and ( n78137 , n78040 , n78136 );
buf ( n78138 , n78136 );
buf ( n78139 , n78040 );
or ( n78140 , n78137 , n78138 , n78139 );
and ( n78141 , n78037 , n78140 );
and ( n78142 , n78035 , n78140 );
or ( n78143 , n78038 , n78141 , n78142 );
and ( n78144 , n77974 , n78143 );
xor ( n78145 , n77974 , n78143 );
xor ( n78146 , n78035 , n78037 );
xor ( n78147 , n78146 , n78140 );
not ( n78148 , n78147 );
xor ( n78149 , n78040 , n78136 );
not ( n78150 , n78149 );
not ( n78151 , n78150 );
xor ( n78152 , n78042 , n78044 );
xor ( n78153 , n78152 , n78133 );
buf ( n78154 , n78153 );
xor ( n78155 , n78090 , n78092 );
xor ( n78156 , n78155 , n78130 );
buf ( n78157 , n78156 );
xor ( n78158 , n78095 , n78124 );
xor ( n78159 , n78158 , n78127 );
buf ( n78160 , n78159 );
xor ( n78161 , n78097 , n78099 );
xor ( n78162 , n78161 , n78121 );
xor ( n78163 , n78052 , n78057 );
xor ( n78164 , n78163 , n78084 );
buf ( n78165 , n78164 );
and ( n78166 , n78162 , n78165 );
xor ( n78167 , n78162 , n78165 );
xor ( n78168 , n78113 , n78115 );
xor ( n78169 , n78168 , n78118 );
buf ( n78170 , n78169 );
buf ( n78171 , n78101 );
xor ( n78172 , n78171 , n78111 );
xor ( n78173 , n78067 , n78070 );
xor ( n78174 , n78173 , n78075 );
buf ( n78175 , n78174 );
and ( n78176 , n78172 , n78175 );
and ( n78177 , n78170 , n78176 );
and ( n78178 , n78167 , n78177 );
or ( n78179 , n78166 , n78178 );
and ( n78180 , n78160 , n78179 );
and ( n78181 , n78157 , n78180 );
and ( n78182 , n78154 , n78181 );
and ( n78183 , n78151 , n78182 );
or ( n78184 , n78150 , n78183 );
and ( n78185 , n78148 , n78184 );
or ( n78186 , n78147 , n78185 );
and ( n78187 , n78145 , n78186 );
or ( n78188 , n78144 , n78187 );
and ( n78189 , n77972 , n78188 );
and ( n78190 , n77970 , n78189 );
and ( n78191 , n77969 , n78190 );
and ( n78192 , n77967 , n78191 );
and ( n78193 , n77965 , n78192 );
or ( n78194 , n77964 , n78193 );
and ( n78195 , n77539 , n78194 );
and ( n78196 , n77538 , n78195 );
and ( n78197 , n77537 , n78196 );
and ( n78198 , n77535 , n78197 );
and ( n78199 , n77534 , n78198 );
or ( n78200 , n77533 , n78199 );
and ( n78201 , n77210 , n78200 );
and ( n78202 , n77208 , n78201 );
and ( n78203 , n77207 , n78202 );
and ( n78204 , n77205 , n78203 );
or ( n78205 , n77204 , n78204 );
and ( n78206 , n77202 , n78205 );
or ( n78207 , n77201 , n78206 );
and ( n78208 , n75943 , n78207 );
or ( n78209 , n75942 , n78208 );
and ( n78210 , n75403 , n78209 );
or ( n78211 , n75402 , n78210 );
and ( n78212 , n75398 , n78211 );
or ( n78213 , n75397 , n78212 );
and ( n78214 , n75127 , n78213 );
or ( n78215 , n75126 , n78214 );
and ( n78216 , n74518 , n78215 );
and ( n78217 , n74516 , n78216 );
or ( n78218 , n74515 , n78217 );
and ( n78219 , n74513 , n78218 );
or ( n78220 , n74512 , n78219 );
and ( n78221 , n73854 , n78220 );
and ( n78222 , n73852 , n78221 );
and ( n78223 , n73850 , n78222 );
or ( n78224 , n73849 , n78223 );
and ( n78225 , n73847 , n78224 );
and ( n78226 , n73845 , n78225 );
and ( n78227 , n73844 , n78226 );
and ( n78228 , n73842 , n78227 );
and ( n78229 , n73840 , n78228 );
and ( n78230 , n73838 , n78229 );
or ( n78231 , n73837 , n78230 );
and ( n78232 , n70382 , n78231 );
and ( n78233 , n70380 , n78232 );
or ( n78234 , n70379 , n78233 );
and ( n78235 , n70377 , n78234 );
or ( n78236 , n70376 , n78235 );
and ( n78237 , n69049 , n78236 );
or ( n78238 , n69048 , n78237 );
and ( n78239 , n68590 , n78238 );
or ( n78240 , n68589 , n78239 );
and ( n78241 , n68177 , n78240 );
and ( n78242 , n68176 , n78241 );
or ( n78243 , n68175 , n78242 );
and ( n78244 , n68173 , n78243 );
and ( n78245 , n68172 , n78244 );
or ( n78246 , n68171 , n78245 );
and ( n78247 , n68169 , n78246 );
or ( n78248 , n68168 , n78247 );
and ( n78249 , n66383 , n78248 );
or ( n78250 , n66382 , n78249 );
and ( n78251 , n66380 , n78250 );
and ( n78252 , n66378 , n78251 );
and ( n78253 , n66376 , n78252 );
and ( n78254 , n66375 , n78253 );
and ( n78255 , n66374 , n78254 );
or ( n78256 , n66373 , n78255 );
and ( n78257 , n66371 , n78256 );
or ( n78258 , n66370 , n78257 );
and ( n78259 , n66368 , n78258 );
or ( n78260 , n66367 , n78259 );
and ( n78261 , n62836 , n78260 );
or ( n78262 , n62835 , n78261 );
and ( n78263 , n62833 , n78262 );
and ( n78264 , n62832 , n78263 );
or ( n78265 , n62831 , n78264 );
and ( n78266 , n61730 , n78265 );
or ( n78267 , n61729 , n78266 );
and ( n78268 , n61727 , n78267 );
or ( n78269 , n61726 , n78268 );
and ( n78270 , n61724 , n78269 );
and ( n78271 , n61723 , n78270 );
or ( n78272 , n61722 , n78271 );
and ( n78273 , n61720 , n78272 );
and ( n78274 , n61718 , n78273 );
or ( n78275 , n61717 , n78274 );
and ( n78276 , n59479 , n78275 );
or ( n78277 , n59478 , n78276 );
and ( n78278 , n58698 , n78277 );
or ( n78279 , n58697 , n78278 );
and ( n78280 , n58695 , n78279 );
or ( n78281 , n58694 , n78280 );
and ( n78282 , n58028 , n78281 );
and ( n78283 , n58027 , n78282 );
or ( n78284 , n58026 , n78283 );
and ( n78285 , n58024 , n78284 );
or ( n78286 , n58023 , n78285 );
and ( n78287 , n57027 , n78286 );
or ( n78288 , n57026 , n78287 );
and ( n78289 , n56704 , n78288 );
and ( n78290 , n56703 , n78289 );
and ( n78291 , n56701 , n78290 );
or ( n78292 , n56700 , n78291 );
and ( n78293 , n56698 , n78292 );
and ( n78294 , n56697 , n78293 );
or ( n78295 , n56696 , n78294 );
and ( n78296 , n55370 , n78295 );
and ( n78297 , n55369 , n78296 );
and ( n78298 , n55368 , n78297 );
or ( n78299 , n55367 , n78298 );
and ( n78300 , n54703 , n78299 );
or ( n78301 , n54702 , n78300 );
and ( n78302 , n54700 , n78301 );
and ( n78303 , n54698 , n78302 );
and ( n78304 , n54697 , n78303 );
or ( n78305 , n54696 , n78304 );
and ( n78306 , n53239 , n78305 );
or ( n78307 , n53238 , n78306 );
and ( n78308 , n52417 , n78307 );
or ( n78309 , n52416 , n78308 );
and ( n78310 , n52170 , n78309 );
or ( n78311 , n52169 , n78310 );
and ( n78312 , n51904 , n78311 );
and ( n78313 , n51903 , n78312 );
and ( n78314 , n51902 , n78313 );
or ( n78315 , n51901 , n78314 );
and ( n78316 , n51411 , n78315 );
and ( n78317 , n51409 , n78316 );
or ( n78318 , n51408 , n78317 );
and ( n78319 , n51406 , n78318 );
and ( n78320 , n51404 , n78319 );
or ( n78321 , n51403 , n78320 );
and ( n78322 , n51401 , n78321 );
and ( n78323 , n51400 , n78322 );
or ( n78324 , n51399 , n78323 );
and ( n78325 , n51397 , n78324 );
or ( n78326 , n51396 , n78325 );
and ( n78327 , n49629 , n78326 );
or ( n78328 , n49628 , n78327 );
and ( n78329 , n49244 , n78328 );
or ( n78330 , n49243 , n78329 );
and ( n78331 , n49241 , n78330 );
or ( n78332 , n49240 , n78331 );
and ( n78333 , n48869 , n78332 );
or ( n78334 , n48868 , n78333 );
and ( n78335 , n48866 , n78334 );
or ( n78336 , n48865 , n78335 );
and ( n78337 , n48511 , n78336 );
and ( n78338 , n48510 , n78337 );
and ( n78339 , n48509 , n78338 );
and ( n78340 , n48507 , n78339 );
or ( n78341 , n48506 , n78340 );
and ( n78342 , n47910 , n78341 );
or ( n78343 , n47909 , n78342 );
and ( n78344 , n47907 , n78343 );
or ( n78345 , n47906 , n78344 );
and ( n78346 , n47525 , n78345 );
and ( n78347 , n47523 , n78346 );
and ( n78348 , n47522 , n78347 );
and ( n78349 , n47520 , n78348 );
or ( n78350 , n47519 , n78349 );
and ( n78351 , n47517 , n78350 );
or ( n78352 , n47516 , n78351 );
and ( n78353 , n46891 , n78352 );
and ( n78354 , n46890 , n78353 );
or ( n78355 , n46889 , n78354 );
and ( n78356 , n46668 , n78355 );
and ( n78357 , n46667 , n78356 );
or ( n78358 , n46666 , n78357 );
and ( n78359 , n46387 , n78358 );
and ( n78360 , n46386 , n78359 );
or ( n78361 , n46385 , n78360 );
and ( n78362 , n46212 , n78361 );
and ( n78363 , n46211 , n78362 );
or ( n78364 , n46210 , n78363 );
and ( n78365 , n46026 , n78364 );
and ( n78366 , n46025 , n78365 );
or ( n78367 , n46024 , n78366 );
and ( n78368 , n45876 , n78367 );
xor ( n78369 , n45875 , n78368 );
buf ( n78370 , n78369 );
xor ( n78371 , n45876 , n78367 );
buf ( n78372 , n78371 );
xor ( n78373 , n46025 , n78365 );
buf ( n78374 , n78373 );
xor ( n78375 , n46026 , n78364 );
buf ( n78376 , n78375 );
xor ( n78377 , n46211 , n78362 );
buf ( n78378 , n78377 );
xor ( n78379 , n46212 , n78361 );
buf ( n78380 , n78379 );
xor ( n78381 , n46386 , n78359 );
buf ( n78382 , n78381 );
xor ( n78383 , n46387 , n78358 );
buf ( n78384 , n78383 );
xor ( n78385 , n46667 , n78356 );
buf ( n78386 , n78385 );
xor ( n78387 , n46668 , n78355 );
buf ( n78388 , n78387 );
xor ( n78389 , n46890 , n78353 );
buf ( n78390 , n78389 );
xor ( n78391 , n46891 , n78352 );
buf ( n78392 , n78391 );
xor ( n78393 , n47517 , n78350 );
buf ( n78394 , n78393 );
xor ( n78395 , n47520 , n78348 );
buf ( n78396 , n78395 );
xor ( n78397 , n47522 , n78347 );
buf ( n78398 , n78397 );
xor ( n78399 , n47523 , n78346 );
buf ( n78400 , n78399 );
xor ( n78401 , n47525 , n78345 );
buf ( n78402 , n78401 );
xor ( n78403 , n47907 , n78343 );
buf ( n78404 , n78403 );
xor ( n78405 , n47910 , n78341 );
buf ( n78406 , n78405 );
xor ( n78407 , n48507 , n78339 );
buf ( n78408 , n78407 );
xor ( n78409 , n48509 , n78338 );
buf ( n78410 , n78409 );
xor ( n78411 , n48510 , n78337 );
buf ( n78412 , n78411 );
xor ( n78413 , n48511 , n78336 );
buf ( n78414 , n78413 );
xor ( n78415 , n48866 , n78334 );
buf ( n78416 , n78415 );
xor ( n78417 , n48869 , n78332 );
buf ( n78418 , n78417 );
xor ( n78419 , n49241 , n78330 );
buf ( n78420 , n78419 );
xor ( n78421 , n49244 , n78328 );
buf ( n78422 , n78421 );
xor ( n78423 , n49629 , n78326 );
buf ( n78424 , n78423 );
xor ( n78425 , n51397 , n78324 );
buf ( n78426 , n78425 );
xor ( n78427 , n51400 , n78322 );
buf ( n78428 , n78427 );
xor ( n78429 , n51401 , n78321 );
buf ( n78430 , n78429 );
xor ( n78431 , n51404 , n78319 );
buf ( n78432 , n78431 );
xor ( n78433 , n51406 , n78318 );
buf ( n78434 , n78433 );
xor ( n78435 , n51409 , n78316 );
buf ( n78436 , n78435 );
xor ( n78437 , n51411 , n78315 );
buf ( n78438 , n78437 );
xor ( n78439 , n51902 , n78313 );
buf ( n78440 , n78439 );
xor ( n78441 , n51903 , n78312 );
buf ( n78442 , n78441 );
xor ( n78443 , n51904 , n78311 );
buf ( n78444 , n78443 );
xor ( n78445 , n52170 , n78309 );
buf ( n78446 , n78445 );
xor ( n78447 , n52417 , n78307 );
buf ( n78448 , n78447 );
xor ( n78449 , n53239 , n78305 );
buf ( n78450 , n78449 );
xor ( n78451 , n54697 , n78303 );
buf ( n78452 , n78451 );
xor ( n78453 , n54698 , n78302 );
buf ( n78454 , n78453 );
xor ( n78455 , n54700 , n78301 );
buf ( n78456 , n78455 );
xor ( n78457 , n54703 , n78299 );
buf ( n78458 , n78457 );
xor ( n78459 , n55368 , n78297 );
buf ( n78460 , n78459 );
xor ( n78461 , n55369 , n78296 );
buf ( n78462 , n78461 );
xor ( n78463 , n55370 , n78295 );
buf ( n78464 , n78463 );
xor ( n78465 , n56697 , n78293 );
buf ( n78466 , n78465 );
xor ( n78467 , n56698 , n78292 );
buf ( n78468 , n78467 );
xor ( n78469 , n56701 , n78290 );
buf ( n78470 , n78469 );
xor ( n78471 , n56703 , n78289 );
buf ( n78472 , n78471 );
xor ( n78473 , n56704 , n78288 );
buf ( n78474 , n78473 );
xor ( n78475 , n57027 , n78286 );
buf ( n78476 , n78475 );
xor ( n78477 , n58024 , n78284 );
buf ( n78478 , n78477 );
xor ( n78479 , n58027 , n78282 );
buf ( n78480 , n78479 );
xor ( n78481 , n58028 , n78281 );
buf ( n78482 , n78481 );
xor ( n78483 , n58695 , n78279 );
buf ( n78484 , n78483 );
xor ( n78485 , n58698 , n78277 );
buf ( n78486 , n78485 );
xor ( n78487 , n59479 , n78275 );
buf ( n78488 , n78487 );
xor ( n78489 , n61718 , n78273 );
buf ( n78490 , n78489 );
xor ( n78491 , n61720 , n78272 );
buf ( n78492 , n78491 );
xor ( n78493 , n61723 , n78270 );
buf ( n78494 , n78493 );
xor ( n78495 , n61724 , n78269 );
buf ( n78496 , n78495 );
xor ( n78497 , n61727 , n78267 );
buf ( n78498 , n78497 );
xor ( n78499 , n61730 , n78265 );
buf ( n78500 , n78499 );
xor ( n78501 , n62832 , n78263 );
buf ( n78502 , n78501 );
xor ( n78503 , n62833 , n78262 );
buf ( n78504 , n78503 );
xor ( n78505 , n62836 , n78260 );
buf ( n78506 , n78505 );
xor ( n78507 , n66368 , n78258 );
buf ( n78508 , n78507 );
xor ( n78509 , n66371 , n78256 );
buf ( n78510 , n78509 );
xor ( n78511 , n66374 , n78254 );
buf ( n78512 , n78511 );
xor ( n78513 , n66375 , n78253 );
buf ( n78514 , n78513 );
xor ( n78515 , n66376 , n78252 );
buf ( n78516 , n78515 );
xor ( n78517 , n66378 , n78251 );
buf ( n78518 , n78517 );
xor ( n78519 , n66380 , n78250 );
buf ( n78520 , n78519 );
xor ( n78521 , n66383 , n78248 );
buf ( n78522 , n78521 );
xor ( n78523 , n68169 , n78246 );
buf ( n78524 , n78523 );
xor ( n78525 , n68172 , n78244 );
buf ( n78526 , n78525 );
xor ( n78527 , n68173 , n78243 );
buf ( n78528 , n78527 );
xor ( n78529 , n68176 , n78241 );
buf ( n78530 , n78529 );
xor ( n78531 , n68177 , n78240 );
buf ( n78532 , n78531 );
xor ( n78533 , n68590 , n78238 );
buf ( n78534 , n78533 );
xor ( n78535 , n69049 , n78236 );
buf ( n78536 , n78535 );
xor ( n78537 , n70377 , n78234 );
buf ( n78538 , n78537 );
xor ( n78539 , n70380 , n78232 );
buf ( n78540 , n78539 );
xor ( n78541 , n70382 , n78231 );
buf ( n78542 , n78541 );
xor ( n78543 , n73838 , n78229 );
buf ( n78544 , n78543 );
xor ( n78545 , n73840 , n78228 );
buf ( n78546 , n78545 );
xor ( n78547 , n73842 , n78227 );
buf ( n78548 , n78547 );
xor ( n78549 , n73844 , n78226 );
buf ( n78550 , n78549 );
xor ( n78551 , n73845 , n78225 );
buf ( n78552 , n78551 );
xor ( n78553 , n73847 , n78224 );
buf ( n78554 , n78553 );
xor ( n78555 , n73850 , n78222 );
buf ( n78556 , n78555 );
xor ( n78557 , n73852 , n78221 );
buf ( n78558 , n78557 );
xor ( n78559 , n73854 , n78220 );
buf ( n78560 , n78559 );
xor ( n78561 , n74513 , n78218 );
buf ( n78562 , n78561 );
xor ( n78563 , n74516 , n78216 );
buf ( n78564 , n78563 );
xor ( n78565 , n74518 , n78215 );
buf ( n78566 , n78565 );
xor ( n78567 , n75127 , n78213 );
buf ( n78568 , n78567 );
xor ( n78569 , n75398 , n78211 );
buf ( n78570 , n78569 );
xor ( n78571 , n75403 , n78209 );
buf ( n78572 , n78571 );
xor ( n78573 , n75943 , n78207 );
buf ( n78574 , n78573 );
xor ( n78575 , n77202 , n78205 );
buf ( n78576 , n78575 );
xor ( n78577 , n77205 , n78203 );
buf ( n78578 , n78577 );
xor ( n78579 , n77207 , n78202 );
buf ( n78580 , n78579 );
xor ( n78581 , n77208 , n78201 );
buf ( n78582 , n78581 );
xor ( n78583 , n77210 , n78200 );
buf ( n78584 , n78583 );
xor ( n78585 , n77534 , n78198 );
buf ( n78586 , n78585 );
xor ( n78587 , n77535 , n78197 );
buf ( n78588 , n78587 );
xor ( n78589 , n77537 , n78196 );
buf ( n78590 , n78589 );
xor ( n78591 , n77538 , n78195 );
buf ( n78592 , n78591 );
xor ( n78593 , n77539 , n78194 );
buf ( n78594 , n78593 );
xor ( n78595 , n77965 , n78192 );
buf ( n78596 , n78595 );
xor ( n78597 , n77967 , n78191 );
buf ( n78598 , n78597 );
xor ( n78599 , n77969 , n78190 );
buf ( n78600 , n78599 );
xor ( n78601 , n77970 , n78189 );
buf ( n78602 , n78601 );
xor ( n78603 , n77972 , n78188 );
buf ( n78604 , n78603 );
xor ( n78605 , n78145 , n78186 );
buf ( n78606 , n78605 );
xor ( n78607 , n78148 , n78184 );
buf ( n78608 , n78607 );
xor ( n78609 , n78151 , n78182 );
buf ( n78610 , n78609 );
xor ( n78611 , n78154 , n78181 );
buf ( n78612 , n78611 );
xor ( n78613 , n78157 , n78180 );
buf ( n78614 , n78613 );
xor ( n78615 , n78160 , n78179 );
buf ( n78616 , n78615 );
xor ( n78617 , n78167 , n78177 );
buf ( n78618 , n78617 );
xor ( n78619 , n78170 , n78176 );
buf ( n78620 , n78619 );
xor ( n78621 , n78172 , n78175 );
buf ( n78622 , n78621 );
xor ( n78623 , n78068 , n78105 );
xor ( n78624 , n78623 , n78108 );
buf ( n78625 , n78624 );
buf ( n78626 , n78625 );
not ( C0n , n0 );
and ( C0 , C0n , n0 );
endmodule
