//NOTE: no-implementation module stub

module dmux (
    input wire SYSCLK,
    input wire TMODE,
    input wire SEN,
    input wire RESET_D1_R_N,
    input wire CLMI_RHOLD,
    input wire REGA_S,
    input wire REGB_S,
    input wire IMMED_S,
    input wire SELA_S,
    input wire SELBR_S,
    input wire SELBI_S,
    input wire ALURES_E,
    input wire SELC_M,
    input wire RDBUSINM,
    input wire REGC_W_R,
    input wire REGA_E_R,
    input wire REGBI_E_R,
    input wire REGBR_E_R,
    input wire CP0_PCREL_S,
    input wire CINA_E_R,
    input wire CINBI_E_R,
    input wire Z_E
);

endmodule
