// IWLS benchmark module "i8" printed on Wed May 29 17:27:06 2002
module i8(\V133(3) , \V133(1) , \V133(2) , \V133(0) , \V133(5) , \V133(10) , \V133(6) , \V133(7) , \V133(8) , \V47(31) , \V47(30) , \V47(29) , \V47(28) , \V47(27) , \V47(26) , \V47(25) , \V47(24) , \V47(23) , \V47(22) , \V47(21) , \V47(20) , \V47(19) , \V47(18) , \V47(17) , \V47(16) , \V47(15) , \V47(14) , \V47(13) , \V47(12) , \V47(11) , \V47(10) , \V47(9) , \V47(8) , \V47(7) , \V47(6) , \V47(5) , \V47(4) , \V47(3) , \V47(2) , \V47(1) , \V47(0) , \V84(11) , \V84(10) , \V84(9) , \V84(8) , \V84(7) , \V84(6) , \V84(5) , \V84(4) , \V84(3) , \V84(2) , \V84(1) , \V15(14) , \V15(13) , \V15(12) , \V15(11) , \V15(10) , \V15(9) , \V15(8) , \V15(7) , \V15(6) , \V15(5) , \V15(4) , \V15(3) , \V15(2) , \V15(1) , \V15(0) , \V84(31) , \V84(30) , \V84(29) , \V84(28) , \V84(27) , \V84(26) , \V84(25) , \V84(24) , \V84(23) , \V84(22) , \V84(21) , \V84(20) , \V84(19) , \V84(18) , \V84(17) , \V84(16) , \V84(15) , \V84(14) , \V84(13) , \V84(12) , \V84(0) , \V48(0) , \V49(0) , \V116(0) , \V50(0) , \V52(0) , \V51(0) , \V116(2) , \V133(9) , \V116(1) , \V116(8) , \V116(7) , \V116(6) , \V116(5) , \V116(4) , \V116(3) , \V116(9) , \V116(11) , \V116(10) , \V116(12) , \V116(15) , \V116(14) , \V116(13) , \V116(16) , \V116(31) , \V116(30) , \V116(29) , \V116(28) , \V116(27) , \V116(26) , \V116(25) , \V116(24) , \V116(23) , \V116(22) , \V116(21) , \V116(20) , \V116(19) , \V116(18) , \V116(17) , \V121(16) , \V119(0) , \V121(17) , \V122(0) , \V133(4) , \V118(0) , \V118(1) , \V134(0) , \V136(1) , \V136(0) , \V142(5) , \V142(4) , \V142(3) , \V142(2) , \V142(1) , \V142(0) , \V143(0) , \V145(1) , \V145(0) , \V146(0) , \V149(2) , \V149(1) , \V149(0) , \V150(0) , \V165(14) , \V165(13) , \V165(12) , \V165(11) , \V165(10) , \V165(9) , \V165(8) , \V165(7) , \V165(6) , \V165(5) , \V165(4) , \V165(3) , \V165(2) , \V165(1) , \V165(0) , \V197(31) , \V197(30) , \V197(29) , \V197(28) , \V197(27) , \V197(26) , \V197(25) , \V197(24) , \V197(23) , \V197(22) , \V197(21) , \V197(20) , \V197(19) , \V197(18) , \V197(17) , \V197(16) , \V197(15) , \V197(14) , \V197(13) , \V197(12) , \V197(11) , \V197(10) , \V197(9) , \V197(8) , \V197(7) , \V197(6) , \V197(5) , \V197(4) , \V197(3) , \V197(2) , \V197(1) , \V197(0) , \V212(14) , \V212(13) , \V212(12) , \V212(11) , \V212(10) , \V212(9) , \V212(8) , \V212(7) , \V212(6) , \V212(5) , \V212(4) , \V212(3) , \V212(2) , \V212(1) , \V212(0) , \V213(0) , \V214(0) );
input
  \V47(24) ,
  \V84(31) ,
  \V15(14) ,
  \V84(30) ,
  \V47(21) ,
  \V47(20) ,
  \V15(11) ,
  \V15(10) ,
  \V47(27) ,
  \V47(26) ,
  \V47(29) ,
  \V47(28) ,
  \V47(31) ,
  \V133(10) ,
  \V47(30) ,
  \V116(27) ,
  \V116(26) ,
  \V116(29) ,
  \V116(28) ,
  \V116(3) ,
  \V116(2) ,
  \V116(5) ,
  \V116(4) ,
  \V116(21) ,
  \V116(1) ,
  \V116(20) ,
  \V116(0) ,
  \V47(0) ,
  \V116(23) ,
  \V47(1) ,
  \V116(22) ,
  \V47(2) ,
  \V116(25) ,
  \V121(17) ,
  \V47(3) ,
  \V116(24) ,
  \V121(16) ,
  \V47(4) ,
  \V116(17) ,
  \V116(7) ,
  \V47(5) ,
  \V116(16) ,
  \V116(6) ,
  \V47(6) ,
  \V116(19) ,
  \V48(0) ,
  \V116(9) ,
  \V47(7) ,
  \V116(18) ,
  \V116(8) ,
  \V47(8) ,
  \V47(9) ,
  \V118(1) ,
  \V118(0) ,
  \V49(0) ,
  \V116(11) ,
  \V84(0) ,
  \V116(10) ,
  \V84(1) ,
  \V116(13) ,
  \V84(2) ,
  \V116(12) ,
  \V84(3) ,
  \V116(15) ,
  \V84(4) ,
  \V119(0) ,
  \V116(14) ,
  \V84(5) ,
  \V84(6) ,
  \V84(7) ,
  \V84(8) ,
  \V84(9) ,
  \V84(13) ,
  \V116(31) ,
  \V84(12) ,
  \V116(30) ,
  \V84(15) ,
  \V84(14) ,
  \V84(11) ,
  \V84(10) ,
  \V133(3) ,
  \V133(2) ,
  \V133(5) ,
  \V15(0) ,
  \V133(4) ,
  \V15(1) ,
  \V84(17) ,
  \V50(0) ,
  \V15(2) ,
  \V84(16) ,
  \V15(3) ,
  \V133(1) ,
  \V84(19) ,
  \V15(4) ,
  \V133(0) ,
  \V84(18) ,
  \V15(5) ,
  \V84(23) ,
  \V15(6) ,
  \V84(22) ,
  \V15(7) ,
  \V84(25) ,
  \V15(8) ,
  \V51(0) ,
  \V47(13) ,
  \V84(24) ,
  \V15(9) ,
  \V47(12) ,
  \V133(7) ,
  \V47(15) ,
  \V133(6) ,
  \V47(14) ,
  \V133(9) ,
  \V84(21) ,
  \V133(8) ,
  \V84(20) ,
  \V47(11) ,
  \V52(0) ,
  \V47(10) ,
  \V84(27) ,
  \V84(26) ,
  \V84(29) ,
  \V47(17) ,
  \V84(28) ,
  \V122(0) ,
  \V47(16) ,
  \V47(19) ,
  \V47(18) ,
  \V47(23) ,
  \V47(22) ,
  \V15(13) ,
  \V47(25) ,
  \V15(12) ;
output
  \V165(11) ,
  \V165(10) ,
  \V165(13) ,
  \V165(12) ,
  \V165(14) ,
  \V197(31) ,
  \V197(30) ,
  \V212(3) ,
  \V212(2) ,
  \V212(5) ,
  \V212(4) ,
  \V212(1) ,
  \V212(0) ,
  \V212(7) ,
  \V212(6) ,
  \V213(0) ,
  \V212(9) ,
  \V212(8) ,
  \V150(0) ,
  \V214(0) ,
  \V165(3) ,
  \V165(2) ,
  \V165(5) ,
  \V165(4) ,
  \V165(1) ,
  \V165(0) ,
  \V212(11) ,
  \V212(10) ,
  \V212(13) ,
  \V165(7) ,
  \V212(12) ,
  \V165(6) ,
  \V165(9) ,
  \V212(14) ,
  \V165(8) ,
  \V142(3) ,
  \V142(2) ,
  \V142(5) ,
  \V142(4) ,
  \V142(1) ,
  \V142(0) ,
  \V143(0) ,
  \V197(27) ,
  \V197(26) ,
  \V197(29) ,
  \V197(28) ,
  \V145(1) ,
  \V145(0) ,
  \V197(21) ,
  \V197(20) ,
  \V197(23) ,
  \V197(22) ,
  \V197(25) ,
  \V197(24) ,
  \V146(0) ,
  \V197(17) ,
  \V197(16) ,
  \V197(19) ,
  \V197(18) ,
  \V134(0) ,
  \V197(3) ,
  \V197(11) ,
  \V197(2) ,
  \V197(10) ,
  \V197(5) ,
  \V197(13) ,
  \V149(2) ,
  \V197(4) ,
  \V197(12) ,
  \V197(15) ,
  \V197(14) ,
  \V197(1) ,
  \V197(0) ,
  \V149(1) ,
  \V149(0) ,
  \V136(1) ,
  \V197(7) ,
  \V136(0) ,
  \V197(6) ,
  \V197(9) ,
  \V197(8) ;
wire
  \[60] ,
  V831,
  \[61] ,
  \[62] ,
  \[63] ,
  \[64] ,
  \[65] ,
  \[66] ,
  \[67] ,
  \[68] ,
  \[69] ,
  \[0] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  \[70] ,
  \[5] ,
  \[71] ,
  \[6] ,
  \[72] ,
  \[7] ,
  \[73] ,
  V967,
  \[8] ,
  \[74] ,
  \[9] ,
  \[75] ,
  \[76] ,
  \[77] ,
  \[78] ,
  \[79] ,
  \[80] ,
  \[82] ,
  \[83] ,
  \[84] ,
  \[85] ,
  \[86] ,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[90] ,
  \[14] ,
  \[91] ,
  \[15] ,
  \[92] ,
  \[16] ,
  \[93] ,
  \[17] ,
  \[94] ,
  \[18] ,
  \[95] ,
  \[19] ,
  \[96] ,
  \[97] ,
  \[98] ,
  \[100] ,
  \[99] ,
  \[101] ,
  V1117,
  \[104] ,
  \[20] ,
  \[105] ,
  \[21] ,
  \[106] ,
  \[22] ,
  V1146,
  \[23] ,
  V1153,
  \[108] ,
  \[24] ,
  \[109] ,
  \[25] ,
  \[26] ,
  \[27] ,
  \[28] ,
  \[29] ,
  \[110] ,
  \[111] ,
  \[112] ,
  \[113] ,
  \[114] ,
  \[30] ,
  \[31] ,
  \[32] ,
  V553,
  V554,
  \[117] ,
  \[33] ,
  V560,
  \[118] ,
  V569,
  \[34] ,
  \[119] ,
  \[35] ,
  \[36] ,
  \[37] ,
  \[38] ,
  \[39] ,
  \[120] ,
  \[121] ,
  \[122] ,
  \[123] ,
  V622,
  \[124] ,
  \[40] ,
  V631,
  \[125] ,
  \[41] ,
  \[126] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[129] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \[130] ,
  \[131] ,
  V715,
  \[134] ,
  \[50] ,
  V732,
  \[135] ,
  \[51] ,
  V749,
  \[52] ,
  \[53] ,
  V766,
  \[138] ,
  \[54] ,
  \[139] ,
  \[55] ,
  \[56] ,
  V799,
  \[57] ,
  \[58] ,
  \[59] ,
  \V235(2) ,
  \[140] ,
  \V235(1) ,
  \V235(0) ;
assign
  \[60]  = (\[94]  & (\[93]  & \V47(27) )) | ((\[93]  & (\[92]  & \V47(24) )) | ((\[93]  & (\[91]  & \V47(20) )) | ((\[93]  & (\V235(0)  & \V84(3) )) | ((\[97]  & \V116(3) ) | (\[93]  & V553))))),
  V831 = V715 & ~\V133(5) ,
  \[61]  = (\[94]  & (\[93]  & \V47(26) )) | ((\[93]  & (\[92]  & \V47(23) )) | ((\[93]  & (\[91]  & \V47(19) )) | ((\[93]  & (\V235(0)  & \V84(2) )) | ((\[97]  & \V116(2) ) | (\[93]  & V553))))),
  \V165(11)  = \[20] ,
  \[62]  = (\[94]  & (\[93]  & \V47(25) )) | ((\[93]  & (\[92]  & \V47(22) )) | ((\[93]  & (\[91]  & \V47(18) )) | ((\[93]  & (\V235(0)  & \V84(1) )) | ((\[97]  & \V116(1) ) | (\[93]  & V553))))),
  \V165(10)  = \[21] ,
  \[63]  = (\[94]  & (\[93]  & \V47(24) )) | ((\[93]  & (\[92]  & \V47(21) )) | ((\[93]  & (\[91]  & \V47(17) )) | ((\[93]  & (\V235(0)  & \V84(0) )) | ((\[97]  & \V116(0) ) | (\[93]  & V553))))),
  \V165(13)  = \[18] ,
  \[64]  = (\[114]  & \V116(14) ) | ((\[98]  & \V84(31) ) | V1117),
  \V165(12)  = \[19] ,
  \[65]  = (\[114]  & \V116(13) ) | ((\[98]  & \V84(30) ) | V1117),
  \[66]  = (\[114]  & \V116(12) ) | ((\[98]  & \V84(29) ) | V1117),
  \V165(14)  = \[17] ,
  \[67]  = (\[114]  & \V116(11) ) | ((\[98]  & \V84(28) ) | V1117),
  \[68]  = (\[114]  & \V116(10) ) | ((\[98]  & \V84(27) ) | V1117),
  \[69]  = (\[114]  & \V116(9) ) | ((\[98]  & \V84(26) ) | V1117),
  \[0]  = (\[131]  & (\[85]  & (~V554 & \V84(0) ))) | ((\[131]  & (\[85]  & (~V554 & ~\V133(10) ))) | ((\[85]  & (\V48(0)  & ~\V133(10) )) | ((V799 & \V116(0) ) | (V560 & \V49(0) )))),
  \[1]  = (\[129]  & (\[91]  & \V15(1) )) | ((\[129]  & (\V235(0)  & \V47(2) )) | ((\[117]  & (\[100]  & \V52(0) )) | ((\[134]  & \[129] ) | (V799 & \V116(2) )))),
  \[2]  = (\[138]  & (~V799 & \V50(0) )) | ((\[129]  & (\[91]  & \V15(0) )) | ((\[129]  & (\V235(0)  & \V47(1) )) | ((\[117]  & (\[100]  & \V51(0) )) | ((\[135]  & \[129] ) | (V799 & \V116(1) ))))),
  \[3]  = (\[140]  & \V47(0) ) | ((\[123]  & \V15(7) ) | ((\[121]  & \V116(8) ) | ((\[120]  & \V47(8) ) | ((\[119]  & \V84(8) ) | \[122] )))),
  \[4]  = (\[123]  & \V15(6) ) | ((\[121]  & \V116(7) ) | ((\[120]  & \V47(7) ) | ((\[119]  & \V84(7) ) | \[122] ))),
  \[70]  = (\[114]  & \V116(8) ) | ((\[98]  & \V84(25) ) | V1117),
  \V197(31)  = \[32] ,
  \[5]  = (\[123]  & \V15(5) ) | ((\[121]  & \V116(6) ) | ((\[120]  & \V47(6) ) | ((\[119]  & \V84(6) ) | \[122] ))),
  \[71]  = (\[114]  & \V116(7) ) | ((\[98]  & \V84(24) ) | V1117),
  \V197(30)  = \[33] ,
  \[6]  = (\[123]  & \V15(4) ) | ((\[121]  & \V116(5) ) | ((\[120]  & \V47(5) ) | ((\[119]  & \V84(5) ) | \[122] ))),
  \[72]  = (\[114]  & \V116(6) ) | ((\[98]  & \V84(23) ) | V1117),
  \[7]  = (\[123]  & \V15(3) ) | ((\[121]  & \V116(4) ) | ((\[120]  & \V47(4) ) | ((\[119]  & \V84(4) ) | \[122] ))),
  \[73]  = (\[114]  & \V116(5) ) | ((\[98]  & \V84(22) ) | V1117),
  \V212(3)  = \[75] ,
  V967 = V766 & ~\V133(1) ,
  \[8]  = (\[123]  & \V15(2) ) | ((\[121]  & \V116(3) ) | ((\[120]  & \V47(3) ) | ((\[119]  & \V84(3) ) | \[122] ))),
  \[74]  = (\[114]  & \V116(4) ) | ((\[98]  & \V84(21) ) | V1117),
  \V212(2)  = \[76] ,
  \[9]  = (\[94]  & (\[85]  & \V47(1) )) | ((\[94]  & (V622 & \V47(1) )) | ((\[91]  & (\[85]  & \V15(8) )) | ((\[91]  & (V622 & \V15(8) )) | ((\[85]  & (\V235(0)  & \V47(9) )) | ((V622 & (\V235(0)  & \V47(9) )) | ((\[126]  & \[85] ) | ((\[126]  & V622) | (\[118]  & \V116(9) )))))))),
  \[75]  = (\[114]  & \V116(3) ) | ((\[98]  & \V84(20) ) | V1117),
  \V212(5)  = \[73] ,
  \[76]  = (\[114]  & \V116(2) ) | ((\[98]  & \V84(19) ) | V1117),
  \V212(4)  = \[74] ,
  \[77]  = (\[114]  & \V116(1) ) | ((\[98]  & \V84(18) ) | V1117),
  \[78]  = (\[114]  & \V116(0) ) | ((\[98]  & \V84(17) ) | V1117),
  \[79]  = (\[138]  & (~V1153 & ~V799)) | ((~\[101]  & (\V121(16)  & ~\V133(8) )) | ((~\[85]  & (~V1153 & ~V799)) | (\V119(0)  & \V133(10) ))),
  \V212(1)  = \[77] ,
  \V212(0)  = \[78] ,
  \V212(7)  = \[71] ,
  \[80]  = (~\[101]  & \V121(17) ) | ((\[101]  & V1153) | (\V122(0)  & \V133(10) )),
  \V212(6)  = \[72] ,
  \V213(0)  = \[79] ,
  \V212(9)  = \[69] ,
  \[82]  = (~V799 & ~V560) | (V749 | V732),
  \V212(8)  = \[70] ,
  \[83]  = \[82]  | V715,
  \[84]  = ~\V235(1)  & ~\V235(0) ,
  \[85]  = V766 | \V133(10) ,
  \V150(0)  = \[16] ,
  \[86]  = \[85]  | V631,
  \V214(0)  = \[80] ,
  \V165(3)  = \[28] ,
  \V165(2)  = \[29] ,
  \V165(5)  = \[26] ,
  \V165(4)  = \[27] ,
  \[10]  = (\[140]  & \V47(3) ) | ((\[123]  & \V15(10) ) | ((\[121]  & \V116(11) ) | ((\[120]  & \V47(11) ) | ((\[119]  & \V84(11) ) | \[122] )))),
  \V165(1)  = \[30] ,
  \[11]  = (\[140]  & \V47(2) ) | ((\[123]  & \V15(9) ) | ((\[121]  & \V116(10) ) | ((\[120]  & \V47(10) ) | ((\[119]  & \V84(10) ) | \[122] )))),
  \V165(0)  = \[31] ,
  \[12]  = (\[139]  & (\[94]  & \V47(4) )) | ((\[139]  & (\[92]  & \V47(1) )) | ((\[139]  & (\[91]  & \V15(11) )) | ((\[139]  & (\V235(0)  & \V47(12) )) | ((\[104]  & (~V732 & \V84(12) )) | ((\[94]  & (\[82]  & \V47(4) )) | ((\[92]  & (\[82]  & \V47(1) )) | ((\[91]  & (\[82]  & \V15(11) )) | ((\[82]  & (\V235(0)  & \V47(12) )) | ((V799 & (~V732 & \V116(12) )) | ((\[139]  & V553) | (\[82]  & V553))))))))))),
  \[13]  = (\[112]  & \V47(7) ) | ((\[110]  & \V15(14) ) | ((\[109]  & \V47(15) ) | ((\[108]  & \V47(4) ) | ((\[106]  & \V116(15) ) | ((\[105]  & \V84(15) ) | \[111] ))))),
  \[90]  = (~\V118(0)  & (~\V133(9)  & (\V133(5)  & ~\V133(1) ))) | ((~\V133(9)  & (\V133(5)  & (~\V133(0)  & ~\V133(1) ))) | ((\[96]  & (V749 & V631)) | (V967 | V831))),
  \[14]  = (\[112]  & \V47(6) ) | ((\[110]  & \V15(13) ) | ((\[109]  & \V47(14) ) | ((\[108]  & \V47(3) ) | ((\[106]  & \V116(14) ) | ((\[105]  & \V84(14) ) | \[111] ))))),
  \[91]  = \[84]  & ~\V235(2) ,
  \V212(11)  = \[67] ,
  \[15]  = (\[112]  & \V47(5) ) | ((\[110]  & \V15(12) ) | ((\[109]  & \V47(13) ) | ((\[108]  & \V47(2) ) | ((\[106]  & \V116(13) ) | ((\[105]  & \V84(13) ) | \[111] ))))),
  \[92]  = \[84]  & \V235(2) ,
  \V212(10)  = \[68] ,
  \[16]  = (\[139]  & (\[94]  & (\V47(8)  & ~\V133(2) ))) | ((\[139]  & (\[92]  & (\V47(5)  & ~\V133(2) ))) | ((\[139]  & (\[91]  & (\V47(1)  & ~\V133(2) ))) | ((\[139]  & (\V235(0)  & (\V47(16)  & ~\V133(2) ))) | ((\[139]  & (V553 & ~\V133(2) )) | ((\[94]  & (\[83]  & \V47(8) )) | ((\[92]  & (\[83]  & \V47(5) )) | ((\[91]  & (\[83]  & \V47(1) )) | ((\[83]  & (\V235(0)  & \V47(16) )) | ((\[106]  & \V116(16) ) | ((\[105]  & \V84(16) ) | (\[83]  & V553))))))))))),
  \[93]  = \[90]  | \V133(10) ,
  \V212(13)  = \[65] ,
  \V165(7)  = \[24] ,
  \[17]  = (\[112]  & \V47(23) ) | ((\[110]  & \V47(16) ) | ((\[109]  & \V47(31) ) | ((\[108]  & \V47(20) ) | ((\[106]  & \V116(31) ) | ((\[105]  & \V84(31) ) | \[111] ))))),
  \[94]  = \V235(1)  & ~\V235(0) ,
  \V212(12)  = \[66] ,
  \V165(6)  = \[25] ,
  \[18]  = (\[112]  & \V47(22) ) | ((\[110]  & \V47(15) ) | ((\[109]  & \V47(30) ) | ((\[108]  & \V47(19) ) | ((\[106]  & \V116(30) ) | ((\[105]  & \V84(30) ) | \[111] ))))),
  \[95]  = (V967 & ~\V133(2) ) | (V831 & V732),
  \V165(9)  = \[22] ,
  \[19]  = (\[112]  & \V47(21) ) | ((\[110]  & \V47(14) ) | ((\[109]  & \V47(29) ) | ((\[108]  & \V47(18) ) | ((\[106]  & \V116(29) ) | ((\[105]  & \V84(29) ) | \[111] ))))),
  \[96]  = ~V732 & ~V715,
  \V212(14)  = \[64] ,
  \V165(8)  = \[23] ,
  \[97]  = V799,
  \[98]  = \[95]  | \V133(10) ,
  \[100]  = ~\[99]  | V1146,
  \[99]  = ~V560 | \V133(2) ,
  \[101]  = ~V766 | \V133(10) ,
  V1117 = ~\[99]  & (V1146 & (~\V118(1)  & (~\V118(0)  & \V133(5) ))),
  \[104]  = V1153 & (V622 & (V560 & ~\V235(0) )),
  \[20]  = (\[112]  & \V47(20) ) | ((\[110]  & \V47(13) ) | ((\[109]  & \V47(28) ) | ((\[108]  & \V47(17) ) | ((\[106]  & \V116(28) ) | ((\[105]  & \V84(28) ) | \[111] ))))),
  \[105]  = \[104] ,
  \[21]  = (\[112]  & \V47(19) ) | ((\[110]  & \V47(12) ) | ((\[109]  & \V47(27) ) | ((\[108]  & \V47(16) ) | ((\[106]  & \V116(27) ) | ((\[105]  & \V84(27) ) | \[111] ))))),
  \[106]  = V799,
  \[22]  = (\[112]  & \V47(18) ) | ((\[110]  & \V47(11) ) | ((\[109]  & \V47(26) ) | ((\[108]  & \V47(15) ) | ((\[106]  & \V116(26) ) | ((\[105]  & \V84(26) ) | \[111] ))))),
  V1146 = V560 & ~\V133(1) ,
  \[23]  = (\[112]  & \V47(17) ) | ((\[110]  & \V47(10) ) | ((\[109]  & \V47(25) ) | ((\[108]  & \V47(14) ) | ((\[106]  & \V116(25) ) | ((\[105]  & \V84(25) ) | \[111] ))))),
  V1153 = \[130]  & (~\V133(9)  & ~\V133(10) ),
  \[108]  = \[92]  & \[83] ,
  \[24]  = (\[112]  & \V47(16) ) | ((\[110]  & \V47(9) ) | ((\[109]  & \V47(24) ) | ((\[108]  & \V47(13) ) | ((\[106]  & \V116(24) ) | ((\[105]  & \V84(24) ) | \[111] ))))),
  \[109]  = \[83]  & \V235(0) ,
  \[25]  = (\[112]  & \V47(15) ) | ((\[110]  & \V47(8) ) | ((\[109]  & \V47(23) ) | ((\[108]  & \V47(12) ) | ((\[106]  & \V116(23) ) | ((\[105]  & \V84(23) ) | \[111] ))))),
  \V142(3)  = \[5] ,
  \[26]  = (\[112]  & \V47(14) ) | ((\[110]  & \V47(7) ) | ((\[109]  & \V47(22) ) | ((\[108]  & \V47(11) ) | ((\[106]  & \V116(22) ) | ((\[105]  & \V84(22) ) | \[111] ))))),
  \V142(2)  = \[6] ,
  \[27]  = (\[112]  & \V47(13) ) | ((\[110]  & \V47(6) ) | ((\[109]  & \V47(21) ) | ((\[108]  & \V47(10) ) | ((\[106]  & \V116(21) ) | ((\[105]  & \V84(21) ) | \[111] ))))),
  \V142(5)  = \[3] ,
  \[28]  = (\[112]  & \V47(12) ) | ((\[110]  & \V47(5) ) | ((\[109]  & \V47(20) ) | ((\[108]  & \V47(9) ) | ((\[106]  & \V116(20) ) | ((\[105]  & \V84(20) ) | \[111] ))))),
  \V142(4)  = \[4] ,
  \[29]  = (\[112]  & \V47(11) ) | ((\[110]  & \V47(4) ) | ((\[109]  & \V47(19) ) | ((\[108]  & \V47(8) ) | ((\[106]  & \V116(19) ) | ((\[105]  & \V84(19) ) | \[111] ))))),
  \V142(1)  = \[7] ,
  \[110]  = \[91]  & \[83] ,
  \V142(0)  = \[8] ,
  \[111]  = \[83]  & V553,
  \[112]  = \[94]  & \[83] ,
  \[113]  = 0,
  \[114]  = V799,
  \[30]  = (\[112]  & \V47(10) ) | ((\[110]  & \V47(3) ) | ((\[109]  & \V47(18) ) | ((\[108]  & \V47(7) ) | ((\[106]  & \V116(18) ) | ((\[105]  & \V84(18) ) | \[111] ))))),
  \[31]  = (\[112]  & \V47(9) ) | ((\[110]  & \V47(2) ) | ((\[109]  & \V47(17) ) | ((\[108]  & \V47(6) ) | ((\[106]  & \V116(17) ) | ((\[105]  & \V84(17) ) | \[111] ))))),
  \[32]  = (\[94]  & (\[93]  & \V84(23) )) | ((\[93]  & (\[92]  & \V84(20) )) | ((\[93]  & (\[91]  & \V84(16) )) | ((\[93]  & (\V235(0)  & \V84(31) )) | ((\[97]  & \V116(31) ) | (\[93]  & V553))))),
  V553 = (\[125]  & (\[91]  & ~\V133(7) )) | ((\[131]  & \[91] ) | (\[91]  & \V133(1) )),
  V554 = ~\[101]  & V967,
  \V143(0)  = \[9] ,
  \[117]  = (~\[85]  & ~\V133(8) ) | V799,
  \[33]  = (\[94]  & (\[93]  & \V84(22) )) | ((\[93]  & (\[92]  & \V84(19) )) | ((\[93]  & (\[91]  & \V84(15) )) | ((\[93]  & (\V235(0)  & \V84(30) )) | ((\[97]  & \V116(30) ) | (\[93]  & V553))))),
  V560 = ~\V133(9)  & (~\V133(7)  & ~\V133(10) ),
  \[118]  = V799,
  V569 = \[130]  & (V622 & ~\V133(8) ),
  \[34]  = (\[94]  & (\[93]  & \V84(21) )) | ((\[93]  & (\[92]  & \V84(18) )) | ((\[93]  & (\[91]  & \V84(14) )) | ((\[93]  & (\V235(0)  & \V84(29) )) | ((\[97]  & \V116(29) ) | (\[93]  & V553))))),
  \[119]  = \[92]  & \[86] ,
  \[35]  = (\[94]  & (\[93]  & \V84(20) )) | ((\[93]  & (\[92]  & \V84(17) )) | ((\[93]  & (\[91]  & \V84(13) )) | ((\[93]  & (\V235(0)  & \V84(28) )) | ((\[97]  & \V116(28) ) | (\[93]  & V553))))),
  \[36]  = (\[94]  & (\[93]  & \V84(19) )) | ((\[93]  & (\[92]  & \V84(16) )) | ((\[93]  & (\[91]  & \V84(12) )) | ((\[93]  & (\V235(0)  & \V84(27) )) | ((\[97]  & \V116(27) ) | (\[93]  & V553))))),
  \V197(27)  = \[36] ,
  \[37]  = (\[94]  & (\[93]  & \V84(18) )) | ((\[93]  & (\[92]  & \V84(15) )) | ((\[93]  & (\[91]  & \V84(11) )) | ((\[93]  & (\V235(0)  & \V84(26) )) | ((\[97]  & \V116(26) ) | (\[93]  & V553))))),
  \V197(26)  = \[37] ,
  \[38]  = (\[94]  & (\[93]  & \V84(17) )) | ((\[93]  & (\[92]  & \V84(14) )) | ((\[93]  & (\[91]  & \V84(10) )) | ((\[93]  & (\V235(0)  & \V84(25) )) | ((\[97]  & \V116(25) ) | (\[93]  & V553))))),
  \V197(29)  = \[34] ,
  \[39]  = (\[94]  & (\[93]  & \V84(16) )) | ((\[93]  & (\[92]  & \V84(13) )) | ((\[93]  & (\[91]  & \V84(9) )) | ((\[93]  & (\V235(0)  & \V84(24) )) | ((\[97]  & \V116(24) ) | (\[93]  & V553))))),
  \V197(28)  = \[35] ,
  \[120]  = \[86]  & \V235(0) ,
  \[121]  = \[118] ,
  \[122]  = \[86]  & V553,
  \V145(1)  = \[10] ,
  \[123]  = \[91]  & \[86] ,
  \V145(0)  = \[11] ,
  V622 = ~\V133(4)  & ~\V133(9) ,
  \[124]  = (V766 & ~\V133(8) ) | V569,
  \[40]  = (\[94]  & (\[93]  & \V84(15) )) | ((\[93]  & (\[92]  & \V84(12) )) | ((\[93]  & (\[91]  & \V84(8) )) | ((\[93]  & (\V235(0)  & \V84(23) )) | ((\[97]  & \V116(23) ) | (\[93]  & V553))))),
  V631 = V622 & ~\V133(6) ,
  \V197(21)  = \[42] ,
  \[125]  = \V133(6)  | \V133(5) ,
  \[41]  = (\[94]  & (\[93]  & \V84(14) )) | ((\[93]  & (\[92]  & \V84(11) )) | ((\[93]  & (\[91]  & \V84(7) )) | ((\[93]  & (\V235(0)  & \V84(22) )) | ((\[97]  & \V116(22) ) | (\[93]  & V553))))),
  \V197(20)  = \[43] ,
  \[126]  = (\[92]  & \V84(9) ) | V553,
  \[42]  = (\[94]  & (\[93]  & \V84(13) )) | ((\[93]  & (\[92]  & \V84(10) )) | ((\[93]  & (\[91]  & \V84(6) )) | ((\[93]  & (\V235(0)  & \V84(21) )) | ((\[97]  & \V116(21) ) | (\[93]  & V553))))),
  \V197(23)  = \[40] ,
  \[43]  = (\[94]  & (\[93]  & \V84(12) )) | ((\[93]  & (\[91]  & \V84(5) )) | ((\[93]  & (\V235(0)  & \V84(20) )) | ((\[126]  & \[93] ) | (\[97]  & \V116(20) )))),
  \V197(22)  = \[41] ,
  \[44]  = (\[94]  & (\[93]  & \V84(11) )) | ((\[93]  & (\[92]  & \V84(8) )) | ((\[93]  & (\[91]  & \V84(4) )) | ((\[93]  & (\V235(0)  & \V84(19) )) | ((\[97]  & \V116(19) ) | (\[93]  & V553))))),
  \V197(25)  = \[38] ,
  \[129]  = \[124]  | \V133(10) ,
  \[45]  = (\[94]  & (\[93]  & \V84(10) )) | ((\[93]  & (\[92]  & \V84(7) )) | ((\[93]  & (\[91]  & \V84(3) )) | ((\[93]  & (\V235(0)  & \V84(18) )) | ((\[97]  & \V116(18) ) | (\[93]  & V553))))),
  \V197(24)  = \[39] ,
  \V146(0)  = \[12] ,
  \[46]  = (\[94]  & (\[93]  & \V84(9) )) | ((\[93]  & (\[92]  & \V84(6) )) | ((\[93]  & (\[91]  & \V84(2) )) | ((\[93]  & (\V235(0)  & \V84(17) )) | ((\[97]  & \V116(17) ) | (\[93]  & V553))))),
  \V197(17)  = \[46] ,
  \[47]  = (\[94]  & (\[93]  & \V84(8) )) | ((\[93]  & (\[92]  & \V84(5) )) | ((\[93]  & (\[91]  & \V84(1) )) | ((\[93]  & (\V235(0)  & \V84(16) )) | ((\[97]  & \V116(16) ) | (\[93]  & V553))))),
  \V197(16)  = \[47] ,
  \[48]  = (\[94]  & (\[93]  & \V84(7) )) | ((\[93]  & (\[92]  & \V84(4) )) | ((\[93]  & (\[91]  & \V84(0) )) | ((\[93]  & (\V235(0)  & \V84(15) )) | ((\[97]  & \V116(15) ) | (\[93]  & V553))))),
  \V197(19)  = \[44] ,
  \[49]  = (\[94]  & (\[93]  & \V84(6) )) | ((\[93]  & (\[92]  & \V84(3) )) | ((\[93]  & (\[91]  & \V47(31) )) | ((\[93]  & (\V235(0)  & \V84(14) )) | ((\[97]  & \V116(14) ) | (\[93]  & V553))))),
  \V197(18)  = \[45] ,
  \[130]  = \V133(2)  & \V133(1) ,
  \[131]  = \V133(10)  | \V133(2) ,
  V715 = \[139]  & V631,
  \[134]  = (\[92]  & \V84(2) ) | V553,
  \V134(0)  = \[0] ,
  \V197(3)  = \[60] ,
  \[50]  = (\[94]  & (\[93]  & \V84(5) )) | ((\[93]  & (\[91]  & \V47(30) )) | ((\[93]  & (\V235(0)  & \V84(13) )) | ((\[134]  & \[93] ) | (\[97]  & \V116(13) )))),
  \V197(11)  = \[52] ,
  V732 = V631 & ~\V133(2) ,
  \[135]  = (\[92]  & \V84(1) ) | V553,
  \V197(2)  = \[61] ,
  \[51]  = (\[94]  & (\[93]  & \V84(4) )) | ((\[93]  & (\[91]  & \V47(29) )) | ((\[93]  & (\V235(0)  & \V84(12) )) | ((\[135]  & \[93] ) | (\[97]  & \V116(12) )))),
  \V197(10)  = \[53] ,
  \V197(5)  = \[58] ,
  V749 = V622 & \V133(3) ,
  \[52]  = (\[94]  & (\[93]  & \V84(3) )) | ((\[93]  & (\[92]  & \V84(0) )) | ((\[93]  & (\[91]  & \V47(28) )) | ((\[93]  & (\V235(0)  & \V84(11) )) | ((\[97]  & \V116(11) ) | (\[93]  & V553))))),
  \V197(13)  = \[50] ,
  \V149(2)  = \[13] ,
  \V197(4)  = \[59] ,
  \[53]  = (\[94]  & (\[93]  & \V84(2) )) | ((\[93]  & (\[92]  & \V47(31) )) | ((\[93]  & (\[91]  & \V47(27) )) | ((\[93]  & (\V235(0)  & \V84(10) )) | ((\[97]  & \V116(10) ) | (\[93]  & V553))))),
  \V197(12)  = \[51] ,
  V766 = ~\V133(9)  & \V133(7) ,
  \[138]  = \V133(8)  & ~\V133(10) ,
  \[54]  = (\[94]  & (\[93]  & \V84(1) )) | ((\[93]  & (\[92]  & \V47(30) )) | ((\[93]  & (\[91]  & \V47(26) )) | ((\[93]  & (\V235(0)  & \V84(9) )) | ((\[97]  & \V116(9) ) | (\[93]  & V553))))),
  \V197(15)  = \[48] ,
  \[139]  = V622 & ~\V133(1) ,
  \[55]  = (\[94]  & (\[93]  & \V84(0) )) | ((\[93]  & (\[92]  & \V47(29) )) | ((\[93]  & (\[91]  & \V47(25) )) | ((\[93]  & (\V235(0)  & \V84(8) )) | ((\[97]  & \V116(8) ) | (\[93]  & V553))))),
  \V197(14)  = \[49] ,
  \V197(1)  = \[62] ,
  \[56]  = (\[94]  & (\[93]  & \V47(31) )) | ((\[93]  & (\[92]  & \V47(28) )) | ((\[93]  & (\[91]  & \V47(24) )) | ((\[93]  & (\V235(0)  & \V84(7) )) | ((\[97]  & \V116(7) ) | (\[93]  & V553))))),
  \V197(0)  = \[63] ,
  V799 = \V133(9)  & ~\V133(10) ,
  \[57]  = (\[94]  & (\[93]  & \V47(30) )) | ((\[93]  & (\[92]  & \V47(27) )) | ((\[93]  & (\[91]  & \V47(23) )) | ((\[93]  & (\V235(0)  & \V84(6) )) | ((\[97]  & \V116(6) ) | (\[93]  & V553))))),
  \V149(1)  = \[14] ,
  \[58]  = (\[94]  & (\[93]  & \V47(29) )) | ((\[93]  & (\[92]  & \V47(26) )) | ((\[93]  & (\[91]  & \V47(22) )) | ((\[93]  & (\V235(0)  & \V84(5) )) | ((\[97]  & \V116(5) ) | (\[93]  & V553))))),
  \V149(0)  = \[15] ,
  \[59]  = (\[94]  & (\[93]  & \V47(28) )) | ((\[93]  & (\[92]  & \V47(25) )) | ((\[93]  & (\[91]  & \V47(21) )) | ((\[93]  & (\V235(0)  & \V84(4) )) | ((\[97]  & \V116(4) ) | (\[93]  & V553))))),
  \V235(2)  = (~\[125]  & \V133(2) ) | ((\V133(8)  & \V133(2) ) | \[130] ),
  \V136(1)  = \[1] ,
  \[140]  = \[94]  & \[86] ,
  \V197(7)  = \[56] ,
  \V136(0)  = \[2] ,
  \V197(6)  = \[57] ,
  \V197(9)  = \[54] ,
  \V235(1)  = (~\[131]  & (~\[125]  & \V133(1) )) | ((\[138]  & \V133(1) ) | ((\V133(7)  & ~\V133(0) ) | (~\V133(5)  & ~\V133(0) ))),
  \V197(8)  = \[55] ,
  \V235(0)  = (\[130]  & \V133(3) ) | \V133(10) ;
endmodule

