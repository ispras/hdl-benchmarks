//NOTE: no-implementation module stub

module REG16LC (
    input wire DSPCLK,
    input wire MMR_web,
    input wire FSDIV_we_PSET,
    input wire [15:0] DMD_FSDIV,
    output reg [15:0] FSDIV,
    input wire RST
);

endmodule
