--------------------------------------------------------------------
--       Actel Axcelerator VITAL Library
--       NAME: axcelerator.vhd
--       DATE: July 20, 2004
---------------------------------------------------------------------/

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.VITAL_Timing.all;

package COMPONENTS is

constant DefaultTimingChecksOn : Boolean := True;
constant DefaultXGenerationOn : Boolean := False;
constant DefaultXon : Boolean := False;
constant DefaultMsgOn : Boolean := True;



------ Component ADD1 ------
 component ADD1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		FCI		: in    STD_ULOGIC;
		S		: out    STD_ULOGIC;
		FCO		: out    STD_ULOGIC);
 end component;


------ Component AND2 ------
 component AND2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND2A ------
 component AND2A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND2B ------
 component AND2B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND3 ------
 component AND3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND3A ------
 component AND3A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND3B ------
 component AND3B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND3C ------
 component AND3C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND4 ------
 component AND4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND4A ------
 component AND4A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND4B ------
 component AND4B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND4C ------
 component AND4C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND4D ------
 component AND4D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND5A ------
 component AND5A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND5B ------
 component AND5B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND5C ------
 component AND5C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO1 ------
 component AO1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO10 ------
 component AO10
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO11 ------
 component AO11
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO12 ------
 component AO12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO13 ------
 component AO13
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO14 ------
 component AO14
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO15 ------
 component AO15
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO16 ------
 component AO16
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO17 ------
 component AO17
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO18 ------
 component AO18
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO1A ------
 component AO1A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO1B ------
 component AO1B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO1C ------
 component AO1C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO1D ------
 component AO1D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO1E ------
 component AO1E
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO2 ------
 component AO2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO2A ------
 component AO2A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO2B ------
 component AO2B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO2C ------
 component AO2C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO2D ------
 component AO2D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO2E ------
 component AO2E
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO3 ------
 component AO3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO3A ------
 component AO3A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO3B ------
 component AO3B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO3C ------
 component AO3C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO4A ------
 component AO4A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO5A ------
 component AO5A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO6 ------
 component AO6
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO6A ------
 component AO6A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO7 ------
 component AO7
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO8 ------
 component AO8
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO9 ------
 component AO9
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI1 ------
 component AOI1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI1A ------
 component AOI1A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI1B ------
 component AOI1B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI1C ------
 component AOI1C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI1D ------
 component AOI1D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI2A ------
 component AOI2A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI2B ------
 component AOI2B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI3A ------
 component AOI3A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI4 ------
 component AOI4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI4A ------
 component AOI4A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI5 ------
 component AOI5
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AFCNTECP1 ------
 component AFCNTECP1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_UD_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_Q_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_UD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		Q		:  out STD_ULOGIC;
		UD		:  in    STD_ULOGIC;
		FCI		:  in    STD_ULOGIC;
		FCO		:  out    STD_ULOGIC);

 end component;


------ Component ARCNTECP1 ------
 component ARCNTECP1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_UD_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_Q_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_UD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		Q		:  out STD_ULOGIC;
		UD		:  in    STD_ULOGIC;
		FCI		:  in    STD_ULOGIC;
		FCO		:  out    STD_ULOGIC);

 end component;


------ Component AFCNTELDCP1 ------
 component AFCNTELDCP1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_UD_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_LD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_LD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_LD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_LD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_LD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_UD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		LD		:  in    STD_ULOGIC;
		Q		:  out STD_ULOGIC;
		UD		:  in    STD_ULOGIC;
		FCI		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		FCO		:  out    STD_ULOGIC);

 end component;


------ Component ARCNTELDCP1 ------
 component ARCNTELDCP1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_UD_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_LD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_LD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_LD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_LD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_LD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_UD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		LD		:  in    STD_ULOGIC;
		Q		:  out STD_ULOGIC;
		UD		:  in    STD_ULOGIC;
		FCI		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		FCO		:  out    STD_ULOGIC);

 end component;


------ Component AX1 ------
 component AX1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AX1A ------
 component AX1A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AX1B ------
 component AX1B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AX1C ------
 component AX1C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AX1D ------
 component AX1D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AX1E ------
 component AX1E
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXO1 ------
 component AXO1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXO2 ------
 component AXO2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXO3 ------
 component AXO3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXO5 ------
 component AXO5
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXO6 ------
 component AXO6
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXO7 ------
 component AXO7
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXOI1 ------
 component AXOI1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXOI2 ------
 component AXOI2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXOI3 ------
 component AXOI3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXOI4 ------
 component AXOI4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXOI5 ------
 component AXOI5
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXOI7 ------
 component AXOI7
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF ------
 component BIBUF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_8 ------
 component BIBUF_S_8
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_8D ------
 component BIBUF_S_8D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_8U ------
 component BIBUF_S_8U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_12 ------
 component BIBUF_S_12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_12D ------
 component BIBUF_S_12D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_12U ------
 component BIBUF_S_12U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_16 ------
 component BIBUF_S_16
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_16D ------
 component BIBUF_S_16D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_16U ------
 component BIBUF_S_16U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_24 ------
 component BIBUF_S_24
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_24D ------
 component BIBUF_S_24D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_24U ------
 component BIBUF_S_24U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_8 ------
 component BIBUF_F_8
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_8D ------
 component BIBUF_F_8D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_8U ------
 component BIBUF_F_8U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_12 ------
 component BIBUF_F_12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_12D ------
 component BIBUF_F_12D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_12U ------
 component BIBUF_F_12U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_16 ------
 component BIBUF_F_16
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_16D ------
 component BIBUF_F_16D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_16U ------
 component BIBUF_F_16U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_24 ------
 component BIBUF_F_24
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_24D ------
 component BIBUF_F_24D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_24U ------
 component BIBUF_F_24U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS25 ------
 component BIBUF_LVCMOS25
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS25D ------
 component BIBUF_LVCMOS25D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS25U ------
 component BIBUF_LVCMOS25U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS18 ------
 component BIBUF_LVCMOS18
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS18D ------
 component BIBUF_LVCMOS18D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS18U ------
 component BIBUF_LVCMOS18U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS15 ------
 component BIBUF_LVCMOS15
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS15D ------
 component BIBUF_LVCMOS15D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS15U ------
 component BIBUF_LVCMOS15U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_PCI ------
 component BIBUF_PCI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_PCIX ------
 component BIBUF_PCIX
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_GTLP33 ------
 component BIBUF_GTLP33
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_GTLP25 ------
 component BIBUF_GTLP25
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BUFA ------
 component BUFA
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BUFD ------
 component BUFD
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBIBUF ------
 component CLKBIBUF
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;
                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_D_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_D                  : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E                  : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                PAD             : inout  STD_ULOGIC;
                D               : in     STD_ULOGIC;
                E               : in     STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 end component;


------ Component CLKBUF ------
 component CLKBUF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF_LVCMOS25 ------
 component CLKBUF_LVCMOS25
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF_LVCMOS18 ------
 component CLKBUF_LVCMOS18
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF_LVCMOS15 ------
 component CLKBUF_LVCMOS15
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF_PCI ------
 component CLKBUF_PCI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF_PCIX ------
 component CLKBUF_PCIX
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF_GTLP33 ------
 component CLKBUF_GTLP33
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF_GTLP25 ------
 component CLKBUF_GTLP25
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF_HSTL_I ------
 component CLKBUF_HSTL_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF_SSTL3_I ------
 component CLKBUF_SSTL3_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF_SSTL3_II ------
 component CLKBUF_SSTL3_II
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF_SSTL2_I ------
 component CLKBUF_SSTL2_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF_SSTL2_II ------
 component CLKBUF_SSTL2_II
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CM7 ------
 component CM7
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S0		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CM8 ------
 component CM8
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CM8BUFF ------
 component CM8BUFF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
                tpw_A_posedge   : VitalDelayType := 0.000 ns;
                tpw_A_negedge   : VitalDelayType := 0.000 ns;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CM8INV ------
 component CM8INV
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMA9 ------
 component CMA9
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMAF ------
 component CMAF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMB3 ------
 component CMB3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMB7 ------
 component CMB7
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMBB ------
 component CMBB
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMBF ------
 component CMBF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMEA ------
 component CMEA
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMEB ------
 component CMEB
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMEE ------
 component CMEE
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMEF ------
 component CMEF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMF1 ------
 component CMF1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMF2 ------
 component CMF2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMF3 ------
 component CMF3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMF4 ------
 component CMF4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMF5 ------
 component CMF5
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMF6 ------
 component CMF6
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMF7 ------
 component CMF7
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMF8 ------
 component CMF8
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMF9 ------
 component CMF9
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMFA ------
 component CMFA
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMFB ------
 component CMFB
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMFC ------
 component CMFC
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMFD ------
 component CMFD
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CMFE ------
 component CMFE
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CS1 ------
 component CS1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CS2 ------
 component CS2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CY2A ------
 component CY2A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B0		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A1		: in    STD_ULOGIC;
		B1		: in    STD_ULOGIC;
		A0		: in    STD_ULOGIC;
		B0		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CY2B ------
 component CY2B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B0		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A1		: in    STD_ULOGIC;
		B1		: in    STD_ULOGIC;
		A0		: in    STD_ULOGIC;
		B0		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component DF1 ------
 component DF1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DF1_CC ------
 component DF1_CC
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DF1B ------
 component DF1B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFC1B ------
 component DFC1B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFC1B_CC ------
 component DFC1B_CC
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFC1D ------
 component DFC1D
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFE1C ------
 component DFE1C
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFE1B ------
 component DFE1B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFE3C ------
 component DFE3C
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFE3D ------
 component DFE3D
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFE4F ------
 component DFE4F
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFE4G ------
 component DFE4G
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFEG ------
 component DFEG
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFEH ------
 component DFEH
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFP1 ------
 component DFP1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFP1A ------
 component DFP1A
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFP1B ------
 component DFP1B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFP1B_CC ------
 component DFP1B_CC
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFP1D ------
 component DFP1D
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFPC ------
 component DFPC
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFPCB ------
 component DFPCB
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFPCC ------
 component DFPCC
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DL1 ------
 component DL1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DL1A ------
 component DL1A
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DL1B ------
 component DL1B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DL1C ------
 component DL1C
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DL2A ------
 component DL2A
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DL2C ------
 component DL2C
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLC ------
 component DLC
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLC1 ------
 component DLC1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLC1A ------
 component DLC1A
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLC1F ------
 component DLC1F
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DLC1G ------
 component DLC1G
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DLCA ------
 component DLCA
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLE ------
 component DLE
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_E_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLE1D ------
 component DLE1D
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_E_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DLE2B ------
 component DLE2B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_E_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLE2C ------
 component DLE2C
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_E_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLE3B ------
 component DLE3B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_E_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLE3C ------
 component DLE3C
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_E_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLEA ------
 component DLEA
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_E_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLEB ------
 component DLEB
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_E_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLEC ------
 component DLEC
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_E_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLM ------
 component DLM
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_A_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		A		:  in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLM2 ------
 component DLM2
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_A_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		A		:  in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLM2B ------
 component DLM2B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_A_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		A		:  in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLM3 ------
 component DLM3
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D0_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S0_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S1_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D0_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D0_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D0_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D0_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S0_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S0_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S0_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S0_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D1_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D1_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D1_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D1_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S1_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S1_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S1_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S1_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D2_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D2_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D2_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D2_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D3_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D3_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D3_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D3_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D0		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S0		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S1		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D0		:  in    STD_ULOGIC;
		S0		:  in    STD_ULOGIC;
		D1		:  in    STD_ULOGIC;
		S1		:  in    STD_ULOGIC;
		D2		:  in    STD_ULOGIC;
		D3		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLM3A ------
 component DLM3A
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D0_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S0_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S1_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D0_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D0_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D0_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D0_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S0_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S0_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S0_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S0_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D1_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D1_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D1_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D1_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S1_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S1_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S1_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S1_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D2_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D2_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D2_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D2_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D3_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D3_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D3_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D3_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D0		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S0		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S1		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D0		:  in    STD_ULOGIC;
		S0		:  in    STD_ULOGIC;
		D1		:  in    STD_ULOGIC;
		S1		:  in    STD_ULOGIC;
		D2		:  in    STD_ULOGIC;
		D3		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLM4 ------
 component DLM4
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S0_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D0_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S10_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S10_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S10_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S10_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S11_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S11_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S11_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S11_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S0_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S0_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S0_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S0_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D0_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D0_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D0_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D0_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D1_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D1_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D1_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D1_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D2_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D2_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D2_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D2_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D3_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D3_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D3_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D3_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S0		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D0		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		S10		:  in    STD_ULOGIC;
		S11		:  in    STD_ULOGIC;
		S0		:  in    STD_ULOGIC;
		D0		:  in    STD_ULOGIC;
		D1		:  in    STD_ULOGIC;
		D2		:  in    STD_ULOGIC;
		D3		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLM4A ------
 component DLM4A
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S0_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D0_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S10_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S10_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S10_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S10_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S11_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S11_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S11_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S11_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S0_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S0_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S0_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S0_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D0_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D0_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D0_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D0_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D1_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D1_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D1_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D1_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D2_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D2_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D2_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D2_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D3_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D3_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D3_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D3_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S0		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D0		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		S10		:  in    STD_ULOGIC;
		S11		:  in    STD_ULOGIC;
		S0		:  in    STD_ULOGIC;
		D0		:  in    STD_ULOGIC;
		D1		:  in    STD_ULOGIC;
		D2		:  in    STD_ULOGIC;
		D3		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLMA ------
 component DLMA
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_A_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		A		:  in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLME1A ------
 component DLME1A
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_A_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_E_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		A		:  in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLP1 ------
 component DLP1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLP1A ------
 component DLP1A
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLP1B ------
 component DLP1B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLP1C ------
 component DLP1C
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLP1D ------
 component DLP1D
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DLP1E ------
 component DLP1E
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component FA1 ------
 component FA1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CI_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CI_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CI		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		CI		: in    STD_ULOGIC;
		S		: out    STD_ULOGIC;
		CO		: out    STD_ULOGIC);
 end component;


------ Component FCEND_BUFF ------
 component FCEND_BUFF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_FCI_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_FCI		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		FCI		: in    STD_ULOGIC;
		CO		: out    STD_ULOGIC);
 end component;


------ Component FCEND_INV ------
 component FCEND_INV
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_FCI_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_FCI		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		FCI		: in    STD_ULOGIC;
		CO		: out    STD_ULOGIC);
 end component;


------ Component FCINIT_BUFF ------
 component FCINIT_BUFF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		FCO		: out    STD_ULOGIC);
 end component;


------ Component FCINIT_GND ------
 component FCINIT_GND
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True		);
    port(
		FCO		: out    STD_ULOGIC);
 end component;


------ Component FCINIT_INV ------
 component FCINIT_INV
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		FCO		: out    STD_ULOGIC);
 end component;


------ Component FCINIT_VCC ------
 component FCINIT_VCC
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True		);
    port(
		FCO		: out    STD_ULOGIC);
 end component;


------ Component GAND2 ------
 component GAND2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		G		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component GMX4 ------
 component GMX4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S0		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		G		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component GNAND2 ------
 component GNAND2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		G		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component GND ------
 component GND
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True		);
    port(
		Y		: out    STD_ULOGIC);
 end component;


------ Component GNOR2 ------
 component GNOR2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		G		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component GOR2 ------
 component GOR2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		G		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component GXOR2 ------
 component GXOR2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		G		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component HA1 ------
 component HA1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		S		: out    STD_ULOGIC;
		CO		: out    STD_ULOGIC);
 end component;


------ Component HA1A ------
 component HA1A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		S		: out    STD_ULOGIC;
		CO		: out    STD_ULOGIC);
 end component;


------ Component HA1B ------
 component HA1B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		S		: out    STD_ULOGIC;
		CO		: out    STD_ULOGIC);
 end component;


------ Component HA1C ------
 component HA1C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		S		: out    STD_ULOGIC;
		CO		: out    STD_ULOGIC);
 end component;


------ Component HCLKBIBUF ------
 component HCLKBIBUF
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;
                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_D_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_D                  : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E                  : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                PAD             : inout  STD_ULOGIC;
                D               : in     STD_ULOGIC;
                E               : in     STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 end component;


------ Component HCLKBUF ------
 component HCLKBUF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component HCLKBUF_LVCMOS25 ------
 component HCLKBUF_LVCMOS25
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component HCLKBUF_LVCMOS18 ------
 component HCLKBUF_LVCMOS18
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component HCLKBUF_LVCMOS15 ------
 component HCLKBUF_LVCMOS15
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component HCLKBUF_PCI ------
 component HCLKBUF_PCI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component HCLKBUF_PCIX ------
 component HCLKBUF_PCIX
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component HCLKBUF_GTLP33 ------
 component HCLKBUF_GTLP33
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component HCLKBUF_GTLP25 ------
 component HCLKBUF_GTLP25
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component HCLKBUF_HSTL_I ------
 component HCLKBUF_HSTL_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component HCLKBUF_SSTL3_I ------
 component HCLKBUF_SSTL3_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component HCLKBUF_SSTL3_II ------
 component HCLKBUF_SSTL3_II
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component HCLKBUF_SSTL2_I ------
 component HCLKBUF_SSTL2_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component HCLKBUF_SSTL2_II ------
 component HCLKBUF_SSTL2_II
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component HCLKINT ------
 component HCLKINT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF ------
 component INBUF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS25 ------
 component INBUF_LVCMOS25
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS25D ------
 component INBUF_LVCMOS25D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS25U ------
 component INBUF_LVCMOS25U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS18 ------
 component INBUF_LVCMOS18
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS18D ------
 component INBUF_LVCMOS18D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS18U ------
 component INBUF_LVCMOS18U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS15 ------
 component INBUF_LVCMOS15
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS15D ------
 component INBUF_LVCMOS15D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS15U ------
 component INBUF_LVCMOS15U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_PCI ------
 component INBUF_PCI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_PCIX ------
 component INBUF_PCIX
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_GTLP33 ------
 component INBUF_GTLP33
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_GTLP25 ------
 component INBUF_GTLP25
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_HSTL_I ------
 component INBUF_HSTL_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_SSTL3_I ------
 component INBUF_SSTL3_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_SSTL3_II ------
 component INBUF_SSTL3_II
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_SSTL2_I ------
 component INBUF_SSTL2_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_SSTL2_II ------
 component INBUF_SSTL2_II
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INV ------
 component INV
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INVA ------
 component INVA
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INVD ------
 component INVD
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOI_DFEG ------
 component IOI_DFEG
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component IOI_DFEH ------
 component IOI_DFEH
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component IOI_BUFF ------
 component IOI_BUFF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOOE_BUFF ------
 component IOOE_BUFF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOOE_DFEG ------
 component IOOE_DFEG
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_YOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_YOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_YOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tperiod_CLK_negedge        :  VitalDelayType := 0.000 ns;
		tpw_CLK_posedge        :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge        :  VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                CLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                Q                : out    STD_ULOGIC;
                YOUT                : out    STD_ULOGIC);
 end component;


------ Component IOOE_DFEH ------
 component IOOE_DFEH
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_YOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_YOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_YOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge   :   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge	:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge       :   VitalDelayType := 0.000 ns;
		tperiod_CLK_negedge        :  VitalDelayType := 0.000 ns;
		tpw_CLK_posedge        :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge        :  VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge   :   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge	:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                CLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                Q                : out    STD_ULOGIC;
                YOUT                : out    STD_ULOGIC);
 end component;


------ Component IOPAD_IN ------
 component IOPAD_IN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
-- DNW: Add the following 2 lines
		tpw_PAD_posedge		: VitalDelayType := 0.000 ns;
		tpw_PAD_negedge		: VitalDelayType := 0.000 ns;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOPAD_TRI ------
 component IOPAD_TRI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_D_posedge	: VitalDelayType := 0.000 ns;
		tpw_D_negedge	: VitalDelayType := 0.000 ns;
		tpw_E_posedge   : VitalDelayType := 0.000 ns;
		tpw_E_negedge	: VitalDelayType := 0.000 ns;

		tpd_D_PAD       : VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component IOPAD_BI ------
 component IOPAD_BI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		
                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;
  
                tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component JKF ------
 component JKF
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_J_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_J_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_J_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		thold_J_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_K_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		thold_K_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge		:  VitalDelayType := 0.000 ns;
		tipd_J      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_K      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK	:   VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		J	:  in    STD_ULOGIC;
		K	:  in    STD_ULOGIC;
	        CLK	:  in    STD_ULOGIC;
		Q	:  out    STD_ULOGIC);

 end component;


------ Component JKF1B ------
 component JKF1B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_J_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_J_CLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
		tsetup_J_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		thold_J_CLK_negedge_negedge   :   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_K_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		thold_K_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge		:  VitalDelayType := 0.000 ns;
		tipd_J      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_K      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK	:   VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		J	:  in    STD_ULOGIC;
		K	:  in    STD_ULOGIC;
	        CLK	:  in    STD_ULOGIC;
		Q	:  out    STD_ULOGIC);

 end component;


------ Component JKF2A ------
 component JKF2A
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_J_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_J_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_J_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		thold_J_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_K_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		thold_K_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge	:  VitalDelayType := 0.000 ns;
		tipd_CLR	:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_J      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_K      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK	:   VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		J	:  in    STD_ULOGIC;
		K	:  in    STD_ULOGIC;
	        CLR	:  in    STD_ULOGIC;
	        CLK	:  in    STD_ULOGIC;
		Q	:  out    STD_ULOGIC);

 end component;


------ Component JKF2B ------
 component JKF2B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_J_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_J_CLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
		tsetup_J_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		thold_J_CLK_negedge_negedge   :   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_K_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		thold_K_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge           :   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge	:  VitalDelayType := 0.000 ns;
		tipd_CLR	:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_J      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_K      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK	:   VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		J	:  in    STD_ULOGIC;
		K	:  in    STD_ULOGIC;
	        CLR	:  in    STD_ULOGIC;
	        CLK	:  in    STD_ULOGIC;
		Q	:  out    STD_ULOGIC);

 end component;


------ Component JKF3A ------
 component JKF3A
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_J_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_J_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_J_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		thold_J_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_K_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		thold_K_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge   	:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE	:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_J      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_K      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK	:   VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		J	:  in    STD_ULOGIC;
		K	:  in    STD_ULOGIC;
	        PRE	:  in    STD_ULOGIC;
	        CLK	:  in    STD_ULOGIC;
		Q	:  out    STD_ULOGIC);

 end component;


------ Component JKF3B ------
 component JKF3B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_J_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_J_CLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
		tsetup_J_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		thold_J_CLK_negedge_negedge   :   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_K_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		thold_K_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge   	:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE	:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_J      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_K      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK	:   VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		J	:  in    STD_ULOGIC;
		K	:  in    STD_ULOGIC;
	        PRE	:  in    STD_ULOGIC;
	        CLK	:  in    STD_ULOGIC;
		Q	:  out    STD_ULOGIC);

 end component;


------ Component MAJ3 ------
 component MAJ3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MAJ3X ------
 component MAJ3X
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MAJ3XI ------
 component MAJ3XI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MIN3 ------
 component MIN3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MIN3X ------
 component MIN3X
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MIN3XI ------
 component MIN3XI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MULT1 ------
 component MULT1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_PO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_PO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PI_PO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_PO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PI_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PI		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		PI		: in    STD_ULOGIC;
		FCI		: in    STD_ULOGIC;
		PO		: out    STD_ULOGIC;
		FCO		: out    STD_ULOGIC);
 end component;


------ Component MX2 ------
 component MX2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MX2A ------
 component MX2A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MX2B ------
 component MX2B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MX2C ------
 component MX2C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MX4 ------
 component MX4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S0		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S1		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND2 ------
 component NAND2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND2A ------
 component NAND2A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND2B ------
 component NAND2B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND3 ------
 component NAND3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND3A ------
 component NAND3A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND3B ------
 component NAND3B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND3C ------
 component NAND3C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND4 ------
 component NAND4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND4A ------
 component NAND4A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND4B ------
 component NAND4B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND4C ------
 component NAND4C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND4D ------
 component NAND4D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND5B ------
 component NAND5B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND5C ------
 component NAND5C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR2 ------
 component NOR2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR2A ------
 component NOR2A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR2B ------
 component NOR2B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR3 ------
 component NOR3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR3A ------
 component NOR3A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR3B ------
 component NOR3B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR3C ------
 component NOR3C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR4 ------
 component NOR4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR4A ------
 component NOR4A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR4B ------
 component NOR4B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR4C ------
 component NOR4C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR4D ------
 component NOR4D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR5B ------
 component NOR5B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR5C ------
 component NOR5C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA1 ------
 component OA1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA1A ------
 component OA1A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA1B ------
 component OA1B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		C		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA1C ------
 component OA1C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		C		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA2 ------
 component OA2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA2A ------
 component OA2A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA3 ------
 component OA3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA3A ------
 component OA3A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA3B ------
 component OA3B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA4 ------
 component OA4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA4A ------
 component OA4A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA5 ------
 component OA5
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OAI1 ------
 component OAI1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OAI2A ------
 component OAI2A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OAI3 ------
 component OAI3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OAI3A ------
 component OAI3A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR2 ------
 component OR2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR2A ------
 component OR2A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR2B ------
 component OR2B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR3 ------
 component OR3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR3A ------
 component OR3A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR3B ------
 component OR3B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR3C ------
 component OR3C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR4 ------
 component OR4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR4A ------
 component OR4A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR4B ------
 component OR4B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR4C ------
 component OR4C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR4D ------
 component OR4D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR5A ------
 component OR5A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR5B ------
 component OR5B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR5C ------
 component OR5C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF ------
 component OUTBUF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_S_8 ------
 component OUTBUF_S_8
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_S_12 ------
 component OUTBUF_S_12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_S_16 ------
 component OUTBUF_S_16
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_S_24 ------
 component OUTBUF_S_24
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_F_8 ------
 component OUTBUF_F_8
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_F_12 ------
 component OUTBUF_F_12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_F_16 ------
 component OUTBUF_F_16
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_F_24 ------
 component OUTBUF_F_24
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_LVCMOS25 ------
 component OUTBUF_LVCMOS25
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_LVCMOS18 ------
 component OUTBUF_LVCMOS18
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_LVCMOS15 ------
 component OUTBUF_LVCMOS15
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_PCI ------
 component OUTBUF_PCI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_PCIX ------
 component OUTBUF_PCIX
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_GTLP33 ------
 component OUTBUF_GTLP33
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_GTLP25 ------
 component OUTBUF_GTLP25
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_HSTL_I ------
 component OUTBUF_HSTL_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_SSTL3_I ------
 component OUTBUF_SSTL3_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_SSTL3_II ------
 component OUTBUF_SSTL3_II
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_SSTL2_I ------
 component OUTBUF_SSTL2_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_SSTL2_II ------
 component OUTBUF_SSTL2_II
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component PLLHCLK ------
 component PLLHCLK
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component PLLRCLK ------
 component PLLRCLK
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component SFCNTECP1 ------
 component SFCNTECP1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_UD_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_Q_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_UD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		Q		:  out STD_ULOGIC;
		UD		:  in    STD_ULOGIC;
		FCI		:  in    STD_ULOGIC;
		FCO		:  out    STD_ULOGIC);

 end component;


------ Component SRCNTECP1 ------
 component SRCNTECP1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_UD_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_Q_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_UD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		Q		:  out STD_ULOGIC;
		UD		:  in    STD_ULOGIC;
		FCI		:  in    STD_ULOGIC;
		FCO		:  out    STD_ULOGIC);

 end component;


------ Component SFCNTELDCP1 ------
 component SFCNTELDCP1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_UD_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_Q_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_LD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_LD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_LD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_LD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_UD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_LD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		Q		:  out STD_ULOGIC;
		UD		:  in    STD_ULOGIC;
		FCI		:  in    STD_ULOGIC;
		LD		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		FCO		:  out    STD_ULOGIC);

 end component;


------ Component SRCNTELDCP1 ------
 component SRCNTELDCP1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_UD_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_Q_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_LD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_LD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_LD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_LD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_UD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_LD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		Q		:  out STD_ULOGIC;
		UD		:  in    STD_ULOGIC;
		FCI		:  in    STD_ULOGIC;
		LD		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		FCO		:  out    STD_ULOGIC);

 end component;


------ Component SUB1 ------
 component SUB1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		FCI		: in    STD_ULOGIC;
		S		: out    STD_ULOGIC;
		FCO		: out    STD_ULOGIC);
 end component;


------ Component TF1A ------
 component TF1A
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_T_CLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_T_CLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_T_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_T_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge	:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge	:  VitalDelayType := 0.000 ns;
		tipd_CLK	:  VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR	:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_T	:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		T	:  in    STD_ULOGIC;
		CLR	:  in    STD_ULOGIC;
	        CLK	:  in    STD_ULOGIC;
		Q	:  out    STD_ULOGIC);

 end component;


------ Component TF1B ------
 component TF1B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_T_CLK_negedge_negedge	:   VitalDelayType := 0.000 ns;
		thold_T_CLK_negedge_negedge	:   VitalDelayType := 0.000 ns;
		tsetup_T_CLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
		thold_T_CLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge	:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge	:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge	:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge	:  VitalDelayType := 0.000 ns;
		tipd_CLK	:  VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR	:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_T	:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		T	:  in    STD_ULOGIC;
		CLR	:  in    STD_ULOGIC;
	        CLK	:  in    STD_ULOGIC;
		Q	:  out    STD_ULOGIC);

 end component;


------ Component TRIBUFF ------
 component TRIBUFF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_8 ------
 component TRIBUFF_S_8
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_8D ------
 component TRIBUFF_S_8D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_8U ------
 component TRIBUFF_S_8U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_12 ------
 component TRIBUFF_S_12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_12D ------
 component TRIBUFF_S_12D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_12U ------
 component TRIBUFF_S_12U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_16 ------
 component TRIBUFF_S_16
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_16D ------
 component TRIBUFF_S_16D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_16U ------
 component TRIBUFF_S_16U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_24 ------
 component TRIBUFF_S_24
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_24D ------
 component TRIBUFF_S_24D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_24U ------
 component TRIBUFF_S_24U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_8 ------
 component TRIBUFF_F_8
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_8D ------
 component TRIBUFF_F_8D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_8U ------
 component TRIBUFF_F_8U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_12 ------
 component TRIBUFF_F_12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_12D ------
 component TRIBUFF_F_12D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_12U ------
 component TRIBUFF_F_12U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_16 ------
 component TRIBUFF_F_16
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_16D ------
 component TRIBUFF_F_16D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_16U ------
 component TRIBUFF_F_16U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_24 ------
 component TRIBUFF_F_24
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_24D ------
 component TRIBUFF_F_24D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_24U ------
 component TRIBUFF_F_24U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS25 ------
 component TRIBUFF_LVCMOS25
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS25D ------
 component TRIBUFF_LVCMOS25D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS25U ------
 component TRIBUFF_LVCMOS25U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS18 ------
 component TRIBUFF_LVCMOS18
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS18D ------
 component TRIBUFF_LVCMOS18D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS18U ------
 component TRIBUFF_LVCMOS18U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS15 ------
 component TRIBUFF_LVCMOS15
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS15D ------
 component TRIBUFF_LVCMOS15D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS15U ------
 component TRIBUFF_LVCMOS15U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_PCI ------
 component TRIBUFF_PCI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_PCIX ------
 component TRIBUFF_PCIX
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_GTLP33 ------
 component TRIBUFF_GTLP33
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_GTLP25 ------
 component TRIBUFF_GTLP25
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component VCC ------
 component VCC
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True		);
    port(
		Y		: out    STD_ULOGIC);
 end component;


------ Component XA1 ------
 component XA1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XA1A ------
 component XA1A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XA1B ------
 component XA1B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XA1C ------
 component XA1C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XAI1 ------
 component XAI1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XAI1A ------
 component XAI1A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XNOR2 ------
 component XNOR2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XNOR3 ------
 component XNOR3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XNOR4 ------
 component XNOR4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XO1 ------
 component XO1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XO1A ------
 component XO1A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XOR2 ------
 component XOR2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XOR3 ------
 component XOR3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XOR4 ------
 component XOR4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XOR4_FCI ------
 component XOR4_FCI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		FCI		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component ZOR3 ------
 component ZOR3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component ZOR3I ------
 component ZOR3I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOFIFO_BIBUF ------
 component IOFIFO_BIBUF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_AIN_YIN		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_AOUT_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_AIN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_AOUT		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		AIN		: in    STD_ULOGIC;
		AOUT		: in    STD_ULOGIC;
		YIN		: out    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC);
 end component;


------ Component IOI_FCLK_EN_BUFF ------
 component IOI_FCLK_EN_BUFF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_ENOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		ENOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 end component;


------ Component IOI_FCLK_BUFF ------
 component IOI_FCLK_BUFF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 end component;


------ Component IOI_RCLK_EN_BUFF ------
 component IOI_RCLK_EN_BUFF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_ENOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		ENOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 end component;


------ Component IOI_RCLK_BUFF ------
 component IOI_RCLK_BUFF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 end component;


------ Component IOOE_FCLK_EN_BUFF ------
 component IOOE_FCLK_EN_BUFF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_ENOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC;
		ENOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 end component;


------ Component IOOE_FCLK ------
 component IOOE_FCLK
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		: in    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 end component;


------ Component IOOE_RCLK_EN_BUFF ------
 component IOOE_RCLK_EN_BUFF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_ENOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC;
		ENOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 end component;


------ Component IOOE_RCLK_CLR_EN ------
 component IOOE_RCLK_CLR_EN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_CLR_CLROUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_ENOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_CLR		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		CLROUT		: out    STD_ULOGIC;
		ENOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 end component;


------ Component IOOE_RCLK_BUFF ------
 component IOOE_RCLK_BUFF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 end component;


------ Component IOOE_RCLK ------
 component IOOE_RCLK
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		: in    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 end component;


------ Component PLLINT ------
 component PLLINT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component PLLOUT ------
 component PLLOUT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_HSTL_I ------
 component BIBUF_HSTL_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_SSTL3_I ------
 component BIBUF_SSTL3_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_SSTL3_II ------
 component BIBUF_SSTL3_II
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_SSTL2_I ------
 component BIBUF_SSTL2_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_SSTL2_II ------
 component BIBUF_SSTL2_II
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BUFF ------
 component BUFF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKINT ------
 component CLKINT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKINT_W ------
 component CLKINT_W
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKOUT_E ------
 component CLKOUT_E
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKOUT_W ------
 component CLKOUT_W
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component DFM ------
 component DFM
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFM3B ------
 component DFM3B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFM4A ------
 component DFM4A
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFM4B ------
 component DFM4B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFMA ------
 component DFMA
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFMB ------
 component DFMB
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFME1A ------
 component DFME1A
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFME1B ------
 component DFME1B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFME2A ------
 component DFME2A
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFME2B ------
 component DFME2B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFME3A ------
 component DFME3A
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFME3B ------
 component DFME3B
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFMEG ------
 component DFMEG
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFMEH ------
 component DFMEH
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFMPCA ------
 component DFMPCA
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFMPCB ------
 component DFMPCB
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component HCLKMUX ------
 component HCLKMUX
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		
                tpw_A_posedge   : VitalDelayType := 0.000 ns;
                tpw_A_negedge   : VitalDelayType := 0.000 ns;    
                tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOFIFO_INBUF ------
 component IOFIFO_INBUF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOFIFO_OUTBUF ------
 component IOFIFO_OUTBUF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOOE_FCLK_BUFF ------
 component IOOE_FCLK_BUFF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 end component;


------ Component IOOE_OUT_FCLK ------
 component IOOE_OUT_FCLK
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 end component;


------ Component IOOE_OUT_FCLK_CLR_EN ------
 component IOOE_OUT_FCLK_CLR_EN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_ENOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_CLROUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		CLR		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC;
		ENOUT		: out    STD_ULOGIC;
		CLROUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 end component;


------ Component IOOE_OUT_RCLK ------
 component IOOE_OUT_RCLK
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 end component;


------ Component IOOE_OUT_RCLK_CLR_EN ------
 component IOOE_OUT_RCLK_CLR_EN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_ENOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_CLROUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		CLR		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC;
		ENOUT		: out    STD_ULOGIC;
		CLROUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 end component;


------ Component IOOE_FCLK_CLR_EN ------
 component IOOE_FCLK_CLR_EN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_EN_ENOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_CLROUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		EN		: in    STD_ULOGIC;
		CLR		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		ENOUT		: out    STD_ULOGIC;
		CLROUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 end component;


------ Component IOPAD_IN_U ------
 component IOPAD_IN_U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_PAD_posedge		: VitalDelayType := 0.000 ns;
		tpw_PAD_negedge		: VitalDelayType := 0.000 ns;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOPAD_IN_D ------
 component IOPAD_IN_D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_PAD_posedge		: VitalDelayType := 0.000 ns;
		tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOPAD_TRI_U ------
 component IOPAD_TRI_U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_D_posedge	: VitalDelayType := 0.000 ns;
		tpw_D_negedge	: VitalDelayType := 0.000 ns;
		tpw_E_posedge	: VitalDelayType := 0.000 ns;
		tpw_E_negedge       : VitalDelayType := 0.000 ns;
		
                tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component IOPAD_TRI_D ------
 component IOPAD_TRI_D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_D_posedge	: VitalDelayType := 0.000 ns;
	        tpw_D_negedge   : VitalDelayType := 0.000 ns;
		tpw_E_posedge   : VitalDelayType := 0.000 ns;
                tpw_E_negedge 	: VitalDelayType := 0.000 ns;

                tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component IOPAD_BI_U ------
 component IOPAD_BI_U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

		tpw_D_posedge	    : VitalDelayType := 0.000 ns;
	        tpw_D_negedge       : VitalDelayType := 0.000 ns;
		tpw_E_posedge       : VitalDelayType := 0.000 ns;
                tpw_E_negedge 	    : VitalDelayType := 0.000 ns;
		tpw_PAD_posedge     : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge     : VitalDelayType := 0.000 ns;

                tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);

		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOPAD_BI_D ------
 component IOPAD_BI_D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
	
		tpw_E_posedge       : VitalDelayType := 0.000 ns;
                tpw_E_negedge 	    : VitalDelayType := 0.000 ns;
		tpw_D_posedge       : VitalDelayType := 0.000 ns;
                tpw_D_negedge 	    : VitalDelayType := 0.000 ns;
		tpw_PAD_posedge     : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge     : VitalDelayType := 0.000 ns;

        	tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component RCLKMUX ------
 component RCLKMUX
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
	   
                tpw_A_posedge   : VitalDelayType := 0.000 ns;
                tpw_A_negedge   : VitalDelayType := 0.000 ns;
         	tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_HSTL_I ------
 component TRIBUFF_HSTL_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		
                tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_SSTL3_I ------
 component TRIBUFF_SSTL3_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_SSTL3_II ------
 component TRIBUFF_SSTL3_II
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_SSTL2_I ------
 component TRIBUFF_SSTL2_I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_SSTL2_II ------
 component TRIBUFF_SSTL2_II
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;

component BIOFIFO_BIDIRINFIFO 
  GENERIC (
        tipd_A       : VitalDelayType01 := (0.00 ns, 0.00 ns);
        tipd_D       : VitalDelayType01 := (0.00 ns, 0.00 ns);
        tipd_WENB       : VitalDelayType01 := (0.00 ns, 0.00 ns);
        tipd_WCLK     : VitalDelayType01 := (0.00 ns, 0.00 ns);
        tipd_RENB       : VitalDelayType01 := (0.00 ns, 0.00 ns);
        tipd_RCLK     : VitalDelayType01 := (0.00 ns, 0.00 ns);
        tipd_CLRB      : VitalDelayType01 := (0.00 ns, 0.00 ns);
        tpd_A_Y   : VitalDelayType01 := (0.1000 ns, 0.1000 ns);
        tpd_RCLK_Q   : VitalDelayType01 := (0.1000 ns, 0.1000 ns);
        tpd_CLRB_Q    : VitalDelayType01 := (0.1000 ns, 0.1000 ns);
        tsetup_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_D_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_negedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLRB_WCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLRB_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True
        );
  PORT (
        A     : IN STD_ULOGIC ;
        D     : IN STD_ULOGIC ;
        WENB     : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RENB     : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        CLRB    : IN STD_ULOGIC ;
        Q     : OUT STD_ULOGIC ;
        Y     : OUT STD_ULOGIC
        );

  
end component;


component BIOFIFO_BIDIROUTFIFO 
  GENERIC (
        tipd_A       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_D       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_CLRB      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_A_Y   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_Q   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLRB_Q    : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tsetup_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_D_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_negedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLRB_WCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLRB_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True
        );
  PORT (
        A     : IN STD_ULOGIC ;
        D     : IN STD_ULOGIC ;
        WENB     : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RENB     : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        CLRB    : IN STD_ULOGIC ;
        Q     : OUT STD_ULOGIC ;
        Y     : OUT STD_ULOGIC
        );

  
end component;


component BIOFIFO_INFIFO 
  GENERIC (
        tipd_D       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_CLRB      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_Q   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLRB_Q    : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tsetup_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_negedge_posedge     :   VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLRB_WCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLRB_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True
        );
  PORT (
        D     : IN STD_ULOGIC ;
        WENB     : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RENB     : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        CLRB    : IN STD_ULOGIC ;
        Q     : OUT STD_ULOGIC
        );

  
end component;

component BIOFIFO_OUTFIFO 
  GENERIC (
        tipd_D       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_CLRB      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_Q   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLRB_Q    : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tsetup_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_negedge_posedge     :   VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLRB_WCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLRB_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True
        );
  PORT (
        D     : IN STD_ULOGIC ;
        WENB     : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RENB     : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        CLRB    : IN STD_ULOGIC ;
        Q     : OUT STD_ULOGIC
        );


end component;


component IOFIFO_BIDIRINFIFO 
  GENERIC (
        tipd_A       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_D       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_CLRB      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_A_Y   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_Q   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLRB_Q    : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tsetup_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_D_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_negedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLRB_WCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLRB_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True
        );
  PORT (
        A     : IN STD_ULOGIC ;
        D     : IN STD_ULOGIC ;
        WENB     : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RENB     : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        CLRB    : IN STD_ULOGIC ;
        Q     : OUT STD_ULOGIC ;
        Y     : OUT STD_ULOGIC
        );


  
end component;


component IOFIFO_BIDIROUTFIFO 
  GENERIC (
        tipd_A       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_D       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_CLRB      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_A_Y   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_Q   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLRB_Q    : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tsetup_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_D_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_negedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLRB_WCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLRB_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True
        );
  PORT (
        A     : IN STD_ULOGIC ;
        D     : IN STD_ULOGIC ;
        WENB     : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RENB     : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        CLRB    : IN STD_ULOGIC ;
        Q     : OUT STD_ULOGIC ;
        Y     : OUT STD_ULOGIC
        );

  
end component;


component IOFIFO_INFIFO 
  GENERIC (
        tipd_D       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_CLRB      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_Q   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLRB_Q    : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tsetup_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_negedge_posedge     :   VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLRB_WCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLRB_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True
        );
  PORT (
        D     : IN STD_ULOGIC ;
        WENB     : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RENB     : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        CLRB    : IN STD_ULOGIC ;
        Q     : OUT STD_ULOGIC
        );

  
end component;

component IOFIFO_OUTFIFO 
  GENERIC (
        tipd_D       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_CLRB      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_Q   : VitalDelayType01 := (0.1000 ns, 0.100 ns);
        tpd_CLRB_Q    : VitalDelayType01 := (0.1000 ns, 0.1000 ns);
        tsetup_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_negedge_posedge     :   VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLRB_WCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLRB_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True
        );
  PORT (
        D     : IN STD_ULOGIC ;
        WENB     : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RENB     : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        CLRB    : IN STD_ULOGIC ;
        Q     : OUT STD_ULOGIC
        );

  
end component;

component IOPADP_IN
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      
      tpw_PAD_posedge 		: VitalDelayType := 0.000 ns;
      tpw_PAD_negedge           : VitalDelayType := 0.000 ns;
      tpw_N2PIN_posedge 	: VitalDelayType := 0.000 ns;
      tpw_N2PIN_negedge         : VitalDelayType := 0.000 ns;   

      tpd_PAD_Y                 :        VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_N2PIN_Y               :        VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PAD         	     :        VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_N2PIN       	     :        VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :        in    STD_ULOGIC;
      N2PIN                          :        in    STD_ULOGIC;
      Y                              :        out   STD_ULOGIC);

end component;


component IOPADN_IN 
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      
      tpw_PAD_posedge 		: VitalDelayType := 0.000 ns;
      tpw_PAD_negedge           : VitalDelayType := 0.000 ns;
 
      tpd_PAD_N2POUT                 :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PAD                       	     :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      N2POUT                         :	out   STD_ULOGIC);

end component;

component IOPADP_TRI 
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpw_E_posedge           : VitalDelayType := 0.000 ns;
      tpw_E_negedge           : VitalDelayType := 0.000 ns;
      tpw_D_posedge           : VitalDelayType := 0.000 ns;
      tpw_D_negedge           : VitalDelayType := 0.000 ns;
      
tpd_E_PAD                      :	VitalDelayType01z := 
               (0.100 ns, 0.100 ns, 0.100 ns, 0.000 ns, 0.100 ns, 0.100 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);

end component;

component IOPADN_TRI 
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      
      tpw_DB_posedge 	    :   VitalDelayType := 0.000 ns;
      tpw_DB_negedge            :   VitalDelayType := 0.000 ns;
      tpw_E_posedge 		: VitalDelayType := 0.000 ns;
      tpw_E_negedge           : VitalDelayType := 0.000 ns;

      tpd_E_PAD                     :	VitalDelayType01z := 
               (0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns);
      tpd_DB_PAD                      :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_DB                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      DB                             :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);

end component;


component CLKBUF_LVDS 
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                             :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);

end component;

component CLKBUF_LVPECL 
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                             :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);

end component;

component HCLKBUF_LVDS 
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                             :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);

end component;

component HCLKBUF_LVPECL 
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                             :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);

end component;

component INBUF_LVDS 
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                             :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);

end component;

component INBUF_LVPECL 
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                             :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);

end component;

component OUTBUF_LVDS 
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_PADP                     :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D_PADN                     :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_D                                 :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      PADP                           :	out   STD_ULOGIC;
      PADN                           :	out   STD_ULOGIC);

end component;

component OUTBUF_LVPECL 
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_PADP                     :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D_PADN                     :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      PADP                           :	out   STD_ULOGIC;
      PADN                           :	out   STD_ULOGIC);

end component;


component CM8F
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S11_Y                      :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_S10_Y                      :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_S01_Y                      :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_S00_Y                      :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_S11_FY                     :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_S10_FY                     :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_S01_FY                     :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_S00_FY                     :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D3_FY                      :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D2_FY                      :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D1_FY                      :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D0_FY                      :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S00                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S01                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S00                            :	in    STD_ULOGIC;
      S01                            :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      FY                             :	out   STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component FIFO64K36 
  GENERIC (
        tipd_DEPTH3   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH2   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH1   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH0   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WIDTH2   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WIDTH1   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WIDTH0   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AEVAL7   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AEVAL6   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AEVAL5   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AEVAL4   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AEVAL3   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AEVAL2   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AEVAL1   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AEVAL0   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AFVAL7   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AFVAL6   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AFVAL5   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AFVAL4   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AFVAL3   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AFVAL2   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AFVAL1   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AFVAL0   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_REN      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD35     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD34     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD33     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD32     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD31     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD30     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD29     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD28     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD27     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD26     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD25     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD24     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD23     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD22     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD21     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD20     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD19     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD18     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD17     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD16     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD15     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD14     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD13     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD12     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD11     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD10     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD9      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD8      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD7      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD6      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD5      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD4      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD3      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WEN      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_CLR      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD1  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD2  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD3  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD4  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD5  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD6  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD7  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD8  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD9  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD10 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD11 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD12 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD13 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD14 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD15 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD16 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD17 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD18 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD19 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD20 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD21 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD22 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD23 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD24 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD25 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD26 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD27 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD28 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD29 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD30 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD31 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD32 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD33 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD34 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD35 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_FULL   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_AFULL  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_EMPTY  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_AEMPTY : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD0  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD1  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD2  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD3  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD4  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD5  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD6  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD7  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD8  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD9  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD10 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD11 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD12 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD13 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD14 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD15 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD16 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD17 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD18 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD19 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD20 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD21 : VitalDelayType01 := (0.100 ns, 0.10 ns);
        tpd_CLR_RD22 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD23 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD24 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD25 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD26 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD27 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD28 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD29 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD30 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD31 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD32 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD33 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD34 : VitalDelayType01 := (0.1000 ns, 0.100 ns);
        tpd_CLR_RD35 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_FULL   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_AFULL  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_EMPTY  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_AEMPTY : VitalDelayType01 := (0.100 ns, 0.100 ns);


        tsetup_WD35_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD34_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD33_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD32_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD31_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD30_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD29_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD28_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD27_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD26_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD25_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD24_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD23_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD22_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD21_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD20_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD19_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD18_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD17_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD16_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD15_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD14_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD13_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD12_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD11_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD10_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD9_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD8_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD35_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD34_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD33_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD32_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD31_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD30_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD29_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD28_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD27_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD26_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD25_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD24_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD23_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD22_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD21_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD20_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD19_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD18_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD17_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD16_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD15_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD14_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD13_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD12_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD11_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD10_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD9_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD8_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;

        tsetup_WEN_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

        tsetup_DEPTH3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        tsetup_WIDTH2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_AEVAL7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_AFVAL7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_DEPTH3_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH3_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        tsetup_WIDTH2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        tsetup_AEVAL7_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL6_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL5_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL4_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL3_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL7_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL6_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL5_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL4_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL3_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_AFVAL7_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL6_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL5_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL4_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL3_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL7_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL6_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL5_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL4_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL3_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_REN_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

        thold_WD35_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD34_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD33_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD32_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD31_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD30_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD29_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD28_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD27_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD26_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD25_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD24_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD23_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD22_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD21_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD20_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD19_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD18_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD17_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD16_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD15_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD14_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD13_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD12_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD11_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD10_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD9_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD8_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD35_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD34_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD33_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD32_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD31_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD30_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD29_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD28_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD27_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD26_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD25_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD24_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD23_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD22_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD21_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD20_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD19_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD18_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD17_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD16_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD15_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD14_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD13_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD12_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD11_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD10_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD9_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD8_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;


        thold_WEN_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

        thold_DEPTH3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        thold_WIDTH2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        thold_AEVAL7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        thold_AFVAL7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;



        thold_DEPTH3_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH3_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        thold_WIDTH2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        thold_AEVAL7_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL6_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL5_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL4_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL3_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL7_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL6_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL5_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL4_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL3_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        thold_AFVAL7_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL6_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL5_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL4_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL3_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL7_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL6_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL5_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL4_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL3_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        thold_REN_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

        trecovery_CLR_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLR_RCLK_posedge_posedge      :  VitalDelayType := 0.000 ns;

        trecovery_CLR_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLR_WCLK_posedge_posedge      :  VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLR_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True
        );
  PORT (
        DEPTH3 : IN STD_ULOGIC ;
        DEPTH2 : IN STD_ULOGIC ;
        DEPTH1 : IN STD_ULOGIC ;
        DEPTH0 : IN STD_ULOGIC ;
        WIDTH2 : IN STD_ULOGIC ;
        WIDTH1 : IN STD_ULOGIC ;
        WIDTH0 : IN STD_ULOGIC ;
        AEVAL7 : IN STD_ULOGIC ;
        AEVAL6 : IN STD_ULOGIC ;
        AEVAL5 : IN STD_ULOGIC ;
        AEVAL4 : IN STD_ULOGIC ;
        AEVAL3 : IN STD_ULOGIC ;
        AEVAL2 : IN STD_ULOGIC ;
        AEVAL1 : IN STD_ULOGIC ;
        AEVAL0 : IN STD_ULOGIC ;
        AFVAL7 : IN STD_ULOGIC ;
        AFVAL6 : IN STD_ULOGIC ;
        AFVAL5 : IN STD_ULOGIC ;
        AFVAL4 : IN STD_ULOGIC ;
        AFVAL3 : IN STD_ULOGIC ;
        AFVAL2 : IN STD_ULOGIC ;
        AFVAL1 : IN STD_ULOGIC ;
        AFVAL0 : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        WD35   : IN STD_ULOGIC ;
        WD34   : IN STD_ULOGIC ;
        WD33   : IN STD_ULOGIC ;
        WD32   : IN STD_ULOGIC ;
        WD31   : IN STD_ULOGIC ;
        WD30   : IN STD_ULOGIC ;
        WD29   : IN STD_ULOGIC ;
        WD28   : IN STD_ULOGIC ;
        WD27   : IN STD_ULOGIC ;
        WD26   : IN STD_ULOGIC ;
        WD25   : IN STD_ULOGIC ;
        WD24   : IN STD_ULOGIC ;
        WD23   : IN STD_ULOGIC ;
        WD22   : IN STD_ULOGIC ;
        WD21   : IN STD_ULOGIC ;
        WD20   : IN STD_ULOGIC ;
        WD19   : IN STD_ULOGIC ;
        WD18   : IN STD_ULOGIC ;
        WD17   : IN STD_ULOGIC ;
        WD16   : IN STD_ULOGIC ;
        WD15   : IN STD_ULOGIC ;
        WD14   : IN STD_ULOGIC ;
        WD13   : IN STD_ULOGIC ;
        WD12   : IN STD_ULOGIC ;
        WD11   : IN STD_ULOGIC ;
        WD10   : IN STD_ULOGIC ;
        WD9    : IN STD_ULOGIC ;
        WD8    : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        CLR    : IN STD_ULOGIC ;
        RD35   : OUT STD_ULOGIC ;
        RD34   : OUT STD_ULOGIC ;
        RD33   : OUT STD_ULOGIC ;
        RD32   : OUT STD_ULOGIC ;
        RD31   : OUT STD_ULOGIC ;
        RD30   : OUT STD_ULOGIC ;
        RD29   : OUT STD_ULOGIC ;
        RD28   : OUT STD_ULOGIC ;
        RD27   : OUT STD_ULOGIC ;
        RD26   : OUT STD_ULOGIC ;
        RD25   : OUT STD_ULOGIC ;
        RD24   : OUT STD_ULOGIC ;
        RD23   : OUT STD_ULOGIC ;
        RD22   : OUT STD_ULOGIC ;
        RD21   : OUT STD_ULOGIC ;
        RD20   : OUT STD_ULOGIC ;
        RD19   : OUT STD_ULOGIC ;
        RD18   : OUT STD_ULOGIC ;
        RD17   : OUT STD_ULOGIC ;
        RD16   : OUT STD_ULOGIC ;
        RD15   : OUT STD_ULOGIC ;
        RD14   : OUT STD_ULOGIC ;
        RD13   : OUT STD_ULOGIC ;
        RD12   : OUT STD_ULOGIC ;
        RD11   : OUT STD_ULOGIC ;
        RD10   : OUT STD_ULOGIC ;
        RD9    : OUT STD_ULOGIC ;
        RD8    : OUT STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC ;
        RD6    : OUT STD_ULOGIC ;
        RD5    : OUT STD_ULOGIC ;
        RD4    : OUT STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC ;
        RD2    : OUT STD_ULOGIC ;
        RD1    : OUT STD_ULOGIC ;
        RD0    : OUT STD_ULOGIC ;
        FULL   : OUT STD_ULOGIC ;
        AFULL  : OUT STD_ULOGIC ;
        EMPTY  : OUT STD_ULOGIC ;
        AEMPTY : OUT STD_ULOGIC
        );


  
end component;

component RAM64K36 
  GENERIC (
        tipd_DEPTH3   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH2   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH1   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH0   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD15   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD14   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD13   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD12   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD11   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD10   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD9    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD8    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD7    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD6    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD5    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD35     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD34     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD33     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD32     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD31     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD30     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD29     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD28     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD27     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD26     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD25     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD24     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD23     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD22     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD21     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD20     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD19     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD18     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD17     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD16     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD15     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD14     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD13     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD12     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD11     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD10     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD9      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD8      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD7      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD6      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD5      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD4      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD3      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WW2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WW1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WW0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WEN      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD15   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD14   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD13   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD12   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD11   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD10   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD9    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD8    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD7    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD6    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD5    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD4    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RW2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RW1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RW0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_REN      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);


        tpd_RCLK_RD0  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD1  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD2  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD3  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD4  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD5  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD6  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD7  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD8  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD9  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD10 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD11 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD12 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD13 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD14 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD15 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD16 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD17 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD18 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD19 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD20 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD21 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD22 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD23 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD24 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD25 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD26 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD27 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD28 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD29 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD30 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD31 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD32 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD33 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD34 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD35 : VitalDelayType01 := (0.100 ns, 0.100 ns);


        tsetup_RDAD15_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD14_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD13_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD12_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD11_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD10_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD9_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD8_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD7_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD6_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD5_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD4_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_RDAD15_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD14_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD13_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD12_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD11_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD10_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD9_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD8_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD7_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD6_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD5_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD4_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        tsetup_RW2_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW1_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW0_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW2_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW1_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW0_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;


        tsetup_DEPTH3_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH2_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH1_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH0_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH3_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH2_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH1_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH0_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;



        tsetup_WRAD15_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD14_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD13_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD12_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD11_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD10_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD9_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD8_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_WRAD15_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD14_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD13_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD12_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD11_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD10_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD9_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD8_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_WD35_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD34_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD33_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD32_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD31_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD30_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD29_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD28_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD27_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD26_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD25_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD24_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD23_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD22_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD21_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD20_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD19_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD18_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD17_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD16_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD15_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD14_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD13_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD12_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD11_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD10_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD9_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD8_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD35_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD34_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD33_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD32_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD31_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD30_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD29_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD28_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD27_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD26_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD25_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD24_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD23_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD22_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD21_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD20_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD19_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD18_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD17_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD16_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD15_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD14_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD13_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD12_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD11_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD10_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD9_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD8_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;


        tsetup_WW2_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW2_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;


        thold_RDAD15_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD14_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD13_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD12_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD11_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD10_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD9_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD8_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD7_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD6_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD5_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;

        thold_RDAD15_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD14_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD13_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD12_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD11_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD10_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD9_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD8_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD7_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD6_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD5_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;



        thold_RW2_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW1_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW0_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW2_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW1_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW0_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

        thold_DEPTH3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        thold_WRAD15_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD14_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD13_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD12_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD11_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD10_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD9_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD8_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;

        thold_WRAD15_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD14_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD13_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD12_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD11_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD10_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD9_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD8_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        thold_WD35_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD34_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD33_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD32_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD31_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD30_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD29_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD28_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD27_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD26_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD25_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD24_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD23_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD22_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD21_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD20_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD19_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD18_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD17_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD16_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD15_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD14_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD13_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD12_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD11_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD10_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD9_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD8_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD35_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD34_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD33_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD32_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD31_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD30_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD29_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD28_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD27_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD26_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD25_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD24_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD23_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD22_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD21_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD20_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD19_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD18_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD17_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD16_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD15_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD14_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD13_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD12_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD11_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD10_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD9_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD8_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;


        thold_WW2_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW1_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW0_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW2_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW1_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW0_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

        tsetup_REN_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True
        );
  PORT (
        DEPTH3 : IN STD_ULOGIC ;
        DEPTH2 : IN STD_ULOGIC ;
        DEPTH1 : IN STD_ULOGIC ;
        DEPTH0 : IN STD_ULOGIC ;
        WRAD15 : IN STD_ULOGIC ;
        WRAD14 : IN STD_ULOGIC ;
        WRAD13 : IN STD_ULOGIC ;
        WRAD12 : IN STD_ULOGIC ;
        WRAD11 : IN STD_ULOGIC ;
        WRAD10 : IN STD_ULOGIC ;
        WRAD9  : IN STD_ULOGIC ;
        WRAD8  : IN STD_ULOGIC ;
        WRAD7  : IN STD_ULOGIC ;
        WRAD6  : IN STD_ULOGIC ;
        WRAD5  : IN STD_ULOGIC ;
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD35   : IN STD_ULOGIC ;
        WD34   : IN STD_ULOGIC ;
        WD33   : IN STD_ULOGIC ;
        WD32   : IN STD_ULOGIC ;
        WD31   : IN STD_ULOGIC ;
        WD30   : IN STD_ULOGIC ;
        WD29   : IN STD_ULOGIC ;
        WD28   : IN STD_ULOGIC ;
        WD27   : IN STD_ULOGIC ;
        WD26   : IN STD_ULOGIC ;
        WD25   : IN STD_ULOGIC ;
        WD24   : IN STD_ULOGIC ;
        WD23   : IN STD_ULOGIC ;
        WD22   : IN STD_ULOGIC ;
        WD21   : IN STD_ULOGIC ;
        WD20   : IN STD_ULOGIC ;
        WD19   : IN STD_ULOGIC ;
        WD18   : IN STD_ULOGIC ;
        WD17   : IN STD_ULOGIC ;
        WD16   : IN STD_ULOGIC ;
        WD15   : IN STD_ULOGIC ;
        WD14   : IN STD_ULOGIC ;
        WD13   : IN STD_ULOGIC ;
        WD12   : IN STD_ULOGIC ;
        WD11   : IN STD_ULOGIC ;
        WD10   : IN STD_ULOGIC ;
        WD9    : IN STD_ULOGIC ;
        WD8    : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        WW2    : IN STD_ULOGIC ;
        WW1    : IN STD_ULOGIC ;
        WW0    : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RDAD15 : IN STD_ULOGIC ;
        RDAD14 : IN STD_ULOGIC ;
        RDAD13 : IN STD_ULOGIC ;
        RDAD12 : IN STD_ULOGIC ;
        RDAD11 : IN STD_ULOGIC ;
        RDAD10 : IN STD_ULOGIC ;
        RDAD9  : IN STD_ULOGIC ;
        RDAD8  : IN STD_ULOGIC ;
        RDAD7  : IN STD_ULOGIC ;
        RDAD6  : IN STD_ULOGIC ;
        RDAD5  : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        RW2    : IN STD_ULOGIC ;
        RW1    : IN STD_ULOGIC ;
        RW0    : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD35   : OUT STD_ULOGIC ;
        RD34   : OUT STD_ULOGIC ;
        RD33   : OUT STD_ULOGIC ;
        RD32   : OUT STD_ULOGIC ;
        RD31   : OUT STD_ULOGIC ;
        RD30   : OUT STD_ULOGIC ;
        RD29   : OUT STD_ULOGIC ;
        RD28   : OUT STD_ULOGIC ;
        RD27   : OUT STD_ULOGIC ;
        RD26   : OUT STD_ULOGIC ;
        RD25   : OUT STD_ULOGIC ;
        RD24   : OUT STD_ULOGIC ;
        RD23   : OUT STD_ULOGIC ;
        RD22   : OUT STD_ULOGIC ;
        RD21   : OUT STD_ULOGIC ;
        RD20   : OUT STD_ULOGIC ;
        RD19   : OUT STD_ULOGIC ;
        RD18   : OUT STD_ULOGIC ;
        RD17   : OUT STD_ULOGIC ;
        RD16   : OUT STD_ULOGIC ;
        RD15   : OUT STD_ULOGIC ;
        RD14   : OUT STD_ULOGIC ;
        RD13   : OUT STD_ULOGIC ;
        RD12   : OUT STD_ULOGIC ;
        RD11   : OUT STD_ULOGIC ;
        RD10   : OUT STD_ULOGIC ;
        RD9    : OUT STD_ULOGIC ;
        RD8    : OUT STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC ;
        RD6    : OUT STD_ULOGIC ;
        RD5    : OUT STD_ULOGIC ;
        RD4    : OUT STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC ;
        RD2    : OUT STD_ULOGIC ;
        RD1    : OUT STD_ULOGIC ;
        RD0    : OUT STD_ULOGIC
        );


end component;


component RAM64K36P 
  GENERIC (
        tipd_DEPTH3   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH2   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH1   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH0   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD15   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD14   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD13   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD12   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD11   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD10   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD9    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD8    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD7    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD6    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD5    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD35     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD34     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD33     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD32     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD31     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD30     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD29     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD28     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD27     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD26     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD25     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD24     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD23     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD22     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD21     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD20     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD19     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD18     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD17     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD16     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD15     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD14     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD13     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD12     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD11     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD10     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD9      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD8      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD7      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD6      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD5      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD4      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD3      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WW2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WW1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WW0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WEN      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD15   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD14   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD13   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD12   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD11   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD10   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD9    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD8    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD7    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD6    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD5    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD4    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RW2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RW1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RW0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_REN      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);


        tpd_RCLK_RD0  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD1  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD2  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD3  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD4  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD5  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD6  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD7  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD8  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD9  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD10 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD11 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD12 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD13 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD14 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD15 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD16 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD17 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD18 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD19 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD20 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD21 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD22 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD23 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD24 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD25 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD26 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD27 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD28 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD29 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD30 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD31 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD32 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD33 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD34 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD35 : VitalDelayType01 := (0.100 ns, 0.100 ns);


        tsetup_RDAD15_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD14_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD13_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD12_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD11_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD10_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD9_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD8_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD7_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD6_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD5_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD4_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_RDAD15_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD14_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD13_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD12_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD11_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD10_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD9_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD8_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD7_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD6_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD5_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD4_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;



        tsetup_RW2_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW1_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW0_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW2_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW1_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW0_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;


        tsetup_DEPTH3_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH2_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH1_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH0_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH3_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH2_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH1_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH0_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;



        tsetup_WRAD15_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD14_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD13_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD12_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD11_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD10_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD9_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD8_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_WRAD15_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD14_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD13_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD12_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD11_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD10_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD9_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD8_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        tsetup_WD35_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD34_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD33_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD32_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD31_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD30_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD29_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD28_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD27_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD26_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD25_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD24_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD23_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD22_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD21_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD20_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD19_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD18_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD17_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD16_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD15_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD14_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD13_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD12_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD11_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD10_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD9_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD8_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD35_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD34_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD33_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD32_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD31_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD30_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD29_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD28_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD27_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD26_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD25_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD24_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD23_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD22_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD21_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD20_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD19_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD18_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD17_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD16_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD15_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD14_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD13_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD12_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD11_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD10_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD9_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD8_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;



        tsetup_WW2_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW2_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;


        thold_RDAD15_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD14_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD13_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD12_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD11_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD10_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD9_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD8_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD7_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD6_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD5_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;

        thold_RDAD15_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD14_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD13_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD12_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD11_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD10_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD9_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD8_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD7_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD6_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD5_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;

        thold_RW2_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW1_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW0_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW2_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW1_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW0_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

        thold_DEPTH3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        thold_WRAD15_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD14_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD13_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD12_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD11_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD10_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD9_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD8_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;

        thold_WRAD15_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD14_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD13_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD12_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD11_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD10_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD9_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD8_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        thold_WD35_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD34_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD33_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD32_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD31_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD30_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD29_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD28_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD27_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD26_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD25_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD24_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD23_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD22_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD21_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD20_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD19_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD18_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD17_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD16_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD15_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD14_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD13_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD12_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD11_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD10_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD9_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD8_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD35_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD34_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD33_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD32_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD31_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD30_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD29_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD28_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD27_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD26_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD25_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD24_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD23_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD22_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD21_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD20_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD19_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD18_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD17_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD16_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD15_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD14_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD13_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD12_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD11_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD10_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD9_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD8_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;


        thold_WW2_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW1_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW0_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW2_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW1_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW0_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

        tsetup_REN_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;



        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True
        );
  PORT (
        DEPTH3 : IN STD_ULOGIC ;
        DEPTH2 : IN STD_ULOGIC ;
        DEPTH1 : IN STD_ULOGIC ;
        DEPTH0 : IN STD_ULOGIC ;
        WRAD15 : IN STD_ULOGIC ;
        WRAD14 : IN STD_ULOGIC ;
        WRAD13 : IN STD_ULOGIC ;
        WRAD12 : IN STD_ULOGIC ;
        WRAD11 : IN STD_ULOGIC ;
        WRAD10 : IN STD_ULOGIC ;
        WRAD9  : IN STD_ULOGIC ;
        WRAD8  : IN STD_ULOGIC ;
        WRAD7  : IN STD_ULOGIC ;
        WRAD6  : IN STD_ULOGIC ;
        WRAD5  : IN STD_ULOGIC ;
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD35   : IN STD_ULOGIC ;
        WD34   : IN STD_ULOGIC ;
        WD33   : IN STD_ULOGIC ;
        WD32   : IN STD_ULOGIC ;
        WD31   : IN STD_ULOGIC ;
        WD30   : IN STD_ULOGIC ;
        WD29   : IN STD_ULOGIC ;
        WD28   : IN STD_ULOGIC ;
        WD27   : IN STD_ULOGIC ;
        WD26   : IN STD_ULOGIC ;
        WD25   : IN STD_ULOGIC ;
        WD24   : IN STD_ULOGIC ;
        WD23   : IN STD_ULOGIC ;
        WD22   : IN STD_ULOGIC ;
        WD21   : IN STD_ULOGIC ;
        WD20   : IN STD_ULOGIC ;
        WD19   : IN STD_ULOGIC ;
        WD18   : IN STD_ULOGIC ;
        WD17   : IN STD_ULOGIC ;
        WD16   : IN STD_ULOGIC ;
        WD15   : IN STD_ULOGIC ;
        WD14   : IN STD_ULOGIC ;
        WD13   : IN STD_ULOGIC ;
        WD12   : IN STD_ULOGIC ;
        WD11   : IN STD_ULOGIC ;
        WD10   : IN STD_ULOGIC ;
        WD9    : IN STD_ULOGIC ;
        WD8    : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        WW2    : IN STD_ULOGIC ;
        WW1    : IN STD_ULOGIC ;
        WW0    : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RDAD15 : IN STD_ULOGIC ;
        RDAD14 : IN STD_ULOGIC ;
        RDAD13 : IN STD_ULOGIC ;
        RDAD12 : IN STD_ULOGIC ;
        RDAD11 : IN STD_ULOGIC ;
        RDAD10 : IN STD_ULOGIC ;
        RDAD9  : IN STD_ULOGIC ;
        RDAD8  : IN STD_ULOGIC ;
        RDAD7  : IN STD_ULOGIC ;
        RDAD6  : IN STD_ULOGIC ;
        RDAD5  : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        RW2    : IN STD_ULOGIC ;
        RW1    : IN STD_ULOGIC ;
        RW0    : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD35   : OUT STD_ULOGIC ;
        RD34   : OUT STD_ULOGIC ;
        RD33   : OUT STD_ULOGIC ;
        RD32   : OUT STD_ULOGIC ;
        RD31   : OUT STD_ULOGIC ;
        RD30   : OUT STD_ULOGIC ;
        RD29   : OUT STD_ULOGIC ;
        RD28   : OUT STD_ULOGIC ;
        RD27   : OUT STD_ULOGIC ;
        RD26   : OUT STD_ULOGIC ;
        RD25   : OUT STD_ULOGIC ;
        RD24   : OUT STD_ULOGIC ;
        RD23   : OUT STD_ULOGIC ;
        RD22   : OUT STD_ULOGIC ;
        RD21   : OUT STD_ULOGIC ;
        RD20   : OUT STD_ULOGIC ;
        RD19   : OUT STD_ULOGIC ;
        RD18   : OUT STD_ULOGIC ;
        RD17   : OUT STD_ULOGIC ;
        RD16   : OUT STD_ULOGIC ;
        RD15   : OUT STD_ULOGIC ;
        RD14   : OUT STD_ULOGIC ;
        RD13   : OUT STD_ULOGIC ;
        RD12   : OUT STD_ULOGIC ;
        RD11   : OUT STD_ULOGIC ;
        RD10   : OUT STD_ULOGIC ;
        RD9    : OUT STD_ULOGIC ;
        RD8    : OUT STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC ;
        RD6    : OUT STD_ULOGIC ;
        RD5    : OUT STD_ULOGIC ;
        RD4    : OUT STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC ;
        RD2    : OUT STD_ULOGIC ;
        RD1    : OUT STD_ULOGIC ;
        RD0    : OUT STD_ULOGIC
        );

 
  
end component;

component DDR_OUT
    port(DR, DF, E, CLK, PRE, CLR : in std_logic;  Q : out std_logic) ;
end component; 

component DDR_REG
    port(D, E, CLK, CLR, PRE : in std_logic;  QR, QF : out std_logic) ;
end component; 

component PLL
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;

      f_REFCLK_LOCK          :	Integer := 3; -- Number of REFCLK pulses after which LOCK is raised

      tipd_PWRDWN            :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_REFCLK            :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_LOWFREQ           :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OSC2              :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OSC1              :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OSC0              :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI5             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI4             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI3             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI2             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI1             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI0             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ5             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ4             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ3             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ2             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ1             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ0             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE4        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE3        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE2        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE1        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE0        :	VitalDelayType01 := (0.000 ns, 0.000 ns);

      tpd_REFCLK_CLK1        :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_REFCLK_CLK2        :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_REFCLK_LOCK        :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PWRDWN                  :	in    STD_ULOGIC; -- Active high
      REFCLK                  :	in    STD_ULOGIC;
      LOWFREQ                 : in    STD_ULOGIC; 
      OSC2                    : in    STD_ULOGIC; 
      OSC1                    : in    STD_ULOGIC; 
      OSC0                    : in    STD_ULOGIC; 
      DIVI5                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI4                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI3                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI2                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI1                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI0                   : in    STD_ULOGIC; -- Clock multiplier
      DIVJ5                   : in    STD_ULOGIC; -- Clock divider
      DIVJ4                   : in    STD_ULOGIC; -- Clock divider
      DIVJ3                   : in    STD_ULOGIC; -- Clock divider
      DIVJ2                   : in    STD_ULOGIC; -- Clock divider
      DIVJ1                   : in    STD_ULOGIC; -- Clock divider
      DIVJ0                   : in    STD_ULOGIC; -- Clock divider
      DELAYLINE4              : in    STD_ULOGIC; -- Delay Value
      DELAYLINE3              : in    STD_ULOGIC; -- Delay Value
      DELAYLINE2              : in    STD_ULOGIC; -- Delay Value
      DELAYLINE1              : in    STD_ULOGIC; -- Delay Value
      DELAYLINE0              : in    STD_ULOGIC; -- Delay Value
      LOCK                    :	out   STD_ULOGIC;
      CLK1                    :	out   STD_ULOGIC;
      CLK2                    :	out   STD_ULOGIC);

end component; 

component PLLFB
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;

      f_REFCLK_LOCK          :	Integer := 3; -- Number of REFCLK pulses after which LOCK is raised

      tipd_PWRDWN            :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_REFCLK            :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_FB                :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_LOWFREQ           :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OSC2              :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OSC1              :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OSC0              :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI5             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI4             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI3             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI2             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI1             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI0             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ5             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ4             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ3             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ2             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ1             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ0             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE4        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE3        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE2        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE1        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE0        :	VitalDelayType01 := (0.000 ns, 0.000 ns);

      tpd_REFCLK_CLK1        :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_REFCLK_CLK2        :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_REFCLK_LOCK        :  VitalDelayType01 := (0.000 ns, 0.000 ns));


   port(
      PWRDWN                  :	in    STD_ULOGIC; -- Active high
      REFCLK                  :	in    STD_ULOGIC;
      FB                      :	in    STD_ULOGIC;
      LOWFREQ                 : in    STD_ULOGIC; 
      OSC2                    : in    STD_ULOGIC; 
      OSC1                    : in    STD_ULOGIC; 
      OSC0                    : in    STD_ULOGIC; 
      DIVI5                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI4                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI3                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI2                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI1                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI0                   : in    STD_ULOGIC; -- Clock multiplier
      DIVJ5                   : in    STD_ULOGIC; -- Clock divider
      DIVJ4                   : in    STD_ULOGIC; -- Clock divider
      DIVJ3                   : in    STD_ULOGIC; -- Clock divider
      DIVJ2                   : in    STD_ULOGIC; -- Clock divider
      DIVJ1                   : in    STD_ULOGIC; -- Clock divider
      DIVJ0                   : in    STD_ULOGIC; -- Clock divider
      DELAYLINE4              : in    STD_ULOGIC; -- Delay Value
      DELAYLINE3              : in    STD_ULOGIC; -- Delay Value
      DELAYLINE2              : in    STD_ULOGIC; -- Delay Value
      DELAYLINE1              : in    STD_ULOGIC; -- Delay Value
      DELAYLINE0              : in    STD_ULOGIC; -- Delay Value
      LOCK                    :	out   STD_ULOGIC;
      CLK1                    :	out   STD_ULOGIC;
      CLK2                    :	out   STD_ULOGIC);

end component; 


---------------- CELL:NOR5D ---------------

COMPONENT NOR5D
   port(
          A     : in std_logic;
          B     : in std_logic;
          C     : in std_logic;
          D     : in std_logic;
          E     : in std_logic;
          Y             : out std_logic);
END COMPONENT;




------ Component ADDSUB1 ------
 component ADDSUB1
    generic(
                TimingChecksOn:Boolean :=True;
                Xon: Boolean :=False;
                InstancePath: STRING :="*";
                MsgOn: Boolean :=True;
                tpd_A_S         : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_FCI_S               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_B_S         : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_A_FCO               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_B_FCO               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_AS_FCO              : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_FCI_FCO             : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_A          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_FCI                : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_B          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_AS         : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                A               : in    STD_ULOGIC;
                FCI             : in    STD_ULOGIC;
                B               : in    STD_ULOGIC;
                AS              : in    STD_ULOGIC;
                S               : out    STD_ULOGIC;
                FCO             : out    STD_ULOGIC);
 end component;



---------------- CELL:NAND5D ---------------

COMPONENT NAND5D
   port(
          A     : in std_logic;
          B     : in std_logic;
          C     : in std_logic;
          D     : in std_logic;
          E     : in std_logic;
          Y             : out std_logic);
END COMPONENT;



------ Component FA1A ------
 component FA1A
    generic(
                TimingChecksOn:Boolean :=True;
                Xon: Boolean :=False;
                InstancePath: STRING :="*";
                MsgOn: Boolean :=True;
                tpd_CI_CO               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_B_CO                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_A_CO                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CI_S                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_A_S         : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_B_S         : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_CI         : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_B          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_A          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                CI              : in    STD_ULOGIC;
                B               : in    STD_ULOGIC;
                A               : in    STD_ULOGIC;
                CO              : out    STD_ULOGIC;
                S               : out    STD_ULOGIC);
 end component;



------ Component FA1B ------
 component FA1B
    generic(
                TimingChecksOn:Boolean :=True;
                Xon: Boolean :=False;
                InstancePath: STRING :="*";
                MsgOn: Boolean :=True;
                tpd_A_CO                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_B_CO                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CI_CO               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CI_S                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_A_S         : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_B_S         : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_A          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_B          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CI         : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                A               : in    STD_ULOGIC;
                B               : in    STD_ULOGIC;
                CI              : in    STD_ULOGIC;
                CO              : out    STD_ULOGIC;
                S               : out    STD_ULOGIC);
 end component;



------ Component FA2A ------
 component FA2A
    generic(
                TimingChecksOn:Boolean :=True;
                Xon: Boolean :=False;
                InstancePath: STRING :="*";
                MsgOn: Boolean :=True;
                tpd_CI_CO               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_B_CO                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_A0_CO               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_A1_CO               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_A0_S                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_A1_S                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_B_S         : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CI_S                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_CI         : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_B          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_A0         : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_A1         : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                CI              : in    STD_ULOGIC;
                B               : in    STD_ULOGIC;
                A0              : in    STD_ULOGIC;
                A1              : in    STD_ULOGIC;
                CO              : out    STD_ULOGIC;
                S               : out    STD_ULOGIC);
 end component;

 END COMPONENTS;
--------------------- END OF COMPONENTS PACKAGE SECTION  ----------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;

use IEEE.VITAL_Timing.all;
use IEEE.VITAL_Primitives.all;

package VTABLES is

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

-- CLR_ipd, CLK_delayed, Q_zd, D, E_delayed, PRE_ipd, CLK_ipd
CONSTANT DFEG_Q_tab : VitalStateTableType := (
( L,  x,  x,  x,  x,  x,  x,  x,  L ),
( H,  L,  H,  H,  x,  x,  H,  x,  H ),
( H,  L,  H,  x,  H,  x,  H,  x,  H ),
( H,  L,  x,  H,  L,  x,  H,  x,  H ),
( H,  H,  x,  x,  x,  H,  x,  x,  S ),
( H,  x,  x,  x,  x,  L,  x,  x,  H ),
( H,  x,  x,  x,  x,  H,  L,  x,  S ),
( x,  L,  L,  L,  x,  H,  H,  x,  L ),
( x,  L,  L,  x,  H,  H,  H,  x,  L ),
( x,  L,  x,  L,  L,  H,  H,  x,  L ),
( U,  x,  L,  x,  x,  H,  x,  x,  L ),
( H,  x,  H,  x,  x,  U,  x,  x,  H )); 

-- CLR_ipd, CLK_delayed, T_delayed, Q_zd, CLK_ipd
CONSTANT tflipflop_Q_tab : VitalStateTableType := (
( L,  x,  x,  x,  x,  x,  L ),
( H,  L,  L,  H,  H,  x,  H ),
( H,  L,  H,  L,  H,  x,  H ),
( H,  H,  x,  x,  x,  x,  S ),
( H,  x,  x,  x,  L,  x,  S ),
( x,  L,  L,  L,  H,  x,  L ),
( x,  L,  H,  H,  H,  x,  L ));

-- CLR_ipd, CLK_delayed, PRE_delayed,K_delayed,J_delayed, Q_zd, CLK_ipd
CONSTANT jkflipflop_Q_tab : VitalStateTableType := (
( L,  x,  H,  x,  x,  x,  x,  x,  U ),
( L,  x,  L,  x,  x,  x,  x,  x,  L ),
( H,  L,  x,  L,  H,  x,  H,  x,  H ),
( H,  L,  x,  L,  x,  H,  H,  x,  H ),
( H,  L,  x,  x,  H,  L,  H,  x,  H ),
( H,  H,  L,  x,  x,  x,  x,  x,  S ),
( H,  x,  L,  x,  x,  x,  L,  x,  S ),
( H,  x,  H,  x,  x,  x,  x,  x,  H ),
( x,  L,  L,  H,  L,  x,  H,  x,  L ),
( x,  L,  L,  H,  x,  H,  H,  x,  L ),
( x,  L,  L,  x,  L,  L,  H,  x,  L ),
( U,  x,  L,  x,  x,  L,  x,  x,  L ),
( H,  x,  U,  x,  x,  H,  x,  x,  H ));

CONSTANT JKF2A_Q_tab : VitalStateTableType := (
( L,  x,  x,  x,  x,  x,  x,  L ),
( H,  L,  L,  H,  x,  H,  x,  H ),
( H,  L,  L,  x,  H,  H,  x,  H ),
( H,  L,  x,  H,  L,  H,  x,  H ),
( H,  H,  x,  x,  x,  x,  x,  S ),
( H,  x,  x,  x,  x,  L,  x,  S ),
( x,  L,  H,  L,  x,  H,  x,  L ),
( x,  L,  H,  x,  H,  H,  x,  L ),
( x,  L,  x,  L,  L,  H,  x,  L ),
( U,  x,  x,  x,  L,  x,  x,  L ));

CONSTANT JKF3A_Q_tab : VitalStateTableType := (
( L,  H,  L,  x,  H,  H,  x,  L ),
( L,  H,  x,  H,  H,  H,  x,  L ),
( L,  L,  H,  x,  x,  H,  x,  H ),
( L,  L,  x,  H,  x,  H,  x,  H ),
( L,  x,  L,  L,  H,  H,  x,  L ),
( L,  x,  H,  L,  x,  H,  x,  H ),
( H,  x,  x,  x,  H,  x,  x,  S ),
( x,  x,  x,  x,  L,  x,  x,  H ),
( x,  x,  x,  x,  H,  L,  x,  S ),
( x,  x,  x,  H,  U,  x,  x,  H ));

CONSTANT dlatch_DLE3B_Q_tab : VitalStateTableType := (
( x,  x,  x,  H,  x,  H ),   --active high preset

( H,  x,  x,  L,  x,  S ),   --latch
( x,  H,  x,  L,  x,  S ),   --latch

( L,  L,  H,  L,  x,  H ),   --transparent
( L,  L,  L,  L,  x,  L ),   --transparent

( U,  x,  H,  L,  H,  H ),   --o/p mux pessimism
( x,  U,  H,  L,  H,  H ),   --o/p mux pessimism
( U,  x,  L,  L,  L,  L ),   --o/p mux pessimism
( x,  U,  L,  L,  L,  L ),   --o/p mux pessimism

( L,  L,  H,  U,  x,  H ),   --PRE==X
( H,  x,  x,  U,  H,  H ),   --PRE==X
( x,  H,  x,  U,  H,  H ),   --PRE==X
( L,  U,  H,  U,  H,  H ),   --PRE==X
( U,  L,  H,  U,  H,  H ),   --PRE==X
( U,  U,  H,  U,  H,  H ));  --PRE==X
--G, E, D, P, Qn, Qn+1

CONSTANT dlatch_DLE2B_Q_tab : VitalStateTableType := (
( L,  x,  x,  x,  x,  L ),   --active low clear

( H,  H,  x,  x,  x,  S ),   --latch
( H,  x,  H,  x,  x,  S ),   --latch

( H,  L,  L,  H,  x,  H ),   --transparent
( H,  L,  L,  L,  x,  L ),   --transparent

( H,  x,  x,  L,  L,  L ),   --o/p mux pessimism
( H,  x,  x,  H,  H,  H ),   --o/p mux pessimism

( U,  x,  x,  L,  L,  L ),   --CLR==X, o/p mux pessimism
( U,  H,  x,  x,  L,  L ),   --CLR==X, o/p mux pessimism, latch
( U,  x,  H,  x,  L,  L ),   --CLR==X, o/p mux pessimism, latch
( U,  L,  L,  L,  x,  L ));  --CLR==X, i/p mux pessimism
--C, G, E, D, Qn, Qn+1


CONSTANT dlatch_DL2C_Q_tab : VitalStateTableType := (
( L,  x,  x,  x,  x,  L ),   --active low clear
( H,  x,  x,  H,  x,  H ),   --active high preset

( H,  H,  x,  L,  x,  S ),   --latch
( H,  L,  L,  L,  x,  L ),   --transparent

( U,  L,  L,  L,  x,  L ),   --CLR==U
( U,  H,  x,  L,  L,  L ),   --CLR==U
( x,  U,  L,  L,  L,  L ),   --CLR,G==U

( H,  U,  H,  x,  H,  H ),   --PRE==U/x,G==U
( H,  L,  H,  x,  x,  H ),   --PRE==U/x
( H,  H,  x,  U,  H,  H ));  --PRE==U
--CLR, G, D, PRE, Qn, Qn+1

end VTABLES;



--------------------- END OF VITABLE TABLE SECTION  ----------------



 ---- CELL ADD1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity ADD1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		FCI		: in    STD_ULOGIC;
		S		: out    STD_ULOGIC;
		FCO		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of ADD1 :  entity is TRUE;
 end ADD1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of ADD1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL FCI_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (FCI_ipd, FCI, tipd_FCI);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, FCI_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS S_zd : STD_LOGIC is Results(1);
	ALIAS FCO_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE S_GlitchData  : VitalGlitchDataType;
	VARIABLE FCO_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       S_zd := ( VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) XOR  FCI_ipd );
       FCO_zd := ((( A_ipd  AND  B_ipd ) OR ( A_ipd  AND  FCI_ipd )) OR ( B_ipd  AND  FCI_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => S,
	   GlitchData => S_GlitchData,
	   OutSignalName => "S",
	   OutTemp => S_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_S, true),
	             1 => (B_ipd'last_event,tpd_B_S, true),
	             2 => (FCI_ipd'last_event,tpd_FCI_S, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => FCO,
	   GlitchData => FCO_GlitchData,
	   OutSignalName => "FCO",
	   OutTemp => FCO_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_FCO, true),
	             1 => (B_ipd'last_event,tpd_B_FCO, true),
	             2 => (FCI_ipd'last_event,tpd_FCI_FCO, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_ADD1_VITAL of ADD1 is 
    for VITAL_ACT
    end for;
 end CFG_ADD1_VITAL;



 ---- CELL AND2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND2 :  entity is TRUE;
 end AND2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AND2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( A_ipd  AND  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND2_VITAL of AND2 is 
    for VITAL_ACT
    end for;
 end CFG_AND2_VITAL;



 ---- CELL AND2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND2A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND2A :  entity is TRUE;
 end AND2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AND2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( (NOT A_ipd)  AND  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND2A_VITAL of AND2A is 
    for VITAL_ACT
    end for;
 end CFG_AND2A_VITAL;



 ---- CELL AND2B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND2B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND2B :  entity is TRUE;
 end AND2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AND2B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( (NOT A_ipd)  AND  (NOT B_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND2B_VITAL of AND2B is 
    for VITAL_ACT
    end for;
 end CFG_AND2B_VITAL;



 ---- CELL AND3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND3 :  entity is TRUE;
 end AND3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AND3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  B_ipd ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND3_VITAL of AND3 is 
    for VITAL_ACT
    end for;
 end CFG_AND3_VITAL;



 ---- CELL AND3A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND3A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND3A :  entity is TRUE;
 end AND3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AND3A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  B_ipd ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND3A_VITAL of AND3A is 
    for VITAL_ACT
    end for;
 end CFG_AND3A_VITAL;



 ---- CELL AND3B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND3B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND3B :  entity is TRUE;
 end AND3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AND3B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND3B_VITAL of AND3B is 
    for VITAL_ACT
    end for;
 end CFG_AND3B_VITAL;



 ---- CELL AND3C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND3C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND3C :  entity is TRUE;
 end AND3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AND3C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND3C_VITAL of AND3C is 
    for VITAL_ACT
    end for;
 end CFG_AND3C_VITAL;



 ---- CELL AND4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND4 :  entity is TRUE;
 end AND4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AND4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A_ipd  AND  B_ipd ) AND  C_ipd ) AND  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND4_VITAL of AND4 is 
    for VITAL_ACT
    end for;
 end CFG_AND4_VITAL;



 ---- CELL AND4A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND4A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND4A :  entity is TRUE;
 end AND4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AND4A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  AND  B_ipd ) AND  C_ipd ) AND  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND4A_VITAL of AND4A is 
    for VITAL_ACT
    end for;
 end CFG_AND4A_VITAL;



 ---- CELL AND4B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND4B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND4B :  entity is TRUE;
 end AND4B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AND4B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  C_ipd ) AND  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND4B_VITAL of AND4B is 
    for VITAL_ACT
    end for;
 end CFG_AND4B_VITAL;



 ---- CELL AND4C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND4C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND4C :  entity is TRUE;
 end AND4C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AND4C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  (NOT C_ipd) ) AND  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND4C_VITAL of AND4C is 
    for VITAL_ACT
    end for;
 end CFG_AND4C_VITAL;



 ---- CELL AND4D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND4D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND4D :  entity is TRUE;
 end AND4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AND4D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  (NOT C_ipd) ) AND  (NOT D_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND4D_VITAL of AND4D is 
    for VITAL_ACT
    end for;
 end CFG_AND4D_VITAL;



 ---- CELL AND5A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND5A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND5A :  entity is TRUE;
 end AND5A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AND5A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (((( (NOT A_ipd)  AND  B_ipd ) AND  C_ipd ) AND  D_ipd ) AND  E_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true),
	             4 => (E_ipd'last_event,tpd_E_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND5A_VITAL of AND5A is 
    for VITAL_ACT
    end for;
 end CFG_AND5A_VITAL;



 ---- CELL AND5B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND5B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND5B :  entity is TRUE;
 end AND5B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AND5B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (((( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  C_ipd ) AND  D_ipd ) AND  E_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true),
	             4 => (E_ipd'last_event,tpd_E_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND5B_VITAL of AND5B is 
    for VITAL_ACT
    end for;
 end CFG_AND5B_VITAL;



 ---- CELL AND5C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND5C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND5C :  entity is TRUE;
 end AND5C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AND5C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (((( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  (NOT C_ipd) ) AND  D_ipd ) AND  E_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true),
	             4 => (E_ipd'last_event,tpd_E_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND5C_VITAL of AND5C is 
    for VITAL_ACT
    end for;
 end CFG_AND5C_VITAL;



 ---- CELL AO1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO1 :  entity is TRUE;
 end AO1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO1_VITAL of AO1 is 
    for VITAL_ACT
    end for;
 end CFG_AO1_VITAL;



 ---- CELL AO10 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO10 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO10 :  entity is TRUE;
 end AO10;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO10 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A_ipd  AND  B_ipd ) OR  C_ipd ) AND ( D_ipd  OR  E_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true),
	             4 => (E_ipd'last_event,tpd_E_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO10_VITAL of AO10 is 
    for VITAL_ACT
    end for;
 end CFG_AO10_VITAL;



 ---- CELL AO11 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO11 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO11 :  entity is TRUE;
 end AO11;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO11 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  B_ipd ) OR (( A_ipd  OR  B_ipd ) AND  C_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO11_VITAL of AO11 is 
    for VITAL_ACT
    end for;
 end CFG_AO11_VITAL;



 ---- CELL AO12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO12 :  entity is TRUE;
 end AO12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2( B_ipd ,( A_ipd  AND  (NOT B_ipd) ), (NOT C_ipd) ) OR (( (NOT A_ipd)  AND  B_ipd ) OR ( (NOT A_ipd)  AND  (NOT C_ipd) )));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO12_VITAL of AO12 is 
    for VITAL_ACT
    end for;
 end CFG_AO12_VITAL;



 ---- CELL AO13 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO13 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO13 :  entity is TRUE;
 end AO13;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO13 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A_ipd  AND  B_ipd ) OR ( A_ipd  AND  (NOT C_ipd) )) OR ( B_ipd  AND  (NOT C_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO13_VITAL of AO13 is 
    for VITAL_ACT
    end for;
 end CFG_AO13_VITAL;



 ---- CELL AO14 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO14 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO14 :  entity is TRUE;
 end AO14;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO14 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2(( (NOT A_ipd)  AND  (NOT B_ipd) ), B_ipd , C_ipd ) OR (( A_ipd  AND  B_ipd ) OR ( A_ipd  AND  (NOT C_ipd) )));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO14_VITAL of AO14 is 
    for VITAL_ACT
    end for;
 end CFG_AO14_VITAL;



 ---- CELL AO15 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO15 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO15 :  entity is TRUE;
 end AO15;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO15 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2(( A_ipd  AND  (NOT B_ipd) ),( (NOT A_ipd)  AND  (NOT B_ipd) ), C_ipd ) OR (( (NOT A_ipd)  AND  B_ipd ) AND  C_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO15_VITAL of AO15 is 
    for VITAL_ACT
    end for;
 end CFG_AO15_VITAL;



 ---- CELL AO16 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO16 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO16 :  entity is TRUE;
 end AO16;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO16 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2(( A_ipd  AND  B_ipd ),( (NOT A_ipd)  AND  (NOT B_ipd) ), (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO16_VITAL of AO16 is 
    for VITAL_ACT
    end for;
 end CFG_AO16_VITAL;



 ---- CELL AO17 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO17 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO17 :  entity is TRUE;
 end AO17;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO17 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2(( (NOT A_ipd)  AND  (NOT B_ipd) ),( (NOT A_ipd)  AND  B_ipd ), C_ipd ) OR (( A_ipd  AND  B_ipd ) AND  C_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO17_VITAL of AO17 is 
    for VITAL_ACT
    end for;
 end CFG_AO17_VITAL;



 ---- CELL AO18 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO18 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO18 :  entity is TRUE;
 end AO18;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO18 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  AND  B_ipd ) OR ( (NOT A_ipd)  AND  (NOT C_ipd) )) OR ( B_ipd  AND  (NOT C_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO18_VITAL of AO18 is 
    for VITAL_ACT
    end for;
 end CFG_AO18_VITAL;



 ---- CELL AO1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO1A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO1A :  entity is TRUE;
 end AO1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO1A_VITAL of AO1A is 
    for VITAL_ACT
    end for;
 end CFG_AO1A_VITAL;



 ---- CELL AO1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO1B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO1B :  entity is TRUE;
 end AO1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  B_ipd ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO1B_VITAL of AO1B is 
    for VITAL_ACT
    end for;
 end CFG_AO1B_VITAL;



 ---- CELL AO1C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO1C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO1C :  entity is TRUE;
 end AO1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO1C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  B_ipd ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO1C_VITAL of AO1C is 
    for VITAL_ACT
    end for;
 end CFG_AO1C_VITAL;



 ---- CELL AO1D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO1D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO1D :  entity is TRUE;
 end AO1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO1D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  (NOT B_ipd) ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO1D_VITAL of AO1D is 
    for VITAL_ACT
    end for;
 end CFG_AO1D_VITAL;



 ---- CELL AO1E ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO1E is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO1E :  entity is TRUE;
 end AO1E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO1E is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  (NOT B_ipd) ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO1E_VITAL of AO1E is 
    for VITAL_ACT
    end for;
 end CFG_AO1E_VITAL;



 ---- CELL AO2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO2 :  entity is TRUE;
 end AO2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A_ipd  AND  B_ipd ) OR  C_ipd ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO2_VITAL of AO2 is 
    for VITAL_ACT
    end for;
 end CFG_AO2_VITAL;



 ---- CELL AO2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO2A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO2A :  entity is TRUE;
 end AO2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  AND  B_ipd ) OR  C_ipd ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO2A_VITAL of AO2A is 
    for VITAL_ACT
    end for;
 end CFG_AO2A_VITAL;



 ---- CELL AO2B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO2B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO2B :  entity is TRUE;
 end AO2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO2B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  AND  (NOT B_ipd) ) OR  C_ipd ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO2B_VITAL of AO2B is 
    for VITAL_ACT
    end for;
 end CFG_AO2B_VITAL;



 ---- CELL AO2C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO2C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO2C :  entity is TRUE;
 end AO2C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO2C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  AND  B_ipd ) OR  (NOT C_ipd) ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO2C_VITAL of AO2C is 
    for VITAL_ACT
    end for;
 end CFG_AO2C_VITAL;



 ---- CELL AO2D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO2D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO2D :  entity is TRUE;
 end AO2D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO2D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  AND  (NOT B_ipd) ) OR  (NOT C_ipd) ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO2D_VITAL of AO2D is 
    for VITAL_ACT
    end for;
 end CFG_AO2D_VITAL;



 ---- CELL AO2E ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO2E is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO2E :  entity is TRUE;
 end AO2E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO2E is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  AND  (NOT B_ipd) ) OR  (NOT C_ipd) ) OR  (NOT D_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO2E_VITAL of AO2E is 
    for VITAL_ACT
    end for;
 end CFG_AO2E_VITAL;



 ---- CELL AO3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO3 :  entity is TRUE;
 end AO3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  AND  B_ipd ) AND  C_ipd ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO3_VITAL of AO3 is 
    for VITAL_ACT
    end for;
 end CFG_AO3_VITAL;



 ---- CELL AO3A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO3A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO3A :  entity is TRUE;
 end AO3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO3A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A_ipd  AND  B_ipd ) AND  C_ipd ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO3A_VITAL of AO3A is 
    for VITAL_ACT
    end for;
 end CFG_AO3A_VITAL;



 ---- CELL AO3B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO3B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO3B :  entity is TRUE;
 end AO3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO3B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  C_ipd ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO3B_VITAL of AO3B is 
    for VITAL_ACT
    end for;
 end CFG_AO3B_VITAL;



 ---- CELL AO3C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO3C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO3C :  entity is TRUE;
 end AO3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO3C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  (NOT C_ipd) ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO3C_VITAL of AO3C is 
    for VITAL_ACT
    end for;
 end CFG_AO3C_VITAL;



 ---- CELL AO4A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO4A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO4A :  entity is TRUE;
 end AO4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO4A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2(( B_ipd  AND  C_ipd ),( C_ipd  AND  D_ipd ), (NOT A_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO4A_VITAL of AO4A is 
    for VITAL_ACT
    end for;
 end CFG_AO4A_VITAL;



 ---- CELL AO5A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO5A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO5A :  entity is TRUE;
 end AO5A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO5A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2( B_ipd , C_ipd , (NOT A_ipd) ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO5A_VITAL of AO5A is 
    for VITAL_ACT
    end for;
 end CFG_AO5A_VITAL;



 ---- CELL AO6 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO6 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO6 :  entity is TRUE;
 end AO6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO6 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  B_ipd ) OR ( C_ipd  AND  D_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO6_VITAL of AO6 is 
    for VITAL_ACT
    end for;
 end CFG_AO6_VITAL;



 ---- CELL AO6A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO6A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO6A :  entity is TRUE;
 end AO6A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO6A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  B_ipd ) OR ( C_ipd  AND  (NOT D_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO6A_VITAL of AO6A is 
    for VITAL_ACT
    end for;
 end CFG_AO6A_VITAL;



 ---- CELL AO7 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO7 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO7 :  entity is TRUE;
 end AO7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO7 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (((( A_ipd  AND  B_ipd ) AND  C_ipd ) OR  D_ipd ) OR  E_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true),
	             4 => (E_ipd'last_event,tpd_E_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO7_VITAL of AO7 is 
    for VITAL_ACT
    end for;
 end CFG_AO7_VITAL;



 ---- CELL AO8 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO8 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO8 :  entity is TRUE;
 end AO8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO8 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A_ipd  AND  B_ipd ) OR ( (NOT C_ipd)  AND  (NOT D_ipd) )) OR  E_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true),
	             4 => (E_ipd'last_event,tpd_E_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO8_VITAL of AO8 is 
    for VITAL_ACT
    end for;
 end CFG_AO8_VITAL;



 ---- CELL AO9 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO9 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO9 :  entity is TRUE;
 end AO9;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AO9 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (((( A_ipd  AND  B_ipd ) OR  C_ipd ) OR  D_ipd ) OR  E_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true),
	             4 => (E_ipd'last_event,tpd_E_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO9_VITAL of AO9 is 
    for VITAL_ACT
    end for;
 end CFG_AO9_VITAL;



 ---- CELL AOI1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI1 :  entity is TRUE;
 end AOI1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AOI1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( A_ipd  AND  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI1_VITAL of AOI1 is 
    for VITAL_ACT
    end for;
 end CFG_AOI1_VITAL;



 ---- CELL AOI1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI1A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI1A :  entity is TRUE;
 end AOI1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AOI1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  AND  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI1A_VITAL of AOI1A is 
    for VITAL_ACT
    end for;
 end CFG_AOI1A_VITAL;



 ---- CELL AOI1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI1B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI1B :  entity is TRUE;
 end AOI1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AOI1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( A_ipd  AND  B_ipd ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI1B_VITAL of AOI1B is 
    for VITAL_ACT
    end for;
 end CFG_AOI1B_VITAL;



 ---- CELL AOI1C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI1C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI1C :  entity is TRUE;
 end AOI1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AOI1C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  AND  (NOT B_ipd) ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI1C_VITAL of AOI1C is 
    for VITAL_ACT
    end for;
 end CFG_AOI1C_VITAL;



 ---- CELL AOI1D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI1D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI1D :  entity is TRUE;
 end AOI1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AOI1D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  AND  (NOT B_ipd) ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI1D_VITAL of AOI1D is 
    for VITAL_ACT
    end for;
 end CFG_AOI1D_VITAL;



 ---- CELL AOI2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI2A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI2A :  entity is TRUE;
 end AOI2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AOI2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( (( (NOT A_ipd)  AND  B_ipd ) OR  C_ipd ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI2A_VITAL of AOI2A is 
    for VITAL_ACT
    end for;
 end CFG_AOI2A_VITAL;



 ---- CELL AOI2B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI2B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI2B :  entity is TRUE;
 end AOI2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AOI2B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( (( (NOT A_ipd)  AND  B_ipd ) OR  (NOT C_ipd) ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI2B_VITAL of AOI2B is 
    for VITAL_ACT
    end for;
 end CFG_AOI2B_VITAL;



 ---- CELL AOI3A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI3A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI3A :  entity is TRUE;
 end AOI3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AOI3A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A_ipd  OR  B_ipd ) OR  C_ipd ) AND ( A_ipd  OR  D_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI3A_VITAL of AOI3A is 
    for VITAL_ACT
    end for;
 end CFG_AOI3A_VITAL;



 ---- CELL AOI4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI4 :  entity is TRUE;
 end AOI4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AOI4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( A_ipd  AND  B_ipd ) OR ( C_ipd  AND  D_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI4_VITAL of AOI4 is 
    for VITAL_ACT
    end for;
 end CFG_AOI4_VITAL;



 ---- CELL AOI4A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI4A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI4A :  entity is TRUE;
 end AOI4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AOI4A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( A_ipd  AND  B_ipd ) OR ( (NOT C_ipd)  AND  D_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI4A_VITAL of AOI4A is 
    for VITAL_ACT
    end for;
 end CFG_AOI4A_VITAL;



 ---- CELL AOI5 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI5 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI5 :  entity is TRUE;
 end AOI5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AOI5 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT VitalMUX2(( (NOT A_ipd)  AND  B_ipd ),( A_ipd  AND  (NOT B_ipd) ), C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI5_VITAL of AOI5 is 
    for VITAL_ACT
    end for;
 end CFG_AOI5_VITAL;



 ---- CELL AFCNTECP1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AFCNTECP1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_UD_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_Q_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_UD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		Q		:  out STD_ULOGIC;
		UD		:  in    STD_ULOGIC;
		FCI		:  in    STD_ULOGIC;
		FCO		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of AFCNTECP1 :  entity is TRUE;
 end AFCNTECP1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AFCNTECP1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL UD_ipd  : STD_ULOGIC := 'X';
	SIGNAL FCI_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (UD_ipd, UD, tipd_UD);
	  VitalWireDelay (FCI_ipd, FCI, tipd_FCI);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (UD_ipd, FCI_ipd, PRE_ipd,CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_UD_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_UD_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_FCI_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_FCI_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_1	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);
	ALIAS FCO_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;
	VARIABLE FCO_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_UD_CLK_negedge, 
	 TimingData		=> Tmkr_UD_CLK_negedge, 
	 TestSignal		=> UD_ipd,
	 TestSignalName		=> "UD",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_UD_CLK_posedge_negedge,
	 SetupLow		=> tsetup_UD_CLK_negedge_negedge,
	 HoldHigh		=> thold_UD_CLK_posedge_negedge,
	 HoldLow		=> thold_UD_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/AFCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_FCI_CLK_negedge, 
	 TimingData		=> Tmkr_FCI_CLK_negedge, 
	 TestSignal		=> FCI_ipd,
	 TestSignalName		=> "FCI",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_FCI_CLK_posedge_negedge,
	 SetupLow		=> tsetup_FCI_CLK_negedge_negedge,
	 HoldHigh		=> thold_FCI_CLK_posedge_negedge,
	 HoldLow		=> thold_FCI_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/AFCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (CLR_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "AFCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "AFCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "AFCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "AFCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "AFCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "AFCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_UD_CLK_negedge or 
	 Tviol_FCI_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, Q_zd, NET_0_1, E_delayed, PRE_ipd, CLK_delayed));
   Q_zd := Violation XOR Q_zd;
    --- combinatorial output logic. 
   FCO_zd := ((( Q_zd  AND  UD_ipd ) OR ( Q_zd  AND  FCI_ipd )) OR ( FCI_ipd  AND  UD_ipd ));
         --- now combinatorial logic input to the DFF 
   NET_0_1 := (( Q_zd  XOR  UD_ipd ) XOR  FCI_ipd );
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => FCO,
	 GlitchData => FCO_GlitchData,
	 OutSignalName => "FCO",
	 OutTemp => FCO_zd,
	 Paths => (
	         0 => (UD_ipd'last_event, tpd_UD_FCO, true),
	         1 => (FCI_ipd'last_event, tpd_FCI_FCO, true),
		 2 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		 3 => (CLR_ipd'last_event, tpd_CLR_Q, true),
	           4 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_AFCNTECP1_VITAL of AFCNTECP1 is
   for VITAL_ACT
   end for;
end CFG_AFCNTECP1_VITAL;



 ---- CELL ARCNTECP1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity ARCNTECP1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_UD_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_Q_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_UD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		Q		:  out STD_ULOGIC;
		UD		:  in    STD_ULOGIC;
		FCI		:  in    STD_ULOGIC;
		FCO		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of ARCNTECP1 :  entity is TRUE;
 end ARCNTECP1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of ARCNTECP1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL UD_ipd  : STD_ULOGIC := 'X';
	SIGNAL FCI_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (UD_ipd, UD, tipd_UD);
	  VitalWireDelay (FCI_ipd, FCI, tipd_FCI);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (UD_ipd, FCI_ipd, PRE_ipd,CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_UD_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_UD_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_FCI_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_FCI_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_1	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);
	ALIAS FCO_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;
	VARIABLE FCO_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_UD_CLK_posedge,
	 TimingData		=> Tmkr_UD_CLK_posedge,
	 TestSignal		=> UD_ipd,
	 TestSignalName		=> "UD",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_UD_CLK_posedge_posedge,
	 SetupLow		=> tsetup_UD_CLK_negedge_posedge,
	 HoldHigh		=> thold_UD_CLK_posedge_posedge,
	 HoldLow		=> thold_UD_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/ARCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_FCI_CLK_posedge,
	 TimingData		=> Tmkr_FCI_CLK_posedge,
	 TestSignal		=> FCI_ipd,
	 TestSignalName		=> "FCI",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_FCI_CLK_posedge_posedge,
	 SetupLow		=> tsetup_FCI_CLK_negedge_posedge,
	 HoldHigh		=> thold_FCI_CLK_posedge_posedge,
	 HoldLow		=> thold_FCI_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/ARCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "ARCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "ARCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "ARCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "ARCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "ARCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "ARCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_UD_CLK_posedge or 
	 Tviol_FCI_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, NET_0_1, E_delayed, PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;
    --- combinatorial output logic. 
   FCO_zd := ((( Q_zd  AND  UD_ipd ) OR ( Q_zd  AND  FCI_ipd )) OR ( FCI_ipd  AND  UD_ipd ));
         --- now combinatorial logic input to the DFF 
   NET_0_1 := (( Q_zd  XOR  UD_ipd ) XOR  FCI_ipd );
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => FCO,
	 GlitchData => FCO_GlitchData,
	 OutSignalName => "FCO",
	 OutTemp => FCO_zd,
	 Paths => (
	         0 => (UD_ipd'last_event, tpd_UD_FCO, true),
	         1 => (FCI_ipd'last_event, tpd_FCI_FCO, true),
		 2 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		 3 => (CLR_ipd'last_event, tpd_CLR_Q, true),
	           4 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_ARCNTECP1_VITAL of ARCNTECP1 is
   for VITAL_ACT
   end for;
end CFG_ARCNTECP1_VITAL;



 ---- CELL AFCNTELDCP1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AFCNTELDCP1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_UD_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_LD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_LD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_LD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_LD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_LD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_UD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		LD		:  in    STD_ULOGIC;
		Q		:  out STD_ULOGIC;
		UD		:  in    STD_ULOGIC;
		FCI		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		FCO		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of AFCNTELDCP1 :  entity is TRUE;
 end AFCNTELDCP1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AFCNTELDCP1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL LD_ipd  : STD_ULOGIC := 'X';
	SIGNAL UD_ipd  : STD_ULOGIC := 'X';
	SIGNAL FCI_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (LD_ipd, LD, tipd_LD);
	  VitalWireDelay (UD_ipd, UD, tipd_UD);
	  VitalWireDelay (FCI_ipd, FCI, tipd_FCI);
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (LD_ipd, UD_ipd, FCI_ipd, D_ipd, PRE_ipd,CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_LD_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_LD_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_UD_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_UD_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_FCI_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_FCI_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_4	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);
	ALIAS FCO_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;
	VARIABLE FCO_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_LD_CLK_negedge, 
	 TimingData		=> Tmkr_LD_CLK_negedge, 
	 TestSignal		=> LD_ipd,
	 TestSignalName		=> "LD",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_LD_CLK_posedge_negedge,
	 SetupLow		=> tsetup_LD_CLK_negedge_negedge,
	 HoldHigh		=> thold_LD_CLK_posedge_negedge,
	 HoldLow		=> thold_LD_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/AFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_UD_CLK_negedge, 
	 TimingData		=> Tmkr_UD_CLK_negedge, 
	 TestSignal		=> UD_ipd,
	 TestSignalName		=> "UD",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_UD_CLK_posedge_negedge,
	 SetupLow		=> tsetup_UD_CLK_negedge_negedge,
	 HoldHigh		=> thold_UD_CLK_posedge_negedge,
	 HoldLow		=> thold_UD_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/AFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_FCI_CLK_negedge, 
	 TimingData		=> Tmkr_FCI_CLK_negedge, 
	 TestSignal		=> FCI_ipd,
	 TestSignalName		=> "FCI",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_FCI_CLK_posedge_negedge,
	 SetupLow		=> tsetup_FCI_CLK_negedge_negedge,
	 HoldHigh		=> thold_FCI_CLK_posedge_negedge,
	 HoldLow		=> thold_FCI_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/AFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/AFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (CLR_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "AFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "AFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "AFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "AFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "AFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "AFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_LD_CLK_negedge or 
	 Tviol_UD_CLK_negedge or 
	 Tviol_FCI_CLK_negedge or Tviol_D_CLK_negedge or Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, Q_zd, NET_0_4, E_delayed, PRE_ipd, CLK_delayed));
   Q_zd := Violation XOR Q_zd;
    --- combinatorial output logic. 
   FCO_zd := ((( Q_zd  AND  UD_ipd ) OR ( Q_zd  AND  FCI_ipd )) OR ( FCI_ipd  AND  UD_ipd ));
         --- now combinatorial logic input to the DFF 
   NET_0_4 :=  VitalMUX2((( Q_zd  XOR  UD_ipd ) XOR  FCI_ipd ), D_ipd , (NOT LD_ipd) );
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => FCO,
	 GlitchData => FCO_GlitchData,
	 OutSignalName => "FCO",
	 OutTemp => FCO_zd,
	 Paths => (
	         0 => (UD_ipd'last_event, tpd_UD_FCO, true),
	         1 => (FCI_ipd'last_event, tpd_FCI_FCO, true),
		 2 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		 3 => (CLR_ipd'last_event, tpd_CLR_Q, true),
	           4 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_AFCNTELDCP1_VITAL of AFCNTELDCP1 is
   for VITAL_ACT
   end for;
end CFG_AFCNTELDCP1_VITAL;



 ---- CELL ARCNTELDCP1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity ARCNTELDCP1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_UD_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_LD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_LD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_LD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_LD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_LD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_UD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		LD		:  in    STD_ULOGIC;
		Q		:  out STD_ULOGIC;
		UD		:  in    STD_ULOGIC;
		FCI		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		FCO		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of ARCNTELDCP1 :  entity is TRUE;
 end ARCNTELDCP1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of ARCNTELDCP1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL LD_ipd  : STD_ULOGIC := 'X';
	SIGNAL UD_ipd  : STD_ULOGIC := 'X';
	SIGNAL FCI_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (LD_ipd, LD, tipd_LD);
	  VitalWireDelay (UD_ipd, UD, tipd_UD);
	  VitalWireDelay (FCI_ipd, FCI, tipd_FCI);
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (LD_ipd, UD_ipd, FCI_ipd, D_ipd, PRE_ipd,CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_LD_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_LD_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_UD_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_UD_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_FCI_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_FCI_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_4	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);
	ALIAS FCO_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;
	VARIABLE FCO_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_LD_CLK_posedge,
	 TimingData		=> Tmkr_LD_CLK_posedge,
	 TestSignal		=> LD_ipd,
	 TestSignalName		=> "LD",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_LD_CLK_posedge_posedge,
	 SetupLow		=> tsetup_LD_CLK_negedge_posedge,
	 HoldHigh		=> thold_LD_CLK_posedge_posedge,
	 HoldLow		=> thold_LD_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/ARCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_UD_CLK_posedge,
	 TimingData		=> Tmkr_UD_CLK_posedge,
	 TestSignal		=> UD_ipd,
	 TestSignalName		=> "UD",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_UD_CLK_posedge_posedge,
	 SetupLow		=> tsetup_UD_CLK_negedge_posedge,
	 HoldHigh		=> thold_UD_CLK_posedge_posedge,
	 HoldLow		=> thold_UD_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/ARCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_FCI_CLK_posedge,
	 TimingData		=> Tmkr_FCI_CLK_posedge,
	 TestSignal		=> FCI_ipd,
	 TestSignalName		=> "FCI",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_FCI_CLK_posedge_posedge,
	 SetupLow		=> tsetup_FCI_CLK_negedge_posedge,
	 HoldHigh		=> thold_FCI_CLK_posedge_posedge,
	 HoldLow		=> thold_FCI_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/ARCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/ARCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "ARCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "ARCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "ARCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "ARCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "ARCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "ARCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_LD_CLK_posedge or 
	 Tviol_UD_CLK_posedge or 
	 Tviol_FCI_CLK_posedge or Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, NET_0_4, E_delayed, PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;
    --- combinatorial output logic. 
   FCO_zd := ((( Q_zd  AND  UD_ipd ) OR ( Q_zd  AND  FCI_ipd )) OR ( FCI_ipd  AND  UD_ipd ));
         --- now combinatorial logic input to the DFF 
   NET_0_4 :=  VitalMUX2((( Q_zd  XOR  UD_ipd ) XOR  FCI_ipd ), D_ipd , (NOT LD_ipd) );
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => FCO,
	 GlitchData => FCO_GlitchData,
	 OutSignalName => "FCO",
	 OutTemp => FCO_zd,
	 Paths => (
	         0 => (UD_ipd'last_event, tpd_UD_FCO, true),
	         1 => (FCI_ipd'last_event, tpd_FCI_FCO, true),
		 2 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		 3 => (CLR_ipd'last_event, tpd_CLR_Q, true),
	           4 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_ARCNTELDCP1_VITAL of ARCNTELDCP1 is
   for VITAL_ACT
   end for;
end CFG_ARCNTELDCP1_VITAL;



 ---- CELL AX1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AX1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AX1 :  entity is TRUE;
 end AX1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AX1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  B_ipd ) XOR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AX1_VITAL of AX1 is 
    for VITAL_ACT
    end for;
 end CFG_AX1_VITAL;



 ---- CELL AX1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AX1A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AX1A :  entity is TRUE;
 end AX1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AX1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  AND  B_ipd ) XOR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AX1A_VITAL of AX1A is 
    for VITAL_ACT
    end for;
 end CFG_AX1A_VITAL;



 ---- CELL AX1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AX1B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AX1B :  entity is TRUE;
 end AX1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AX1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  (NOT B_ipd) ) XOR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AX1B_VITAL of AX1B is 
    for VITAL_ACT
    end for;
 end CFG_AX1B_VITAL;



 ---- CELL AX1C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AX1C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AX1C :  entity is TRUE;
 end AX1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AX1C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  B_ipd ) XOR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AX1C_VITAL of AX1C is 
    for VITAL_ACT
    end for;
 end CFG_AX1C_VITAL;



 ---- CELL AX1D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AX1D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AX1D :  entity is TRUE;
 end AX1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AX1D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  AND  (NOT B_ipd) ) XOR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AX1D_VITAL of AX1D is 
    for VITAL_ACT
    end for;
 end CFG_AX1D_VITAL;



 ---- CELL AX1E ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AX1E is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AX1E :  entity is TRUE;
 end AX1E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AX1E is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( A_ipd  AND  B_ipd ) XOR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AX1E_VITAL of AX1E is 
    for VITAL_ACT
    end for;
 end CFG_AX1E_VITAL;



 ---- CELL AXO1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXO1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXO1 :  entity is TRUE;
 end AXO1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AXO1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( B_ipd  AND  (NOT C_ipd) ) OR  VitalMUX2( C_ipd , A_ipd , (NOT B_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXO1_VITAL of AXO1 is 
    for VITAL_ACT
    end for;
 end CFG_AXO1_VITAL;



 ---- CELL AXO2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXO2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXO2 :  entity is TRUE;
 end AXO2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AXO2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( B_ipd  AND  (NOT C_ipd) ) OR  VitalMUX2( C_ipd , (NOT A_ipd) , (NOT B_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXO2_VITAL of AXO2 is 
    for VITAL_ACT
    end for;
 end CFG_AXO2_VITAL;



 ---- CELL AXO3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXO3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXO3 :  entity is TRUE;
 end AXO3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AXO3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT B_ipd)  AND  C_ipd ) OR  VitalMUX2( A_ipd , (NOT C_ipd) , (NOT B_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXO3_VITAL of AXO3 is 
    for VITAL_ACT
    end for;
 end CFG_AXO3_VITAL;



 ---- CELL AXO5 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXO5 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXO5 :  entity is TRUE;
 end AXO5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AXO5 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( B_ipd  AND  C_ipd ) OR  VitalMUX2( (NOT A_ipd) , (NOT C_ipd) , B_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXO5_VITAL of AXO5 is 
    for VITAL_ACT
    end for;
 end CFG_AXO5_VITAL;



 ---- CELL AXO6 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXO6 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXO6 :  entity is TRUE;
 end AXO6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AXO6 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT B_ipd)  AND  (NOT C_ipd) ) OR  VitalMUX2( C_ipd , A_ipd , B_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXO6_VITAL of AXO6 is 
    for VITAL_ACT
    end for;
 end CFG_AXO6_VITAL;



 ---- CELL AXO7 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXO7 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXO7 :  entity is TRUE;
 end AXO7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AXO7 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT B_ipd)  AND  C_ipd ) OR  VitalMUX2( (NOT A_ipd) , (NOT C_ipd) , (NOT B_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXO7_VITAL of AXO7 is 
    for VITAL_ACT
    end for;
 end CFG_AXO7_VITAL;



 ---- CELL AXOI1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXOI1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXOI1 :  entity is TRUE;
 end AXOI1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AXOI1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( B_ipd  AND  (NOT C_ipd) ) OR  VitalMUX2( C_ipd , A_ipd , (NOT B_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXOI1_VITAL of AXOI1 is 
    for VITAL_ACT
    end for;
 end CFG_AXOI1_VITAL;



 ---- CELL AXOI2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXOI2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXOI2 :  entity is TRUE;
 end AXOI2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AXOI2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( B_ipd  AND  (NOT C_ipd) ) OR  VitalMUX2( C_ipd , (NOT A_ipd) , (NOT B_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXOI2_VITAL of AXOI2 is 
    for VITAL_ACT
    end for;
 end CFG_AXOI2_VITAL;



 ---- CELL AXOI3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXOI3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXOI3 :  entity is TRUE;
 end AXOI3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AXOI3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT B_ipd)  AND  C_ipd ) OR  VitalMUX2( A_ipd , (NOT C_ipd) , (NOT B_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXOI3_VITAL of AXOI3 is 
    for VITAL_ACT
    end for;
 end CFG_AXOI3_VITAL;



 ---- CELL AXOI4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXOI4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXOI4 :  entity is TRUE;
 end AXOI4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AXOI4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( B_ipd  AND  C_ipd ) OR  VitalMUX2( A_ipd , (NOT C_ipd) , B_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXOI4_VITAL of AXOI4 is 
    for VITAL_ACT
    end for;
 end CFG_AXOI4_VITAL;



 ---- CELL AXOI5 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXOI5 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXOI5 :  entity is TRUE;
 end AXOI5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AXOI5 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( B_ipd  AND  C_ipd ) OR  VitalMUX2( (NOT A_ipd) , (NOT C_ipd) , B_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXOI5_VITAL of AXOI5 is 
    for VITAL_ACT
    end for;
 end CFG_AXOI5_VITAL;



 ---- CELL AXOI7 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXOI7 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXOI7 :  entity is TRUE;
 end AXOI7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of AXOI7 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT B_ipd)  AND  C_ipd ) OR  VitalMUX2( (NOT A_ipd) , (NOT C_ipd) , (NOT B_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXOI7_VITAL of AXOI7 is 
    for VITAL_ACT
    end for;
 end CFG_AXOI7_VITAL;



 ---- CELL BIBUF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF :  entity is TRUE;
 end BIBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_VITAL of BIBUF is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_VITAL;



 ---- CELL BIBUF_S_8 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_8 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_8 :  entity is TRUE;
 end BIBUF_S_8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_8 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_8_VITAL of BIBUF_S_8 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_8_VITAL;



 ---- CELL BIBUF_S_8D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_8D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_8D :  entity is TRUE;
 end BIBUF_S_8D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_8D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_8D_VITAL of BIBUF_S_8D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_8D_VITAL;



 ---- CELL BIBUF_S_8U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_8U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_8U :  entity is TRUE;
 end BIBUF_S_8U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_8U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_8U_VITAL of BIBUF_S_8U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_8U_VITAL;



 ---- CELL BIBUF_S_12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_12 :  entity is TRUE;
 end BIBUF_S_12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_12_VITAL of BIBUF_S_12 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_12_VITAL;



 ---- CELL BIBUF_S_12D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_12D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_12D :  entity is TRUE;
 end BIBUF_S_12D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_12D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_12D_VITAL of BIBUF_S_12D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_12D_VITAL;



 ---- CELL BIBUF_S_12U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_12U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_12U :  entity is TRUE;
 end BIBUF_S_12U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_12U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_12U_VITAL of BIBUF_S_12U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_12U_VITAL;



 ---- CELL BIBUF_S_16 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_16 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_16 :  entity is TRUE;
 end BIBUF_S_16;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_16 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_16_VITAL of BIBUF_S_16 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_16_VITAL;



 ---- CELL BIBUF_S_16D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_16D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_16D :  entity is TRUE;
 end BIBUF_S_16D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_16D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_16D_VITAL of BIBUF_S_16D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_16D_VITAL;



 ---- CELL BIBUF_S_16U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_16U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_16U :  entity is TRUE;
 end BIBUF_S_16U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_16U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_16U_VITAL of BIBUF_S_16U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_16U_VITAL;



 ---- CELL BIBUF_S_24 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_24 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_24 :  entity is TRUE;
 end BIBUF_S_24;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_24 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_24_VITAL of BIBUF_S_24 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_24_VITAL;



 ---- CELL BIBUF_S_24D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_24D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_24D :  entity is TRUE;
 end BIBUF_S_24D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_24D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_24D_VITAL of BIBUF_S_24D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_24D_VITAL;



 ---- CELL BIBUF_S_24U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_24U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_24U :  entity is TRUE;
 end BIBUF_S_24U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_24U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_24U_VITAL of BIBUF_S_24U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_24U_VITAL;



 ---- CELL BIBUF_F_8 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_8 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_8 :  entity is TRUE;
 end BIBUF_F_8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_8 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_8_VITAL of BIBUF_F_8 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_8_VITAL;



 ---- CELL BIBUF_F_8D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_8D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_8D :  entity is TRUE;
 end BIBUF_F_8D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_8D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_8D_VITAL of BIBUF_F_8D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_8D_VITAL;



 ---- CELL BIBUF_F_8U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_8U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_8U :  entity is TRUE;
 end BIBUF_F_8U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_8U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_8U_VITAL of BIBUF_F_8U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_8U_VITAL;



 ---- CELL BIBUF_F_12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_12 :  entity is TRUE;
 end BIBUF_F_12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_12_VITAL of BIBUF_F_12 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_12_VITAL;



 ---- CELL BIBUF_F_12D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_12D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_12D :  entity is TRUE;
 end BIBUF_F_12D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_12D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_12D_VITAL of BIBUF_F_12D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_12D_VITAL;



 ---- CELL BIBUF_F_12U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_12U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_12U :  entity is TRUE;
 end BIBUF_F_12U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_12U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_12U_VITAL of BIBUF_F_12U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_12U_VITAL;



 ---- CELL BIBUF_F_16 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_16 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_16 :  entity is TRUE;
 end BIBUF_F_16;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_16 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_16_VITAL of BIBUF_F_16 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_16_VITAL;



 ---- CELL BIBUF_F_16D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_16D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_16D :  entity is TRUE;
 end BIBUF_F_16D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_16D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_16D_VITAL of BIBUF_F_16D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_16D_VITAL;



 ---- CELL BIBUF_F_16U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_16U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_16U :  entity is TRUE;
 end BIBUF_F_16U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_16U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_16U_VITAL of BIBUF_F_16U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_16U_VITAL;



 ---- CELL BIBUF_F_24 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_24 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_24 :  entity is TRUE;
 end BIBUF_F_24;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_24 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_24_VITAL of BIBUF_F_24 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_24_VITAL;



 ---- CELL BIBUF_F_24D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_24D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_24D :  entity is TRUE;
 end BIBUF_F_24D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_24D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_24D_VITAL of BIBUF_F_24D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_24D_VITAL;



 ---- CELL BIBUF_F_24U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_24U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_24U :  entity is TRUE;
 end BIBUF_F_24U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_24U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_24U_VITAL of BIBUF_F_24U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_24U_VITAL;



 ---- CELL BIBUF_LVCMOS25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS25 :  entity is TRUE;
 end BIBUF_LVCMOS25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS25_VITAL of BIBUF_LVCMOS25 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS25_VITAL;



 ---- CELL BIBUF_LVCMOS25D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS25D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS25D :  entity is TRUE;
 end BIBUF_LVCMOS25D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS25D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS25D_VITAL of BIBUF_LVCMOS25D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS25D_VITAL;



 ---- CELL BIBUF_LVCMOS25U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS25U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS25U :  entity is TRUE;
 end BIBUF_LVCMOS25U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS25U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS25U_VITAL of BIBUF_LVCMOS25U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS25U_VITAL;



 ---- CELL BIBUF_LVCMOS18 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS18 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS18 :  entity is TRUE;
 end BIBUF_LVCMOS18;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS18 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS18_VITAL of BIBUF_LVCMOS18 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS18_VITAL;



 ---- CELL BIBUF_LVCMOS18D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS18D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS18D :  entity is TRUE;
 end BIBUF_LVCMOS18D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS18D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS18D_VITAL of BIBUF_LVCMOS18D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS18D_VITAL;



 ---- CELL BIBUF_LVCMOS18U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS18U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS18U :  entity is TRUE;
 end BIBUF_LVCMOS18U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS18U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS18U_VITAL of BIBUF_LVCMOS18U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS18U_VITAL;



 ---- CELL BIBUF_LVCMOS15 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS15 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS15 :  entity is TRUE;
 end BIBUF_LVCMOS15;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS15 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS15_VITAL of BIBUF_LVCMOS15 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS15_VITAL;



 ---- CELL BIBUF_LVCMOS15D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS15D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS15D :  entity is TRUE;
 end BIBUF_LVCMOS15D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS15D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS15D_VITAL of BIBUF_LVCMOS15D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS15D_VITAL;



 ---- CELL BIBUF_LVCMOS15U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS15U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS15U :  entity is TRUE;
 end BIBUF_LVCMOS15U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS15U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS15U_VITAL of BIBUF_LVCMOS15U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS15U_VITAL;



 ---- CELL BIBUF_PCI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_PCI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_PCI :  entity is TRUE;
 end BIBUF_PCI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_PCI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_PCI_VITAL of BIBUF_PCI is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_PCI_VITAL;



 ---- CELL BIBUF_PCIX ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_PCIX is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_PCIX :  entity is TRUE;
 end BIBUF_PCIX;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_PCIX is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_PCIX_VITAL of BIBUF_PCIX is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_PCIX_VITAL;



 ---- CELL BIBUF_GTLP33 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_GTLP33 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_GTLP33 :  entity is TRUE;
 end BIBUF_GTLP33;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_GTLP33 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_GTLP33_VITAL of BIBUF_GTLP33 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_GTLP33_VITAL;



 ---- CELL BIBUF_GTLP25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_GTLP25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_GTLP25 :  entity is TRUE;
 end BIBUF_GTLP25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_GTLP25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_GTLP25_VITAL of BIBUF_GTLP25 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_GTLP25_VITAL;



 ---- CELL BUFA ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BUFA is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BUFA :  entity is TRUE;
 end BUFA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BUFA is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BUFA_VITAL of BUFA is 
    for VITAL_ACT
    end for;
 end CFG_BUFA_VITAL;



 ---- CELL BUFD ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BUFD is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BUFD :  entity is TRUE;
 end BUFD;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BUFD is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BUFD_VITAL of BUFD is 
    for VITAL_ACT
    end for;
 end CFG_BUFD_VITAL;


 ---- CELL CLKBIBUF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBIBUF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D			: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E			: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: inout  STD_ULOGIC;
		D		: in     STD_ULOGIC;
		E		: in     STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBIBUF :  entity is TRUE;
 end CLKBIBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKBIBUF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBIBUF_VITAL of CLKBIBUF is 
    for VITAL_ACT
    end for;
 end CFG_CLKBIBUF_VITAL;


 ---- CELL CLKBUF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF :  entity is TRUE;
 end CLKBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKBUF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_VITAL of CLKBUF is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_VITAL;



 ---- CELL CLKBUF_LVCMOS25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_LVCMOS25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_LVCMOS25 :  entity is TRUE;
 end CLKBUF_LVCMOS25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKBUF_LVCMOS25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_LVCMOS25_VITAL of CLKBUF_LVCMOS25 is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_LVCMOS25_VITAL;



 ---- CELL CLKBUF_LVCMOS18 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_LVCMOS18 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_LVCMOS18 :  entity is TRUE;
 end CLKBUF_LVCMOS18;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKBUF_LVCMOS18 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_LVCMOS18_VITAL of CLKBUF_LVCMOS18 is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_LVCMOS18_VITAL;



 ---- CELL CLKBUF_LVCMOS15 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_LVCMOS15 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_LVCMOS15 :  entity is TRUE;
 end CLKBUF_LVCMOS15;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKBUF_LVCMOS15 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_LVCMOS15_VITAL of CLKBUF_LVCMOS15 is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_LVCMOS15_VITAL;



 ---- CELL CLKBUF_PCI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_PCI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_PCI :  entity is TRUE;
 end CLKBUF_PCI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKBUF_PCI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_PCI_VITAL of CLKBUF_PCI is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_PCI_VITAL;



 ---- CELL CLKBUF_PCIX ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_PCIX is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_PCIX :  entity is TRUE;
 end CLKBUF_PCIX;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKBUF_PCIX is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_PCIX_VITAL of CLKBUF_PCIX is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_PCIX_VITAL;



 ---- CELL CLKBUF_GTLP33 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_GTLP33 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_GTLP33 :  entity is TRUE;
 end CLKBUF_GTLP33;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKBUF_GTLP33 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_GTLP33_VITAL of CLKBUF_GTLP33 is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_GTLP33_VITAL;



 ---- CELL CLKBUF_GTLP25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_GTLP25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_GTLP25 :  entity is TRUE;
 end CLKBUF_GTLP25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKBUF_GTLP25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_GTLP25_VITAL of CLKBUF_GTLP25 is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_GTLP25_VITAL;



 ---- CELL CLKBUF_HSTL_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_HSTL_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_HSTL_I :  entity is TRUE;
 end CLKBUF_HSTL_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKBUF_HSTL_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_HSTL_I_VITAL of CLKBUF_HSTL_I is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_HSTL_I_VITAL;



 ---- CELL CLKBUF_SSTL3_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_SSTL3_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_SSTL3_I :  entity is TRUE;
 end CLKBUF_SSTL3_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKBUF_SSTL3_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_SSTL3_I_VITAL of CLKBUF_SSTL3_I is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_SSTL3_I_VITAL;



 ---- CELL CLKBUF_SSTL3_II ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_SSTL3_II is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_SSTL3_II :  entity is TRUE;
 end CLKBUF_SSTL3_II;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKBUF_SSTL3_II is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_SSTL3_II_VITAL of CLKBUF_SSTL3_II is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_SSTL3_II_VITAL;



 ---- CELL CLKBUF_SSTL2_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_SSTL2_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_SSTL2_I :  entity is TRUE;
 end CLKBUF_SSTL2_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKBUF_SSTL2_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_SSTL2_I_VITAL of CLKBUF_SSTL2_I is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_SSTL2_I_VITAL;



 ---- CELL CLKBUF_SSTL2_II ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_SSTL2_II is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_SSTL2_II :  entity is TRUE;
 end CLKBUF_SSTL2_II;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKBUF_SSTL2_II is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_SSTL2_II_VITAL of CLKBUF_SSTL2_II is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_SSTL2_II_VITAL;



 ---- CELL CM7 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CM7 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S0		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CM7 :  entity is TRUE;
 end CM7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CM7 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL S0_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (S0_ipd, S0, tipd_S0);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, S0_ipd, D1_ipd, S10_ipd, S11_ipd, D2_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( VitalMUX2( D0_ipd , D1_ipd , (NOT S0_ipd) ), VitalMUX2( D2_ipd , D3_ipd , (NOT S0_ipd) ), NOT (  S10_ipd  OR  S11_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (S0_ipd'last_event,tpd_S0_Y, true),
	             2 => (D1_ipd'last_event,tpd_D1_Y, true),
	             3 => (S10_ipd'last_event,tpd_S10_Y, true),
	             4 => (S11_ipd'last_event,tpd_S11_Y, true),
	             5 => (D2_ipd'last_event,tpd_D2_Y, true),
	             6 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CM7_VITAL of CM7 is 
    for VITAL_ACT
    end for;
 end CFG_CM7_VITAL;



 ---- CELL CM8 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CM8 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CM8 :  entity is TRUE;
 end CM8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CM8 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, S00_ipd, S01_ipd, D1_ipd, S10_ipd, S11_ipd, D2_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( VitalMUX2( D0_ipd , D1_ipd , NOT (  S00_ipd  AND  S01_ipd )), VitalMUX2( D2_ipd , D3_ipd , NOT (  S00_ipd  AND  S01_ipd )), NOT (  S10_ipd  OR  S11_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (S00_ipd'last_event,tpd_S00_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (D1_ipd'last_event,tpd_D1_Y, true),
	             4 => (S10_ipd'last_event,tpd_S10_Y, true),
	             5 => (S11_ipd'last_event,tpd_S11_Y, true),
	             6 => (D2_ipd'last_event,tpd_D2_Y, true),
	             7 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CM8_VITAL of CM8 is 
    for VITAL_ACT
    end for;
 end CFG_CM8_VITAL;



 ---- CELL CM8BUFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CM8BUFF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
	
                tpw_A_posedge   : VitalDelayType := 0.000 ns;
                tpw_A_negedge   : VitalDelayType := 0.000 ns;
             	tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CM8BUFF :  entity is TRUE;
 end CM8BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CM8BUFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- timing check results
	VARIABLE Pviol_A       : STD_ULOGIC := '0';
	VARIABLE PeriodData_A  : VitalPeriodDataType := VitalPeriodDataInit;

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_A,
              PeriodData     => PeriodData_A,
              TestSignal     => A_ipd,
              TestSignalName => "A",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_A_posedge,
              PulseWidthLow  => tpw_A_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/CM8BUFF",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CM8BUFF_VITAL of CM8BUFF is 
    for VITAL_ACT
    end for;
 end CFG_CM8BUFF_VITAL;



 ---- CELL CM8INV ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CM8INV is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CM8INV :  entity is TRUE;
 end CM8INV;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CM8INV is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  (NOT A_ipd) ;


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CM8INV_VITAL of CM8INV is 
    for VITAL_ACT
    end for;
 end CFG_CM8INV_VITAL;



 ---- CELL CMA9 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMA9 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMA9 :  entity is TRUE;
 end CMA9;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMA9 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, DB_ipd, S01_ipd, S11_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	CONSTANT CMA9_table : VitalTruthTableType(0 to 10, 0 to 5) :=
	-- Input Pattern                   Response
   -- D0   DB   D3   S01  S11          Y
	(( '-', '0', '-', '0', '-',        '1'), --0
	 ( '-', '1', '-', '-', '1',        '0'),
	 ( '-', '0', '0', '1', '-',        '0'),
	 ( '1', '1', '-', '-', '0',        '1'),
	 ( '1', '-', '1', '-', '0',        '1'),
	 ( '-', '0', '1', '-', '-',        '1'), --5
	 ( '0', '1', '-', '-', '-',        '0'),
	 ( '0', '-', '0', '1', '-',        '0'),
	 ( '1', '-', '-', '0', '0',        '1'),
	 ( '-', '0', '1', '1', '-',        '1'),
	 ( '-', '-', '0', '1', '1',        '0')); --10

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
   Y_zd := VitalTruthTable(
            TruthTable => CMA9_table,
             DataIn => (
              D0_ipd, DB_ipd, D3_ipd, S01_ipd, S11_ipd));



	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (DB_ipd'last_event,tpd_DB_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (S11_ipd'last_event,tpd_S11_Y, true),
	             4 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMA9_VITAL of CMA9 is 
    for VITAL_ACT
    end for;
 end CFG_CMA9_VITAL;



 ---- CELL CMAF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMAF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMAF :  entity is TRUE;
 end CMAF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMAF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, DB_ipd, S11_ipd, D2_ipd, S01_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	CONSTANT CMAF_table : VitalTruthTableType(0 to 25, 0 to 6) :=
	  -- Input Pattern                             Response
	  -- D0   D2   D3   DB   S01  S11       Y
	  (( '0', '0', '0', '-', '-', '-',     '0'), --0
	   ( '1', '1', '1', '-', '-', '-',     '1'),
	   ( '0', '0', '-', '-', '0', '0',     '0'),
	   ( '1', '1', '-', '-', '0', '0',     '1'),
	   ( '0', '0', '-', '1', '-', '-',     '0'),
	   ( '1', '1', '-', '1', '-', '-',     '1'), --5
	   ( '0', '0', '-', '-', '0', '-',     '0'),
	   ( '1', '1', '-', '-', '0', '-',     '1'),
	   ( '-', '0', '0', '-', '1', '1',     '0'),
	   ( '-', '1', '1', '-', '1', '1',     '1'),
	   ( '-', '0', '0', '0', '-', '-',     '0'), --10
	   ( '-', '1', '1', '0', '-', '-',     '1'),
	   ( '-', '0', '0', '-', '-', '1',     '0'),
	   ( '-', '1', '1', '-', '-', '1',     '1'),
	   ( '0', '-', '0', '-', '1', '0',     '0'),
	   ( '1', '-', '1', '-', '1', '0',     '1'), --15
	   ( '-', '0', '-', '0', '0', '-',     '0'),
	   ( '-', '1', '-', '0', '0', '-',     '1'),
	   ( '-', '0', '-', '1', '-', '1',     '0'),
	   ( '-', '1', '-', '1', '-', '1',     '1'),
	   ( '-', '0', '-', '-', '0', '1',     '0'), --20
	   ( '-', '1', '-', '-', '0', '1',     '1'),
	   ( '-', '-', '0', '0', '1', '-',     '0'),
	   ( '-', '-', '1', '0', '1', '-',     '1'),
	   ( '0', '-', '-', '1', '-', '0',     '0'),
  	   ( '1', '-', '-', '1', '-', '0',     '1')); --25

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
      Y_zd := VitalTruthTable(
             TruthTable => CMAF_table,
             DataIn => (
              D0_ipd, D2_ipd, D3_ipd, DB_ipd, S01_ipd, S11_ipd));



	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (DB_ipd'last_event,tpd_DB_Y, true),
	             2 => (S11_ipd'last_event,tpd_S11_Y, true),
	             3 => (D2_ipd'last_event,tpd_D2_Y, true),
	             4 => (S01_ipd'last_event,tpd_S01_Y, true),
	             5 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMAF_VITAL of CMAF is 
    for VITAL_ACT
    end for;
 end CFG_CMAF_VITAL;



 ---- CELL CMB3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMB3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMB3 :  entity is TRUE;
 end CMB3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMB3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, S00_ipd, S01_ipd, D1_ipd, DB_ipd, S11_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( VitalMUX2( D0_ipd , D1_ipd , NOT (  S00_ipd  AND  S01_ipd )), VitalMUX2( (NOT DB_ipd) , (NOT DB_ipd) , NOT (  S00_ipd  AND  S01_ipd )), NOT (  (NOT DB_ipd)  OR  S11_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (S00_ipd'last_event,tpd_S00_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (D1_ipd'last_event,tpd_D1_Y, true),
	             4 => (DB_ipd'last_event,tpd_DB_Y, true),
	             5 => (S11_ipd'last_event,tpd_S11_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMB3_VITAL of CMB3 is 
    for VITAL_ACT
    end for;
 end CFG_CMB3_VITAL;



 ---- CELL CMB7 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMB7 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMB7 :  entity is TRUE;
 end CMB7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMB7 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, S00_ipd, S01_ipd, D1_ipd, DB_ipd, S11_ipd, D2_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

  CONSTANT CMB7_table : VitalTruthTableType(0 to 24, 0 to 7) :=
  -- Input Pattern                             Response
  -- D0   D1   D2   DB   S00  S01  S11          Y
  (( '0', '0', '0', '1', '-', '-', '-',        '0'), --0
   ( '-', '-', '1', '0', '-', '-', '-',        '1'),
   ( '-', '0', '-', '1', '1', '1', '0',        '0'),
   ( '-', '1', '-', '-', '1', '1', '0',        '1'),
   ( '0', '-', '-', '1', '0', '-', '0',        '0'),
   ( '0', '-', '-', '1', '-', '0', '0',        '0'), --5
   ( '1', '-', '-', '1', '0', '-', '0',        '1'),
   ( '1', '-', '-', '1', '-', '0', '0',        '1'),
   ( '-', '-', '-', '1', '1', '1', '1',        '0'),
   ( '-', '-', '-', '0', '1', '1', '-',        '1'),
   ( '-', '-', '0', '0', '0', '-', '-',        '0'), --10
   ( '-', '-', '0', '0', '-', '0', '-',        '0'),
   ( '-', '-', '0', '-', '0', '-', '1',        '0'),
   ( '-', '-', '0', '-', '-', '0', '1',        '0'),
   ( '0', '-', '0', '-', '0', '-', '-',        '0'),
   ( '0', '-', '0', '-', '-', '0', '-',        '0'), --15
   ( '1', '-', '1', '-', '0', '-', '-',        '1'),
   ( '1', '-', '1', '-', '-', '0', '-',        '1'),
   ( '-', '-', '1', '-', '0', '-', '1',        '1'),
   ( '-', '-', '1', '-', '-', '0', '1',        '1'),
   ( '-', '0', '-', '1', '1', '1', '-',        '0'), --20
   ( '0', '0', '-', '1', '-', '-', '0',        '0'),
   ( '1', '1', '-', '1', '-', '-', '0',        '1'),
   ( '-', '-', '0', '1', '-', '-', '1',        '0'),
   ( '1', '1', '1', '-', '-', '-', '0',        '1'));

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
    Y_zd := VitalTruthTable (
             TruthTable => CMB7_table,
             DataIn => (
              D0_ipd, D1_ipd, D2_ipd, DB_ipd, S00_ipd, S01_ipd, S11_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (S00_ipd'last_event,tpd_S00_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (D1_ipd'last_event,tpd_D1_Y, true),
	             4 => (DB_ipd'last_event,tpd_DB_Y, true),
	             5 => (S11_ipd'last_event,tpd_S11_Y, true),
	             6 => (D2_ipd'last_event,tpd_D2_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMB7_VITAL of CMB7 is 
    for VITAL_ACT
    end for;
 end CFG_CMB7_VITAL;



 ---- CELL CMBB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMBB is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMBB :  entity is TRUE;
 end CMBB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMBB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, S00_ipd, S01_ipd, D1_ipd, DB_ipd, S11_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

 CONSTANT CMBB_table : VitalTruthTableType(0 to 23, 0 to 7) :=
  -- Input Pattern                             Response
  -- D0   D1   DB   D3   S00  S01  S11          Y
  (( '0', '0', '1', '0', '-', '-', '-',        '0'), --0
   ( '-', '-', '0', '1', '-', '-', '-',        '1'),
   ( '-', '-', '0', '-', '-', '0', '-',        '1'),
   ( '-', '-', '1', '-', '-', '0', '1',        '0'),
   ( '-', '-', '0', '-', '0', '-', '-',        '1'),
   ( '-', '-', '1', '-', '0', '-', '1',        '0'), --5
   ( '0', '-', '1', '-', '-', '0', '0',        '0'),
   ( '1', '-', '-', '-', '-', '0', '0',        '1'),
   ( '0', '-', '1', '-', '0', '-', '0',        '0'),
   ( '1', '-', '-', '-', '0', '-', '0',        '1'),
   ( '-', '0', '1', '-', '1', '1', '0',        '0'), --10
   ( '-', '1', '1', '-', '1', '1', '0',        '1'),
   ( '-', '-', '-', '0', '1', '1', '1',        '0'),
   ( '-', '-', '-', '1', '1', '1', '1',        '1'),
   ( '-', '-', '0', '0', '1', '1', '-',        '0'),
   ( '-', '-', '0', '1', '1', '1', '-',        '1'), --15
   ( '-', '-', '1', '0', '-', '-', '1',        '0'),
   ( '-', '0', '-', '0', '1', '1', '-',        '0'),
   ( '-', '1', '-', '1', '1', '1', '-',        '1'),
   ( '0', '-', '1', '-', '0', '-', '-',        '0'),
   ( '0', '0', '1', '-', '-', '-', '0',        '0'), --20
   ( '1', '1', '1', '-', '-', '-', '0',        '1'),
   ( '0', '-', '1', '-', '-', '0', '-',        '0'),
   ( '1', '1', '-', '1', '-', '-', '0',        '1'));

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
   Y_zd := VitalTruthTable(
           TruthTable => CMBB_table,
             DataIn => (
              D0_ipd, D1_ipd, DB_ipd, D3_ipd, S00_ipd, S01_ipd, S11_ipd));



	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (S00_ipd'last_event,tpd_S00_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (D1_ipd'last_event,tpd_D1_Y, true),
	             4 => (DB_ipd'last_event,tpd_DB_Y, true),
	             5 => (S11_ipd'last_event,tpd_S11_Y, true),
	             6 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMBB_VITAL of CMBB is 
    for VITAL_ACT
    end for;
 end CFG_CMBB_VITAL;



 ---- CELL CMBF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMBF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMBF :  entity is TRUE;
 end CMBF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMBF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, S00_ipd, S01_ipd, D1_ipd, DB_ipd, S11_ipd, D2_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( VitalMUX2( D0_ipd , D1_ipd , NOT (  S00_ipd  AND  S01_ipd )), VitalMUX2( D2_ipd , D3_ipd , NOT (  S00_ipd  AND  S01_ipd )), NOT (  (NOT DB_ipd)  OR  S11_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (S00_ipd'last_event,tpd_S00_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (D1_ipd'last_event,tpd_D1_Y, true),
	             4 => (DB_ipd'last_event,tpd_DB_Y, true),
	             5 => (S11_ipd'last_event,tpd_S11_Y, true),
	             6 => (D2_ipd'last_event,tpd_D2_Y, true),
	             7 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMBF_VITAL of CMBF is 
    for VITAL_ACT
    end for;
 end CFG_CMBF_VITAL;



 ---- CELL CMEA ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMEA is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMEA :  entity is TRUE;
 end CMEA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMEA is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (DB_ipd, S01_ipd, D1_ipd, S10_ipd, S11_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

   CONSTANT CMEA_table : VitalTruthTableType(0 to 14, 0 to 6) :=
         -- Input Pattern                        Response
         -- DB   D1   D3   S01  S10  S11          Y
         (( '1', '-', '-', '-', '-', '-',        '0'), --0
          ( '0', '1', '1', '-', '-', '-',        '1'),
          ( '0', '0', '-', '1', '0', '0',        '0'),
          ( '0', '1', '-', '-', '0', '0',        '1'),
          ( '-', '0', '-', '1', '0', '0',        '0'),
          ( '0', '-', '0', '1', '1', '-',        '0'),
          ( '0', '-', '0', '1', '-', '1',        '0'), --5
          ( '0', '-', '-', '0', '-', '-',        '1'),
          ( '-', '0', '0', '1', '-', '-',        '0'),
          ( '-', '1', '0', '1', '1', '-',        '0'),
          ( '-', '1', '0', '1', '-', '1',        '0'),
          ( '-', '-', '0', '1', '1', '-',        '0'),
          ( '-', '-', '0', '1', '-', '1',        '0'),
          ( '0', '-', '1', '-', '1', '-',        '1'),
          ( '0', '-', '1', '-', '-', '1',        '1'));

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
      Y_zd := VitalTruthTable(
             TruthTable => CMEA_table,
             DataIn => (
              DB_ipd, D1_ipd, D3_ipd, S01_ipd, S10_ipd, S11_ipd));



	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (DB_ipd'last_event,tpd_DB_Y, true),
	             1 => (S01_ipd'last_event,tpd_S01_Y, true),
	             2 => (D1_ipd'last_event,tpd_D1_Y, true),
	             3 => (S10_ipd'last_event,tpd_S10_Y, true),
	             4 => (S11_ipd'last_event,tpd_S11_Y, true),
	             5 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMEA_VITAL of CMEA is 
    for VITAL_ACT
    end for;
 end CFG_CMEA_VITAL;



 ---- CELL CMEB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMEB is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMEB :  entity is TRUE;
 end CMEB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMEB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, DB_ipd, S01_ipd, D1_ipd, S10_ipd, S11_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	CONSTANT CMEB_table : VitalTruthTableType(0 to 24, 0 to 7) :=
	  -- Input Pattern                             Response
	  -- D0   D1   DB   D3   S01  S10  S11          Y
	  (( '0', '0', '1', '0', '-', '-', '-',        '0'), --0
	   ( '1', '1', '0', '1', '-', '-', '-',        '1'),
	   ( '0', '-', '-', '-', '0', '0', '0',        '0'),
	   ( '1', '-', '-', '-', '0', '0', '0',        '1'),
	   ( '0', '-', '1', '-', '-', '0', '0',        '0'),
	   ( '1', '-', '1', '-', '-', '0', '0',        '1'), --5
	   ( '-', '-', '0', '1', '1', '1', '-',        '1'),
	   ( '-', '-', '0', '1', '1', '-', '1',        '1'),
	   ( '-', '0', '0', '-', '1', '0', '0',        '0'),
	   ( '-', '1', '0', '-', '1', '0', '0',        '1'),
 	   ( '-', '-', '-', '0', '1', '1', '-',        '0'), --10
	   ( '-', '-', '-', '0', '1', '-', '1',        '0'),
	   ( '-', '-', '1', '-', '-', '1', '-',        '0'),
	   ( '-', '-', '1', '-', '-', '-', '1',        '0'),
	   ( '-', '-', '0', '-', '0', '1', '-',        '1'),
	   ( '-', '0', '0', '0', '1', '-', '-',        '0'), --15
	   ( '-', '1', '0', '1', '1', '-', '-',        '1'),
	   ( '0', '0', '-', '-', '-', '0', '0',        '0'),
	   ( '1', '1', '-', '-', '-', '0', '0',        '1'),
	   ( '0', '-', '1', '-', '-', '-', '-',        '0'),
	   ( '1', '-', '0', '-', '0', '-', '-',        '1'), --20
	   ( '-', '-', '0', '1', '-', '1', '-',        '1'),
	   ( '-', '-', '0', '1', '-', '-', '1',        '1'),
	   ( '-', '-', '0', '-', '0', '-', '1',        '1'),
	   ( '0', '0', '-', '0', '1', '-', '-',        '0'));

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
    Y_zd := VitalTruthTable(
     TruthTable => CMEB_table,
             DataIn => (
              D0_ipd, D1_ipd, DB_ipd, D3_ipd, S01_ipd, S10_ipd, S11_ipd));



	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (DB_ipd'last_event,tpd_DB_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (D1_ipd'last_event,tpd_D1_Y, true),
	             4 => (S10_ipd'last_event,tpd_S10_Y, true),
	             5 => (S11_ipd'last_event,tpd_S11_Y, true),
	             6 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMEB_VITAL of CMEB is 
    for VITAL_ACT
    end for;
 end CFG_CMEB_VITAL;



 ---- CELL CMEE ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMEE is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMEE :  entity is TRUE;
 end CMEE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMEE is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (DB_ipd, S01_ipd, D1_ipd, S10_ipd, S11_ipd, D2_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	CONSTANT CMEE_table : VitalTruthTableType(0 to 27, 0 to 7) :=
	  -- Input Pattern                             Response
	  -- DB   D1   D2   D3   S01  S10  S11          Y
	  (( '1', '0', '0', '0', '-', '-', '-',        '0'), --0
	   ( '0', '1', '1', '1', '-', '-', '-',        '1'),
	   ( '-', '0', '-', '-', '1', '0', '0',        '0'),
	   ( '0', '1', '-', '-', '1', '0', '0',        '1'),
	   ( '0', '-', '-', '0', '1', '1', '-',        '0'),
	   ( '0', '-', '-', '1', '1', '1', '-',        '1'), --5
	   ( '0', '-', '-', '0', '1', '-', '1',        '0'),
	   ( '0', '-', '-', '1', '1', '-', '1',        '1'),
	   ( '1', '-', '-', '-', '-', '0', '0',        '0'),
	   ( '0', '-', '-', '-', '0', '0', '0',        '1'),
	   ( '-', '-', '0', '-', '0', '-', '1',        '0'), --10
	   ( '-', '-', '1', '-', '0', '-', '1',        '1'),
	   ( '-', '-', '0', '-', '0', '1', '-',        '0'),
	   ( '-', '-', '1', '-', '0', '1', '-',        '1'),
	   ( '1', '-', '0', '-', '-', '-', '1',        '0'),
	   ( '1', '-', '1', '-', '-', '-', '1',        '1'), --15
	   ( '1', '-', '0', '-', '-', '1', '-',        '0'),
	   ( '1', '-', '1', '-', '-', '1', '-',        '1'),
	   ( '1', '-', '0', '-', '-', '-', '-',        '0'),
	   ( '0', '-', '1', '-', '0', '-', '-',        '1'),
	   ( '-', '-', '0', '0', '-', '1', '-',        '0'), --20
	   ( '-', '-', '1', '1', '-', '1', '-',        '1'),
	   ( '-', '-', '0', '0', '-', '-', '1',        '0'),
	   ( '0', '0', '-', '0', '1', '-', '-',        '0'),
	   ( '0', '1', '-', '1', '1', '-', '-',        '1'),
	   ( '-', '-', '1', '1', '-', '-', '1',        '1'), --25
	   ( '0', '1', '-', '-', '-', '0', '0',        '1'),
	   ( '-', '0', '0', '0', '1', '-', '-',        '0'));

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
          Y_zd := VitalTruthTable(
             TruthTable => CMEE_table,
             DataIn => (
              DB_ipd, D1_ipd, D2_ipd, D3_ipd, S01_ipd, S10_ipd, S11_ipd));



	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (DB_ipd'last_event,tpd_DB_Y, true),
	             1 => (S01_ipd'last_event,tpd_S01_Y, true),
	             2 => (D1_ipd'last_event,tpd_D1_Y, true),
	             3 => (S10_ipd'last_event,tpd_S10_Y, true),
	             4 => (S11_ipd'last_event,tpd_S11_Y, true),
	             5 => (D2_ipd'last_event,tpd_D2_Y, true),
	             6 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMEE_VITAL of CMEE is 
    for VITAL_ACT
    end for;
 end CFG_CMEE_VITAL;



 ---- CELL CMEF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMEF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMEF :  entity is TRUE;
 end CMEF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMEF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, DB_ipd, S01_ipd, D1_ipd, S10_ipd, S11_ipd, D2_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( VitalMUX2( D0_ipd , D1_ipd , NOT (  (NOT DB_ipd)  AND  S01_ipd )), VitalMUX2( D2_ipd , D3_ipd , NOT (  (NOT DB_ipd)  AND  S01_ipd )), NOT (  S10_ipd  OR  S11_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (DB_ipd'last_event,tpd_DB_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (D1_ipd'last_event,tpd_D1_Y, true),
	             4 => (S10_ipd'last_event,tpd_S10_Y, true),
	             5 => (S11_ipd'last_event,tpd_S11_Y, true),
	             6 => (D2_ipd'last_event,tpd_D2_Y, true),
	             7 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMEF_VITAL of CMEF is 
    for VITAL_ACT
    end for;
 end CFG_CMEF_VITAL;



 ---- CELL CMF1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMF1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMF1 :  entity is TRUE;
 end CMF1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMF1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, S00_ipd, S01_ipd, DB_ipd, S10_ipd, S11_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( VitalMUX2( D0_ipd , (NOT DB_ipd) , NOT (  S00_ipd  AND  S01_ipd )), (NOT DB_ipd) , NOT (  S10_ipd  OR  S11_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (S00_ipd'last_event,tpd_S00_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (DB_ipd'last_event,tpd_DB_Y, true),
	             4 => (S10_ipd'last_event,tpd_S10_Y, true),
	             5 => (S11_ipd'last_event,tpd_S11_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMF1_VITAL of CMF1 is 
    for VITAL_ACT
    end for;
 end CFG_CMF1_VITAL;



 ---- CELL CMF2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMF2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMF2 :  entity is TRUE;
 end CMF2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMF2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (DB_ipd, S00_ipd, S01_ipd, D1_ipd, S10_ipd, S11_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( VitalMUX2( (NOT DB_ipd) , D1_ipd , NOT (  S00_ipd  AND  S01_ipd )), (NOT DB_ipd) , NOT (  S10_ipd  OR  S11_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (DB_ipd'last_event,tpd_DB_Y, true),
	             1 => (S00_ipd'last_event,tpd_S00_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (D1_ipd'last_event,tpd_D1_Y, true),
	             4 => (S10_ipd'last_event,tpd_S10_Y, true),
	             5 => (S11_ipd'last_event,tpd_S11_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMF2_VITAL of CMF2 is 
    for VITAL_ACT
    end for;
 end CFG_CMF2_VITAL;



 ---- CELL CMF3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMF3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMF3 :  entity is TRUE;
 end CMF3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMF3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL DB_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, S00_ipd, S01_ipd, D1_ipd, S10_ipd, S11_ipd, DB_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( VitalMUX2( D0_ipd , D1_ipd , NOT (  S00_ipd  AND  S01_ipd )), (NOT DB_ipd) , NOT (  S10_ipd  OR  S11_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (S00_ipd'last_event,tpd_S00_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (D1_ipd'last_event,tpd_D1_Y, true),
	             4 => (S10_ipd'last_event,tpd_S10_Y, true),
	             5 => (S11_ipd'last_event,tpd_S11_Y, true),
	             6 => (DB_ipd'last_event,tpd_DB_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMF3_VITAL of CMF3 is 
    for VITAL_ACT
    end for;
 end CFG_CMF3_VITAL;



 ---- CELL CMF4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMF4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMF4 :  entity is TRUE;
 end CMF4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMF4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (DB_ipd, S10_ipd, S11_ipd, D2_ipd, S00_ipd, S01_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( (NOT DB_ipd) , VitalMUX2( D2_ipd , (NOT DB_ipd) , NOT (  S00_ipd  AND  S01_ipd )), NOT (  S10_ipd  OR  S11_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (DB_ipd'last_event,tpd_DB_Y, true),
	             1 => (S10_ipd'last_event,tpd_S10_Y, true),
	             2 => (S11_ipd'last_event,tpd_S11_Y, true),
	             3 => (D2_ipd'last_event,tpd_D2_Y, true),
	             4 => (S00_ipd'last_event,tpd_S00_Y, true),
	             5 => (S01_ipd'last_event,tpd_S01_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMF4_VITAL of CMF4 is 
    for VITAL_ACT
    end for;
 end CFG_CMF4_VITAL;



 ---- CELL CMF5 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMF5 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMF5 :  entity is TRUE;
 end CMF5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMF5 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL DB_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, S10_ipd, S11_ipd, D2_ipd, S00_ipd, S01_ipd, DB_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( VitalMUX2( D0_ipd , D2_ipd , NOT (  S10_ipd  OR  S11_ipd )), (NOT DB_ipd) , NOT (  S00_ipd  AND  S01_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (S10_ipd'last_event,tpd_S10_Y, true),
	             2 => (S11_ipd'last_event,tpd_S11_Y, true),
	             3 => (D2_ipd'last_event,tpd_D2_Y, true),
	             4 => (S00_ipd'last_event,tpd_S00_Y, true),
	             5 => (S01_ipd'last_event,tpd_S01_Y, true),
	             6 => (DB_ipd'last_event,tpd_DB_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMF5_VITAL of CMF5 is 
    for VITAL_ACT
    end for;
 end CFG_CMF5_VITAL;



 ---- CELL CMF6 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMF6 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMF6 :  entity is TRUE;
 end CMF6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMF6 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (DB_ipd, S00_ipd, S01_ipd, D1_ipd, S10_ipd, S11_ipd, D2_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( VitalMUX2( (NOT DB_ipd) , D1_ipd , NOT (  S00_ipd  AND  S01_ipd )), VitalMUX2( D2_ipd , (NOT DB_ipd) , NOT (  S00_ipd  AND  S01_ipd )), NOT (  S10_ipd  OR  S11_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (DB_ipd'last_event,tpd_DB_Y, true),
	             1 => (S00_ipd'last_event,tpd_S00_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (D1_ipd'last_event,tpd_D1_Y, true),
	             4 => (S10_ipd'last_event,tpd_S10_Y, true),
	             5 => (S11_ipd'last_event,tpd_S11_Y, true),
	             6 => (D2_ipd'last_event,tpd_D2_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMF6_VITAL of CMF6 is 
    for VITAL_ACT
    end for;
 end CFG_CMF6_VITAL;



 ---- CELL CMF7 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMF7 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMF7 :  entity is TRUE;
 end CMF7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMF7 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL DB_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, S00_ipd, S01_ipd, D1_ipd, S10_ipd, S11_ipd, D2_ipd, DB_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( VitalMUX2( D0_ipd , D1_ipd , NOT (  S00_ipd  AND  S01_ipd )), VitalMUX2( D2_ipd , (NOT DB_ipd) , NOT (  S00_ipd  AND  S01_ipd )), NOT (  S10_ipd  OR  S11_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (S00_ipd'last_event,tpd_S00_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (D1_ipd'last_event,tpd_D1_Y, true),
	             4 => (S10_ipd'last_event,tpd_S10_Y, true),
	             5 => (S11_ipd'last_event,tpd_S11_Y, true),
	             6 => (D2_ipd'last_event,tpd_D2_Y, true),
	             7 => (DB_ipd'last_event,tpd_DB_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMF7_VITAL of CMF7 is 
    for VITAL_ACT
    end for;
 end CFG_CMF7_VITAL;



 ---- CELL CMF8 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMF8 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMF8 :  entity is TRUE;
 end CMF8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMF8 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (DB_ipd, S10_ipd, S11_ipd, S00_ipd, S01_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( (NOT DB_ipd) , VitalMUX2( (NOT DB_ipd) , D3_ipd , NOT (  S00_ipd  AND  S01_ipd )), NOT (  S10_ipd  OR  S11_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (DB_ipd'last_event,tpd_DB_Y, true),
	             1 => (S10_ipd'last_event,tpd_S10_Y, true),
	             2 => (S11_ipd'last_event,tpd_S11_Y, true),
	             3 => (S00_ipd'last_event,tpd_S00_Y, true),
	             4 => (S01_ipd'last_event,tpd_S01_Y, true),
	             5 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMF8_VITAL of CMF8 is 
    for VITAL_ACT
    end for;
 end CFG_CMF8_VITAL;



 ---- CELL CMF9 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMF9 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMF9 :  entity is TRUE;
 end CMF9;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMF9 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, S00_ipd, S01_ipd, DB_ipd, S10_ipd, S11_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( VitalMUX2( D0_ipd , (NOT DB_ipd) , NOT (  S00_ipd  AND  S01_ipd )), VitalMUX2( (NOT DB_ipd) , D3_ipd , NOT (  S00_ipd  AND  S01_ipd )), NOT (  S10_ipd  OR  S11_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (S00_ipd'last_event,tpd_S00_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (DB_ipd'last_event,tpd_DB_Y, true),
	             4 => (S10_ipd'last_event,tpd_S10_Y, true),
	             5 => (S11_ipd'last_event,tpd_S11_Y, true),
	             6 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMF9_VITAL of CMF9 is 
    for VITAL_ACT
    end for;
 end CFG_CMF9_VITAL;



 ---- CELL CMFA ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMFA is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMFA :  entity is TRUE;
 end CMFA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMFA is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (DB_ipd, S00_ipd, S01_ipd, D1_ipd, S10_ipd, S11_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( (NOT DB_ipd) , VitalMUX2( D1_ipd , D3_ipd , NOT (  S10_ipd  OR  S11_ipd )), NOT (  S00_ipd  AND  S01_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (DB_ipd'last_event,tpd_DB_Y, true),
	             1 => (S00_ipd'last_event,tpd_S00_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (D1_ipd'last_event,tpd_D1_Y, true),
	             4 => (S10_ipd'last_event,tpd_S10_Y, true),
	             5 => (S11_ipd'last_event,tpd_S11_Y, true),
	             6 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMFA_VITAL of CMFA is 
    for VITAL_ACT
    end for;
 end CFG_CMFA_VITAL;



 ---- CELL CMFB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMFB is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMFB :  entity is TRUE;
 end CMFB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMFB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, S00_ipd, S01_ipd, D1_ipd, S10_ipd, S11_ipd, DB_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( VitalMUX2( D0_ipd , D1_ipd , NOT (  S00_ipd  AND  S01_ipd )), VitalMUX2( (NOT DB_ipd) , D3_ipd , NOT (  S00_ipd  AND  S01_ipd )), NOT (  S10_ipd  OR  S11_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (S00_ipd'last_event,tpd_S00_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (D1_ipd'last_event,tpd_D1_Y, true),
	             4 => (S10_ipd'last_event,tpd_S10_Y, true),
	             5 => (S11_ipd'last_event,tpd_S11_Y, true),
	             6 => (DB_ipd'last_event,tpd_DB_Y, true),
	             7 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMFB_VITAL of CMFB is 
    for VITAL_ACT
    end for;
 end CFG_CMFB_VITAL;



 ---- CELL CMFC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMFC is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMFC :  entity is TRUE;
 end CMFC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMFC is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (DB_ipd, S10_ipd, S11_ipd, D2_ipd, S00_ipd, S01_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( (NOT DB_ipd) , VitalMUX2( D2_ipd , D3_ipd , NOT (  S00_ipd  AND  S01_ipd )), NOT (  S10_ipd  OR  S11_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (DB_ipd'last_event,tpd_DB_Y, true),
	             1 => (S10_ipd'last_event,tpd_S10_Y, true),
	             2 => (S11_ipd'last_event,tpd_S11_Y, true),
	             3 => (D2_ipd'last_event,tpd_D2_Y, true),
	             4 => (S00_ipd'last_event,tpd_S00_Y, true),
	             5 => (S01_ipd'last_event,tpd_S01_Y, true),
	             6 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMFC_VITAL of CMFC is 
    for VITAL_ACT
    end for;
 end CFG_CMFC_VITAL;



 ---- CELL CMFD ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMFD is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		DB		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMFD :  entity is TRUE;
 end CMFD;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMFD is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, S00_ipd, S01_ipd, DB_ipd, S10_ipd, S11_ipd, D2_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( VitalMUX2( D0_ipd , (NOT DB_ipd) , NOT (  S00_ipd  AND  S01_ipd )), VitalMUX2( D2_ipd , D3_ipd , NOT (  S00_ipd  AND  S01_ipd )), NOT (  S10_ipd  OR  S11_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (S00_ipd'last_event,tpd_S00_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (DB_ipd'last_event,tpd_DB_Y, true),
	             4 => (S10_ipd'last_event,tpd_S10_Y, true),
	             5 => (S11_ipd'last_event,tpd_S11_Y, true),
	             6 => (D2_ipd'last_event,tpd_D2_Y, true),
	             7 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMFD_VITAL of CMFD is 
    for VITAL_ACT
    end for;
 end CFG_CMFD_VITAL;



 ---- CELL CMFE ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CMFE is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_DB_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S00_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S01_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S00		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S01		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		S00		: in    STD_ULOGIC;
		S01		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S10		: in    STD_ULOGIC;
		S11		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CMFE :  entity is TRUE;
 end CMFE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CMFE is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL DB_ipd  : STD_ULOGIC := 'X';
	SIGNAL S00_ipd  : STD_ULOGIC := 'X';
	SIGNAL S01_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	VitalWireDelay (S00_ipd, S00, tipd_S00);
	VitalWireDelay (S01_ipd, S01, tipd_S01);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (DB_ipd, S00_ipd, S01_ipd, D1_ipd, S10_ipd, S11_ipd, D2_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( VitalMUX2( (NOT DB_ipd) , D1_ipd , NOT (  S00_ipd  AND  S01_ipd )), VitalMUX2( D2_ipd , D3_ipd , NOT (  S00_ipd  AND  S01_ipd )), NOT (  S10_ipd  OR  S11_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (DB_ipd'last_event,tpd_DB_Y, true),
	             1 => (S00_ipd'last_event,tpd_S00_Y, true),
	             2 => (S01_ipd'last_event,tpd_S01_Y, true),
	             3 => (D1_ipd'last_event,tpd_D1_Y, true),
	             4 => (S10_ipd'last_event,tpd_S10_Y, true),
	             5 => (S11_ipd'last_event,tpd_S11_Y, true),
	             6 => (D2_ipd'last_event,tpd_D2_Y, true),
	             7 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CMFE_VITAL of CMFE is 
    for VITAL_ACT
    end for;
 end CFG_CMFE_VITAL;



 ---- CELL CS1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CS1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CS1 :  entity is TRUE;
 end CS1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CS1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( C_ipd , D_ipd , NOT (  A_ipd  OR ( S_ipd  AND  B_ipd )));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (S_ipd'last_event,tpd_S_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true),
	             3 => (C_ipd'last_event,tpd_C_Y, true),
	             4 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CS1_VITAL of CS1 is 
    for VITAL_ACT
    end for;
 end CFG_CS1_VITAL;



 ---- CELL CS2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CS2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CS2 :  entity is TRUE;
 end CS2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CS2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( C_ipd , D_ipd , NOT ( ( A_ipd  OR  S_ipd ) AND  B_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (S_ipd'last_event,tpd_S_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true),
	             3 => (C_ipd'last_event,tpd_C_Y, true),
	             4 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CS2_VITAL of CS2 is 
    for VITAL_ACT
    end for;
 end CFG_CS2_VITAL;



 ---- CELL CY2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CY2A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B0		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A1		: in    STD_ULOGIC;
		B1		: in    STD_ULOGIC;
		A0		: in    STD_ULOGIC;
		B0		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CY2A :  entity is TRUE;
 end CY2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CY2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A1_ipd  : STD_ULOGIC := 'X';
	SIGNAL B1_ipd  : STD_ULOGIC := 'X';
	SIGNAL A0_ipd  : STD_ULOGIC := 'X';
	SIGNAL B0_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A1_ipd, A1, tipd_A1);
	VitalWireDelay (B1_ipd, B1, tipd_B1);
	VitalWireDelay (A0_ipd, A0, tipd_A0);
	VitalWireDelay (B0_ipd, B0, tipd_B0);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A1_ipd, B1_ipd, A0_ipd, B0_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A1_ipd  AND  B1_ipd ) OR (( A0_ipd  AND  B0_ipd ) AND  A1_ipd )) OR (( A0_ipd  AND  B0_ipd ) AND  B1_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A1_ipd'last_event,tpd_A1_Y, true),
	             1 => (B1_ipd'last_event,tpd_B1_Y, true),
	             2 => (A0_ipd'last_event,tpd_A0_Y, true),
	             3 => (B0_ipd'last_event,tpd_B0_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CY2A_VITAL of CY2A is 
    for VITAL_ACT
    end for;
 end CFG_CY2A_VITAL;



 ---- CELL CY2B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CY2B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B0		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A1		: in    STD_ULOGIC;
		B1		: in    STD_ULOGIC;
		A0		: in    STD_ULOGIC;
		B0		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CY2B :  entity is TRUE;
 end CY2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CY2B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A1_ipd  : STD_ULOGIC := 'X';
	SIGNAL B1_ipd  : STD_ULOGIC := 'X';
	SIGNAL A0_ipd  : STD_ULOGIC := 'X';
	SIGNAL B0_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A1_ipd, A1, tipd_A1);
	VitalWireDelay (B1_ipd, B1, tipd_B1);
	VitalWireDelay (A0_ipd, A0, tipd_A0);
	VitalWireDelay (B0_ipd, B0, tipd_B0);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A1_ipd, B1_ipd, A0_ipd, B0_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A1_ipd  AND  B1_ipd ) OR (( A0_ipd  OR  B0_ipd ) AND  A1_ipd )) OR (( A0_ipd  OR  B0_ipd ) AND  B1_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A1_ipd'last_event,tpd_A1_Y, true),
	             1 => (B1_ipd'last_event,tpd_B1_Y, true),
	             2 => (A0_ipd'last_event,tpd_A0_Y, true),
	             3 => (B0_ipd'last_event,tpd_B0_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CY2B_VITAL of CY2B is 
    for VITAL_ACT
    end for;
 end CFG_CY2B_VITAL;



 ---- CELL DF1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DF1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DF1 :  entity is TRUE;
 end DF1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DF1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DF1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DF1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed, '0', '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DF1_VITAL of DF1 is
   for VITAL_ACT
   end for;
end CFG_DF1_VITAL;



 ---- CELL DF1_CC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DF1_CC is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DF1_CC :  entity is TRUE;
 end DF1_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DF1_CC is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DF1_CC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DF1_CC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed, '0', '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DF1_CC_VITAL of DF1_CC is
   for VITAL_ACT
   end for;
end CFG_DF1_CC_VITAL;



 ---- CELL DF1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DF1B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DF1B :  entity is TRUE;
 end DF1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DF1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DF1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DF1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, D_delayed, '0', '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DF1B_VITAL of DF1B is
   for VITAL_ACT
   end for;
end CFG_DF1B_VITAL;



 ---- CELL DFC1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFC1B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFC1B :  entity is TRUE;
 end DFC1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFC1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFC1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>    TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFC1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFC1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFC1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, D_delayed, '0', '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFC1B_VITAL of DFC1B is
   for VITAL_ACT
   end for;
end CFG_DFC1B_VITAL;



 ---- CELL DFC1B_CC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFC1B_CC is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFC1B_CC :  entity is TRUE;
 end DFC1B_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFC1B_CC is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFC1B_CC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>    TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFC1B_CC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFC1B_CC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFC1B_CC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, D_delayed, '0', '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFC1B_CC_VITAL of DFC1B_CC is
   for VITAL_ACT
   end for;
end CFG_DFC1B_CC_VITAL;



 ---- CELL DFC1D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFC1D is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFC1D :  entity is TRUE;
 end DFC1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFC1D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFC1D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>    TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFC1D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFC1D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFC1D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, Q_zd, D_delayed, '0', '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFC1D_VITAL of DFC1D is
   for VITAL_ACT
   end for;
end CFG_DFC1D_VITAL;



 ---- CELL DFE1C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFE1C is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFE1C :  entity is TRUE;
 end DFE1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFE1C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFE1C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TRUE,	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFE1C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFE1C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, D_delayed, E_delayed, '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFE1C_VITAL of DFE1C is
   for VITAL_ACT
   end for;
end CFG_DFE1C_VITAL;



 ---- CELL DFE1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFE1B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFE1B :  entity is TRUE;
 end DFE1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFE1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFE1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TRUE,	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFE1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFE1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed, E_delayed, '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFE1B_VITAL of DFE1B is
   for VITAL_ACT
   end for;
end CFG_DFE1B_VITAL;



 ---- CELL DFE3C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFE3C is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFE3C :  entity is TRUE;
 end DFE3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFE3C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFE3C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFE3C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFE3C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFE3C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFE3C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, D_delayed, E_delayed, '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFE3C_VITAL of DFE3C is
   for VITAL_ACT
   end for;
end CFG_DFE3C_VITAL;



 ---- CELL DFE3D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFE3D is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFE3D :  entity is TRUE;
 end DFE3D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFE3D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFE3D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFE3D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFE3D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFE3D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFE3D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, Q_zd, D_delayed, E_delayed, '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFE3D_VITAL of DFE3D is
   for VITAL_ACT
   end for;
end CFG_DFE3D_VITAL;



 ---- CELL DFE4F ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFE4F is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFE4F :  entity is TRUE;
 end DFE4F;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFE4F is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFE4F",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFE4F",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFE4F",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFE4F",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFE4F",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed, E_delayed, PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFE4F_VITAL of DFE4F is
   for VITAL_ACT
   end for;
end CFG_DFE4F_VITAL;



 ---- CELL DFE4G ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFE4G is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFE4G :  entity is TRUE;
 end DFE4G;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFE4G is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFE4G",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFE4G",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFE4G",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFE4G",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFE4G",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or 
	 Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, D_delayed, E_delayed, PRE_ipd, CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFE4G_VITAL of DFE4G is
   for VITAL_ACT
   end for;
end CFG_DFE4G_VITAL;



 ---- CELL DFEG ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFEG is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFEG :  entity is TRUE;
 end DFEG;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFEG is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DFEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, D_delayed, E_delayed, PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFEG_VITAL of DFEG is
   for VITAL_ACT
   end for;
end CFG_DFEG_VITAL;



 ---- CELL DFEH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFEH is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFEH :  entity is TRUE;
 end DFEH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFEH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (CLR_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DFEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or 
	 Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, Q_zd, D_delayed, E_delayed, PRE_ipd, CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFEH_VITAL of DFEH is
   for VITAL_ACT
   end for;
end CFG_DFEH_VITAL;



 ---- CELL DFP1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFP1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFP1 :  entity is TRUE;
 end DFP1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFP1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_posedge,
	 Removal		=> thold_PRE_CLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed, '0', (NOT PRE_ipd), CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFP1_VITAL of DFP1 is
   for VITAL_ACT
   end for;
end CFG_DFP1_VITAL;



 ---- CELL DFP1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFP1A is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFP1A :  entity is TRUE;
 end DFP1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFP1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFP1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_negedge,
	 Removal		=> thold_PRE_CLK_negedge_negedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFP1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFP1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFP1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, D_delayed, '0', (NOT PRE_ipd), CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFP1A_VITAL of DFP1A is
   for VITAL_ACT
   end for;
end CFG_DFP1A_VITAL;



 ---- CELL DFP1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFP1B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFP1B :  entity is TRUE;
 end DFP1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFP1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFP1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFP1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFP1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFP1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed, '0', PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFP1B_VITAL of DFP1B is
   for VITAL_ACT
   end for;
end CFG_DFP1B_VITAL;



 ---- CELL DFP1B_CC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFP1B_CC is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFP1B_CC :  entity is TRUE;
 end DFP1B_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFP1B_CC is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFP1B_CC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFP1B_CC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFP1B_CC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFP1B_CC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed, '0', PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFP1B_CC_VITAL of DFP1B_CC is
   for VITAL_ACT
   end for;
end CFG_DFP1B_CC_VITAL;



 ---- CELL DFP1D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFP1D is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFP1D :  entity is TRUE;
 end DFP1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFP1D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFP1D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFP1D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFP1D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFP1D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or 
	 Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, D_delayed, '0', PRE_ipd, CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFP1D_VITAL of DFP1D is
   for VITAL_ACT
   end for;
end CFG_DFP1D_VITAL;



 ---- CELL DFPC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFPC is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFPC :  entity is TRUE;
 end DFPC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFPC is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (NOT PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFPC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_posedge,
	 Removal		=> thold_PRE_CLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01((CLR_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFPC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01(( NOT PRE_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFPC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFPC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFPC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DFPC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, D_delayed, '0', (NOT PRE_ipd), CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFPC_VITAL of DFPC is
   for VITAL_ACT
   end for;
end CFG_DFPC_VITAL;



 ---- CELL DFPCB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFPCB is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFPCB :  entity is TRUE;
 end DFPCB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFPCB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFPCB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFPCB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFPCB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFPCB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFPCB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DFPCB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, D_delayed, '0', PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFPCB_VITAL of DFPCB is
   for VITAL_ACT
   end for;
end CFG_DFPCB_VITAL;



 ---- CELL DFPCC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFPCC is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFPCC :  entity is TRUE;
 end DFPCC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFPCC is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFPCC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFPCC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFPCC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFPCC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFPCC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DFPCC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or 
	 Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, Q_zd, D_delayed, '0', PRE_ipd, CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFPCC_VITAL of DFPCC is
   for VITAL_ACT
   end for;
end CFG_DFPCC_VITAL;



 ---- CELL DL1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DL1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DL1 :  entity is TRUE;
 end DL1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DL1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DL1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TRUE, 
	 HeaderMsg		=> InstancePath & "DL1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT G_ipd),D_ipd,'0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		    1 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DL1_VITAL of DL1 is
   for VITAL_ACT
   end for;
end CFG_DL1_VITAL;



 ---- CELL DL1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DL1A is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DL1A :  entity is TRUE;
 end DL1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DL1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DL1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TRUE, 
	 HeaderMsg		=> InstancePath & "DL1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT G_ipd),D_ipd,'0'));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		    1 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DL1A_VITAL of DL1A is
   for VITAL_ACT
   end for;
end CFG_DL1A_VITAL;



 ---- CELL DL1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DL1B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DL1B :  entity is TRUE;
 end DL1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DL1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DL1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TRUE, 
	 HeaderMsg		=> InstancePath & "DL1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',G_ipd,D_ipd,'0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		    1 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DL1B_VITAL of DL1B is
   for VITAL_ACT
   end for;
end CFG_DL1B_VITAL;



 ---- CELL DL1C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DL1C is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DL1C :  entity is TRUE;
 end DL1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DL1C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DL1C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TRUE, 
	 HeaderMsg		=> InstancePath & "DL1C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',G_ipd,D_ipd,'0'));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		    1 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DL1C_VITAL of DL1C is
   for VITAL_ACT
   end for;
end CFG_DL1C_VITAL;



 ---- CELL DL2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DL2A is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DL2A :  entity is TRUE;
 end DL2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DL2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_negedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) OR (PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DL2A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_negedge,
	 TimingData		=> Tmkr_CLR_G_negedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_posedge_negedge,
	 Removal                => thold_CLR_G_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TO_X01(( NOT PRE_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DL2A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_negedge,
	 TimingData		=> Tmkr_PRE_G_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_negedge_negedge,
	 Removal		=> thold_PRE_G_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01((CLR_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DL2A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (NOT PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DL2A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DL2A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DL2A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or 
		       Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		CLR_ipd,(NOT G_ipd),D_ipd,PRE_ipd));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		    2 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    3 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DL2A_VITAL of DL2A is
   for VITAL_ACT
   end for;
end CFG_DL2A_VITAL;



 ---- CELL DL2C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DL2C is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DL2C :  entity is TRUE;
 end DL2C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DL2C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_posedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) OR (PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DL2C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_posedge,
	 TimingData		=> Tmkr_CLR_G_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_posedge_posedge,
	 Removal                => thold_CLR_G_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TO_X01(( NOT PRE_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DL2C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_posedge,
	 TimingData		=> Tmkr_PRE_G_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_negedge_posedge,
	 Removal		=> thold_PRE_G_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01((CLR_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DL2C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (NOT PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DL2C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DL2C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DL2C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_PRE or 
		       Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		CLR_ipd,G_ipd,D_ipd,PRE_ipd));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		    2 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    3 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DL2C_VITAL of DL2C is
   for VITAL_ACT
   end for;
end CFG_DL2C_VITAL;



 ---- CELL DLC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLC is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLC :  entity is TRUE;
 end DLC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLC is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_negedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_negedge,
	 TimingData		=> Tmkr_CLR_G_negedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_posedge_negedge,
	 Removal                => thold_CLR_G_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		CLR_ipd,(NOT G_ipd),D_ipd,'0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLC_VITAL of DLC is
   for VITAL_ACT
   end for;
end CFG_DLC_VITAL;



 ---- CELL DLC1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLC1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLC1 :  entity is TRUE;
 end DLC1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLC1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_negedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLC1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_negedge,
	 TimingData		=> Tmkr_CLR_G_negedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_negedge_negedge,
	 Removal		=> thold_CLR_G_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLC1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLC1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLC1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),(NOT G_ipd),D_ipd,'0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLC1_VITAL of DLC1 is
   for VITAL_ACT
   end for;
end CFG_DLC1_VITAL;



 ---- CELL DLC1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLC1A is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLC1A :  entity is TRUE;
 end DLC1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLC1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_posedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLC1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_posedge,
	 TimingData		=> Tmkr_CLR_G_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_negedge_posedge,
	 Removal		=> thold_CLR_G_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLC1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLC1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLC1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),G_ipd,D_ipd,'0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLC1A_VITAL of DLC1A is
   for VITAL_ACT
   end for;
end CFG_DLC1A_VITAL;



 ---- CELL DLC1F ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLC1F is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLC1F :  entity is TRUE;
 end DLC1F;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLC1F is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_negedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLC1F",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_negedge,
	 TimingData		=> Tmkr_CLR_G_negedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_negedge_negedge,
	 Removal		=> thold_CLR_G_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLC1F",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLC1F",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLC1F",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),(NOT G_ipd),D_ipd,'0'));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_QN, true),
		    2 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLC1F_VITAL of DLC1F is
   for VITAL_ACT
   end for;
end CFG_DLC1F_VITAL;



 ---- CELL DLC1G ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLC1G is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLC1G :  entity is TRUE;
 end DLC1G;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLC1G is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_posedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLC1G",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_posedge,
	 TimingData		=> Tmkr_CLR_G_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_negedge_posedge,
	 Removal		=> thold_CLR_G_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLC1G",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLC1G",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLC1G",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),G_ipd,D_ipd,'0'));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_QN, true),
		    2 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLC1G_VITAL of DLC1G is
   for VITAL_ACT
   end for;
end CFG_DLC1G_VITAL;



 ---- CELL DLCA ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLCA is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLCA :  entity is TRUE;
 end DLCA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLCA is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_posedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLCA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_posedge,
	 TimingData		=> Tmkr_CLR_G_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_posedge_posedge,
	 Removal                => thold_CLR_G_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLCA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLCA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLCA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		CLR_ipd,G_ipd,D_ipd,'0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLCA_VITAL of DLCA is
   for VITAL_ACT
   end for;
end CFG_DLCA_VITAL;



 ---- CELL DLE ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLE is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_E_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLE :  entity is TRUE;
 end DLE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLE is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd,E, tipd_E);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, E_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D_E_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_E_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tviol_E_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_E_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tmkr_E_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_E		: STD_ULOGIC := '0';
	VARIABLE PInfo_E		: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLE",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_E_negedge,
	 TimingData		=> Tmkr_D_E_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> E_ipd,
	 RefSignalName		=> "E",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_E_posedge_negedge,
	 SetupLow		=> tsetup_D_E_negedge_negedge,
	 HoldHigh               => thold_D_E_posedge_negedge,
	 HoldLow		=> thold_D_E_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT G_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLE",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_negedge,
	 TimingData             => Tmkr_E_G_negedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,
	 SetupLow               => 0 ns,
	 HoldHigh               => thold_E_G_negedge_negedge,
	 HoldLow                => 0 ns,
	 CheckEnabled           =>  TRUE, 
	 RefTransition          => 'F',
	 HeaderMsg              => InstancePath & "/DLE",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_posedge,
	 TimingData             => Tmkr_E_G_posedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => tsetup_E_G_posedge_posedge,
	 SetupLow              => 0 ns,
	 HoldHigh               => 0 ns,
	 HoldLow                => 0 ns,
	 CheckEnabled           =>  TRUE, 
	 RefTransition          => 'R',
	 HeaderMsg              => InstancePath & "/DLE",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((E_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLE",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_E,
	 PeriodData		=> PInfo_E,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 Period	        	=> 0 ns,
         PulseWidthLow          => 0 ns,
	 PulseWidthHigh		=> tpw_E_posedge,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLE",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Tviol_D_E_negedge or Pviol_E or 
		      Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DLE3B_Q_tab,
	 DataIn => (
		  (NOT G_ipd),(NOT E_ipd),D_ipd,'0'));

	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 =>(E_ipd'last_event, tpd_E_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLE_VITAL of DLE is
   for VITAL_ACT
   end for;
end CFG_DLE_VITAL;



 ---- CELL DLE1D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLE1D is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_E_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLE1D :  entity is TRUE;
 end DLE1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLE1D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd,E, tipd_E);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, E_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D_E_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_E_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tviol_E_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_E_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tmkr_E_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_E		: STD_ULOGIC := '0';
	VARIABLE PInfo_E		: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((E_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLE1D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_E_posedge,
	 TimingData		=> Tmkr_D_E_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> E_ipd,
	 RefSignalName		=> "E",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_E_posedge_posedge,
	 SetupLow		=> tsetup_D_E_negedge_posedge,
	 HoldHigh               => thold_D_E_posedge_posedge,
	 HoldLow		=> thold_D_E_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((G_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLE1D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_posedge,
	 TimingData             => Tmkr_E_G_posedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,
	 SetupLow               => 0 ns,
	 HoldHigh               => 0 ns,
	 HoldLow                => thold_E_G_posedge_posedge,
	 CheckEnabled           =>  TRUE, 
	 RefTransition          => 'R',
	 HeaderMsg              => InstancePath & "/DLE1D",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_negedge,
	 TimingData             => Tmkr_E_G_negedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,
	 SetupLow              => tsetup_E_G_negedge_negedge,
	 HoldHigh               => 0 ns,
	 HoldLow                => 0 ns,
	 CheckEnabled           =>  TRUE, 
	 RefTransition          => 'F',
	 HeaderMsg              => InstancePath & "/DLE1D",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLE1D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_E,
	 PeriodData		=> PInfo_E,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 Period	        	=> 0 ns,
         PulseWidthLow          => tpw_E_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLE1D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Tviol_D_E_posedge or Pviol_E or 
		      Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DLE3B_Q_tab,
	 DataIn => (
		  G_ipd,E_ipd,D_ipd,'0'));

	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		     1 =>(E_ipd'last_event, tpd_E_QN, true),
		    2 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLE1D_VITAL of DLE1D is
   for VITAL_ACT
   end for;
end CFG_DLE1D_VITAL;



 ---- CELL DLE2B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLE2B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_E_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLE2B :  entity is TRUE;
 end DLE2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLE2B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (E_ipd,E, tipd_E);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D_E_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_E_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tviol_E_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_E_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tmkr_E_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_posedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Tviol_CLR_E_posedge : STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_E_posedge         : VitalTimingDataType   := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_E		: STD_ULOGIC := '0';
	VARIABLE PInfo_E		: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) OR (E_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLE2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_E_posedge,
	 TimingData		=> Tmkr_D_E_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> E_ipd,
	 RefSignalName		=> "E",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_E_posedge_posedge,
	 SetupLow		=> tsetup_D_E_negedge_posedge,
	 HoldHigh               => thold_D_E_posedge_posedge,
	 HoldLow		=> thold_D_E_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) OR (G_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLE2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_posedge,
	 TimingData             => Tmkr_E_G_posedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,
	 SetupLow               => 0 ns,
	 HoldHigh               => 0 ns,
	 HoldLow                => thold_E_G_posedge_posedge,
	 CheckEnabled           =>  TO_X01(((NOT CLR_ipd) ) ) /= '1', 
	 RefTransition          => 'R',
	 HeaderMsg              => InstancePath & "/DLE2B",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_negedge,
	 TimingData             => Tmkr_E_G_negedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,
	 SetupLow              => tsetup_E_G_negedge_negedge,
	 HoldHigh               => 0 ns,
	 HoldLow                => 0 ns,
	 CheckEnabled           =>  TO_X01(((NOT CLR_ipd) ) ) /= '1', 
	 RefTransition          => 'F',
	 HeaderMsg              => InstancePath & "/DLE2B",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_posedge,
	 TimingData		=> Tmkr_CLR_G_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_posedge_posedge,
	 Removal                => thold_CLR_G_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLE2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_E_posedge,
	 TimingData		=> Tmkr_CLR_E_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> E_ipd,
	 RefSignalName		=> "E",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_E_posedge_posedge,
	 Removal                => thold_CLR_E_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>  TO_X01((NOT G_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLE2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLE2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_E,
	 PeriodData		=> PInfo_E,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 Period	        	=> 0 ns,
         PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_E_negedge,
	 CheckEnabled		=> TO_X01((NOT CLR_ipd)) /= '1',
	 HeaderMsg		=> InstancePath & "DLE2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLE2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Tviol_D_E_posedge or Pviol_CLR or 
		      Pviol_E or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DLE2B_Q_tab,
	 DataIn => (
		    CLR_ipd,G_ipd,E_ipd,D_ipd));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 =>(E_ipd'last_event, tpd_E_Q, true),
		    2 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    3 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLE2B_VITAL of DLE2B is
   for VITAL_ACT
   end for;
end CFG_DLE2B_VITAL;



 ---- CELL DLE2C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLE2C is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_E_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLE2C :  entity is TRUE;
 end DLE2C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLE2C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (E_ipd,E, tipd_E);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D_E_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_E_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tviol_E_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_E_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tmkr_E_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_posedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Tviol_CLR_E_posedge : STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_E_posedge         : VitalTimingDataType   := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_E		: STD_ULOGIC := '0';
	VARIABLE PInfo_E		: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) OR (E_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLE2C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_E_posedge,
	 TimingData		=> Tmkr_D_E_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> E_ipd,
	 RefSignalName		=> "E",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_E_posedge_posedge,
	 SetupLow		=> tsetup_D_E_negedge_posedge,
	 HoldHigh               => thold_D_E_posedge_posedge,
	 HoldLow		=> thold_D_E_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) OR (G_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLE2C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_posedge,
	 TimingData             => Tmkr_E_G_posedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,
	 SetupLow               => 0 ns,
	 HoldHigh               => 0 ns,
	 HoldLow                => thold_E_G_posedge_posedge,
	 CheckEnabled           =>  TO_X01(((CLR_ipd) ) ) /= '1', 
	 RefTransition          => 'R',
	 HeaderMsg              => InstancePath & "/DLE2C",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_negedge,
	 TimingData             => Tmkr_E_G_negedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,
	 SetupLow              => tsetup_E_G_negedge_negedge,
	 HoldHigh               => 0 ns,
	 HoldLow                => 0 ns,
	 CheckEnabled           =>  TO_X01(((CLR_ipd) ) ) /= '1', 
	 RefTransition          => 'F',
	 HeaderMsg              => InstancePath & "/DLE2C",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_posedge,
	 TimingData		=> Tmkr_CLR_G_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_negedge_posedge,
	 Removal		=> thold_CLR_G_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLE2C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_E_posedge,
	 TimingData		=> Tmkr_CLR_E_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> E_ipd,
	 RefSignalName		=> "E",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_E_negedge_posedge,
	 Removal		=> thold_CLR_E_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>  TO_X01((NOT G_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLE2C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLE2C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_E,
	 PeriodData		=> PInfo_E,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 Period	        	=> 0 ns,
         PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_E_negedge,
	 CheckEnabled		=> TO_X01((CLR_ipd)) /= '1',
	 HeaderMsg		=> InstancePath & "DLE2C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLE2C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Tviol_D_E_posedge or Pviol_CLR or 
		      Pviol_E or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DLE2B_Q_tab,
	 DataIn => (
		    (NOT CLR_ipd),G_ipd,E_ipd,D_ipd));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 =>(E_ipd'last_event, tpd_E_Q, true),
		    2 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    3 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLE2C_VITAL of DLE2C is
   for VITAL_ACT
   end for;
end CFG_DLE2C_VITAL;



 ---- CELL DLE3B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLE3B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_E_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLE3B :  entity is TRUE;
 end DLE3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLE3B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (E_ipd,E, tipd_E);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D_E_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_E_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tviol_E_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_E_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tmkr_E_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_E_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_E_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_E		: STD_ULOGIC := '0';
	VARIABLE PInfo_E		: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) OR (E_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLE3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_E_posedge,
	 TimingData		=> Tmkr_D_E_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> E_ipd,
	 RefSignalName		=> "E",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_E_posedge_posedge,
	 SetupLow		=> tsetup_D_E_negedge_posedge,
	 HoldHigh               => thold_D_E_posedge_posedge,
	 HoldLow		=> thold_D_E_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) OR (G_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLE3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_posedge,
	 TimingData             => Tmkr_E_G_posedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,
	 SetupLow               => thold_E_G_posedge_posedge,
	 HoldHigh               => 0 ns,
	 HoldLow                => 0 ns,
	 CheckEnabled           =>  TO_X01(((PRE_ipd) ) ) /= '1', 
	 RefTransition          => 'R',
	 HeaderMsg              => InstancePath & "/DLE3B",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_negedge,
	 TimingData             => Tmkr_E_G_negedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,
	 SetupLow              => tsetup_E_G_negedge_negedge,
	 HoldHigh               => 0 ns,
	 HoldLow                => 0 ns,
	 CheckEnabled           =>  TO_X01(((PRE_ipd) ) ) /= '1', 
	 RefTransition          => 'F',
	 HeaderMsg              => InstancePath & "/DLE3B",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_posedge,
	 TimingData		=> Tmkr_PRE_G_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_negedge_posedge,
	 Removal		=> thold_PRE_G_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLE3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_E_posedge,
	 TimingData		=> Tmkr_PRE_E_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> E_ipd,
	 RefSignalName		=> "E",
	 RefDelay	 => 0 ns,
	 Recovery	 => trecovery_PRE_E_negedge_posedge,
	 Removal		=> thold_PRE_E_negedge_posedge,
	 ActiveLow		=> FALSE,
   CheckEnabled		=>  TO_X01((NOT G_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLE3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLE3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_E,
	 PeriodData		=> PInfo_E,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 Period	        	=> 0 ns,
         PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_E_negedge,
	 CheckEnabled		=> TO_X01( (PRE_ipd)) /= '1',
	 HeaderMsg		=> InstancePath & "DLE3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 	TRUE,
	 HeaderMsg		=> InstancePath & "DLE3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Tviol_D_E_posedge or Tviol_PRE_G_posedge or 
		      Pviol_PRE or Pviol_E or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DLE3B_Q_tab,
	 DataIn => (
		  G_ipd,E_ipd,D_ipd,PRE_ipd));

	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 =>(E_ipd'last_event, tpd_E_Q, true),
		     2 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		    3 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLE3B_VITAL of DLE3B is
   for VITAL_ACT
   end for;
end CFG_DLE3B_VITAL;



 ---- CELL DLE3C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLE3C is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_E_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLE3C :  entity is TRUE;
 end DLE3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLE3C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (E_ipd,E, tipd_E);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D_E_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_E_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tviol_E_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_E_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tmkr_E_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_E_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_E_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_E		: STD_ULOGIC := '0';
	VARIABLE PInfo_E		: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) OR (E_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLE3C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_E_posedge,
	 TimingData		=> Tmkr_D_E_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> E_ipd,
	 RefSignalName		=> "E",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_E_posedge_posedge,
	 SetupLow		=> tsetup_D_E_negedge_posedge,
	 HoldHigh               => thold_D_E_posedge_posedge,
	 HoldLow		=> thold_D_E_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) OR (G_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLE3C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_posedge,
	 TimingData             => Tmkr_E_G_posedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,	 
         SetupLow               => 0 ns,
	 HoldHigh               => 0 ns,
	 HoldLow                => thold_E_G_posedge_posedge,
	 CheckEnabled           =>  TO_X01(((NOT PRE_ipd) ) ) /= '1', 
	 RefTransition          => 'R',
	 HeaderMsg              => InstancePath & "/DLE3C",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_negedge,
	 TimingData             => Tmkr_E_G_negedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,
	 SetupLow              => tsetup_E_G_negedge_negedge,
	 HoldHigh               => 0 ns,
	 HoldLow                => 0 ns,
	 CheckEnabled           =>  TO_X01(((NOT PRE_ipd) ) ) /= '1', 
	 RefTransition          => 'F',
	 HeaderMsg              => InstancePath & "/DLE3C",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_posedge,
	 TimingData		=> Tmkr_PRE_G_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_posedge_posedge,
	 Removal                => thold_PRE_G_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLE3C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_E_posedge,
	 TimingData		=> Tmkr_PRE_E_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> E_ipd,
	 RefSignalName		=> "E",
	 RefDelay	 => 0 ns,
	 Recovery	 => trecovery_PRE_E_posedge_posedge,
	 Removal                => thold_PRE_E_posedge_posedge,
	 ActiveLow		=> TRUE,
         CheckEnabled		=>  TO_X01((NOT G_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLE3C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLE3C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_E,
	 PeriodData		=> PInfo_E,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 Period	        	=> 0 ns,
         PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_E_negedge,
	 CheckEnabled		=> TO_X01( (NOT PRE_ipd)) /= '1',
	 HeaderMsg		=> InstancePath & "DLE3C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 	TRUE,
	 HeaderMsg		=> InstancePath & "DLE3C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Tviol_D_E_posedge or Tviol_PRE_G_posedge or 
		      Pviol_PRE or Pviol_E or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DLE3B_Q_tab,
	 DataIn => (
		  G_ipd,E_ipd,D_ipd,(NOT PRE_ipd)));

	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 =>(E_ipd'last_event, tpd_E_Q, true),
		     2 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		    3 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLE3C_VITAL of DLE3C is
   for VITAL_ACT
   end for;
end CFG_DLE3C_VITAL;



 ---- CELL DLEA ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLEA is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_E_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLEA :  entity is TRUE;
 end DLEA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLEA is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd,E, tipd_E);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, E_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D_E_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_E_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tviol_E_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_E_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tmkr_E_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_E		: STD_ULOGIC := '0';
	VARIABLE PInfo_E		: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((E_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLEA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_E_posedge,
	 TimingData		=> Tmkr_D_E_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> E_ipd,
	 RefSignalName		=> "E",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_E_posedge_posedge,
	 SetupLow		=> tsetup_D_E_negedge_posedge,
	 HoldHigh               => thold_D_E_posedge_posedge,
	 HoldLow		=> thold_D_E_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT G_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLEA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_negedge,
	 TimingData             => Tmkr_E_G_negedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,	 SetupLow               => 0 ns,
	 HoldHigh               => 0 ns,
	 HoldLow                => thold_E_G_posedge_negedge,
	 CheckEnabled           =>  TRUE, 
	 RefTransition          => 'F',
	 HeaderMsg              => InstancePath & "/DLEA",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_posedge,
	 TimingData             => Tmkr_E_G_posedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,
	 SetupLow              => tsetup_E_G_negedge_posedge,
	 HoldHigh               => 0 ns,
	 HoldLow                => 0 ns,
	 CheckEnabled           =>  TRUE, 
	 RefTransition          => 'R',
	 HeaderMsg              => InstancePath & "/DLEA",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLEA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_E,
	 PeriodData		=> PInfo_E,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 Period	        	=> 0 ns,
         PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_E_negedge,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLEA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Tviol_D_E_posedge or Pviol_E or 
		      Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DLE3B_Q_tab,
	 DataIn => (
		  (NOT G_ipd),E_ipd,D_ipd,'0'));

	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 =>(E_ipd'last_event, tpd_E_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLEA_VITAL of DLEA is
   for VITAL_ACT
   end for;
end CFG_DLEA_VITAL;



 ---- CELL DLEB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLEB is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_E_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLEB :  entity is TRUE;
 end DLEB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLEB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd,E, tipd_E);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, E_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D_E_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_E_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tviol_E_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_E_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tmkr_E_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_E		: STD_ULOGIC := '0';
	VARIABLE PInfo_E		: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLEB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_E_negedge,
	 TimingData		=> Tmkr_D_E_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> E_ipd,
	 RefSignalName		=> "E",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_E_posedge_negedge,
	 SetupLow		=> tsetup_D_E_negedge_negedge,
	 HoldHigh               => thold_D_E_posedge_negedge,
	 HoldLow		=> thold_D_E_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((G_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLEB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_posedge,
	 TimingData             => Tmkr_E_G_posedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,	 SetupLow               => 0 ns,
	 HoldHigh               => thold_E_G_negedge_posedge,
	 HoldLow                =>  0 ns,
	 CheckEnabled           =>  TRUE, 
	 RefTransition          => 'R',
	 HeaderMsg              => InstancePath & "/DLEB",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_negedge,
	 TimingData             => Tmkr_E_G_negedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => tsetup_E_G_posedge_negedge,
	 SetupLow              => 0 ns,
	 HoldHigh               => 0 ns,
	 HoldLow                => 0 ns,
	 CheckEnabled           =>  TRUE, 
	 RefTransition          => 'F',
	 HeaderMsg              => InstancePath & "/DLEB",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((E_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLEB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_E,
	 PeriodData		=> PInfo_E,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 Period	        	=> 0 ns,
         PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_E_posedge,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLEB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Tviol_D_E_negedge or Pviol_E or 
		      Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DLE3B_Q_tab,
	 DataIn => (
		  G_ipd,(NOT E_ipd),D_ipd,'0'));

	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 =>(E_ipd'last_event, tpd_E_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLEB_VITAL of DLEB is
   for VITAL_ACT
   end for;
end CFG_DLEB_VITAL;



 ---- CELL DLEC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLEC is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_E_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLEC :  entity is TRUE;
 end DLEC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLEC is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd,E, tipd_E);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, E_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D_E_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_E_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tviol_E_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_E_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tmkr_E_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_E		: STD_ULOGIC := '0';
	VARIABLE PInfo_E		: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((E_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLEC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_E_posedge,
	 TimingData		=> Tmkr_D_E_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> E_ipd,
	 RefSignalName		=> "E",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_E_posedge_posedge,
	 SetupLow		=> tsetup_D_E_negedge_posedge,
	 HoldHigh               => thold_D_E_posedge_posedge,
	 HoldLow		=> thold_D_E_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((G_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLEC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_posedge,
	 TimingData             => Tmkr_E_G_posedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,	 SetupLow               => 0 ns,
	 HoldHigh               => 0 ns,
	 HoldLow                => thold_E_G_posedge_posedge,
	 CheckEnabled           => TRUE, 
	 RefTransition          => 'R',
	 HeaderMsg              => InstancePath & "/DLEC",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_negedge,
	 TimingData             => Tmkr_E_G_negedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,
	 SetupLow              => tsetup_E_G_negedge_negedge,
	 HoldHigh               => 0 ns,
	 HoldLow                => 0 ns,
	 CheckEnabled           =>  TRUE, 
	 RefTransition          => 'F',
	 HeaderMsg              => InstancePath & "/DLEC",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLEC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_E,
	 PeriodData		=> PInfo_E,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 Period	        	=> 0 ns,
         PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_E_negedge,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLEC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Tviol_D_E_posedge or Pviol_E or 
		      Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DLE3B_Q_tab,
	 DataIn => (
		  G_ipd,E_ipd,D_ipd,'0'));

	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 =>(E_ipd'last_event, tpd_E_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLEC_VITAL of DLEC is
   for VITAL_ACT
   end for;
end CFG_DLEC_VITAL;



 ---- CELL DLM ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLM is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_A_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		A		:  in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLM :  entity is TRUE;
 end DLM;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLM is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd, G_ipd)

	-- timing check results
	VARIABLE Tviol_A_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_A_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_S_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_S_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_B_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_G_negedge,
	 TimingData		=> Tmkr_A_G_negedge,
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_G_posedge_negedge,
	 SetupLow		=> tsetup_A_G_negedge_negedge,
	 HoldHigh		=> thold_A_G_posedge_negedge,
	 HoldLow		=> thold_A_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_G_negedge,
	 TimingData		=> Tmkr_S_G_negedge,
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_G_posedge_negedge,
	 SetupLow		=> tsetup_S_G_negedge_negedge,
	 HoldHigh		=> thold_S_G_posedge_negedge,
	 HoldLow		=> thold_S_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_G_negedge,
	 TimingData		=> Tmkr_B_G_negedge,
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_G_posedge_negedge,
	 SetupLow		=> tsetup_B_G_negedge_negedge,
	 HoldHigh		=> thold_B_G_posedge_negedge,
	 HoldLow		=> thold_B_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TRUE, 
	 HeaderMsg		=> InstancePath & "DLM",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_A_G_negedge or Tviol_S_G_negedge or Tviol_B_G_negedge or 
		      Pviol_G;
	 --- now combinatorial logic input to the DFF 
	 NET_0_2 := 
 VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT G_ipd),NET_0_2, '0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (A_ipd'last_event, tpd_A_Q, true),
		    1 => (S_ipd'last_event, tpd_S_Q, true),
		    2 => (B_ipd'last_event, tpd_B_Q, true),
		    3 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLM_VITAL of DLM is
   for VITAL_ACT
   end for;
end CFG_DLM_VITAL;



 ---- CELL DLM2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLM2 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_A_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		A		:  in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLM2 :  entity is TRUE;
 end DLM2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLM2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd, CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_A_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_A_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_S_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_S_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_B_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_negedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_G_negedge,
	 TimingData		=> Tmkr_A_G_negedge,
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_G_posedge_negedge,
	 SetupLow		=> tsetup_A_G_negedge_negedge,
	 HoldHigh		=> thold_A_G_posedge_negedge,
	 HoldLow		=> thold_A_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM2",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_G_negedge,
	 TimingData		=> Tmkr_S_G_negedge,
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_G_posedge_negedge,
	 SetupLow		=> tsetup_S_G_negedge_negedge,
	 HoldHigh		=> thold_S_G_posedge_negedge,
	 HoldLow		=> thold_S_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM2",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_G_negedge,
	 TimingData		=> Tmkr_B_G_negedge,
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_G_posedge_negedge,
	 SetupLow		=> tsetup_B_G_negedge_negedge,
	 HoldHigh		=> thold_B_G_posedge_negedge,
	 HoldLow		=> thold_B_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM2",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_negedge,
	 TimingData		=> Tmkr_CLR_G_negedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_posedge_negedge,
	 Removal                => thold_CLR_G_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLM2",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLM2",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLM2",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_A_G_negedge or Tviol_S_G_negedge or Tviol_B_G_negedge or 
		      Pviol_CLR or Pviol_G;
	 --- now combinatorial logic input to the DFF 
	 NET_0_2 := 
 VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		CLR_ipd,(NOT G_ipd),NET_0_2, '0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (A_ipd'last_event, tpd_A_Q, true),
		    1 => (S_ipd'last_event, tpd_S_Q, true),
		    2 => (B_ipd'last_event, tpd_B_Q, true),
		    3 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    4 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLM2_VITAL of DLM2 is
   for VITAL_ACT
   end for;
end CFG_DLM2_VITAL;



 ---- CELL DLM2B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLM2B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_A_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		A		:  in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLM2B :  entity is TRUE;
 end DLM2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLM2B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd, CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_A_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_A_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_S_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_S_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_B_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_posedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_G_posedge,
	 TimingData		=> Tmkr_A_G_posedge,
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_G_posedge_posedge,
	 SetupLow		=> tsetup_A_G_negedge_posedge,
	 HoldHigh		=> thold_A_G_posedge_posedge,
	 HoldLow		=> thold_A_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLM2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_G_posedge,
	 TimingData		=> Tmkr_S_G_posedge,
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_G_posedge_posedge,
	 SetupLow		=> tsetup_S_G_negedge_posedge,
	 HoldHigh		=> thold_S_G_posedge_posedge,
	 HoldLow		=> thold_S_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLM2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_G_posedge,
	 TimingData		=> Tmkr_B_G_posedge,
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_G_posedge_posedge,
	 SetupLow		=> tsetup_B_G_negedge_posedge,
	 HoldHigh		=> thold_B_G_posedge_posedge,
	 HoldLow		=> thold_B_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLM2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_posedge,
	 TimingData		=> Tmkr_CLR_G_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_posedge_posedge,
	 Removal                => thold_CLR_G_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLM2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLM2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLM2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_A_G_posedge or Tviol_S_G_posedge or Tviol_B_G_posedge or 
		      Pviol_CLR or Pviol_G;
	 --- now combinatorial logic input to the DFF 
	 NET_0_2 := 
 VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		CLR_ipd,G_ipd,NET_0_2, '0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (A_ipd'last_event, tpd_A_Q, true),
		    1 => (S_ipd'last_event, tpd_S_Q, true),
		    2 => (B_ipd'last_event, tpd_B_Q, true),
		    3 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    4 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLM2B_VITAL of DLM2B is
   for VITAL_ACT
   end for;
end CFG_DLM2B_VITAL;



 ---- CELL DLM3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLM3 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D0_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S0_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S1_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D0_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D0_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D0_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D0_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S0_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S0_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S0_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S0_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D1_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D1_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D1_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D1_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S1_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S1_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S1_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S1_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D2_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D2_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D2_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D2_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D3_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D3_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D3_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D3_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D0		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S0		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S1		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D0		:  in    STD_ULOGIC;
		S0		:  in    STD_ULOGIC;
		D1		:  in    STD_ULOGIC;
		S1		:  in    STD_ULOGIC;
		D2		:  in    STD_ULOGIC;
		D3		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLM3 :  entity is TRUE;
 end DLM3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLM3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL S0_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL S1_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (S0_ipd, S0, tipd_S0);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (S1_ipd, S1, tipd_S1);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D0_ipd, S0_ipd, D1_ipd, S1_ipd, D2_ipd, D3_ipd, G_ipd)

	-- timing check results
	VARIABLE Tviol_D0_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D0_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_S0_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_S0_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D1_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D1_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_S1_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_S1_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D2_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D2_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D3_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D3_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE NET_0_8	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D0_G_negedge,
	 TimingData		=> Tmkr_D0_G_negedge,
	 TestSignal		=> D0_ipd,
	 TestSignalName		=> "D0",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D0_G_posedge_negedge,
	 SetupLow		=> tsetup_D0_G_negedge_negedge,
	 HoldHigh		=> thold_D0_G_posedge_negedge,
	 HoldLow		=> thold_D0_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM3",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_S0_G_negedge,
	 TimingData		=> Tmkr_S0_G_negedge,
	 TestSignal		=> S0_ipd,
	 TestSignalName		=> "S0",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S0_G_posedge_negedge,
	 SetupLow		=> tsetup_S0_G_negedge_negedge,
	 HoldHigh		=> thold_S0_G_posedge_negedge,
	 HoldLow		=> thold_S0_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM3",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D1_G_negedge,
	 TimingData		=> Tmkr_D1_G_negedge,
	 TestSignal		=> D1_ipd,
	 TestSignalName		=> "D1",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D1_G_posedge_negedge,
	 SetupLow		=> tsetup_D1_G_negedge_negedge,
	 HoldHigh		=> thold_D1_G_posedge_negedge,
	 HoldLow		=> thold_D1_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM3",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_S1_G_negedge,
	 TimingData		=> Tmkr_S1_G_negedge,
	 TestSignal		=> S1_ipd,
	 TestSignalName		=> "S1",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S1_G_posedge_negedge,
	 SetupLow		=> tsetup_S1_G_negedge_negedge,
	 HoldHigh		=> thold_S1_G_posedge_negedge,
	 HoldLow		=> thold_S1_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM3",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D2_G_negedge,
	 TimingData		=> Tmkr_D2_G_negedge,
	 TestSignal		=> D2_ipd,
	 TestSignalName		=> "D2",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D2_G_posedge_negedge,
	 SetupLow		=> tsetup_D2_G_negedge_negedge,
	 HoldHigh		=> thold_D2_G_posedge_negedge,
	 HoldLow		=> thold_D2_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM3",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D3_G_negedge,
	 TimingData		=> Tmkr_D3_G_negedge,
	 TestSignal		=> D3_ipd,
	 TestSignalName		=> "D3",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D3_G_posedge_negedge,
	 SetupLow		=> tsetup_D3_G_negedge_negedge,
	 HoldHigh		=> thold_D3_G_posedge_negedge,
	 HoldLow		=> thold_D3_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM3",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TRUE, 
	 HeaderMsg		=> InstancePath & "DLM3",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D0_G_negedge or Tviol_S0_G_negedge or Tviol_D1_G_negedge or 
		      Tviol_S1_G_negedge or Tviol_D2_G_negedge or Tviol_D3_G_negedge or 
		      Pviol_G;
	 --- now combinatorial logic input to the DFF 
	 NET_0_8 := 
 VitalMUX2( VitalMUX2( D0_ipd , D1_ipd , (NOT S0_ipd) ), VitalMUX2( D2_ipd , D3_ipd , (NOT S0_ipd) ), (NOT S1_ipd) );

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT G_ipd),NET_0_8, '0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D0_ipd'last_event, tpd_D0_Q, true),
		    1 => (S0_ipd'last_event, tpd_S0_Q, true),
		    2 => (D1_ipd'last_event, tpd_D1_Q, true),
		    3 => (S1_ipd'last_event, tpd_S1_Q, true),
		    4 => (D2_ipd'last_event, tpd_D2_Q, true),
		    5 => (D3_ipd'last_event, tpd_D3_Q, true),
		    6 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLM3_VITAL of DLM3 is
   for VITAL_ACT
   end for;
end CFG_DLM3_VITAL;



 ---- CELL DLM3A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLM3A is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D0_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S0_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S1_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D0_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D0_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D0_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D0_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S0_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S0_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S0_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S0_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D1_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D1_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D1_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D1_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S1_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S1_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S1_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S1_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D2_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D2_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D2_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D2_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D3_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D3_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D3_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D3_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D0		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S0		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S1		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D0		:  in    STD_ULOGIC;
		S0		:  in    STD_ULOGIC;
		D1		:  in    STD_ULOGIC;
		S1		:  in    STD_ULOGIC;
		D2		:  in    STD_ULOGIC;
		D3		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLM3A :  entity is TRUE;
 end DLM3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLM3A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL S0_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL S1_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (S0_ipd, S0, tipd_S0);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (S1_ipd, S1, tipd_S1);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D0_ipd, S0_ipd, D1_ipd, S1_ipd, D2_ipd, D3_ipd, G_ipd)

	-- timing check results
	VARIABLE Tviol_D0_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D0_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_S0_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_S0_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D1_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D1_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_S1_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_S1_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D2_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D2_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D3_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D3_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE NET_0_8	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D0_G_posedge,
	 TimingData		=> Tmkr_D0_G_posedge,
	 TestSignal		=> D0_ipd,
	 TestSignalName		=> "D0",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D0_G_posedge_posedge,
	 SetupLow		=> tsetup_D0_G_negedge_posedge,
	 HoldHigh		=> thold_D0_G_posedge_posedge,
	 HoldLow		=> thold_D0_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLM3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_S0_G_posedge,
	 TimingData		=> Tmkr_S0_G_posedge,
	 TestSignal		=> S0_ipd,
	 TestSignalName		=> "S0",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S0_G_posedge_posedge,
	 SetupLow		=> tsetup_S0_G_negedge_posedge,
	 HoldHigh		=> thold_S0_G_posedge_posedge,
	 HoldLow		=> thold_S0_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLM3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D1_G_posedge,
	 TimingData		=> Tmkr_D1_G_posedge,
	 TestSignal		=> D1_ipd,
	 TestSignalName		=> "D1",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D1_G_posedge_posedge,
	 SetupLow		=> tsetup_D1_G_negedge_posedge,
	 HoldHigh		=> thold_D1_G_posedge_posedge,
	 HoldLow		=> thold_D1_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLM3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_S1_G_posedge,
	 TimingData		=> Tmkr_S1_G_posedge,
	 TestSignal		=> S1_ipd,
	 TestSignalName		=> "S1",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S1_G_posedge_posedge,
	 SetupLow		=> tsetup_S1_G_negedge_posedge,
	 HoldHigh		=> thold_S1_G_posedge_posedge,
	 HoldLow		=> thold_S1_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLM3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D2_G_posedge,
	 TimingData		=> Tmkr_D2_G_posedge,
	 TestSignal		=> D2_ipd,
	 TestSignalName		=> "D2",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D2_G_posedge_posedge,
	 SetupLow		=> tsetup_D2_G_negedge_posedge,
	 HoldHigh		=> thold_D2_G_posedge_posedge,
	 HoldLow		=> thold_D2_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLM3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D3_G_posedge,
	 TimingData		=> Tmkr_D3_G_posedge,
	 TestSignal		=> D3_ipd,
	 TestSignalName		=> "D3",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D3_G_posedge_posedge,
	 SetupLow		=> tsetup_D3_G_negedge_posedge,
	 HoldHigh		=> thold_D3_G_posedge_posedge,
	 HoldLow		=> thold_D3_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLM3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TRUE, 
	 HeaderMsg		=> InstancePath & "DLM3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D0_G_posedge or Tviol_S0_G_posedge or Tviol_D1_G_posedge or 
		      Tviol_S1_G_posedge or Tviol_D2_G_posedge or Tviol_D3_G_posedge or 
		      Pviol_G;
	 --- now combinatorial logic input to the DFF 
	 NET_0_8 := 
 VitalMUX2( VitalMUX2( D0_ipd , D1_ipd , (NOT S0_ipd) ), VitalMUX2( D2_ipd , D3_ipd , (NOT S0_ipd) ), (NOT S1_ipd) );

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',G_ipd,NET_0_8, '0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D0_ipd'last_event, tpd_D0_Q, true),
		    1 => (S0_ipd'last_event, tpd_S0_Q, true),
		    2 => (D1_ipd'last_event, tpd_D1_Q, true),
		    3 => (S1_ipd'last_event, tpd_S1_Q, true),
		    4 => (D2_ipd'last_event, tpd_D2_Q, true),
		    5 => (D3_ipd'last_event, tpd_D3_Q, true),
		    6 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLM3A_VITAL of DLM3A is
   for VITAL_ACT
   end for;
end CFG_DLM3A_VITAL;



 ---- CELL DLM4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLM4 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S0_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D0_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S10_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S10_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S10_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S10_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S11_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S11_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S11_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S11_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S0_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S0_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S0_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S0_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D0_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D0_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D0_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D0_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D1_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D1_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D1_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D1_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D2_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D2_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D2_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D2_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D3_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D3_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D3_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D3_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S0		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D0		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		S10		:  in    STD_ULOGIC;
		S11		:  in    STD_ULOGIC;
		S0		:  in    STD_ULOGIC;
		D0		:  in    STD_ULOGIC;
		D1		:  in    STD_ULOGIC;
		D2		:  in    STD_ULOGIC;
		D3		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLM4 :  entity is TRUE;
 end DLM4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLM4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL S0_ipd  : STD_ULOGIC := 'X';
	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (S0_ipd, S0, tipd_S0);
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (S10_ipd, S11_ipd, S0_ipd, D0_ipd, D1_ipd, D2_ipd, D3_ipd, G_ipd)

	-- timing check results
	VARIABLE Tviol_S10_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_S10_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_S11_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_S11_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_S0_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_S0_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D0_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D0_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D1_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D1_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D2_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D2_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D3_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D3_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE NET_0_20	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S10_G_negedge,
	 TimingData		=> Tmkr_S10_G_negedge,
	 TestSignal		=> S10_ipd,
	 TestSignalName		=> "S10",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S10_G_posedge_negedge,
	 SetupLow		=> tsetup_S10_G_negedge_negedge,
	 HoldHigh		=> thold_S10_G_posedge_negedge,
	 HoldLow		=> thold_S10_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM4",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_S11_G_negedge,
	 TimingData		=> Tmkr_S11_G_negedge,
	 TestSignal		=> S11_ipd,
	 TestSignalName		=> "S11",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S11_G_posedge_negedge,
	 SetupLow		=> tsetup_S11_G_negedge_negedge,
	 HoldHigh		=> thold_S11_G_posedge_negedge,
	 HoldLow		=> thold_S11_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM4",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_S0_G_negedge,
	 TimingData		=> Tmkr_S0_G_negedge,
	 TestSignal		=> S0_ipd,
	 TestSignalName		=> "S0",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S0_G_posedge_negedge,
	 SetupLow		=> tsetup_S0_G_negedge_negedge,
	 HoldHigh		=> thold_S0_G_posedge_negedge,
	 HoldLow		=> thold_S0_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM4",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D0_G_negedge,
	 TimingData		=> Tmkr_D0_G_negedge,
	 TestSignal		=> D0_ipd,
	 TestSignalName		=> "D0",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D0_G_posedge_negedge,
	 SetupLow		=> tsetup_D0_G_negedge_negedge,
	 HoldHigh		=> thold_D0_G_posedge_negedge,
	 HoldLow		=> thold_D0_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM4",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D1_G_negedge,
	 TimingData		=> Tmkr_D1_G_negedge,
	 TestSignal		=> D1_ipd,
	 TestSignalName		=> "D1",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D1_G_posedge_negedge,
	 SetupLow		=> tsetup_D1_G_negedge_negedge,
	 HoldHigh		=> thold_D1_G_posedge_negedge,
	 HoldLow		=> thold_D1_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM4",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D2_G_negedge,
	 TimingData		=> Tmkr_D2_G_negedge,
	 TestSignal		=> D2_ipd,
	 TestSignalName		=> "D2",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D2_G_posedge_negedge,
	 SetupLow		=> tsetup_D2_G_negedge_negedge,
	 HoldHigh		=> thold_D2_G_posedge_negedge,
	 HoldLow		=> thold_D2_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM4",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D3_G_negedge,
	 TimingData		=> Tmkr_D3_G_negedge,
	 TestSignal		=> D3_ipd,
	 TestSignalName		=> "D3",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D3_G_posedge_negedge,
	 SetupLow		=> tsetup_D3_G_negedge_negedge,
	 HoldHigh		=> thold_D3_G_posedge_negedge,
	 HoldLow		=> thold_D3_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLM4",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TRUE, 
	 HeaderMsg		=> InstancePath & "DLM4",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S10_G_negedge or Tviol_S11_G_negedge or Tviol_S0_G_negedge or 
		      Tviol_D0_G_negedge or Tviol_D1_G_negedge or Tviol_D2_G_negedge or 
		      Tviol_D3_G_negedge or Pviol_G;
	 --- now combinatorial logic input to the DFF 
	 NET_0_20 := 
 VitalMUX2( VitalMUX2( VitalMUX2( D0_ipd , D1_ipd , (NOT S0_ipd) ), VitalMUX2( D2_ipd , D3_ipd , (NOT S0_ipd) ), (NOT S11_ipd) ), VitalMUX2( VitalMUX2( D2_ipd , D3_ipd , (NOT S0_ipd) ), VitalMUX2( D2_ipd , D3_ipd , (NOT S0_ipd) ), S11_ipd ), (NOT S10_ipd) );

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT G_ipd),NET_0_20, '0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (S10_ipd'last_event, tpd_S10_Q, true),
		    1 => (S11_ipd'last_event, tpd_S11_Q, true),
		    2 => (S0_ipd'last_event, tpd_S0_Q, true),
		    3 => (D0_ipd'last_event, tpd_D0_Q, true),
		    4 => (D1_ipd'last_event, tpd_D1_Q, true),
		    5 => (D2_ipd'last_event, tpd_D2_Q, true),
		    6 => (D3_ipd'last_event, tpd_D3_Q, true),
		    7 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLM4_VITAL of DLM4 is
   for VITAL_ACT
   end for;
end CFG_DLM4_VITAL;



 ---- CELL DLM4A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLM4A is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S10_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S11_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S0_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D0_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S10_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S10_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S10_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S10_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S11_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S11_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S11_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S11_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S0_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S0_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S0_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S0_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D0_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D0_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D0_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D0_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D1_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D1_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D1_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D1_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D2_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D2_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D2_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D2_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D3_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D3_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D3_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D3_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S10		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S11		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S0		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D0		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		S10		:  in    STD_ULOGIC;
		S11		:  in    STD_ULOGIC;
		S0		:  in    STD_ULOGIC;
		D0		:  in    STD_ULOGIC;
		D1		:  in    STD_ULOGIC;
		D2		:  in    STD_ULOGIC;
		D3		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLM4A :  entity is TRUE;
 end DLM4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLM4A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S10_ipd  : STD_ULOGIC := 'X';
	SIGNAL S11_ipd  : STD_ULOGIC := 'X';
	SIGNAL S0_ipd  : STD_ULOGIC := 'X';
	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (S10_ipd, S10, tipd_S10);
	VitalWireDelay (S11_ipd, S11, tipd_S11);
	VitalWireDelay (S0_ipd, S0, tipd_S0);
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (S10_ipd, S11_ipd, S0_ipd, D0_ipd, D1_ipd, D2_ipd, D3_ipd, G_ipd)

	-- timing check results
	VARIABLE Tviol_S10_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_S10_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_S11_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_S11_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_S0_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_S0_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D0_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D0_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D1_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D1_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D2_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D2_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D3_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D3_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE NET_0_20	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S10_G_posedge,
	 TimingData		=> Tmkr_S10_G_posedge,
	 TestSignal		=> S10_ipd,
	 TestSignalName		=> "S10",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S10_G_posedge_posedge,
	 SetupLow		=> tsetup_S10_G_negedge_posedge,
	 HoldHigh		=> thold_S10_G_posedge_posedge,
	 HoldLow		=> thold_S10_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLM4A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_S11_G_posedge,
	 TimingData		=> Tmkr_S11_G_posedge,
	 TestSignal		=> S11_ipd,
	 TestSignalName		=> "S11",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S11_G_posedge_posedge,
	 SetupLow		=> tsetup_S11_G_negedge_posedge,
	 HoldHigh		=> thold_S11_G_posedge_posedge,
	 HoldLow		=> thold_S11_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLM4A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_S0_G_posedge,
	 TimingData		=> Tmkr_S0_G_posedge,
	 TestSignal		=> S0_ipd,
	 TestSignalName		=> "S0",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S0_G_posedge_posedge,
	 SetupLow		=> tsetup_S0_G_negedge_posedge,
	 HoldHigh		=> thold_S0_G_posedge_posedge,
	 HoldLow		=> thold_S0_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLM4A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D0_G_posedge,
	 TimingData		=> Tmkr_D0_G_posedge,
	 TestSignal		=> D0_ipd,
	 TestSignalName		=> "D0",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D0_G_posedge_posedge,
	 SetupLow		=> tsetup_D0_G_negedge_posedge,
	 HoldHigh		=> thold_D0_G_posedge_posedge,
	 HoldLow		=> thold_D0_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLM4A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D1_G_posedge,
	 TimingData		=> Tmkr_D1_G_posedge,
	 TestSignal		=> D1_ipd,
	 TestSignalName		=> "D1",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D1_G_posedge_posedge,
	 SetupLow		=> tsetup_D1_G_negedge_posedge,
	 HoldHigh		=> thold_D1_G_posedge_posedge,
	 HoldLow		=> thold_D1_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLM4A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D2_G_posedge,
	 TimingData		=> Tmkr_D2_G_posedge,
	 TestSignal		=> D2_ipd,
	 TestSignalName		=> "D2",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D2_G_posedge_posedge,
	 SetupLow		=> tsetup_D2_G_negedge_posedge,
	 HoldHigh		=> thold_D2_G_posedge_posedge,
	 HoldLow		=> thold_D2_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLM4A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D3_G_posedge,
	 TimingData		=> Tmkr_D3_G_posedge,
	 TestSignal		=> D3_ipd,
	 TestSignalName		=> "D3",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D3_G_posedge_posedge,
	 SetupLow		=> tsetup_D3_G_negedge_posedge,
	 HoldHigh		=> thold_D3_G_posedge_posedge,
	 HoldLow		=> thold_D3_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLM4A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TRUE, 
	 HeaderMsg		=> InstancePath & "DLM4A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S10_G_posedge or Tviol_S11_G_posedge or Tviol_S0_G_posedge or 
		      Tviol_D0_G_posedge or Tviol_D1_G_posedge or Tviol_D2_G_posedge or 
		      Tviol_D3_G_posedge or Pviol_G;
	 --- now combinatorial logic input to the DFF 
	 NET_0_20 := 
 VitalMUX2( VitalMUX2( VitalMUX2( D0_ipd , D1_ipd , (NOT S0_ipd) ), VitalMUX2( D2_ipd , D3_ipd , (NOT S0_ipd) ), (NOT S11_ipd) ), VitalMUX2( VitalMUX2( D2_ipd , D3_ipd , (NOT S0_ipd) ), VitalMUX2( D2_ipd , D3_ipd , (NOT S0_ipd) ), S11_ipd ), (NOT S10_ipd) );

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',G_ipd,NET_0_20, '0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (S10_ipd'last_event, tpd_S10_Q, true),
		    1 => (S11_ipd'last_event, tpd_S11_Q, true),
		    2 => (S0_ipd'last_event, tpd_S0_Q, true),
		    3 => (D0_ipd'last_event, tpd_D0_Q, true),
		    4 => (D1_ipd'last_event, tpd_D1_Q, true),
		    5 => (D2_ipd'last_event, tpd_D2_Q, true),
		    6 => (D3_ipd'last_event, tpd_D3_Q, true),
		    7 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLM4A_VITAL of DLM4A is
   for VITAL_ACT
   end for;
end CFG_DLM4A_VITAL;



 ---- CELL DLMA ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLMA is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_A_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		A		:  in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLMA :  entity is TRUE;
 end DLMA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLMA is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd, G_ipd)

	-- timing check results
	VARIABLE Tviol_A_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_A_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_S_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_S_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_B_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_G_posedge,
	 TimingData		=> Tmkr_A_G_posedge,
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_G_posedge_posedge,
	 SetupLow		=> tsetup_A_G_negedge_posedge,
	 HoldHigh		=> thold_A_G_posedge_posedge,
	 HoldLow		=> thold_A_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLMA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_G_posedge,
	 TimingData		=> Tmkr_S_G_posedge,
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_G_posedge_posedge,
	 SetupLow		=> tsetup_S_G_negedge_posedge,
	 HoldHigh		=> thold_S_G_posedge_posedge,
	 HoldLow		=> thold_S_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLMA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_G_posedge,
	 TimingData		=> Tmkr_B_G_posedge,
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_G_posedge_posedge,
	 SetupLow		=> tsetup_B_G_negedge_posedge,
	 HoldHigh		=> thold_B_G_posedge_posedge,
	 HoldLow		=> thold_B_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLMA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TRUE, 
	 HeaderMsg		=> InstancePath & "DLMA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_A_G_posedge or Tviol_S_G_posedge or Tviol_B_G_posedge or 
		      Pviol_G;
	 --- now combinatorial logic input to the DFF 
	 NET_0_2 := 
 VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',G_ipd,NET_0_2, '0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (A_ipd'last_event, tpd_A_Q, true),
		    1 => (S_ipd'last_event, tpd_S_Q, true),
		    2 => (B_ipd'last_event, tpd_B_Q, true),
		    3 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLMA_VITAL of DLMA is
   for VITAL_ACT
   end for;
end CFG_DLMA_VITAL;



 ---- CELL DLME1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLME1A is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_A_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_E_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_E_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_E_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		A		:  in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLME1A :  entity is TRUE;
 end DLME1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLME1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (E_ipd,E, tipd_E);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd, E_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_A_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_A_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_A_E_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_A_E_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_S_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_S_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_S_E_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_S_E_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_B_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_E_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_B_E_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tviol_E_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_E_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tmkr_E_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_E		: STD_ULOGIC := '0';
	VARIABLE PInfo_E		: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_G_posedge,
	 TimingData		=> Tmkr_A_G_posedge,
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_G_posedge_posedge,
	 SetupLow		=> tsetup_A_G_negedge_posedge,
	 HoldHigh		=> thold_A_G_posedge_posedge,
	 HoldLow		=> thold_A_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((E_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLME1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_E_posedge,
	 TimingData		=> Tmkr_A_E_posedge,
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> E_ipd,
	 RefSignalName		=> "E",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_E_posedge_posedge,
	 SetupLow		=> tsetup_A_E_negedge_posedge,
	 HoldHigh               => thold_A_E_posedge_posedge,
	 HoldLow		=> thold_A_E_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((G_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLME1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_G_posedge,
	 TimingData		=> Tmkr_S_G_posedge,
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_G_posedge_posedge,
	 SetupLow		=> tsetup_S_G_negedge_posedge,
	 HoldHigh		=> thold_S_G_posedge_posedge,
	 HoldLow		=> thold_S_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((E_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLME1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_E_posedge,
	 TimingData		=> Tmkr_S_E_posedge,
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> E_ipd,
	 RefSignalName		=> "E",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_E_posedge_posedge,
	 SetupLow		=> tsetup_S_E_negedge_posedge,
	 HoldHigh               => thold_S_E_posedge_posedge,
	 HoldLow		=> thold_S_E_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((G_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLME1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_G_posedge,
	 TimingData		=> Tmkr_B_G_posedge,
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_G_posedge_posedge,
	 SetupLow		=> tsetup_B_G_negedge_posedge,
	 HoldHigh		=> thold_B_G_posedge_posedge,
	 HoldLow		=> thold_B_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((E_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLME1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_E_posedge,
	 TimingData		=> Tmkr_B_E_posedge,
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> E_ipd,
	 RefSignalName		=> "E",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_E_posedge_posedge,
	 SetupLow		=> tsetup_B_E_negedge_posedge,
	 HoldHigh               => thold_B_E_posedge_posedge,
	 HoldLow		=> thold_B_E_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((G_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLME1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_posedge,
	 TimingData             => Tmkr_E_G_posedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,	 SetupLow               => 0 ns,
	 HoldHigh               => thold_E_G_posedge_posedge,
	 HoldLow                => 0 ns,
	 CheckEnabled           =>  TRUE, 
	 RefTransition          => 'R',
	 HeaderMsg              => InstancePath & "/DLME1A",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_E_G_negedge,
	 TimingData             => Tmkr_E_G_negedge,
	 TestSignal             => E_ipd,
	 TestSignalName         => "E",
	 TestDelay              => 0 ns,
	 RefSignal              => G_ipd,
	 RefSignalName          => "G",
	 RefDelay               => 0 ns,
	 SetupHigh              => 0 ns,
	 SetupLow              => tsetup_E_G_negedge_negedge,
	 HoldHigh               => 0 ns,
	 HoldLow                => 0 ns,
	 CheckEnabled           =>  TRUE, 
	 RefTransition          => 'F',
	 HeaderMsg              => InstancePath & "/DLME1A",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLME1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_E,
	 PeriodData		=> PInfo_E,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 Period	        	=> 0 ns,
	 PulseWidthHigh		=> tpw_E_negedge,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLME1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_A_G_posedge or Tviol_A_E_posedge or Tviol_S_G_posedge or 
		      Tviol_S_E_posedge or Tviol_B_G_posedge or Tviol_B_E_posedge or 
		      Pviol_E or Pviol_G;
	 --- now combinatorial logic input to the DFF 
	 NET_0_2 := 
 VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DLE3B_Q_tab,
	 DataIn => (
		  G_ipd,E_ipd,NET_0_2, '0'));

	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (A_ipd'last_event, tpd_A_Q, true),
		    1 => (S_ipd'last_event, tpd_S_Q, true),
		    2 => (B_ipd'last_event, tpd_B_Q, true),
		     3 =>(E_ipd'last_event, tpd_E_Q, true),
		    4 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLME1A_VITAL of DLME1A is
   for VITAL_ACT
   end for;
end CFG_DLME1A_VITAL;



 ---- CELL DLP1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLP1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLP1 :  entity is TRUE;
 end DLP1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLP1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_negedge,
	 TimingData		=> Tmkr_PRE_G_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_negedge_negedge,
	 Removal		=> thold_PRE_G_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 	TRUE,
	 HeaderMsg		=> InstancePath & "DLP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or 
		       Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT G_ipd),D_ipd,PRE_ipd));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLP1_VITAL of DLP1 is
   for VITAL_ACT
   end for;
end CFG_DLP1_VITAL;



 ---- CELL DLP1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLP1A is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLP1A :  entity is TRUE;
 end DLP1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLP1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLP1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_posedge,
	 TimingData		=> Tmkr_PRE_G_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_negedge_posedge,
	 Removal		=> thold_PRE_G_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLP1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLP1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 	TRUE,
	 HeaderMsg		=> InstancePath & "DLP1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_PRE or 
		       Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',G_ipd,D_ipd,PRE_ipd));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLP1A_VITAL of DLP1A is
   for VITAL_ACT
   end for;
end CFG_DLP1A_VITAL;



 ---- CELL DLP1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLP1B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLP1B :  entity is TRUE;
 end DLP1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLP1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLP1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_negedge,
	 TimingData		=> Tmkr_PRE_G_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_posedge_negedge,
	 Removal                => thold_PRE_G_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLP1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLP1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 	TRUE,
	 HeaderMsg		=> InstancePath & "DLP1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or 
		       Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT G_ipd),D_ipd,(NOT PRE_ipd)));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLP1B_VITAL of DLP1B is
   for VITAL_ACT
   end for;
end CFG_DLP1B_VITAL;



 ---- CELL DLP1C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLP1C is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLP1C :  entity is TRUE;
 end DLP1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLP1C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLP1C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_posedge,
	 TimingData		=> Tmkr_PRE_G_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_posedge_posedge,
	 Removal                => thold_PRE_G_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLP1C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLP1C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 	TRUE,
	 HeaderMsg		=> InstancePath & "DLP1C",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_PRE or 
		       Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',G_ipd,D_ipd,(NOT PRE_ipd)));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLP1C_VITAL of DLP1C is
   for VITAL_ACT
   end for;
end CFG_DLP1C_VITAL;



 ---- CELL DLP1D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLP1D is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLP1D :  entity is TRUE;
 end DLP1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLP1D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLP1D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_negedge,
	 TimingData		=> Tmkr_PRE_G_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_posedge_negedge,
	 Removal                => thold_PRE_G_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLP1D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLP1D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 	TRUE,
	 HeaderMsg		=> InstancePath & "DLP1D",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or 
		       Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT G_ipd),D_ipd,(NOT PRE_ipd)));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_QN, true),
		    2 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLP1D_VITAL of DLP1D is
   for VITAL_ACT
   end for;
end CFG_DLP1D_VITAL;



 ---- CELL DLP1E ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLP1E is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLP1E :  entity is TRUE;
 end DLP1E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DLP1E is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLP1E",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_posedge,
	 TimingData		=> Tmkr_PRE_G_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_posedge_posedge,
	 Removal                => thold_PRE_G_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLP1E",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLP1E",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 	TRUE,
	 HeaderMsg		=> InstancePath & "DLP1E",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_PRE or 
		       Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',G_ipd,D_ipd,(NOT PRE_ipd)));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_QN, true),
		    2 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLP1E_VITAL of DLP1E is
   for VITAL_ACT
   end for;
end CFG_DLP1E_VITAL;



 ---- CELL FA1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity FA1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CI_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CI_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CI		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		CI		: in    STD_ULOGIC;
		S		: out    STD_ULOGIC;
		CO		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of FA1 :  entity is TRUE;
 end FA1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of FA1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL CI_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (CI_ipd, CI, tipd_CI);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, CI_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS S_zd : STD_LOGIC is Results(1);
	ALIAS CO_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE S_GlitchData  : VitalGlitchDataType;
	VARIABLE CO_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       S_zd := ( VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) XOR  CI_ipd );
       CO_zd := ((( A_ipd  AND  B_ipd ) OR ( A_ipd  AND  CI_ipd )) OR ( B_ipd  AND  CI_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => S,
	   GlitchData => S_GlitchData,
	   OutSignalName => "S",
	   OutTemp => S_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_S, true),
	             1 => (B_ipd'last_event,tpd_B_S, true),
	             2 => (CI_ipd'last_event,tpd_CI_S, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CO,
	   GlitchData => CO_GlitchData,
	   OutSignalName => "CO",
	   OutTemp => CO_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_CO, true),
	             1 => (B_ipd'last_event,tpd_B_CO, true),
	             2 => (CI_ipd'last_event,tpd_CI_CO, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_FA1_VITAL of FA1 is 
    for VITAL_ACT
    end for;
 end CFG_FA1_VITAL;



 ---- CELL FCEND_BUFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity FCEND_BUFF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_FCI_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_FCI		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		FCI		: in    STD_ULOGIC;
		CO		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of FCEND_BUFF :  entity is TRUE;
 end FCEND_BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of FCEND_BUFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL FCI_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (FCI_ipd, FCI, tipd_FCI);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (FCI_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS CO_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE CO_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        CO_zd :=TO_X01(FCI_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => CO,
	   GlitchData => CO_GlitchData,
	   OutSignalName => "CO",
	   OutTemp => CO_zd,
	   Paths => (
	             0 => (FCI_ipd'last_event,tpd_FCI_CO, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_FCEND_BUFF_VITAL of FCEND_BUFF is 
    for VITAL_ACT
    end for;
 end CFG_FCEND_BUFF_VITAL;



 ---- CELL FCEND_INV ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity FCEND_INV is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_FCI_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_FCI		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		FCI		: in    STD_ULOGIC;
		CO		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of FCEND_INV :  entity is TRUE;
 end FCEND_INV;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of FCEND_INV is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL FCI_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (FCI_ipd, FCI, tipd_FCI);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (FCI_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS CO_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE CO_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       CO_zd :=  (NOT FCI_ipd) ;


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => CO,
	   GlitchData => CO_GlitchData,
	   OutSignalName => "CO",
	   OutTemp => CO_zd,
	   Paths => (
	             0 => (FCI_ipd'last_event,tpd_FCI_CO, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_FCEND_INV_VITAL of FCEND_INV is 
    for VITAL_ACT
    end for;
 end CFG_FCEND_INV_VITAL;



 ---- CELL FCINIT_BUFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity FCINIT_BUFF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		FCO		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of FCINIT_BUFF :  entity is TRUE;
 end FCINIT_BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of FCINIT_BUFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS FCO_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE FCO_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        FCO_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => FCO,
	   GlitchData => FCO_GlitchData,
	   OutSignalName => "FCO",
	   OutTemp => FCO_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_FCO, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_FCINIT_BUFF_VITAL of FCINIT_BUFF is 
    for VITAL_ACT
    end for;
 end CFG_FCINIT_BUFF_VITAL;



 ---- CELL FCINIT_GND ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity FCINIT_GND is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True		);
    port(
		FCO		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of FCINIT_GND :  entity is TRUE;
 end FCINIT_GND;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of FCINIT_GND is
	attribute VITAL_LEVEL0 of VITAL_ACT : architecture is TRUE;


begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	--- Empty
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
        FCO<= '0';


end VITAL_ACT;

 configuration CFG_FCINIT_GND_VITAL of FCINIT_GND is 
    for VITAL_ACT
    end for;
 end CFG_FCINIT_GND_VITAL;



 ---- CELL FCINIT_INV ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity FCINIT_INV is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		FCO		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of FCINIT_INV :  entity is TRUE;
 end FCINIT_INV;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of FCINIT_INV is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS FCO_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE FCO_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       FCO_zd :=  (NOT A_ipd) ;


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => FCO,
	   GlitchData => FCO_GlitchData,
	   OutSignalName => "FCO",
	   OutTemp => FCO_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_FCO, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_FCINIT_INV_VITAL of FCINIT_INV is 
    for VITAL_ACT
    end for;
 end CFG_FCINIT_INV_VITAL;



 ---- CELL FCINIT_VCC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity FCINIT_VCC is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True		);
    port(
		FCO		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of FCINIT_VCC :  entity is TRUE;
 end FCINIT_VCC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of FCINIT_VCC is
	attribute VITAL_LEVEL0 of VITAL_ACT : architecture is TRUE;


begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	--- Empty
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
        FCO<= '1';


end VITAL_ACT;

 configuration CFG_FCINIT_VCC_VITAL of FCINIT_VCC is 
    for VITAL_ACT
    end for;
 end CFG_FCINIT_VCC_VITAL;



 ---- CELL GAND2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GAND2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		G		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GAND2 :  entity is TRUE;
 end GAND2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of GAND2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (G_ipd, G, tipd_G);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, G_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( A_ipd  AND  G_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (G_ipd'last_event,tpd_G_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GAND2_VITAL of GAND2 is 
    for VITAL_ACT
    end for;
 end CFG_GAND2_VITAL;



 ---- CELL GMX4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GMX4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S0		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		G		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GMX4 :  entity is TRUE;
 end GMX4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of GMX4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL S0_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (S0_ipd, S0, tipd_S0);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (G_ipd, G, tipd_G);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, S0_ipd, D1_ipd, G_ipd, D2_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( VitalMUX2( D0_ipd , D1_ipd , (NOT S0_ipd) ), VitalMUX2( D2_ipd , D3_ipd , (NOT S0_ipd) ), (NOT G_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (S0_ipd'last_event,tpd_S0_Y, true),
	             2 => (D1_ipd'last_event,tpd_D1_Y, true),
	             3 => (G_ipd'last_event,tpd_G_Y, true),
	             4 => (D2_ipd'last_event,tpd_D2_Y, true),
	             5 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GMX4_VITAL of GMX4 is 
    for VITAL_ACT
    end for;
 end CFG_GMX4_VITAL;



 ---- CELL GNAND2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GNAND2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		G		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GNAND2 :  entity is TRUE;
 end GNAND2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of GNAND2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (G_ipd, G, tipd_G);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, G_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  A_ipd  AND  G_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (G_ipd'last_event,tpd_G_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GNAND2_VITAL of GNAND2 is 
    for VITAL_ACT
    end for;
 end CFG_GNAND2_VITAL;



 ---- CELL GND ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GND is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True		);
    port(
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GND :  entity is TRUE;
 end GND;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of GND is
	attribute VITAL_LEVEL0 of VITAL_ACT : architecture is TRUE;


begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	--- Empty
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
        Y<= '0';


end VITAL_ACT;

 configuration CFG_GND_VITAL of GND is 
    for VITAL_ACT
    end for;
 end CFG_GND_VITAL;



 ---- CELL GNOR2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GNOR2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		G		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GNOR2 :  entity is TRUE;
 end GNOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of GNOR2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (G_ipd, G, tipd_G);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, G_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  A_ipd  OR  G_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (G_ipd'last_event,tpd_G_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GNOR2_VITAL of GNOR2 is 
    for VITAL_ACT
    end for;
 end CFG_GNOR2_VITAL;



 ---- CELL GOR2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GOR2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		G		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GOR2 :  entity is TRUE;
 end GOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of GOR2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (G_ipd, G, tipd_G);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, G_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( A_ipd  OR  G_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (G_ipd'last_event,tpd_G_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GOR2_VITAL of GOR2 is 
    for VITAL_ACT
    end for;
 end CFG_GOR2_VITAL;



 ---- CELL GXOR2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GXOR2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		G		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GXOR2 :  entity is TRUE;
 end GXOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of GXOR2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (G_ipd, G, tipd_G);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, G_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( G_ipd , (NOT G_ipd) , (NOT A_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (G_ipd'last_event,tpd_G_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GXOR2_VITAL of GXOR2 is 
    for VITAL_ACT
    end for;
 end CFG_GXOR2_VITAL;



 ---- CELL HA1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HA1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		S		: out    STD_ULOGIC;
		CO		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HA1 :  entity is TRUE;
 end HA1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HA1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS S_zd : STD_LOGIC is Results(1);
	ALIAS CO_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE S_GlitchData  : VitalGlitchDataType;
	VARIABLE CO_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       S_zd :=  VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) );
       CO_zd := ( A_ipd  AND  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => S,
	   GlitchData => S_GlitchData,
	   OutSignalName => "S",
	   OutTemp => S_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_S, true),
	             1 => (B_ipd'last_event,tpd_B_S, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CO,
	   GlitchData => CO_GlitchData,
	   OutSignalName => "CO",
	   OutTemp => CO_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_CO, true),
	             1 => (B_ipd'last_event,tpd_B_CO, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HA1_VITAL of HA1 is 
    for VITAL_ACT
    end for;
 end CFG_HA1_VITAL;



 ---- CELL HA1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HA1A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		S		: out    STD_ULOGIC;
		CO		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HA1A :  entity is TRUE;
 end HA1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HA1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS S_zd : STD_LOGIC is Results(1);
	ALIAS CO_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE S_GlitchData  : VitalGlitchDataType;
	VARIABLE CO_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       S_zd :=  VitalMUX2( B_ipd , (NOT B_ipd) , A_ipd );
       CO_zd := ( (NOT A_ipd)  AND  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => S,
	   GlitchData => S_GlitchData,
	   OutSignalName => "S",
	   OutTemp => S_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_S, true),
	             1 => (B_ipd'last_event,tpd_B_S, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CO,
	   GlitchData => CO_GlitchData,
	   OutSignalName => "CO",
	   OutTemp => CO_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_CO, true),
	             1 => (B_ipd'last_event,tpd_B_CO, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HA1A_VITAL of HA1A is 
    for VITAL_ACT
    end for;
 end CFG_HA1A_VITAL;



 ---- CELL HA1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HA1B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		S		: out    STD_ULOGIC;
		CO		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HA1B :  entity is TRUE;
 end HA1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HA1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS S_zd : STD_LOGIC is Results(1);
	ALIAS CO_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE S_GlitchData  : VitalGlitchDataType;
	VARIABLE CO_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       S_zd :=  NOT VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) );
       CO_zd :=  NOT (  A_ipd  AND  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => S,
	   GlitchData => S_GlitchData,
	   OutSignalName => "S",
	   OutTemp => S_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_S, true),
	             1 => (B_ipd'last_event,tpd_B_S, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CO,
	   GlitchData => CO_GlitchData,
	   OutSignalName => "CO",
	   OutTemp => CO_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_CO, true),
	             1 => (B_ipd'last_event,tpd_B_CO, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HA1B_VITAL of HA1B is 
    for VITAL_ACT
    end for;
 end CFG_HA1B_VITAL;



 ---- CELL HA1C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HA1C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_CO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		S		: out    STD_ULOGIC;
		CO		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HA1C :  entity is TRUE;
 end HA1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HA1C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS S_zd : STD_LOGIC is Results(1);
	ALIAS CO_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE S_GlitchData  : VitalGlitchDataType;
	VARIABLE CO_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       S_zd :=  VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) );
       CO_zd :=  NOT (  A_ipd  AND  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => S,
	   GlitchData => S_GlitchData,
	   OutSignalName => "S",
	   OutTemp => S_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_S, true),
	             1 => (B_ipd'last_event,tpd_B_S, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CO,
	   GlitchData => CO_GlitchData,
	   OutSignalName => "CO",
	   OutTemp => CO_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_CO, true),
	             1 => (B_ipd'last_event,tpd_B_CO, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HA1C_VITAL of HA1C is 
    for VITAL_ACT
    end for;
 end CFG_HA1C_VITAL;


 ---- CELL HCLKBIBUF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HCLKBIBUF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D			: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E			: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: inout  STD_ULOGIC;
		D		: in     STD_ULOGIC;
		E		: in     STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HCLKBIBUF :  entity is TRUE;
 end HCLKBIBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HCLKBIBUF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HCLKBIBUF_VITAL of HCLKBIBUF is 
    for VITAL_ACT
    end for;
 end CFG_HCLKBIBUF_VITAL;


 ---- CELL HCLKBUF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HCLKBUF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HCLKBUF :  entity is TRUE;
 end HCLKBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HCLKBUF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HCLKBUF_VITAL of HCLKBUF is 
    for VITAL_ACT
    end for;
 end CFG_HCLKBUF_VITAL;



 ---- CELL HCLKBUF_LVCMOS25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HCLKBUF_LVCMOS25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HCLKBUF_LVCMOS25 :  entity is TRUE;
 end HCLKBUF_LVCMOS25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HCLKBUF_LVCMOS25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HCLKBUF_LVCMOS25_VITAL of HCLKBUF_LVCMOS25 is 
    for VITAL_ACT
    end for;
 end CFG_HCLKBUF_LVCMOS25_VITAL;



 ---- CELL HCLKBUF_LVCMOS18 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HCLKBUF_LVCMOS18 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HCLKBUF_LVCMOS18 :  entity is TRUE;
 end HCLKBUF_LVCMOS18;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HCLKBUF_LVCMOS18 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HCLKBUF_LVCMOS18_VITAL of HCLKBUF_LVCMOS18 is 
    for VITAL_ACT
    end for;
 end CFG_HCLKBUF_LVCMOS18_VITAL;



 ---- CELL HCLKBUF_LVCMOS15 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HCLKBUF_LVCMOS15 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HCLKBUF_LVCMOS15 :  entity is TRUE;
 end HCLKBUF_LVCMOS15;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HCLKBUF_LVCMOS15 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HCLKBUF_LVCMOS15_VITAL of HCLKBUF_LVCMOS15 is 
    for VITAL_ACT
    end for;
 end CFG_HCLKBUF_LVCMOS15_VITAL;



 ---- CELL HCLKBUF_PCI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HCLKBUF_PCI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HCLKBUF_PCI :  entity is TRUE;
 end HCLKBUF_PCI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HCLKBUF_PCI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HCLKBUF_PCI_VITAL of HCLKBUF_PCI is 
    for VITAL_ACT
    end for;
 end CFG_HCLKBUF_PCI_VITAL;



 ---- CELL HCLKBUF_PCIX ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HCLKBUF_PCIX is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HCLKBUF_PCIX :  entity is TRUE;
 end HCLKBUF_PCIX;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HCLKBUF_PCIX is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HCLKBUF_PCIX_VITAL of HCLKBUF_PCIX is 
    for VITAL_ACT
    end for;
 end CFG_HCLKBUF_PCIX_VITAL;



 ---- CELL HCLKBUF_GTLP33 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HCLKBUF_GTLP33 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HCLKBUF_GTLP33 :  entity is TRUE;
 end HCLKBUF_GTLP33;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HCLKBUF_GTLP33 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HCLKBUF_GTLP33_VITAL of HCLKBUF_GTLP33 is 
    for VITAL_ACT
    end for;
 end CFG_HCLKBUF_GTLP33_VITAL;



 ---- CELL HCLKBUF_GTLP25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HCLKBUF_GTLP25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HCLKBUF_GTLP25 :  entity is TRUE;
 end HCLKBUF_GTLP25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HCLKBUF_GTLP25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HCLKBUF_GTLP25_VITAL of HCLKBUF_GTLP25 is 
    for VITAL_ACT
    end for;
 end CFG_HCLKBUF_GTLP25_VITAL;



 ---- CELL HCLKBUF_HSTL_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HCLKBUF_HSTL_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HCLKBUF_HSTL_I :  entity is TRUE;
 end HCLKBUF_HSTL_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HCLKBUF_HSTL_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HCLKBUF_HSTL_I_VITAL of HCLKBUF_HSTL_I is 
    for VITAL_ACT
    end for;
 end CFG_HCLKBUF_HSTL_I_VITAL;



 ---- CELL HCLKBUF_SSTL3_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HCLKBUF_SSTL3_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HCLKBUF_SSTL3_I :  entity is TRUE;
 end HCLKBUF_SSTL3_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HCLKBUF_SSTL3_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HCLKBUF_SSTL3_I_VITAL of HCLKBUF_SSTL3_I is 
    for VITAL_ACT
    end for;
 end CFG_HCLKBUF_SSTL3_I_VITAL;



 ---- CELL HCLKBUF_SSTL3_II ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HCLKBUF_SSTL3_II is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HCLKBUF_SSTL3_II :  entity is TRUE;
 end HCLKBUF_SSTL3_II;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HCLKBUF_SSTL3_II is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HCLKBUF_SSTL3_II_VITAL of HCLKBUF_SSTL3_II is 
    for VITAL_ACT
    end for;
 end CFG_HCLKBUF_SSTL3_II_VITAL;



 ---- CELL HCLKBUF_SSTL2_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HCLKBUF_SSTL2_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HCLKBUF_SSTL2_I :  entity is TRUE;
 end HCLKBUF_SSTL2_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HCLKBUF_SSTL2_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HCLKBUF_SSTL2_I_VITAL of HCLKBUF_SSTL2_I is 
    for VITAL_ACT
    end for;
 end CFG_HCLKBUF_SSTL2_I_VITAL;



 ---- CELL HCLKBUF_SSTL2_II ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HCLKBUF_SSTL2_II is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HCLKBUF_SSTL2_II :  entity is TRUE;
 end HCLKBUF_SSTL2_II;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HCLKBUF_SSTL2_II is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HCLKBUF_SSTL2_II_VITAL of HCLKBUF_SSTL2_II is 
    for VITAL_ACT
    end for;
 end CFG_HCLKBUF_SSTL2_II_VITAL;



 ---- CELL HCLKINT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HCLKINT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HCLKINT :  entity is TRUE;
 end HCLKINT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HCLKINT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HCLKINT_VITAL of HCLKINT is 
    for VITAL_ACT
    end for;
 end CFG_HCLKINT_VITAL;



 ---- CELL INBUF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF :  entity is TRUE;
 end INBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_VITAL of INBUF is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_VITAL;



 ---- CELL INBUF_LVCMOS25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS25 :  entity is TRUE;
 end INBUF_LVCMOS25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS25_VITAL of INBUF_LVCMOS25 is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS25_VITAL;



 ---- CELL INBUF_LVCMOS25D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS25D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS25D :  entity is TRUE;
 end INBUF_LVCMOS25D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS25D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','L'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS25D_VITAL of INBUF_LVCMOS25D is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS25D_VITAL;



 ---- CELL INBUF_LVCMOS25U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS25U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS25U :  entity is TRUE;
 end INBUF_LVCMOS25U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS25U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS25U_VITAL of INBUF_LVCMOS25U is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS25U_VITAL;



 ---- CELL INBUF_LVCMOS18 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS18 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS18 :  entity is TRUE;
 end INBUF_LVCMOS18;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS18 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS18_VITAL of INBUF_LVCMOS18 is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS18_VITAL;



 ---- CELL INBUF_LVCMOS18D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS18D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS18D :  entity is TRUE;
 end INBUF_LVCMOS18D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS18D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','L'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS18D_VITAL of INBUF_LVCMOS18D is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS18D_VITAL;



 ---- CELL INBUF_LVCMOS18U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS18U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS18U :  entity is TRUE;
 end INBUF_LVCMOS18U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS18U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS18U_VITAL of INBUF_LVCMOS18U is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS18U_VITAL;



 ---- CELL INBUF_LVCMOS15 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS15 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS15 :  entity is TRUE;
 end INBUF_LVCMOS15;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS15 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS15_VITAL of INBUF_LVCMOS15 is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS15_VITAL;



 ---- CELL INBUF_LVCMOS15D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS15D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS15D :  entity is TRUE;
 end INBUF_LVCMOS15D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS15D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','L'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS15D_VITAL of INBUF_LVCMOS15D is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS15D_VITAL;



 ---- CELL INBUF_LVCMOS15U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS15U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS15U :  entity is TRUE;
 end INBUF_LVCMOS15U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS15U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS15U_VITAL of INBUF_LVCMOS15U is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS15U_VITAL;



 ---- CELL INBUF_PCI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_PCI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_PCI :  entity is TRUE;
 end INBUF_PCI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_PCI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_PCI_VITAL of INBUF_PCI is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_PCI_VITAL;



 ---- CELL INBUF_PCIX ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_PCIX is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_PCIX :  entity is TRUE;
 end INBUF_PCIX;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_PCIX is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_PCIX_VITAL of INBUF_PCIX is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_PCIX_VITAL;



 ---- CELL INBUF_GTLP33 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_GTLP33 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_GTLP33 :  entity is TRUE;
 end INBUF_GTLP33;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_GTLP33 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_GTLP33_VITAL of INBUF_GTLP33 is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_GTLP33_VITAL;



 ---- CELL INBUF_GTLP25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_GTLP25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_GTLP25 :  entity is TRUE;
 end INBUF_GTLP25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_GTLP25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_GTLP25_VITAL of INBUF_GTLP25 is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_GTLP25_VITAL;



 ---- CELL INBUF_HSTL_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_HSTL_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_HSTL_I :  entity is TRUE;
 end INBUF_HSTL_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_HSTL_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_HSTL_I_VITAL of INBUF_HSTL_I is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_HSTL_I_VITAL;



 ---- CELL INBUF_SSTL3_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_SSTL3_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_SSTL3_I :  entity is TRUE;
 end INBUF_SSTL3_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_SSTL3_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_SSTL3_I_VITAL of INBUF_SSTL3_I is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_SSTL3_I_VITAL;



 ---- CELL INBUF_SSTL3_II ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_SSTL3_II is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_SSTL3_II :  entity is TRUE;
 end INBUF_SSTL3_II;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_SSTL3_II is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_SSTL3_II_VITAL of INBUF_SSTL3_II is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_SSTL3_II_VITAL;



 ---- CELL INBUF_SSTL2_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_SSTL2_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_SSTL2_I :  entity is TRUE;
 end INBUF_SSTL2_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_SSTL2_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_SSTL2_I_VITAL of INBUF_SSTL2_I is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_SSTL2_I_VITAL;



 ---- CELL INBUF_SSTL2_II ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_SSTL2_II is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_SSTL2_II :  entity is TRUE;
 end INBUF_SSTL2_II;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INBUF_SSTL2_II is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_SSTL2_II_VITAL of INBUF_SSTL2_II is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_SSTL2_II_VITAL;



 ---- CELL INV ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INV is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INV :  entity is TRUE;
 end INV;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INV is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  (NOT A_ipd) ;


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INV_VITAL of INV is 
    for VITAL_ACT
    end for;
 end CFG_INV_VITAL;



 ---- CELL INVA ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INVA is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INVA :  entity is TRUE;
 end INVA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INVA is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  (NOT A_ipd) ;


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INVA_VITAL of INVA is 
    for VITAL_ACT
    end for;
 end CFG_INVA_VITAL;



 ---- CELL INVD ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INVD is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INVD :  entity is TRUE;
 end INVD;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of INVD is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  (NOT A_ipd) ;


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INVD_VITAL of INVD is 
    for VITAL_ACT
    end for;
 end CFG_INVD_VITAL;



 ---- CELL IOI_DFEG ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOI_DFEG is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOI_DFEG :  entity is TRUE;
 end IOI_DFEG;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOI_DFEG is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOI_DFEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOI_DFEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOI_DFEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOI_DFEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "IOI_DFEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "IOI_DFEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "IOI_DFEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, D_delayed, E_delayed, PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOI_DFEG_VITAL of IOI_DFEG is
   for VITAL_ACT
   end for;
end CFG_IOI_DFEG_VITAL;



 ---- CELL IOI_DFEH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOI_DFEH is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOI_DFEH :  entity is TRUE;
 end IOI_DFEH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOI_DFEH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/IOI_DFEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (CLR_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "IOI_DFEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "IOI_DFEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "IOI_DFEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "IOI_DFEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "IOI_DFEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "IOI_DFEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or 
	 Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, Q_zd, D_delayed, E_delayed, PRE_ipd, CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOI_DFEH_VITAL of IOI_DFEH is
   for VITAL_ACT
   end for;
end CFG_IOI_DFEH_VITAL;



 ---- CELL IOI_BUFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOI_BUFF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOI_BUFF :  entity is TRUE;
 end IOI_BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOI_BUFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOI_BUFF_VITAL of IOI_BUFF is 
    for VITAL_ACT
    end for;
 end CFG_IOI_BUFF_VITAL;



 ---- CELL IOOE_BUFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOOE_BUFF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOOE_BUFF :  entity is TRUE;
 end IOOE_BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOOE_BUFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOOE_BUFF_VITAL of IOOE_BUFF is 
    for VITAL_ACT
    end for;
 end CFG_IOOE_BUFF_VITAL;



 ---- CELL IOOE_DFEG ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOOE_DFEG is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_YOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_YOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_YOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tperiod_CLK_negedge        :  VitalDelayType := 0.000 ns;
		tpw_CLK_posedge        :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge        :  VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                CLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                Q                : out    STD_ULOGIC;
                YOUT                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOOE_DFEG :  entity is TRUE;
 end IOOE_DFEG;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOOE_DFEG is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd, E_ipd, PRE_ipd)


   VARIABLE Tviol_D_CLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_E_CLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_YOUT  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS YOUT_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData  : VitalGlitchDataType;
   VARIABLE YOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_CLK_posedge,
   TimingData             => Tmkr_D_CLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => CLK_ipd,
   RefSignalName          => "CLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_CLK_posedge_posedge,
   SetupLow               => tsetup_D_CLK_negedge_posedge,
   HoldHigh              => thold_D_CLK_posedge_posedge,
   HoldLow                => thold_D_CLK_negedge_posedge,
   CheckEnabled           => TO_X01((NOT E_ipd) AND PRE_ipd AND CLR_ipd) /='0',
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOOE_DFEG",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_CLK_posedge,
   TimingData             => Tmkr_CLR_CLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => CLK_ipd,
   RefSignalName          => "CLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_CLK_posedge_posedge,
   Removal                => thold_CLR_CLK_posedge_posedge,
   ActiveLow               => TRUE,
   CheckEnabled           => TO_X01((NOT E_ipd) AND PRE_ipd) /='0',
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOOE_DFEG",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthLow => tpw_CLR_negedge,
    PulseWidthHigh         => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOOE_DFEG",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_CLK_posedge,
   TimingData             => Tmkr_E_CLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => CLK_ipd,
   RefSignalName          => "CLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_CLK_posedge_posedge,
   SetupLow               => tsetup_E_CLK_negedge_posedge,
   HoldHigh              => thold_E_CLK_posedge_posedge,
   HoldLow                => thold_E_CLK_negedge_posedge,
   CheckEnabled           => TO_X01(PRE_ipd AND CLR_ipd) /='0',
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOOE_DFEG",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_CLK_posedge,
   TimingData             => Tmkr_PRE_CLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => CLK_ipd,
   RefSignalName          => "CLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_CLK_posedge_posedge,
   Removal                => thold_PRE_CLK_posedge_posedge,
   ActiveLow               => TRUE,
   CheckEnabled           => TO_X01((NOT E_ipd) AND CLR_ipd) /='0' ,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOOE_DFEG",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthLow => tpw_PRE_negedge,
    PulseWidthHigh         => 0 ns,
    CheckEnabled           => TO_X01(CLR_ipd) /= '0',
    HeaderMsg              => InstancePath & "IOOE_DFEG",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_CLK_posedge  or Tviol_CLR_CLK_posedge  or Pviol_CLR or Tviol_E_CLK_posedge  or Tviol_PRE_CLK_posedge  or Pviol_PRE;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, D_delayed, E_delayed, PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;

  VitalStateTable(
   Result => YOUT_zd,
   PreviousDataIn => PrevData_YOUT,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, YOUT_zd, D_delayed, E_delayed, PRE_ipd, CLK_ipd));
   YOUT_zd := Violation XOR YOUT_zd;

   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => Q,
    GlitchData => Q_GlitchData,
    OutSignalName => "Q",
    OutTemp => Q_zd,
    Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
              1 => (PRE_ipd'last_event, tpd_PRE_Q, true),
              2 => (CLR_ipd'last_event, tpd_CLR_Q, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => YOUT,
    GlitchData => YOUT_GlitchData,
    OutSignalName => "YOUT",
    OutTemp => YOUT_zd,
    Paths => (0 => (CLK_ipd'last_event, tpd_CLK_YOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_YOUT, true),
              2 => (CLR_ipd'last_event, tpd_CLR_YOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOOE_DFEG_VITAL of IOOE_DFEG is
   for VITAL_ACT
   end for;
end CFG_IOOE_DFEG_VITAL;



 ---- CELL IOOE_DFEH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOOE_DFEH is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_YOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_YOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_YOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge   :   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge	:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge       :   VitalDelayType := 0.000 ns;
		tperiod_CLK_negedge        :  VitalDelayType := 0.000 ns;
		tpw_CLK_posedge        :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge        :  VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge   :   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge	:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                CLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                Q                : out    STD_ULOGIC;
                YOUT                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOOE_DFEH :  entity is TRUE;
 end IOOE_DFEH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOOE_DFEH is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd, E_ipd, PRE_ipd)


   VARIABLE Tviol_D_CLK_negedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_E_CLK_negedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_negedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_YOUT  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS YOUT_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData  : VitalGlitchDataType;
   VARIABLE YOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_CLK_negedge, 
   TimingData             => Tmkr_D_CLK_negedge, 
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => CLK_ipd,
   RefSignalName          => "CLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_CLK_posedge_negedge,
   SetupLow               => tsetup_D_CLK_negedge_negedge,
   HoldHigh              => thold_D_CLK_posedge_negedge,
   HoldLow                => thold_D_CLK_negedge_negedge,
   CheckEnabled           => TO_X01((NOT E_ipd) AND CLR_ipd AND PRE_ipd) /='0',
   RefTransition          => 'F',
   HeaderMsg              => InstancePath & "/IOOE_DFEH",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_CLK_negedge,
   TimingData             => Tmkr_CLR_CLK_negedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => CLK_ipd,
   RefSignalName          => "CLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_CLK_posedge_negedge,
   Removal                => thold_CLR_CLK_posedge_negedge,
   ActiveLow               => TRUE,
   CheckEnabled           => TO_X01((NOT E_ipd) AND PRE_ipd) /= '0',
   RefTransition          => 'F',
   HeaderMsg              => InstancePath & "IOOE_DFEH",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthLow => tpw_CLR_negedge,
    PulseWidthHigh         => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOOE_DFEH",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_CLK_negedge, 
   TimingData             => Tmkr_E_CLK_negedge, 
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => CLK_ipd,
   RefSignalName          => "CLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_CLK_posedge_negedge,
   SetupLow               => tsetup_E_CLK_negedge_negedge,
   HoldHigh              => thold_E_CLK_posedge_negedge,
   HoldLow                => thold_E_CLK_negedge_negedge,
   CheckEnabled           => TO_X01(PRE_ipd AND CLR_ipd) /= '0',
   RefTransition          => 'F',
   HeaderMsg              => InstancePath & "/IOOE_DFEH",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_CLK_negedge,
   TimingData             => Tmkr_PRE_CLK_negedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => CLK_ipd,
   RefSignalName          => "CLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_CLK_posedge_negedge,
   Removal                => thold_PRE_CLK_posedge_negedge,
   ActiveLow              => TRUE,
   CheckEnabled           => TO_X01(CLR_ipd AND (NOT E_ipd)) /='1',
   RefTransition          => 'F',
   HeaderMsg              => InstancePath & "IOOE_DFEH",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthLow => tpw_PRE_negedge,
    PulseWidthHigh         => 0 ns,
    CheckEnabled           => TO_X01(CLR_ipd) /='0',
    HeaderMsg              => InstancePath & "IOOE_DFEH",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_CLK_negedge  or Tviol_CLR_CLK_negedge  or Pviol_CLR or Tviol_E_CLK_negedge  or Tviol_PRE_CLK_negedge  or Pviol_PRE;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, Q_zd, D_delayed, E_delayed, PRE_ipd, CLK_delayed));
   Q_zd := Violation XOR Q_zd;

  VitalStateTable(
   Result => YOUT_zd,
   PreviousDataIn => PrevData_YOUT,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, YOUT_zd, D_delayed, E_delayed, PRE_ipd, CLK_delayed));
   YOUT_zd := Violation XOR YOUT_zd;

   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => Q,
    GlitchData => Q_GlitchData,
    OutSignalName => "Q",
    OutTemp => Q_zd,
    Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
              1 => (PRE_ipd'last_event, tpd_PRE_Q, true),
              2 => (CLR_ipd'last_event, tpd_CLR_Q, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => YOUT,
    GlitchData => YOUT_GlitchData,
    OutSignalName => "YOUT",
    OutTemp => YOUT_zd,
    Paths => (0 => (CLK_ipd'last_event, tpd_CLK_YOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_YOUT, true),
              2 => (CLR_ipd'last_event, tpd_CLR_YOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOOE_DFEH_VITAL of IOOE_DFEH is
   for VITAL_ACT
   end for;
end CFG_IOOE_DFEH_VITAL;



 ---- CELL IOPAD_IN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_IN is
    generic (
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
-- DNW: Add the following 2 lines
		tpw_PAD_posedge		: VitalDelayType := 0.000 ns;
		tpw_PAD_negedge		: VitalDelayType := 0.000 ns;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns)
            );

    port (
		PAD		: in    STD_ULOGIC;
		Y		: out   STD_ULOGIC
         );
 attribute VITAL_LEVEL0 of IOPAD_IN :  entity is TRUE;
 end IOPAD_IN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOPAD_IN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd       : STD_LOGIC is Results(1);

-- DNW: Add the following 4 lines
	-- timing check results
	VARIABLE Pviol_PAD       : STD_ULOGIC := '0';
	VARIABLE PeriodData_PAD  : VitalPeriodDataType := VitalPeriodDataInit;

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

-- DNW: Add the following 20 lines
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_IN",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------

           Y_zd :=TO_X01(PAD_ipd);

	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOPAD_IN_VITAL of IOPAD_IN is 
    for VITAL_ACT
    end for;
 end CFG_IOPAD_IN_VITAL;



 ---- CELL IOPAD_TRI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_TRI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		
                tpw_D_posedge 		: VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge 	 	: VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                
                tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPAD_TRI :  entity is TRUE;
 end IOPAD_TRI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOPAD_TRI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- timing check results
	VARIABLE Pviol_E       : STD_ULOGIC := '0';
	VARIABLE PeriodData_E  : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_D       : STD_ULOGIC := '0';
	VARIABLE PeriodData_D  : VitalPeriodDataType := VitalPeriodDataInit;

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_E, 
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_TRI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

            VitalPeriodPulseCheck (
              Violation      => Pviol_D, 
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_TRI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_IOPAD_TRI_VITAL of IOPAD_TRI is 
    for VITAL_ACT
    end for;
 end CFG_IOPAD_TRI_VITAL;



 ---- CELL IOPAD_BI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_BI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPAD_BI :  entity is TRUE;
 end IOPAD_BI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOPAD_BI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

        -- timing check results
	VARIABLE Pviol_D	:STD_ULOGIC := '0';
        VARIABLE PeriodData_D        :VitalPeriodDataType := VitalPeriodDataInit;
 	VARIABLE Pviol_E	:STD_ULOGIC := '0';
        VARIABLE PeriodData_E        :VitalPeriodDataType := VitalPeriodDataInit;	
        VARIABLE Pviol_PAD	:STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD        :VitalPeriodDataType := VitalPeriodDataInit;     

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin
         
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );
 

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );
          
        end if;
	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOPAD_BI_VITAL of IOPAD_BI is 
    for VITAL_ACT
    end for;
 end CFG_IOPAD_BI_VITAL;



 ---- CELL JKF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity JKF is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_J_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_J_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_J_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		thold_J_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_K_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		thold_K_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge		:  VitalDelayType := 0.000 ns;
		tipd_J      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_K      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK	:   VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		J	:  in    STD_ULOGIC;
		K	:  in    STD_ULOGIC;
	        CLK	:  in    STD_ULOGIC;
		Q	:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of JKF :  entity is FALSE;
 end JKF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of JKF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

	SIGNAL J_ipd  : STD_ULOGIC := 'X';
	SIGNAL K_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (J_ipd, J, tipd_J);
	VitalWireDelay (K_ipd, K, tipd_K);
	VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (J_ipd, K_ipd, CLK_ipd)

	-- timing check results
	VARIABLE Tviol_J_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_J_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_K_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_K_CLK_posedge		:  VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK  : STD_ULOGIC := '0';
	VARIABLE PInfo_CLK  : VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation      : STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 5);
	VARIABLE CLK_delayed        : STD_ULOGIC := 'X';
	VARIABLE J_delayed        : STD_ULOGIC := 'X';
	VARIABLE K_delayed        : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_J_CLK_posedge,
	 TimingData		=> Tmkr_J_CLK_posedge,
	 TestSignal		=> J_ipd,
	 TestSignalName		=> "J",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_J_CLK_posedge_posedge,
	 SetupLow		=> tsetup_J_CLK_negedge_posedge,
	 HoldHigh		=> thold_J_CLK_posedge_posedge,
	 HoldLow		=> thold_J_CLK_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/JKF",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_K_CLK_posedge,
	 TimingData             => Tmkr_K_CLK_posedge,
	 TestSignal             => K_ipd,
	 TestSignalName         => "K",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 SetupHigh              => tsetup_K_CLK_posedge_posedge,
	 SetupLow               => tsetup_K_CLK_negedge_posedge,
	 HoldHigh               => thold_K_CLK_posedge_posedge,
	 HoldLow                => thold_K_CLK_negedge_posedge,
	 CheckEnabled           =>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/JKF",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh => tpw_CLK_posedge,
	 PulseWidthLow => tpw_CLK_negedge,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "JKF",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

	 Violation := Tviol_J_CLK_posedge or 
	 Tviol_K_CLK_posedge or 
   Pviol_CLK;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => JKF2A_Q_tab,
	 DataIn => (
             '1', CLK_delayed, K_delayed, J_delayed, Q_zd, CLK_ipd));
	 Q_zd := Violation XOR Q_zd;
	  --- now combinatorial logic input to the DFF 
	 J_delayed :=  J_ipd ;
          --- now combinatorial logic input to the DFF 
         K_delayed :=  (NOT K_ipd) ;
	 CLK_delayed := CLK_ipd;

	 ----------------------
	 --  Path Delay Section
	 ----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_JKF_VITAL of JKF is
   for VITAL_ACT
   end for;
end CFG_JKF_VITAL;



 ---- CELL JKF1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity JKF1B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_J_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_J_CLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
		tsetup_J_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		thold_J_CLK_negedge_negedge   :   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_K_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		thold_K_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge		:  VitalDelayType := 0.000 ns;
		tipd_J      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_K      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK	:   VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		J	:  in    STD_ULOGIC;
		K	:  in    STD_ULOGIC;
	        CLK	:  in    STD_ULOGIC;
		Q	:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of JKF1B :  entity is FALSE;
 end JKF1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of JKF1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

	SIGNAL J_ipd  : STD_ULOGIC := 'X';
	SIGNAL K_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (J_ipd, J, tipd_J);
	VitalWireDelay (K_ipd, K, tipd_K);
	VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (J_ipd, K_ipd, CLK_ipd)

	-- timing check results
	VARIABLE Tviol_J_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_J_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_K_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_K_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK  : STD_ULOGIC := '0';
	VARIABLE PInfo_CLK  : VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation      : STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 5);
	VARIABLE CLK_delayed        : STD_ULOGIC := 'X';
	VARIABLE J_delayed        : STD_ULOGIC := 'X';
	VARIABLE K_delayed        : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_J_CLK_negedge,
	 TimingData		=> Tmkr_J_CLK_negedge,
	 TestSignal		=> J_ipd,
	 TestSignalName		=> "J",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_J_CLK_posedge_negedge,
	 SetupLow		=> tsetup_J_CLK_negedge_negedge,
	 HoldHigh		=> thold_J_CLK_posedge_negedge,
	 HoldLow		=> thold_J_CLK_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/JKF1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_K_CLK_negedge,
	 TimingData             => Tmkr_K_CLK_negedge,
	 TestSignal             => K_ipd,
	 TestSignalName         => "K",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 SetupHigh              => tsetup_K_CLK_posedge_negedge,
	 SetupLow               => tsetup_K_CLK_negedge_negedge,
	 HoldHigh               => thold_K_CLK_posedge_negedge,
	 HoldLow                => thold_K_CLK_negedge_negedge,
	 CheckEnabled           =>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/JKF1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh => tpw_CLK_negedge,
	 PulseWidthLow => tpw_CLK_posedge,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "JKF1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

	 Violation := Tviol_J_CLK_negedge or 
	 Tviol_K_CLK_negedge or 
   Pviol_CLK;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => JKF2A_Q_tab,
	 DataIn => (
             '1', CLK_ipd, K_delayed, J_delayed, Q_zd, CLK_delayed));
	 Q_zd := Violation XOR Q_zd;
	  --- now combinatorial logic input to the DFF 
	 J_delayed :=  J_ipd ;
          --- now combinatorial logic input to the DFF 
         K_delayed :=  (NOT K_ipd) ;
	 CLK_delayed := CLK_ipd;

	 ----------------------
	 --  Path Delay Section
	 ----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_JKF1B_VITAL of JKF1B is
   for VITAL_ACT
   end for;
end CFG_JKF1B_VITAL;



 ---- CELL JKF2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity JKF2A is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_J_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_J_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_J_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		thold_J_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_K_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		thold_K_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge	:  VitalDelayType := 0.000 ns;
		tipd_CLR	:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_J      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_K      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK	:   VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		J	:  in    STD_ULOGIC;
		K	:  in    STD_ULOGIC;
	        CLR	:  in    STD_ULOGIC;
	        CLK	:  in    STD_ULOGIC;
		Q	:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of JKF2A :  entity is FALSE;
 end JKF2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of JKF2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

	SIGNAL J_ipd  : STD_ULOGIC := 'X';
	SIGNAL K_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (J_ipd, J, tipd_J);
	VitalWireDelay (K_ipd, K, tipd_K);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (J_ipd, K_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_J_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_J_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_K_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_K_CLK_posedge		:  VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK  : STD_ULOGIC := '0';
	VARIABLE PInfo_CLK  : VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
	VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation      : STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 5);
	VARIABLE CLK_delayed        : STD_ULOGIC := 'X';
	VARIABLE J_delayed        : STD_ULOGIC := 'X';
	VARIABLE K_delayed        : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_J_CLK_posedge,
	 TimingData		=> Tmkr_J_CLK_posedge,
	 TestSignal		=> J_ipd,
	 TestSignalName		=> "J",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_J_CLK_posedge_posedge,
	 SetupLow		=> tsetup_J_CLK_negedge_posedge,
	 HoldHigh		=> thold_J_CLK_posedge_posedge,
	 HoldLow		=> thold_J_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01((CLR_ipd)) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/JKF2A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_K_CLK_posedge,
	 TimingData             => Tmkr_K_CLK_posedge,
	 TestSignal             => K_ipd,
	 TestSignalName         => "K",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 SetupHigh              => tsetup_K_CLK_posedge_posedge,
	 SetupLow               => tsetup_K_CLK_negedge_posedge,
	 HoldHigh               => thold_K_CLK_posedge_posedge,
	 HoldLow                => thold_K_CLK_negedge_posedge,
	 CheckEnabled           =>  TO_X01((CLR_ipd)) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/JKF2A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_CLK_posedge,
	 TimingData		=> Tmkr_CLR_CLK_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_CLK_posedge_posedge,
	 Removal		=> thold_CLR_CLK_posedge_posedge,
	 ActiveLow              => TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition          => 'R',
	 HeaderMsg              => InstancePath & "JKF2A",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh => tpw_CLK_posedge,
	 PulseWidthLow => tpw_CLK_negedge,
	 CheckEnabled		=> TO_X01((CLR_ipd)) /= '0',
	 HeaderMsg		=> InstancePath & "JKF2A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "JKF2A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

	 Violation := Tviol_J_CLK_posedge or 
	 Tviol_K_CLK_posedge or 
   Pviol_CLR or 
	 Pviol_CLK;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => JKF2A_Q_tab,
	 DataIn => (
             CLR_ipd, CLK_delayed, K_delayed, J_delayed, Q_zd, CLK_ipd));
	 Q_zd := Violation XOR Q_zd;
	  --- now combinatorial logic input to the DFF 
	 J_delayed :=  J_ipd ;
          --- now combinatorial logic input to the DFF 
         K_delayed :=  (NOT K_ipd) ;
	 CLK_delayed := CLK_ipd;

	 ----------------------
	 --  Path Delay Section
	 ----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1 => (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_JKF2A_VITAL of JKF2A is
   for VITAL_ACT
   end for;
end CFG_JKF2A_VITAL;



 ---- CELL JKF2B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity JKF2B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_J_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_J_CLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
		tsetup_J_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		thold_J_CLK_negedge_negedge   :   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_K_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		thold_K_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge           :   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge	:  VitalDelayType := 0.000 ns;
		tipd_CLR	:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_J      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_K      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK	:   VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		J	:  in    STD_ULOGIC;
		K	:  in    STD_ULOGIC;
	        CLR	:  in    STD_ULOGIC;
	        CLK	:  in    STD_ULOGIC;
		Q	:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of JKF2B :  entity is FALSE;
 end JKF2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of JKF2B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

	SIGNAL J_ipd  : STD_ULOGIC := 'X';
	SIGNAL K_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (J_ipd, J, tipd_J);
	VitalWireDelay (K_ipd, K, tipd_K);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (J_ipd, K_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_J_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_J_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_K_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_K_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK  : STD_ULOGIC := '0';
	VARIABLE PInfo_CLK  : VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
	VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation      : STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 5);
	VARIABLE CLK_delayed        : STD_ULOGIC := 'X';
	VARIABLE J_delayed        : STD_ULOGIC := 'X';
	VARIABLE K_delayed        : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_J_CLK_negedge,
	 TimingData		=> Tmkr_J_CLK_negedge,
	 TestSignal		=> J_ipd,
	 TestSignalName		=> "J",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_J_CLK_posedge_negedge,
	 SetupLow		=> tsetup_J_CLK_negedge_negedge,
	 HoldHigh		=> thold_J_CLK_posedge_negedge,
	 HoldLow		=> thold_J_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01((CLR_ipd)) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/JKF2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_K_CLK_negedge,
	 TimingData             => Tmkr_K_CLK_negedge,
	 TestSignal             => K_ipd,
	 TestSignalName         => "K",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 SetupHigh              => tsetup_K_CLK_posedge_negedge,
	 SetupLow               => tsetup_K_CLK_negedge_negedge,
	 HoldHigh               => thold_K_CLK_posedge_negedge,
	 HoldLow                => thold_K_CLK_negedge_negedge,
	 CheckEnabled           =>  TO_X01((CLR_ipd)) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/JKF2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_CLK_negedge,
	 TimingData		=> Tmkr_CLR_CLK_negedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_CLK_posedge_negedge,
	 Removal		=> thold_CLR_CLK_posedge_negedge,
	 ActiveLow              => TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition          => 'F',
	 HeaderMsg              => InstancePath & "JKF2B",
	 Xon            => Xon,
	 MsgOn          => MsgOn,
	 MsgSeverity            => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh => tpw_CLK_negedge,
	 PulseWidthLow => tpw_CLK_posedge,
	 CheckEnabled		=> TO_X01((CLR_ipd)) /= '0',
	 HeaderMsg		=> InstancePath & "JKF2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "JKF2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

	 Violation := Tviol_J_CLK_negedge or 
	 Tviol_K_CLK_negedge or 
   Pviol_CLR or 
	 Pviol_CLK;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => JKF2A_Q_tab,
	 DataIn => (
             CLR_ipd, CLK_ipd, K_delayed, J_delayed, Q_zd, CLK_delayed));
	 Q_zd := Violation XOR Q_zd;
	  --- now combinatorial logic input to the DFF 
	 J_delayed :=  J_ipd ;
          --- now combinatorial logic input to the DFF 
         K_delayed :=  (NOT K_ipd) ;
	 CLK_delayed := CLK_ipd;

	 ----------------------
	 --  Path Delay Section
	 ----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1 => (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_JKF2B_VITAL of JKF2B is
   for VITAL_ACT
   end for;
end CFG_JKF2B_VITAL;



 ---- CELL JKF3A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity JKF3A is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_J_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_J_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_J_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		thold_J_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_K_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		thold_K_CLK_negedge_posedge           :   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge   	:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE	:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_J      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_K      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK	:   VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		J	:  in    STD_ULOGIC;
		K	:  in    STD_ULOGIC;
	        PRE	:  in    STD_ULOGIC;
	        CLK	:  in    STD_ULOGIC;
		Q	:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of JKF3A :  entity is FALSE;
 end JKF3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of JKF3A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

	SIGNAL J_ipd  : STD_ULOGIC := 'X';
	SIGNAL K_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (J_ipd, J, tipd_J);
	VitalWireDelay (K_ipd, K, tipd_K);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (J_ipd, K_ipd, PRE_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_J_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_J_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_K_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_K_CLK_posedge		:  VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK  : STD_ULOGIC := '0';
	VARIABLE PInfo_CLK  : VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
	VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation      : STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 5);
	VARIABLE CLK_delayed        : STD_ULOGIC := 'X';
	VARIABLE J_delayed        : STD_ULOGIC := 'X';
	VARIABLE K_delayed        : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_J_CLK_posedge,
	 TimingData		=> Tmkr_J_CLK_posedge,
	 TestSignal		=> J_ipd,
	 TestSignalName		=> "J",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_J_CLK_posedge_posedge,
	 SetupLow		=> tsetup_J_CLK_negedge_posedge,
	 HoldHigh		=> thold_J_CLK_posedge_posedge,
	 HoldLow		=> thold_J_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01((PRE_ipd)) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/JKF3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_K_CLK_posedge,
	 TimingData             => Tmkr_K_CLK_posedge,
	 TestSignal             => K_ipd,
	 TestSignalName         => "K",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 SetupHigh              => tsetup_K_CLK_posedge_posedge,
	 SetupLow               => tsetup_K_CLK_negedge_posedge,
	 HoldHigh               => thold_K_CLK_posedge_posedge,
	 HoldLow                => thold_K_CLK_negedge_posedge,
	 CheckEnabled           =>  TO_X01((PRE_ipd)) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/JKF3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay	=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
   CheckEnabled		=>   TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg              => InstancePath & "JKF3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh => tpw_CLK_posedge,
	 PulseWidthLow => tpw_CLK_negedge,
	 CheckEnabled		=> TO_X01((PRE_ipd)) /= '0',
	 HeaderMsg		=> InstancePath & "JKF3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow		=> tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> TRUE, 
	 HeaderMsg		=> InstancePath & "JKF3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

	 Violation := Tviol_J_CLK_posedge or 
	 Tviol_K_CLK_posedge or 
   Tviol_PRE_CLK_posedge or 
	 Pviol_PRE or Pviol_CLK;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
   StateTable => JKF3A_Q_tab,
   DataIn => (
CLK_delayed, K_delayed, J_delayed, Q_zd, PRE_ipd, CLK_ipd));
	 Q_zd := Violation XOR Q_zd;
	  --- now combinatorial logic input to the DFF 
	 J_delayed :=  J_ipd ;
          --- now combinatorial logic input to the DFF 
         K_delayed :=  (NOT K_ipd) ;
	 CLK_delayed := CLK_ipd;

	 ----------------------
	 --  Path Delay Section
	 ----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1 => (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_JKF3A_VITAL of JKF3A is
   for VITAL_ACT
   end for;
end CFG_JKF3A_VITAL;



 ---- CELL JKF3B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity JKF3B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_J_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_J_CLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
		tsetup_J_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		thold_J_CLK_negedge_negedge   :   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_K_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_K_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		thold_K_CLK_negedge_negedge           :   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge   	:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE	:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_J      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_K      :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK	:   VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		J	:  in    STD_ULOGIC;
		K	:  in    STD_ULOGIC;
	        PRE	:  in    STD_ULOGIC;
	        CLK	:  in    STD_ULOGIC;
		Q	:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of JKF3B :  entity is FALSE;
 end JKF3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of JKF3B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

	SIGNAL J_ipd  : STD_ULOGIC := 'X';
	SIGNAL K_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (J_ipd, J, tipd_J);
	VitalWireDelay (K_ipd, K, tipd_K);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (J_ipd, K_ipd, PRE_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_J_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_J_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_K_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_K_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK  : STD_ULOGIC := '0';
	VARIABLE PInfo_CLK  : VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
	VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation      : STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 5);
	VARIABLE CLK_delayed        : STD_ULOGIC := 'X';
	VARIABLE J_delayed        : STD_ULOGIC := 'X';
	VARIABLE K_delayed        : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_J_CLK_negedge,
	 TimingData		=> Tmkr_J_CLK_negedge,
	 TestSignal		=> J_ipd,
	 TestSignalName		=> "J",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_J_CLK_posedge_negedge,
	 SetupLow		=> tsetup_J_CLK_negedge_negedge,
	 HoldHigh		=> thold_J_CLK_posedge_negedge,
	 HoldLow		=> thold_J_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01((PRE_ipd)) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/JKF3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalSetupHoldCheck (
	 Violation              => Tviol_K_CLK_negedge,
	 TimingData             => Tmkr_K_CLK_negedge,
	 TestSignal             => K_ipd,
	 TestSignalName         => "K",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 SetupHigh              => tsetup_K_CLK_posedge_negedge,
	 SetupLow               => tsetup_K_CLK_negedge_negedge,
	 HoldHigh               => thold_K_CLK_posedge_negedge,
	 HoldLow                => thold_K_CLK_negedge_negedge,
	 CheckEnabled           =>  TO_X01((PRE_ipd)) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/JKF3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay	=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
   CheckEnabled		=>   TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg              => InstancePath & "JKF3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh => tpw_CLK_negedge,
	 PulseWidthLow => tpw_CLK_posedge,
	 CheckEnabled		=> TO_X01((PRE_ipd)) /= '0',
	 HeaderMsg		=> InstancePath & "JKF3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow		=> tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> TRUE, 
	 HeaderMsg		=> InstancePath & "JKF3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

	 Violation := Tviol_J_CLK_negedge or 
	 Tviol_K_CLK_negedge or 
   Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLK;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
   StateTable => JKF3A_Q_tab,
   DataIn => (
CLK_ipd, K_delayed, J_delayed, Q_zd, PRE_ipd, CLK_delayed));
	 Q_zd := Violation XOR Q_zd;
	  --- now combinatorial logic input to the DFF 
	 J_delayed :=  J_ipd ;
          --- now combinatorial logic input to the DFF 
         K_delayed :=  (NOT K_ipd) ;
	 CLK_delayed := CLK_ipd;

	 ----------------------
	 --  Path Delay Section
	 ----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1 => (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_JKF3B_VITAL of JKF3B is
   for VITAL_ACT
   end for;
end CFG_JKF3B_VITAL;



 ---- CELL MAJ3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MAJ3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MAJ3 :  entity is TRUE;
 end MAJ3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of MAJ3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A_ipd  AND  B_ipd ) OR ( B_ipd  AND  C_ipd )) OR ( A_ipd  AND  C_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MAJ3_VITAL of MAJ3 is 
    for VITAL_ACT
    end for;
 end CFG_MAJ3_VITAL;



 ---- CELL MAJ3X ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MAJ3X is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MAJ3X :  entity is TRUE;
 end MAJ3X;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of MAJ3X is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2(( A_ipd  AND  B_ipd ),( (NOT A_ipd)  AND  B_ipd ), (NOT C_ipd) ) OR (( A_ipd  AND  (NOT B_ipd) ) AND  C_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MAJ3X_VITAL of MAJ3X is 
    for VITAL_ACT
    end for;
 end CFG_MAJ3X_VITAL;



 ---- CELL MAJ3XI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MAJ3XI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MAJ3XI :  entity is TRUE;
 end MAJ3XI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of MAJ3XI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  VitalMUX2(( A_ipd  AND  B_ipd ),( (NOT A_ipd)  AND  B_ipd ), (NOT C_ipd) ) OR (( A_ipd  AND  (NOT B_ipd) ) AND  C_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MAJ3XI_VITAL of MAJ3XI is 
    for VITAL_ACT
    end for;
 end CFG_MAJ3XI_VITAL;



 ---- CELL MIN3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MIN3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MIN3 :  entity is TRUE;
 end MIN3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of MIN3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  AND  (NOT B_ipd) ) OR ( (NOT A_ipd)  AND  (NOT C_ipd) )) OR ( (NOT B_ipd)  AND  (NOT C_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MIN3_VITAL of MIN3 is 
    for VITAL_ACT
    end for;
 end CFG_MIN3_VITAL;



 ---- CELL MIN3X ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MIN3X is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MIN3X :  entity is TRUE;
 end MIN3X;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of MIN3X is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2(( A_ipd  AND  (NOT B_ipd) ),( (NOT A_ipd)  AND  (NOT B_ipd) ), (NOT C_ipd) ) OR (( (NOT A_ipd)  AND  B_ipd ) AND  (NOT C_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MIN3X_VITAL of MIN3X is 
    for VITAL_ACT
    end for;
 end CFG_MIN3X_VITAL;



 ---- CELL MIN3XI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MIN3XI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MIN3XI :  entity is TRUE;
 end MIN3XI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of MIN3XI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  VitalMUX2(( A_ipd  AND  (NOT B_ipd) ),( (NOT A_ipd)  AND  (NOT B_ipd) ), (NOT C_ipd) ) OR (( (NOT A_ipd)  AND  B_ipd ) AND  (NOT C_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MIN3XI_VITAL of MIN3XI is 
    for VITAL_ACT
    end for;
 end CFG_MIN3XI_VITAL;



 ---- CELL MULT1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MULT1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_PO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_PO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PI_PO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_PO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PI_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PI		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		PI		: in    STD_ULOGIC;
		FCI		: in    STD_ULOGIC;
		PO		: out    STD_ULOGIC;
		FCO		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MULT1 :  entity is TRUE;
 end MULT1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of MULT1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL PI_ipd  : STD_ULOGIC := 'X';
	SIGNAL FCI_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (PI_ipd, PI, tipd_PI);
	VitalWireDelay (FCI_ipd, FCI, tipd_FCI);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, PI_ipd, FCI_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PO_zd : STD_LOGIC is Results(1);
	ALIAS FCO_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PO_GlitchData  : VitalGlitchDataType;
	VARIABLE FCO_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PO_zd := ((( A_ipd  AND  B_ipd ) XOR  PI_ipd ) XOR  FCI_ipd );
       FCO_zd := (((( A_ipd  AND  B_ipd ) AND  PI_ipd ) OR (( A_ipd  AND  B_ipd ) AND  FCI_ipd )) OR ( PI_ipd  AND  FCI_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PO,
	   GlitchData => PO_GlitchData,
	   OutSignalName => "PO",
	   OutTemp => PO_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PO, true),
	             1 => (B_ipd'last_event,tpd_B_PO, true),
	             2 => (PI_ipd'last_event,tpd_PI_PO, true),
	             3 => (FCI_ipd'last_event,tpd_FCI_PO, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => FCO,
	   GlitchData => FCO_GlitchData,
	   OutSignalName => "FCO",
	   OutTemp => FCO_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_FCO, true),
	             1 => (B_ipd'last_event,tpd_B_FCO, true),
	             2 => (PI_ipd'last_event,tpd_PI_FCO, true),
	             3 => (FCI_ipd'last_event,tpd_FCI_FCO, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MULT1_VITAL of MULT1 is 
    for VITAL_ACT
    end for;
 end CFG_MULT1_VITAL;



 ---- CELL MX2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MX2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MX2 :  entity is TRUE;
 end MX2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of MX2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (S_ipd'last_event,tpd_S_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MX2_VITAL of MX2 is 
    for VITAL_ACT
    end for;
 end CFG_MX2_VITAL;



 ---- CELL MX2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MX2A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MX2A :  entity is TRUE;
 end MX2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of MX2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( (NOT A_ipd) , B_ipd , (NOT S_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (S_ipd'last_event,tpd_S_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MX2A_VITAL of MX2A is 
    for VITAL_ACT
    end for;
 end CFG_MX2A_VITAL;



 ---- CELL MX2B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MX2B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MX2B :  entity is TRUE;
 end MX2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of MX2B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( A_ipd , (NOT B_ipd) , (NOT S_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (S_ipd'last_event,tpd_S_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MX2B_VITAL of MX2B is 
    for VITAL_ACT
    end for;
 end CFG_MX2B_VITAL;



 ---- CELL MX2C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MX2C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MX2C :  entity is TRUE;
 end MX2C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of MX2C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( (NOT A_ipd) , (NOT B_ipd) , (NOT S_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (S_ipd'last_event,tpd_S_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MX2C_VITAL of MX2C is 
    for VITAL_ACT
    end for;
 end CFG_MX2C_VITAL;



 ---- CELL MX4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MX4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S0_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S1_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D2_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D3_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S0		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S1		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D2		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D3		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D0		: in    STD_ULOGIC;
		S0		: in    STD_ULOGIC;
		D1		: in    STD_ULOGIC;
		S1		: in    STD_ULOGIC;
		D2		: in    STD_ULOGIC;
		D3		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MX4 :  entity is TRUE;
 end MX4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of MX4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D0_ipd  : STD_ULOGIC := 'X';
	SIGNAL S0_ipd  : STD_ULOGIC := 'X';
	SIGNAL D1_ipd  : STD_ULOGIC := 'X';
	SIGNAL S1_ipd  : STD_ULOGIC := 'X';
	SIGNAL D2_ipd  : STD_ULOGIC := 'X';
	SIGNAL D3_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D0_ipd, D0, tipd_D0);
	VitalWireDelay (S0_ipd, S0, tipd_S0);
	VitalWireDelay (D1_ipd, D1, tipd_D1);
	VitalWireDelay (S1_ipd, S1, tipd_S1);
	VitalWireDelay (D2_ipd, D2, tipd_D2);
	VitalWireDelay (D3_ipd, D3, tipd_D3);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D0_ipd, S0_ipd, D1_ipd, S1_ipd, D2_ipd, D3_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( VitalMUX2( D0_ipd , D1_ipd , (NOT S0_ipd) ), VitalMUX2( D2_ipd , D3_ipd , (NOT S0_ipd) ), (NOT S1_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D0_ipd'last_event,tpd_D0_Y, true),
	             1 => (S0_ipd'last_event,tpd_S0_Y, true),
	             2 => (D1_ipd'last_event,tpd_D1_Y, true),
	             3 => (S1_ipd'last_event,tpd_S1_Y, true),
	             4 => (D2_ipd'last_event,tpd_D2_Y, true),
	             5 => (D3_ipd'last_event,tpd_D3_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MX4_VITAL of MX4 is 
    for VITAL_ACT
    end for;
 end CFG_MX4_VITAL;



 ---- CELL NAND2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND2 :  entity is TRUE;
 end NAND2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NAND2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  A_ipd  AND  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND2_VITAL of NAND2 is 
    for VITAL_ACT
    end for;
 end CFG_NAND2_VITAL;



 ---- CELL NAND2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND2A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND2A :  entity is TRUE;
 end NAND2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NAND2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  (NOT A_ipd)  AND  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND2A_VITAL of NAND2A is 
    for VITAL_ACT
    end for;
 end CFG_NAND2A_VITAL;



 ---- CELL NAND2B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND2B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND2B :  entity is TRUE;
 end NAND2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NAND2B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  (NOT A_ipd)  AND  (NOT B_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND2B_VITAL of NAND2B is 
    for VITAL_ACT
    end for;
 end CFG_NAND2B_VITAL;



 ---- CELL NAND3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND3 :  entity is TRUE;
 end NAND3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NAND3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( A_ipd  AND  B_ipd ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND3_VITAL of NAND3 is 
    for VITAL_ACT
    end for;
 end CFG_NAND3_VITAL;



 ---- CELL NAND3A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND3A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND3A :  entity is TRUE;
 end NAND3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NAND3A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  AND  B_ipd ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND3A_VITAL of NAND3A is 
    for VITAL_ACT
    end for;
 end CFG_NAND3A_VITAL;



 ---- CELL NAND3B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND3B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND3B :  entity is TRUE;
 end NAND3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NAND3B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND3B_VITAL of NAND3B is 
    for VITAL_ACT
    end for;
 end CFG_NAND3B_VITAL;



 ---- CELL NAND3C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND3C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND3C :  entity is TRUE;
 end NAND3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NAND3C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND3C_VITAL of NAND3C is 
    for VITAL_ACT
    end for;
 end CFG_NAND3C_VITAL;



 ---- CELL NAND4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND4 :  entity is TRUE;
 end NAND4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NAND4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  (NOT C_ipd) ) OR  (NOT D_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND4_VITAL of NAND4 is 
    for VITAL_ACT
    end for;
 end CFG_NAND4_VITAL;



 ---- CELL NAND4A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND4A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND4A :  entity is TRUE;
 end NAND4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NAND4A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( (( (NOT A_ipd)  AND  B_ipd ) AND  C_ipd ) AND  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND4A_VITAL of NAND4A is 
    for VITAL_ACT
    end for;
 end CFG_NAND4A_VITAL;



 ---- CELL NAND4B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND4B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND4B :  entity is TRUE;
 end NAND4B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NAND4B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( (( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  C_ipd ) AND  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND4B_VITAL of NAND4B is 
    for VITAL_ACT
    end for;
 end CFG_NAND4B_VITAL;



 ---- CELL NAND4C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND4C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND4C :  entity is TRUE;
 end NAND4C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NAND4C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( (( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  (NOT C_ipd) ) AND  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND4C_VITAL of NAND4C is 
    for VITAL_ACT
    end for;
 end CFG_NAND4C_VITAL;



 ---- CELL NAND4D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND4D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND4D :  entity is TRUE;
 end NAND4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NAND4D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( (( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  (NOT C_ipd) ) AND  (NOT D_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND4D_VITAL of NAND4D is 
    for VITAL_ACT
    end for;
 end CFG_NAND4D_VITAL;



 ---- CELL NAND5B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND5B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND5B :  entity is TRUE;
 end NAND5B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NAND5B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ((( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  C_ipd ) AND  D_ipd ) AND  E_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true),
	             4 => (E_ipd'last_event,tpd_E_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND5B_VITAL of NAND5B is 
    for VITAL_ACT
    end for;
 end CFG_NAND5B_VITAL;



 ---- CELL NAND5C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND5C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND5C :  entity is TRUE;
 end NAND5C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NAND5C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ((( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  (NOT C_ipd) ) AND  D_ipd ) AND  E_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true),
	             4 => (E_ipd'last_event,tpd_E_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND5C_VITAL of NAND5C is 
    for VITAL_ACT
    end for;
 end CFG_NAND5C_VITAL;



 ---- CELL NOR2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR2 :  entity is TRUE;
 end NOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NOR2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  A_ipd  OR  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR2_VITAL of NOR2 is 
    for VITAL_ACT
    end for;
 end CFG_NOR2_VITAL;



 ---- CELL NOR2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR2A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR2A :  entity is TRUE;
 end NOR2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NOR2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  (NOT A_ipd)  OR  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR2A_VITAL of NOR2A is 
    for VITAL_ACT
    end for;
 end CFG_NOR2A_VITAL;



 ---- CELL NOR2B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR2B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR2B :  entity is TRUE;
 end NOR2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NOR2B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  (NOT A_ipd)  OR  (NOT B_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR2B_VITAL of NOR2B is 
    for VITAL_ACT
    end for;
 end CFG_NOR2B_VITAL;



 ---- CELL NOR3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR3 :  entity is TRUE;
 end NOR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NOR3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( A_ipd  OR  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR3_VITAL of NOR3 is 
    for VITAL_ACT
    end for;
 end CFG_NOR3_VITAL;



 ---- CELL NOR3A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR3A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR3A :  entity is TRUE;
 end NOR3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NOR3A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  OR  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR3A_VITAL of NOR3A is 
    for VITAL_ACT
    end for;
 end CFG_NOR3A_VITAL;



 ---- CELL NOR3B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR3B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR3B :  entity is TRUE;
 end NOR3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NOR3B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR3B_VITAL of NOR3B is 
    for VITAL_ACT
    end for;
 end CFG_NOR3B_VITAL;



 ---- CELL NOR3C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR3C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR3C :  entity is TRUE;
 end NOR3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NOR3C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR3C_VITAL of NOR3C is 
    for VITAL_ACT
    end for;
 end CFG_NOR3C_VITAL;



 ---- CELL NOR4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR4 :  entity is TRUE;
 end NOR4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NOR4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  (NOT C_ipd) ) AND  (NOT D_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR4_VITAL of NOR4 is 
    for VITAL_ACT
    end for;
 end CFG_NOR4_VITAL;



 ---- CELL NOR4A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR4A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR4A :  entity is TRUE;
 end NOR4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NOR4A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( (( (NOT A_ipd)  OR  B_ipd ) OR  C_ipd ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR4A_VITAL of NOR4A is 
    for VITAL_ACT
    end for;
 end CFG_NOR4A_VITAL;



 ---- CELL NOR4B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR4B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR4B :  entity is TRUE;
 end NOR4B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NOR4B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( (( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  C_ipd ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR4B_VITAL of NOR4B is 
    for VITAL_ACT
    end for;
 end CFG_NOR4B_VITAL;



 ---- CELL NOR4C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR4C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR4C :  entity is TRUE;
 end NOR4C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NOR4C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( (( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  (NOT C_ipd) ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR4C_VITAL of NOR4C is 
    for VITAL_ACT
    end for;
 end CFG_NOR4C_VITAL;



 ---- CELL NOR4D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR4D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR4D :  entity is TRUE;
 end NOR4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NOR4D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( (( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  (NOT C_ipd) ) OR  (NOT D_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR4D_VITAL of NOR4D is 
    for VITAL_ACT
    end for;
 end CFG_NOR4D_VITAL;



 ---- CELL NOR5B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR5B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR5B :  entity is TRUE;
 end NOR5B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NOR5B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ((( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  C_ipd ) OR  D_ipd ) OR  E_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true),
	             4 => (E_ipd'last_event,tpd_E_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR5B_VITAL of NOR5B is 
    for VITAL_ACT
    end for;
 end CFG_NOR5B_VITAL;



 ---- CELL NOR5C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR5C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR5C :  entity is TRUE;
 end NOR5C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of NOR5C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ((( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  (NOT C_ipd) ) OR  D_ipd ) OR  E_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true),
	             4 => (E_ipd'last_event,tpd_E_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR5C_VITAL of NOR5C is 
    for VITAL_ACT
    end for;
 end CFG_NOR5C_VITAL;



 ---- CELL OA1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA1 :  entity is TRUE;
 end OA1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OA1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  OR  B_ipd ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA1_VITAL of OA1 is 
    for VITAL_ACT
    end for;
 end CFG_OA1_VITAL;



 ---- CELL OA1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA1A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA1A :  entity is TRUE;
 end OA1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OA1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  OR  B_ipd ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA1A_VITAL of OA1A is 
    for VITAL_ACT
    end for;
 end CFG_OA1A_VITAL;



 ---- CELL OA1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA1B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		C		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA1B :  entity is TRUE;
 end OA1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OA1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (C_ipd, A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( (NOT C_ipd)  AND ( A_ipd  OR  B_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (C_ipd'last_event,tpd_C_Y, true),
	             1 => (A_ipd'last_event,tpd_A_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA1B_VITAL of OA1B is 
    for VITAL_ACT
    end for;
 end CFG_OA1B_VITAL;



 ---- CELL OA1C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA1C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		C		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA1C :  entity is TRUE;
 end OA1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OA1C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (C_ipd, A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( (NOT C_ipd)  AND ( (NOT A_ipd)  OR  B_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (C_ipd'last_event,tpd_C_Y, true),
	             1 => (A_ipd'last_event,tpd_A_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA1C_VITAL of OA1C is 
    for VITAL_ACT
    end for;
 end CFG_OA1C_VITAL;



 ---- CELL OA2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA2 :  entity is TRUE;
 end OA2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OA2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  OR  B_ipd ) AND ( C_ipd  OR  D_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA2_VITAL of OA2 is 
    for VITAL_ACT
    end for;
 end CFG_OA2_VITAL;



 ---- CELL OA2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA2A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA2A :  entity is TRUE;
 end OA2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OA2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  OR  B_ipd ) AND ( C_ipd  OR  D_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA2A_VITAL of OA2A is 
    for VITAL_ACT
    end for;
 end CFG_OA2A_VITAL;



 ---- CELL OA3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA3 :  entity is TRUE;
 end OA3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OA3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A_ipd  OR  B_ipd ) AND  C_ipd ) AND  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA3_VITAL of OA3 is 
    for VITAL_ACT
    end for;
 end CFG_OA3_VITAL;



 ---- CELL OA3A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA3A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA3A :  entity is TRUE;
 end OA3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OA3A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A_ipd  OR  B_ipd ) AND  (NOT C_ipd) ) AND  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA3A_VITAL of OA3A is 
    for VITAL_ACT
    end for;
 end CFG_OA3A_VITAL;



 ---- CELL OA3B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA3B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA3B :  entity is TRUE;
 end OA3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OA3B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  OR  B_ipd ) AND  (NOT C_ipd) ) AND  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA3B_VITAL of OA3B is 
    for VITAL_ACT
    end for;
 end CFG_OA3B_VITAL;



 ---- CELL OA4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA4 :  entity is TRUE;
 end OA4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OA4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A_ipd  OR  B_ipd ) OR  C_ipd ) AND  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA4_VITAL of OA4 is 
    for VITAL_ACT
    end for;
 end CFG_OA4_VITAL;



 ---- CELL OA4A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA4A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA4A :  entity is TRUE;
 end OA4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OA4A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A_ipd  OR  B_ipd ) OR  (NOT C_ipd) ) AND  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA4A_VITAL of OA4A is 
    for VITAL_ACT
    end for;
 end CFG_OA4A_VITAL;



 ---- CELL OA5 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA5 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA5 :  entity is TRUE;
 end OA5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OA5 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A_ipd  OR  B_ipd ) OR  C_ipd ) AND ( A_ipd  OR  D_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA5_VITAL of OA5 is 
    for VITAL_ACT
    end for;
 end CFG_OA5_VITAL;



 ---- CELL OAI1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OAI1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OAI1 :  entity is TRUE;
 end OAI1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OAI1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( A_ipd  OR  B_ipd ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OAI1_VITAL of OAI1 is 
    for VITAL_ACT
    end for;
 end CFG_OAI1_VITAL;



 ---- CELL OAI2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OAI2A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OAI2A :  entity is TRUE;
 end OAI2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OAI2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( (( A_ipd  OR  B_ipd ) OR  C_ipd ) AND  (NOT D_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OAI2A_VITAL of OAI2A is 
    for VITAL_ACT
    end for;
 end CFG_OAI2A_VITAL;



 ---- CELL OAI3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OAI3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OAI3 :  entity is TRUE;
 end OAI3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OAI3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( (( A_ipd  OR  B_ipd ) AND  C_ipd ) AND  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OAI3_VITAL of OAI3 is 
    for VITAL_ACT
    end for;
 end CFG_OAI3_VITAL;



 ---- CELL OAI3A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OAI3A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OAI3A :  entity is TRUE;
 end OAI3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OAI3A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( (( A_ipd  OR  B_ipd ) AND  (NOT C_ipd) ) AND  (NOT D_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OAI3A_VITAL of OAI3A is 
    for VITAL_ACT
    end for;
 end CFG_OAI3A_VITAL;



 ---- CELL OR2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR2 :  entity is TRUE;
 end OR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OR2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( A_ipd  OR  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR2_VITAL of OR2 is 
    for VITAL_ACT
    end for;
 end CFG_OR2_VITAL;



 ---- CELL OR2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR2A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR2A :  entity is TRUE;
 end OR2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OR2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( (NOT A_ipd)  OR  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR2A_VITAL of OR2A is 
    for VITAL_ACT
    end for;
 end CFG_OR2A_VITAL;



 ---- CELL OR2B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR2B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR2B :  entity is TRUE;
 end OR2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OR2B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( (NOT A_ipd)  OR  (NOT B_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR2B_VITAL of OR2B is 
    for VITAL_ACT
    end for;
 end CFG_OR2B_VITAL;



 ---- CELL OR3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR3 :  entity is TRUE;
 end OR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OR3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  OR  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR3_VITAL of OR3 is 
    for VITAL_ACT
    end for;
 end CFG_OR3_VITAL;



 ---- CELL OR3A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR3A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR3A :  entity is TRUE;
 end OR3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OR3A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  OR  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR3A_VITAL of OR3A is 
    for VITAL_ACT
    end for;
 end CFG_OR3A_VITAL;



 ---- CELL OR3B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR3B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR3B :  entity is TRUE;
 end OR3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OR3B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR3B_VITAL of OR3B is 
    for VITAL_ACT
    end for;
 end CFG_OR3B_VITAL;



 ---- CELL OR3C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR3C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR3C :  entity is TRUE;
 end OR3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OR3C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR3C_VITAL of OR3C is 
    for VITAL_ACT
    end for;
 end CFG_OR3C_VITAL;



 ---- CELL OR4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR4 :  entity is TRUE;
 end OR4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OR4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A_ipd  OR  B_ipd ) OR  C_ipd ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR4_VITAL of OR4 is 
    for VITAL_ACT
    end for;
 end CFG_OR4_VITAL;



 ---- CELL OR4A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR4A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR4A :  entity is TRUE;
 end OR4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OR4A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  OR  B_ipd ) OR  C_ipd ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR4A_VITAL of OR4A is 
    for VITAL_ACT
    end for;
 end CFG_OR4A_VITAL;



 ---- CELL OR4B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR4B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR4B :  entity is TRUE;
 end OR4B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OR4B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  C_ipd ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR4B_VITAL of OR4B is 
    for VITAL_ACT
    end for;
 end CFG_OR4B_VITAL;



 ---- CELL OR4C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR4C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR4C :  entity is TRUE;
 end OR4C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OR4C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  (NOT C_ipd) ) OR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR4C_VITAL of OR4C is 
    for VITAL_ACT
    end for;
 end CFG_OR4C_VITAL;



 ---- CELL OR4D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR4D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR4D :  entity is TRUE;
 end OR4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OR4D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  (NOT C_ipd) ) OR  (NOT D_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR4D_VITAL of OR4D is 
    for VITAL_ACT
    end for;
 end CFG_OR4D_VITAL;



 ---- CELL OR5A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR5A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR5A :  entity is TRUE;
 end OR5A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OR5A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (((( (NOT A_ipd)  OR  B_ipd ) OR  C_ipd ) OR  D_ipd ) OR  E_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true),
	             4 => (E_ipd'last_event,tpd_E_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR5A_VITAL of OR5A is 
    for VITAL_ACT
    end for;
 end CFG_OR5A_VITAL;



 ---- CELL OR5B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR5B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR5B :  entity is TRUE;
 end OR5B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OR5B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (((( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  C_ipd ) OR  D_ipd ) OR  E_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true),
	             4 => (E_ipd'last_event,tpd_E_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR5B_VITAL of OR5B is 
    for VITAL_ACT
    end for;
 end CFG_OR5B_VITAL;



 ---- CELL OR5C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR5C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR5C :  entity is TRUE;
 end OR5C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OR5C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (((( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  (NOT C_ipd) ) OR  D_ipd ) OR  E_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true),
	             4 => (E_ipd'last_event,tpd_E_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR5C_VITAL of OR5C is 
    for VITAL_ACT
    end for;
 end CFG_OR5C_VITAL;



 ---- CELL OUTBUF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF :  entity is TRUE;
 end OUTBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_VITAL of OUTBUF is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_VITAL;



 ---- CELL OUTBUF_S_8 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_S_8 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_S_8 :  entity is TRUE;
 end OUTBUF_S_8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_S_8 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_S_8_VITAL of OUTBUF_S_8 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_S_8_VITAL;



 ---- CELL OUTBUF_S_12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_S_12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_S_12 :  entity is TRUE;
 end OUTBUF_S_12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_S_12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_S_12_VITAL of OUTBUF_S_12 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_S_12_VITAL;



 ---- CELL OUTBUF_S_16 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_S_16 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_S_16 :  entity is TRUE;
 end OUTBUF_S_16;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_S_16 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_S_16_VITAL of OUTBUF_S_16 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_S_16_VITAL;



 ---- CELL OUTBUF_S_24 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_S_24 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_S_24 :  entity is TRUE;
 end OUTBUF_S_24;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_S_24 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_S_24_VITAL of OUTBUF_S_24 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_S_24_VITAL;



 ---- CELL OUTBUF_F_8 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_F_8 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_F_8 :  entity is TRUE;
 end OUTBUF_F_8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_F_8 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_F_8_VITAL of OUTBUF_F_8 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_F_8_VITAL;



 ---- CELL OUTBUF_F_12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_F_12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_F_12 :  entity is TRUE;
 end OUTBUF_F_12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_F_12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_F_12_VITAL of OUTBUF_F_12 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_F_12_VITAL;



 ---- CELL OUTBUF_F_16 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_F_16 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_F_16 :  entity is TRUE;
 end OUTBUF_F_16;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_F_16 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_F_16_VITAL of OUTBUF_F_16 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_F_16_VITAL;



 ---- CELL OUTBUF_F_24 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_F_24 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_F_24 :  entity is TRUE;
 end OUTBUF_F_24;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_F_24 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_F_24_VITAL of OUTBUF_F_24 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_F_24_VITAL;



 ---- CELL OUTBUF_LVCMOS25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_LVCMOS25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_LVCMOS25 :  entity is TRUE;
 end OUTBUF_LVCMOS25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_LVCMOS25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_LVCMOS25_VITAL of OUTBUF_LVCMOS25 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_LVCMOS25_VITAL;



 ---- CELL OUTBUF_LVCMOS18 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_LVCMOS18 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_LVCMOS18 :  entity is TRUE;
 end OUTBUF_LVCMOS18;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_LVCMOS18 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_LVCMOS18_VITAL of OUTBUF_LVCMOS18 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_LVCMOS18_VITAL;



 ---- CELL OUTBUF_LVCMOS15 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_LVCMOS15 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_LVCMOS15 :  entity is TRUE;
 end OUTBUF_LVCMOS15;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_LVCMOS15 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_LVCMOS15_VITAL of OUTBUF_LVCMOS15 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_LVCMOS15_VITAL;



 ---- CELL OUTBUF_PCI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_PCI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_PCI :  entity is TRUE;
 end OUTBUF_PCI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_PCI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_PCI_VITAL of OUTBUF_PCI is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_PCI_VITAL;



 ---- CELL OUTBUF_PCIX ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_PCIX is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_PCIX :  entity is TRUE;
 end OUTBUF_PCIX;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_PCIX is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_PCIX_VITAL of OUTBUF_PCIX is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_PCIX_VITAL;



 ---- CELL OUTBUF_GTLP33 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_GTLP33 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_GTLP33 :  entity is TRUE;
 end OUTBUF_GTLP33;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_GTLP33 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_GTLP33_VITAL of OUTBUF_GTLP33 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_GTLP33_VITAL;



 ---- CELL OUTBUF_GTLP25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_GTLP25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_GTLP25 :  entity is TRUE;
 end OUTBUF_GTLP25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_GTLP25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_GTLP25_VITAL of OUTBUF_GTLP25 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_GTLP25_VITAL;



 ---- CELL OUTBUF_HSTL_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_HSTL_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_HSTL_I :  entity is TRUE;
 end OUTBUF_HSTL_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_HSTL_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_HSTL_I_VITAL of OUTBUF_HSTL_I is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_HSTL_I_VITAL;



 ---- CELL OUTBUF_SSTL3_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_SSTL3_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_SSTL3_I :  entity is TRUE;
 end OUTBUF_SSTL3_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_SSTL3_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_SSTL3_I_VITAL of OUTBUF_SSTL3_I is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_SSTL3_I_VITAL;



 ---- CELL OUTBUF_SSTL3_II ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_SSTL3_II is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_SSTL3_II :  entity is TRUE;
 end OUTBUF_SSTL3_II;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_SSTL3_II is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_SSTL3_II_VITAL of OUTBUF_SSTL3_II is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_SSTL3_II_VITAL;



 ---- CELL OUTBUF_SSTL2_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_SSTL2_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_SSTL2_I :  entity is TRUE;
 end OUTBUF_SSTL2_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_SSTL2_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_SSTL2_I_VITAL of OUTBUF_SSTL2_I is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_SSTL2_I_VITAL;



 ---- CELL OUTBUF_SSTL2_II ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_SSTL2_II is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_SSTL2_II :  entity is TRUE;
 end OUTBUF_SSTL2_II;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of OUTBUF_SSTL2_II is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_SSTL2_II_VITAL of OUTBUF_SSTL2_II is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_SSTL2_II_VITAL;



 ---- CELL PLLHCLK ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity PLLHCLK is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of PLLHCLK :  entity is TRUE;
 end PLLHCLK;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of PLLHCLK is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_PLLHCLK_VITAL of PLLHCLK is 
    for VITAL_ACT
    end for;
 end CFG_PLLHCLK_VITAL;



 ---- CELL PLLRCLK ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity PLLRCLK is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of PLLRCLK :  entity is TRUE;
 end PLLRCLK;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of PLLRCLK is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_PLLRCLK_VITAL of PLLRCLK is 
    for VITAL_ACT
    end for;
 end CFG_PLLRCLK_VITAL;



 ---- CELL SFCNTECP1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity SFCNTECP1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_UD_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_Q_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_UD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		Q		:  out STD_ULOGIC;
		UD		:  in    STD_ULOGIC;
		FCI		:  in    STD_ULOGIC;
		FCO		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of SFCNTECP1 :  entity is TRUE;
 end SFCNTECP1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of SFCNTECP1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL UD_ipd  : STD_ULOGIC := 'X';
	SIGNAL FCI_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (UD_ipd, UD, tipd_UD);
	  VitalWireDelay (FCI_ipd, FCI, tipd_FCI);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (UD_ipd, FCI_ipd, PRE_ipd,CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_UD_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_UD_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_FCI_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_FCI_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_1	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);
	ALIAS FCO_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;
	VARIABLE FCO_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_UD_CLK_negedge, 
	 TimingData		=> Tmkr_UD_CLK_negedge, 
	 TestSignal		=> UD_ipd,
	 TestSignalName		=> "UD",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_UD_CLK_posedge_negedge,
	 SetupLow		=> tsetup_UD_CLK_negedge_negedge,
	 HoldHigh		=> thold_UD_CLK_posedge_negedge,
	 HoldLow		=> thold_UD_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/SFCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_FCI_CLK_negedge, 
	 TimingData		=> Tmkr_FCI_CLK_negedge, 
	 TestSignal		=> FCI_ipd,
	 TestSignalName		=> "FCI",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_FCI_CLK_posedge_negedge,
	 SetupLow		=> tsetup_FCI_CLK_negedge_negedge,
	 HoldHigh		=> thold_FCI_CLK_posedge_negedge,
	 HoldLow		=> thold_FCI_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/SFCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (CLR_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "SFCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "SFCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "SFCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "SFCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "SFCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "SFCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_UD_CLK_negedge or 
	 Tviol_FCI_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, Q_zd, NET_0_1, E_delayed, PRE_ipd, CLK_delayed));
   Q_zd := Violation XOR Q_zd;
    --- combinatorial output logic. 
   FCO_zd := ((( Q_zd  AND  (NOT UD_ipd) ) OR ( Q_zd  AND  FCI_ipd )) OR ( (NOT UD_ipd)  AND  FCI_ipd ));
         --- now combinatorial logic input to the DFF 
   NET_0_1 := (( Q_zd  XOR  (NOT UD_ipd) ) XOR  FCI_ipd );
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => FCO,
	 GlitchData => FCO_GlitchData,
	 OutSignalName => "FCO",
	 OutTemp => FCO_zd,
	 Paths => (
	         0 => (UD_ipd'last_event, tpd_UD_FCO, true),
	         1 => (FCI_ipd'last_event, tpd_FCI_FCO, true),
		 2 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		 3 => (CLR_ipd'last_event, tpd_CLR_Q, true),
	           4 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_SFCNTECP1_VITAL of SFCNTECP1 is
   for VITAL_ACT
   end for;
end CFG_SFCNTECP1_VITAL;



 ---- CELL SRCNTECP1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity SRCNTECP1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_UD_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_Q_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_UD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		Q		:  out STD_ULOGIC;
		UD		:  in    STD_ULOGIC;
		FCI		:  in    STD_ULOGIC;
		FCO		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of SRCNTECP1 :  entity is TRUE;
 end SRCNTECP1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of SRCNTECP1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL UD_ipd  : STD_ULOGIC := 'X';
	SIGNAL FCI_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (UD_ipd, UD, tipd_UD);
	  VitalWireDelay (FCI_ipd, FCI, tipd_FCI);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (UD_ipd, FCI_ipd, PRE_ipd,CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_UD_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_UD_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_FCI_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_FCI_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_1	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);
	ALIAS FCO_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;
	VARIABLE FCO_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_UD_CLK_posedge,
	 TimingData		=> Tmkr_UD_CLK_posedge,
	 TestSignal		=> UD_ipd,
	 TestSignalName		=> "UD",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_UD_CLK_posedge_posedge,
	 SetupLow		=> tsetup_UD_CLK_negedge_posedge,
	 HoldHigh		=> thold_UD_CLK_posedge_posedge,
	 HoldLow		=> thold_UD_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/SRCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_FCI_CLK_posedge,
	 TimingData		=> Tmkr_FCI_CLK_posedge,
	 TestSignal		=> FCI_ipd,
	 TestSignalName		=> "FCI",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_FCI_CLK_posedge_posedge,
	 SetupLow		=> tsetup_FCI_CLK_negedge_posedge,
	 HoldHigh		=> thold_FCI_CLK_posedge_posedge,
	 HoldLow		=> thold_FCI_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/SRCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "SRCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "SRCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "SRCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "SRCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "SRCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "SRCNTECP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_UD_CLK_posedge or 
	 Tviol_FCI_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, NET_0_1, E_delayed, PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;
    --- combinatorial output logic. 
   FCO_zd := ((( Q_zd  AND  (NOT UD_ipd) ) OR ( Q_zd  AND  FCI_ipd )) OR ( (NOT UD_ipd)  AND  FCI_ipd ));
         --- now combinatorial logic input to the DFF 
   NET_0_1 := (( Q_zd  XOR  (NOT UD_ipd) ) XOR  FCI_ipd );
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => FCO,
	 GlitchData => FCO_GlitchData,
	 OutSignalName => "FCO",
	 OutTemp => FCO_zd,
	 Paths => (
	         0 => (UD_ipd'last_event, tpd_UD_FCO, true),
	         1 => (FCI_ipd'last_event, tpd_FCI_FCO, true),
		 2 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		 3 => (CLR_ipd'last_event, tpd_CLR_Q, true),
	           4 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_SRCNTECP1_VITAL of SRCNTECP1 is
   for VITAL_ACT
   end for;
end CFG_SRCNTECP1_VITAL;



 ---- CELL SFCNTELDCP1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity SFCNTELDCP1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_UD_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_Q_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_LD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_LD_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_LD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_LD_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_UD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_LD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		Q		:  out STD_ULOGIC;
		UD		:  in    STD_ULOGIC;
		FCI		:  in    STD_ULOGIC;
		LD		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		FCO		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of SFCNTELDCP1 :  entity is TRUE;
 end SFCNTELDCP1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of SFCNTELDCP1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL UD_ipd  : STD_ULOGIC := 'X';
	SIGNAL FCI_ipd  : STD_ULOGIC := 'X';
	SIGNAL LD_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (UD_ipd, UD, tipd_UD);
	  VitalWireDelay (FCI_ipd, FCI, tipd_FCI);
	  VitalWireDelay (LD_ipd, LD, tipd_LD);
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (UD_ipd, FCI_ipd, LD_ipd, D_ipd, PRE_ipd,CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_UD_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_UD_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_FCI_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_FCI_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_LD_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_LD_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_4	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);
	ALIAS FCO_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;
	VARIABLE FCO_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_UD_CLK_negedge, 
	 TimingData		=> Tmkr_UD_CLK_negedge, 
	 TestSignal		=> UD_ipd,
	 TestSignalName		=> "UD",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_UD_CLK_posedge_negedge,
	 SetupLow		=> tsetup_UD_CLK_negedge_negedge,
	 HoldHigh		=> thold_UD_CLK_posedge_negedge,
	 HoldLow		=> thold_UD_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/SFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_FCI_CLK_negedge, 
	 TimingData		=> Tmkr_FCI_CLK_negedge, 
	 TestSignal		=> FCI_ipd,
	 TestSignalName		=> "FCI",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_FCI_CLK_posedge_negedge,
	 SetupLow		=> tsetup_FCI_CLK_negedge_negedge,
	 HoldHigh		=> thold_FCI_CLK_posedge_negedge,
	 HoldLow		=> thold_FCI_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/SFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_LD_CLK_negedge, 
	 TimingData		=> Tmkr_LD_CLK_negedge, 
	 TestSignal		=> LD_ipd,
	 TestSignalName		=> "LD",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_LD_CLK_posedge_negedge,
	 SetupLow		=> tsetup_LD_CLK_negedge_negedge,
	 HoldHigh		=> thold_LD_CLK_posedge_negedge,
	 HoldLow		=> thold_LD_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/SFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/SFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (CLR_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "SFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "SFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "SFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "SFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "SFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "SFCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_UD_CLK_negedge or 
	 Tviol_FCI_CLK_negedge or 
	 Tviol_LD_CLK_negedge or Tviol_D_CLK_negedge or Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, Q_zd, NET_0_4, E_delayed, PRE_ipd, CLK_delayed));
   Q_zd := Violation XOR Q_zd;
    --- combinatorial output logic. 
   FCO_zd := ((( Q_zd  AND  (NOT UD_ipd) ) OR ( Q_zd  AND  FCI_ipd )) OR ( (NOT UD_ipd)  AND  FCI_ipd ));
         --- now combinatorial logic input to the DFF 
   NET_0_4 :=  VitalMUX2((( Q_zd  XOR  (NOT UD_ipd) ) XOR  FCI_ipd ), D_ipd , (NOT LD_ipd) );
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => FCO,
	 GlitchData => FCO_GlitchData,
	 OutSignalName => "FCO",
	 OutTemp => FCO_zd,
	 Paths => (
	         0 => (UD_ipd'last_event, tpd_UD_FCO, true),
	         1 => (FCI_ipd'last_event, tpd_FCI_FCO, true),
		 2 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		 3 => (CLR_ipd'last_event, tpd_CLR_Q, true),
	           4 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_SFCNTELDCP1_VITAL of SFCNTELDCP1 is
   for VITAL_ACT
   end for;
end CFG_SFCNTELDCP1_VITAL;



 ---- CELL SRCNTELDCP1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity SRCNTELDCP1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_UD_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_Q_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_LD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_LD_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_Q_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_Q_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_UD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_UD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_FCI_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_FCI_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_LD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_LD_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_UD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_LD		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		Q		:  out STD_ULOGIC;
		UD		:  in    STD_ULOGIC;
		FCI		:  in    STD_ULOGIC;
		LD		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		FCO		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of SRCNTELDCP1 :  entity is TRUE;
 end SRCNTELDCP1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of SRCNTELDCP1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL UD_ipd  : STD_ULOGIC := 'X';
	SIGNAL FCI_ipd  : STD_ULOGIC := 'X';
	SIGNAL LD_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (UD_ipd, UD, tipd_UD);
	  VitalWireDelay (FCI_ipd, FCI, tipd_FCI);
	  VitalWireDelay (LD_ipd, LD, tipd_LD);
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (UD_ipd, FCI_ipd, LD_ipd, D_ipd, PRE_ipd,CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_UD_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_UD_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_FCI_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_FCI_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_LD_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_LD_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_4	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);
	ALIAS FCO_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;
	VARIABLE FCO_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_UD_CLK_posedge,
	 TimingData		=> Tmkr_UD_CLK_posedge,
	 TestSignal		=> UD_ipd,
	 TestSignalName		=> "UD",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_UD_CLK_posedge_posedge,
	 SetupLow		=> tsetup_UD_CLK_negedge_posedge,
	 HoldHigh		=> thold_UD_CLK_posedge_posedge,
	 HoldLow		=> thold_UD_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/SRCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_FCI_CLK_posedge,
	 TimingData		=> Tmkr_FCI_CLK_posedge,
	 TestSignal		=> FCI_ipd,
	 TestSignalName		=> "FCI",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_FCI_CLK_posedge_posedge,
	 SetupLow		=> tsetup_FCI_CLK_negedge_posedge,
	 HoldHigh		=> thold_FCI_CLK_posedge_posedge,
	 HoldLow		=> thold_FCI_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/SRCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_LD_CLK_posedge,
	 TimingData		=> Tmkr_LD_CLK_posedge,
	 TestSignal		=> LD_ipd,
	 TestSignalName		=> "LD",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_LD_CLK_posedge_posedge,
	 SetupLow		=> tsetup_LD_CLK_negedge_posedge,
	 HoldHigh		=> thold_LD_CLK_posedge_posedge,
	 HoldLow		=> thold_LD_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/SRCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/SRCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "SRCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "SRCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "SRCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "SRCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "SRCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "SRCNTELDCP1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_UD_CLK_posedge or 
	 Tviol_FCI_CLK_posedge or 
	 Tviol_LD_CLK_posedge or Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, NET_0_4, E_delayed, PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;
    --- combinatorial output logic. 
   FCO_zd := ((( Q_zd  AND  (NOT UD_ipd) ) OR ( Q_zd  AND  FCI_ipd )) OR ( (NOT UD_ipd)  AND  FCI_ipd ));
         --- now combinatorial logic input to the DFF 
   NET_0_4 :=  VitalMUX2((( Q_zd  XOR  (NOT UD_ipd) ) XOR  FCI_ipd ), D_ipd , (NOT LD_ipd) );
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => FCO,
	 GlitchData => FCO_GlitchData,
	 OutSignalName => "FCO",
	 OutTemp => FCO_zd,
	 Paths => (
	         0 => (UD_ipd'last_event, tpd_UD_FCO, true),
	         1 => (FCI_ipd'last_event, tpd_FCI_FCO, true),
		 2 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		 3 => (CLR_ipd'last_event, tpd_CLR_Q, true),
	           4 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_SRCNTELDCP1_VITAL of SRCNTELDCP1 is
   for VITAL_ACT
   end for;
end CFG_SRCNTELDCP1_VITAL;



 ---- CELL SUB1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity SUB1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_S		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_FCO		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		FCI		: in    STD_ULOGIC;
		S		: out    STD_ULOGIC;
		FCO		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of SUB1 :  entity is TRUE;
 end SUB1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of SUB1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL FCI_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (FCI_ipd, FCI, tipd_FCI);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, FCI_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS S_zd : STD_LOGIC is Results(1);
	ALIAS FCO_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE S_GlitchData  : VitalGlitchDataType;
	VARIABLE FCO_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       S_zd := ( VitalMUX2( (NOT B_ipd) , B_ipd , (NOT A_ipd) ) XOR  FCI_ipd );
       FCO_zd := ((( A_ipd  AND  (NOT B_ipd) ) OR ( A_ipd  AND  FCI_ipd )) OR ( (NOT B_ipd)  AND  FCI_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => S,
	   GlitchData => S_GlitchData,
	   OutSignalName => "S",
	   OutTemp => S_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_S, true),
	             1 => (B_ipd'last_event,tpd_B_S, true),
	             2 => (FCI_ipd'last_event,tpd_FCI_S, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => FCO,
	   GlitchData => FCO_GlitchData,
	   OutSignalName => "FCO",
	   OutTemp => FCO_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_FCO, true),
	             1 => (B_ipd'last_event,tpd_B_FCO, true),
	             2 => (FCI_ipd'last_event,tpd_FCI_FCO, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_SUB1_VITAL of SUB1 is 
    for VITAL_ACT
    end for;
 end CFG_SUB1_VITAL;



 ---- CELL TF1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TF1A is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_T_CLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_T_CLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_T_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_T_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge	:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge	:  VitalDelayType := 0.000 ns;
		tipd_CLK	:  VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR	:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_T	:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		T	:  in    STD_ULOGIC;
		CLR	:  in    STD_ULOGIC;
	        CLK	:  in    STD_ULOGIC;
		Q	:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of TF1A :  entity is TRUE;
 end TF1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TF1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL T_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (T_ipd, T, tipd_T);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (T_ipd, CLR_ipd,CLK_ipd)

   -- timing check results
	VARIABLE Tviol_T_CLK_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_T_CLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK  : STD_ULOGIC := '0';
	VARIABLE PInfo_CLK  : VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
	VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation      : STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 4);
	VARIABLE CLK_delayed        : STD_ULOGIC := 'X';
	VARIABLE T_delayed        : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_T_CLK_posedge,
	 TimingData		=> Tmkr_T_CLK_posedge,
	 TestSignal		=> T_ipd,
	 TestSignalName		=> "T",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_T_CLK_posedge_posedge,
	 SetupLow		=> tsetup_T_CLK_negedge_posedge,
	 HoldHigh		=> thold_T_CLK_posedge_posedge,
	 HoldLow		=> thold_T_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/TF1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_CLK_posedge,
	 TimingData		=> Tmkr_CLR_CLK_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_CLK_posedge_posedge,
 	 Removal                => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	  CheckEnabled		=>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "TF1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled           => TO_X01(( NOT CLR_ipd)) /= '1',
	 HeaderMsg		=> InstancePath & "TF1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled	 => TRUE,
	 HeaderMsg		=> InstancePath & "TF1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

	Violation := Tviol_T_CLK_posedge or 
		      Pviol_CLR or 
		      Pviol_CLK;

	VitalStateTable(
	 Result => Q_zd,
	PreviousDataIn => PrevData_Q,
	StateTable => tflipflop_Q_tab,
	DataIn => (
             CLR_ipd, CLK_delayed, T_delayed, Q_zd, CLK_ipd));
	Q_zd := Violation XOR Q_zd;
	--- now combinatorial logic input to the DFF 
	T_delayed :=  T_ipd ;
	CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	          1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_TF1A_VITAL of TF1A is
   for VITAL_ACT
   end for;
end CFG_TF1A_VITAL;



 ---- CELL TF1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TF1B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_T_CLK_negedge_negedge	:   VitalDelayType := 0.000 ns;
		thold_T_CLK_negedge_negedge	:   VitalDelayType := 0.000 ns;
		tsetup_T_CLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
		thold_T_CLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge	:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge	:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge	:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge	:  VitalDelayType := 0.000 ns;
		tipd_CLK	:  VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR	:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_T	:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		T	:  in    STD_ULOGIC;
		CLR	:  in    STD_ULOGIC;
	        CLK	:  in    STD_ULOGIC;
		Q	:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of TF1B :  entity is TRUE;
 end TF1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TF1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL T_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (T_ipd, T, tipd_T);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (T_ipd, CLR_ipd,CLK_ipd)

   -- timing check results
	VARIABLE Tviol_T_CLK_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_T_CLK_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK  : STD_ULOGIC := '0';
	VARIABLE PInfo_CLK  : VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
	VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation      : STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 4);
	VARIABLE CLK_delayed        : STD_ULOGIC := 'X';
	VARIABLE T_delayed        : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_T_CLK_negedge,
	 TimingData		=> Tmkr_T_CLK_negedge,
	 TestSignal		=> T_ipd,
	 TestSignalName		=> "T",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_T_CLK_posedge_negedge,
	 SetupLow		=> tsetup_T_CLK_negedge_negedge,
	 HoldHigh		=> thold_T_CLK_posedge_negedge,
	 HoldLow		=> thold_T_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/TF1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_CLK_negedge,
	 TimingData		=> Tmkr_CLR_CLK_negedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_CLK_posedge_negedge,
 	 Removal                => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	  CheckEnabled		=>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "TF1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled           => TO_X01(( NOT CLR_ipd)) /= '1',
	 HeaderMsg		=> InstancePath & "TF1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled	 => TRUE,
	 HeaderMsg		=> InstancePath & "TF1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

	Violation := Tviol_T_CLK_negedge or 
		      Pviol_CLR or 
		      Pviol_CLK;

	VitalStateTable(
	 Result => Q_zd,
	PreviousDataIn => PrevData_Q,
	StateTable => tflipflop_Q_tab,
	DataIn => (
             CLR_ipd, CLK_ipd, T_delayed, Q_zd, CLK_delayed));
	Q_zd := Violation XOR Q_zd;
	--- now combinatorial logic input to the DFF 
	T_delayed :=  T_ipd ;
	CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	          1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_TF1B_VITAL of TF1B is
   for VITAL_ACT
   end for;
end CFG_TF1B_VITAL;



 ---- CELL TRIBUFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF :  entity is TRUE;
 end TRIBUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_VITAL of TRIBUFF is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_VITAL;



 ---- CELL TRIBUFF_S_8 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_8 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_8 :  entity is TRUE;
 end TRIBUFF_S_8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_8 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_8_VITAL of TRIBUFF_S_8 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_8_VITAL;



 ---- CELL TRIBUFF_S_8D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_8D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_8D :  entity is TRUE;
 end TRIBUFF_S_8D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_8D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_8D_VITAL of TRIBUFF_S_8D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_8D_VITAL;



 ---- CELL TRIBUFF_S_8U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_8U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_8U :  entity is TRUE;
 end TRIBUFF_S_8U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_8U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_8U_VITAL of TRIBUFF_S_8U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_8U_VITAL;



 ---- CELL TRIBUFF_S_12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_12 :  entity is TRUE;
 end TRIBUFF_S_12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_12_VITAL of TRIBUFF_S_12 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_12_VITAL;



 ---- CELL TRIBUFF_S_12D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_12D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_12D :  entity is TRUE;
 end TRIBUFF_S_12D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_12D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_12D_VITAL of TRIBUFF_S_12D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_12D_VITAL;



 ---- CELL TRIBUFF_S_12U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_12U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_12U :  entity is TRUE;
 end TRIBUFF_S_12U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_12U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_12U_VITAL of TRIBUFF_S_12U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_12U_VITAL;



 ---- CELL TRIBUFF_S_16 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_16 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_16 :  entity is TRUE;
 end TRIBUFF_S_16;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_16 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_16_VITAL of TRIBUFF_S_16 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_16_VITAL;



 ---- CELL TRIBUFF_S_16D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_16D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_16D :  entity is TRUE;
 end TRIBUFF_S_16D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_16D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_16D_VITAL of TRIBUFF_S_16D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_16D_VITAL;



 ---- CELL TRIBUFF_S_16U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_16U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_16U :  entity is TRUE;
 end TRIBUFF_S_16U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_16U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_16U_VITAL of TRIBUFF_S_16U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_16U_VITAL;



 ---- CELL TRIBUFF_S_24 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_24 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_24 :  entity is TRUE;
 end TRIBUFF_S_24;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_24 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_24_VITAL of TRIBUFF_S_24 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_24_VITAL;



 ---- CELL TRIBUFF_S_24D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_24D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_24D :  entity is TRUE;
 end TRIBUFF_S_24D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_24D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_24D_VITAL of TRIBUFF_S_24D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_24D_VITAL;



 ---- CELL TRIBUFF_S_24U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_24U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_24U :  entity is TRUE;
 end TRIBUFF_S_24U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_24U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_24U_VITAL of TRIBUFF_S_24U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_24U_VITAL;



 ---- CELL TRIBUFF_F_8 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_8 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_8 :  entity is TRUE;
 end TRIBUFF_F_8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_8 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_8_VITAL of TRIBUFF_F_8 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_8_VITAL;



 ---- CELL TRIBUFF_F_8D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_8D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_8D :  entity is TRUE;
 end TRIBUFF_F_8D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_8D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_8D_VITAL of TRIBUFF_F_8D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_8D_VITAL;



 ---- CELL TRIBUFF_F_8U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_8U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_8U :  entity is TRUE;
 end TRIBUFF_F_8U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_8U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_8U_VITAL of TRIBUFF_F_8U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_8U_VITAL;



 ---- CELL TRIBUFF_F_12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_12 :  entity is TRUE;
 end TRIBUFF_F_12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_12_VITAL of TRIBUFF_F_12 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_12_VITAL;



 ---- CELL TRIBUFF_F_12D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_12D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_12D :  entity is TRUE;
 end TRIBUFF_F_12D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_12D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_12D_VITAL of TRIBUFF_F_12D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_12D_VITAL;



 ---- CELL TRIBUFF_F_12U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_12U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_12U :  entity is TRUE;
 end TRIBUFF_F_12U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_12U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_12U_VITAL of TRIBUFF_F_12U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_12U_VITAL;



 ---- CELL TRIBUFF_F_16 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_16 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_16 :  entity is TRUE;
 end TRIBUFF_F_16;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_16 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_16_VITAL of TRIBUFF_F_16 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_16_VITAL;



 ---- CELL TRIBUFF_F_16D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_16D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_16D :  entity is TRUE;
 end TRIBUFF_F_16D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_16D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_16D_VITAL of TRIBUFF_F_16D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_16D_VITAL;



 ---- CELL TRIBUFF_F_16U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_16U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_16U :  entity is TRUE;
 end TRIBUFF_F_16U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_16U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_16U_VITAL of TRIBUFF_F_16U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_16U_VITAL;



 ---- CELL TRIBUFF_F_24 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_24 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_24 :  entity is TRUE;
 end TRIBUFF_F_24;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_24 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_24_VITAL of TRIBUFF_F_24 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_24_VITAL;



 ---- CELL TRIBUFF_F_24D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_24D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_24D :  entity is TRUE;
 end TRIBUFF_F_24D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_24D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_24D_VITAL of TRIBUFF_F_24D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_24D_VITAL;



 ---- CELL TRIBUFF_F_24U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_24U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_24U :  entity is TRUE;
 end TRIBUFF_F_24U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_24U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_24U_VITAL of TRIBUFF_F_24U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_24U_VITAL;



 ---- CELL TRIBUFF_LVCMOS25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS25 :  entity is TRUE;
 end TRIBUFF_LVCMOS25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS25_VITAL of TRIBUFF_LVCMOS25 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS25_VITAL;



 ---- CELL TRIBUFF_LVCMOS25D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS25D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS25D :  entity is TRUE;
 end TRIBUFF_LVCMOS25D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS25D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS25D_VITAL of TRIBUFF_LVCMOS25D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS25D_VITAL;



 ---- CELL TRIBUFF_LVCMOS25U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS25U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS25U :  entity is TRUE;
 end TRIBUFF_LVCMOS25U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS25U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS25U_VITAL of TRIBUFF_LVCMOS25U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS25U_VITAL;



 ---- CELL TRIBUFF_LVCMOS18 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS18 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS18 :  entity is TRUE;
 end TRIBUFF_LVCMOS18;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS18 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS18_VITAL of TRIBUFF_LVCMOS18 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS18_VITAL;



 ---- CELL TRIBUFF_LVCMOS18D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS18D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS18D :  entity is TRUE;
 end TRIBUFF_LVCMOS18D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS18D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS18D_VITAL of TRIBUFF_LVCMOS18D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS18D_VITAL;



 ---- CELL TRIBUFF_LVCMOS18U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS18U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS18U :  entity is TRUE;
 end TRIBUFF_LVCMOS18U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS18U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS18U_VITAL of TRIBUFF_LVCMOS18U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS18U_VITAL;



 ---- CELL TRIBUFF_LVCMOS15 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS15 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS15 :  entity is TRUE;
 end TRIBUFF_LVCMOS15;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS15 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS15_VITAL of TRIBUFF_LVCMOS15 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS15_VITAL;



 ---- CELL TRIBUFF_LVCMOS15D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS15D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS15D :  entity is TRUE;
 end TRIBUFF_LVCMOS15D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS15D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS15D_VITAL of TRIBUFF_LVCMOS15D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS15D_VITAL;



 ---- CELL TRIBUFF_LVCMOS15U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS15U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS15U :  entity is TRUE;
 end TRIBUFF_LVCMOS15U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS15U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS15U_VITAL of TRIBUFF_LVCMOS15U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS15U_VITAL;



 ---- CELL TRIBUFF_PCI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_PCI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_PCI :  entity is TRUE;
 end TRIBUFF_PCI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_PCI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_PCI_VITAL of TRIBUFF_PCI is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_PCI_VITAL;



 ---- CELL TRIBUFF_PCIX ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_PCIX is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_PCIX :  entity is TRUE;
 end TRIBUFF_PCIX;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_PCIX is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_PCIX_VITAL of TRIBUFF_PCIX is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_PCIX_VITAL;



 ---- CELL TRIBUFF_GTLP33 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_GTLP33 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_GTLP33 :  entity is TRUE;
 end TRIBUFF_GTLP33;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_GTLP33 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_GTLP33_VITAL of TRIBUFF_GTLP33 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_GTLP33_VITAL;



 ---- CELL TRIBUFF_GTLP25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_GTLP25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_GTLP25 :  entity is TRUE;
 end TRIBUFF_GTLP25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_GTLP25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_GTLP25_VITAL of TRIBUFF_GTLP25 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_GTLP25_VITAL;



 ---- CELL VCC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity VCC is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True		);
    port(
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of VCC :  entity is TRUE;
 end VCC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of VCC is
	attribute VITAL_LEVEL0 of VITAL_ACT : architecture is TRUE;


begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	--- Empty
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
        Y<= '1';


end VITAL_ACT;

 configuration CFG_VCC_VITAL of VCC is 
    for VITAL_ACT
    end for;
 end CFG_VCC_VITAL;



 ---- CELL XA1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XA1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XA1 :  entity is TRUE;
 end XA1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of XA1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XA1_VITAL of XA1 is 
    for VITAL_ACT
    end for;
 end CFG_XA1_VITAL;



 ---- CELL XA1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XA1A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XA1A :  entity is TRUE;
 end XA1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of XA1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( NOT VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XA1A_VITAL of XA1A is 
    for VITAL_ACT
    end for;
 end CFG_XA1A_VITAL;



 ---- CELL XA1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XA1B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XA1B :  entity is TRUE;
 end XA1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of XA1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) AND  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XA1B_VITAL of XA1B is 
    for VITAL_ACT
    end for;
 end CFG_XA1B_VITAL;



 ---- CELL XA1C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XA1C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XA1C :  entity is TRUE;
 end XA1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of XA1C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( NOT VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) AND  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XA1C_VITAL of XA1C is 
    for VITAL_ACT
    end for;
 end CFG_XA1C_VITAL;



 ---- CELL XAI1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XAI1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XAI1 :  entity is TRUE;
 end XAI1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of XAI1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XAI1_VITAL of XAI1 is 
    for VITAL_ACT
    end for;
 end CFG_XAI1_VITAL;



 ---- CELL XAI1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XAI1A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XAI1A :  entity is TRUE;
 end XAI1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of XAI1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  NOT VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XAI1A_VITAL of XAI1A is 
    for VITAL_ACT
    end for;
 end CFG_XAI1A_VITAL;



 ---- CELL XNOR2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XNOR2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XNOR2 :  entity is TRUE;
 end XNOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of XNOR2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XNOR2_VITAL of XNOR2 is 
    for VITAL_ACT
    end for;
 end CFG_XNOR2_VITAL;



 ---- CELL XNOR3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XNOR3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XNOR3 :  entity is TRUE;
 end XNOR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of XNOR3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) XOR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XNOR3_VITAL of XNOR3 is 
    for VITAL_ACT
    end for;
 end CFG_XNOR3_VITAL;



 ---- CELL XNOR4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XNOR4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XNOR4 :  entity is TRUE;
 end XNOR4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of XNOR4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) XOR  C_ipd ) XOR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XNOR4_VITAL of XNOR4 is 
    for VITAL_ACT
    end for;
 end CFG_XNOR4_VITAL;



 ---- CELL XO1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XO1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XO1 :  entity is TRUE;
 end XO1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of XO1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XO1_VITAL of XO1 is 
    for VITAL_ACT
    end for;
 end CFG_XO1_VITAL;



 ---- CELL XO1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XO1A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XO1A :  entity is TRUE;
 end XO1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of XO1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( NOT VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XO1A_VITAL of XO1A is 
    for VITAL_ACT
    end for;
 end CFG_XO1A_VITAL;



 ---- CELL XOR2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XOR2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XOR2 :  entity is TRUE;
 end XOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of XOR2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XOR2_VITAL of XOR2 is 
    for VITAL_ACT
    end for;
 end CFG_XOR2_VITAL;



 ---- CELL XOR3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XOR3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XOR3 :  entity is TRUE;
 end XOR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of XOR3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) XOR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XOR3_VITAL of XOR3 is 
    for VITAL_ACT
    end for;
 end CFG_XOR3_VITAL;



 ---- CELL XOR4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XOR4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		D		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XOR4 :  entity is TRUE;
 end XOR4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of XOR4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) XOR  C_ipd ) XOR  D_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (D_ipd'last_event,tpd_D_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XOR4_VITAL of XOR4 is 
    for VITAL_ACT
    end for;
 end CFG_XOR4_VITAL;



 ---- CELL XOR4_FCI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XOR4_FCI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_FCI_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_FCI		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		FCI		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XOR4_FCI :  entity is TRUE;
 end XOR4_FCI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of XOR4_FCI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL FCI_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (FCI_ipd, FCI, tipd_FCI);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd, FCI_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) XOR  C_ipd ) XOR  FCI_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true),
	             3 => (FCI_ipd'last_event,tpd_FCI_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XOR4_FCI_VITAL of XOR4_FCI is 
    for VITAL_ACT
    end for;
 end CFG_XOR4_FCI_VITAL;



 ---- CELL ZOR3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity ZOR3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of ZOR3 :  entity is TRUE;
 end ZOR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of ZOR3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2(( A_ipd  AND  B_ipd ),( (NOT A_ipd)  AND  (NOT B_ipd) ), C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_ZOR3_VITAL of ZOR3 is 
    for VITAL_ACT
    end for;
 end CFG_ZOR3_VITAL;



 ---- CELL ZOR3I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity ZOR3I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of ZOR3I :  entity is TRUE;
 end ZOR3I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of ZOR3I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT VitalMUX2(( A_ipd  AND  B_ipd ),( (NOT A_ipd)  AND  (NOT B_ipd) ), C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_ZOR3I_VITAL of ZOR3I is 
    for VITAL_ACT
    end for;
 end CFG_ZOR3I_VITAL;



 ---- CELL IOFIFO_BIBUF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOFIFO_BIBUF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_AIN_YIN		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_AOUT_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_AIN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_AOUT		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		AIN		: in    STD_ULOGIC;
		AOUT		: in    STD_ULOGIC;
		YIN		: out    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOFIFO_BIBUF :  entity is TRUE;
 end IOFIFO_BIBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOFIFO_BIBUF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL AIN_ipd  : STD_ULOGIC := 'X';
	SIGNAL AOUT_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (AIN_ipd, AIN, tipd_AIN);
	VitalWireDelay (AOUT_ipd, AOUT, tipd_AOUT);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (AIN_ipd, AOUT_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS YIN_zd : STD_LOGIC is Results(1);
	ALIAS YOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE YIN_GlitchData  : VitalGlitchDataType;
	VARIABLE YOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        YIN_zd :=TO_X01(AIN_ipd);
        YOUT_zd :=TO_X01(AOUT_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => YIN,
	   GlitchData => YIN_GlitchData,
	   OutSignalName => "YIN",
	   OutTemp => YIN_zd,
	   Paths => (
	             0 => (AIN_ipd'last_event,tpd_AIN_YIN, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => YOUT,
	   GlitchData => YOUT_GlitchData,
	   OutSignalName => "YOUT",
	   OutTemp => YOUT_zd,
	   Paths => (
	             0 => (AOUT_ipd'last_event,tpd_AOUT_YOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOFIFO_BIBUF_VITAL of IOFIFO_BIBUF is 
    for VITAL_ACT
    end for;
 end CFG_IOFIFO_BIBUF_VITAL;



 ---- CELL IOI_FCLK_EN_BUFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOI_FCLK_EN_BUFF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_ENOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		ENOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOI_FCLK_EN_BUFF :  entity is TRUE;
 end IOI_FCLK_EN_BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOI_FCLK_EN_BUFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, CLK_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS ENOUT_zd : STD_LOGIC is Results(2);
	ALIAS CLKOUT_zd : STD_LOGIC is Results(3);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE ENOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE CLKOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);
        ENOUT_zd :=TO_X01(EN_ipd);
        CLKOUT_zd :=TO_X01(CLK_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => ENOUT,
	   GlitchData => ENOUT_GlitchData,
	   OutSignalName => "ENOUT",
	   OutTemp => ENOUT_zd,
	   Paths => (
	             0 => (EN_ipd'last_event,tpd_EN_ENOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CLKOUT,
	   GlitchData => CLKOUT_GlitchData,
	   OutSignalName => "CLKOUT",
	   OutTemp => CLKOUT_zd,
	   Paths => (
	             0 => (CLK_ipd'last_event,tpd_CLK_CLKOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOI_FCLK_EN_BUFF_VITAL of IOI_FCLK_EN_BUFF is 
    for VITAL_ACT
    end for;
 end CFG_IOI_FCLK_EN_BUFF_VITAL;



 ---- CELL IOI_FCLK_BUFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOI_FCLK_BUFF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOI_FCLK_BUFF :  entity is TRUE;
 end IOI_FCLK_BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOI_FCLK_BUFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, CLK_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS CLKOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE CLKOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);
        CLKOUT_zd :=TO_X01(CLK_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CLKOUT,
	   GlitchData => CLKOUT_GlitchData,
	   OutSignalName => "CLKOUT",
	   OutTemp => CLKOUT_zd,
	   Paths => (
	             0 => (CLK_ipd'last_event,tpd_CLK_CLKOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOI_FCLK_BUFF_VITAL of IOI_FCLK_BUFF is 
    for VITAL_ACT
    end for;
 end CFG_IOI_FCLK_BUFF_VITAL;



 ---- CELL IOI_RCLK_EN_BUFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOI_RCLK_EN_BUFF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_ENOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		ENOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOI_RCLK_EN_BUFF :  entity is TRUE;
 end IOI_RCLK_EN_BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOI_RCLK_EN_BUFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, CLK_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS ENOUT_zd : STD_LOGIC is Results(2);
	ALIAS CLKOUT_zd : STD_LOGIC is Results(3);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE ENOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE CLKOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);
        ENOUT_zd :=TO_X01(EN_ipd);
        CLKOUT_zd :=TO_X01(CLK_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => ENOUT,
	   GlitchData => ENOUT_GlitchData,
	   OutSignalName => "ENOUT",
	   OutTemp => ENOUT_zd,
	   Paths => (
	             0 => (EN_ipd'last_event,tpd_EN_ENOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CLKOUT,
	   GlitchData => CLKOUT_GlitchData,
	   OutSignalName => "CLKOUT",
	   OutTemp => CLKOUT_zd,
	   Paths => (
	             0 => (CLK_ipd'last_event,tpd_CLK_CLKOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOI_RCLK_EN_BUFF_VITAL of IOI_RCLK_EN_BUFF is 
    for VITAL_ACT
    end for;
 end CFG_IOI_RCLK_EN_BUFF_VITAL;



 ---- CELL IOI_RCLK_BUFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOI_RCLK_BUFF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOI_RCLK_BUFF :  entity is TRUE;
 end IOI_RCLK_BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOI_RCLK_BUFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, CLK_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS CLKOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE CLKOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);
        CLKOUT_zd :=TO_X01(CLK_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CLKOUT,
	   GlitchData => CLKOUT_GlitchData,
	   OutSignalName => "CLKOUT",
	   OutTemp => CLKOUT_zd,
	   Paths => (
	             0 => (CLK_ipd'last_event,tpd_CLK_CLKOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOI_RCLK_BUFF_VITAL of IOI_RCLK_BUFF is 
    for VITAL_ACT
    end for;
 end CFG_IOI_RCLK_BUFF_VITAL;



 ---- CELL IOOE_FCLK_EN_BUFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOOE_FCLK_EN_BUFF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_ENOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC;
		ENOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOOE_FCLK_EN_BUFF :  entity is TRUE;
 end IOOE_FCLK_EN_BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOOE_FCLK_EN_BUFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, CLK_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
	ALIAS YOUT_zd : STD_LOGIC is Results(1);
	ALIAS ENOUT_zd : STD_LOGIC is Results(2);
	ALIAS CLKOUT_zd : STD_LOGIC is Results(3);

	-- output glitch detection variables
	VARIABLE YOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE ENOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE CLKOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        YOUT_zd :=TO_X01(A_ipd);
        ENOUT_zd :=TO_X01(EN_ipd);
        CLKOUT_zd :=TO_X01(CLK_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => YOUT,
	   GlitchData => YOUT_GlitchData,
	   OutSignalName => "YOUT",
	   OutTemp => YOUT_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_YOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => ENOUT,
	   GlitchData => ENOUT_GlitchData,
	   OutSignalName => "ENOUT",
	   OutTemp => ENOUT_zd,
	   Paths => (
	             0 => (EN_ipd'last_event,tpd_EN_ENOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CLKOUT,
	   GlitchData => CLKOUT_GlitchData,
	   OutSignalName => "CLKOUT",
	   OutTemp => CLKOUT_zd,
	   Paths => (
	             0 => (CLK_ipd'last_event,tpd_CLK_CLKOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOOE_FCLK_EN_BUFF_VITAL of IOOE_FCLK_EN_BUFF is 
    for VITAL_ACT
    end for;
 end CFG_IOOE_FCLK_EN_BUFF_VITAL;



 ---- CELL IOOE_FCLK ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOOE_FCLK is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		: in    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOOE_FCLK :  entity is TRUE;
 end IOOE_FCLK;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOOE_FCLK is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL CLK_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (CLK_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS CLKOUT_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE CLKOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        CLKOUT_zd :=TO_X01(CLK_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => CLKOUT,
	   GlitchData => CLKOUT_GlitchData,
	   OutSignalName => "CLKOUT",
	   OutTemp => CLKOUT_zd,
	   Paths => (
	             0 => (CLK_ipd'last_event,tpd_CLK_CLKOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOOE_FCLK_VITAL of IOOE_FCLK is 
    for VITAL_ACT
    end for;
 end CFG_IOOE_FCLK_VITAL;



 ---- CELL IOOE_RCLK_EN_BUFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOOE_RCLK_EN_BUFF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_ENOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC;
		ENOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOOE_RCLK_EN_BUFF :  entity is TRUE;
 end IOOE_RCLK_EN_BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOOE_RCLK_EN_BUFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, CLK_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
	ALIAS YOUT_zd : STD_LOGIC is Results(1);
	ALIAS ENOUT_zd : STD_LOGIC is Results(2);
	ALIAS CLKOUT_zd : STD_LOGIC is Results(3);

	-- output glitch detection variables
	VARIABLE YOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE ENOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE CLKOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        YOUT_zd :=TO_X01(A_ipd);
        ENOUT_zd :=TO_X01(EN_ipd);
        CLKOUT_zd :=TO_X01(CLK_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => YOUT,
	   GlitchData => YOUT_GlitchData,
	   OutSignalName => "YOUT",
	   OutTemp => YOUT_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_YOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => ENOUT,
	   GlitchData => ENOUT_GlitchData,
	   OutSignalName => "ENOUT",
	   OutTemp => ENOUT_zd,
	   Paths => (
	             0 => (EN_ipd'last_event,tpd_EN_ENOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CLKOUT,
	   GlitchData => CLKOUT_GlitchData,
	   OutSignalName => "CLKOUT",
	   OutTemp => CLKOUT_zd,
	   Paths => (
	             0 => (CLK_ipd'last_event,tpd_CLK_CLKOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOOE_RCLK_EN_BUFF_VITAL of IOOE_RCLK_EN_BUFF is 
    for VITAL_ACT
    end for;
 end CFG_IOOE_RCLK_EN_BUFF_VITAL;



 ---- CELL IOOE_RCLK_CLR_EN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOOE_RCLK_CLR_EN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_CLR_CLROUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_ENOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_CLR		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		CLROUT		: out    STD_ULOGIC;
		ENOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOOE_RCLK_CLR_EN :  entity is TRUE;
 end IOOE_RCLK_CLR_EN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOOE_RCLK_CLR_EN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (CLR_ipd, EN_ipd, CLK_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
	ALIAS CLROUT_zd : STD_LOGIC is Results(1);
	ALIAS ENOUT_zd : STD_LOGIC is Results(2);
	ALIAS CLKOUT_zd : STD_LOGIC is Results(3);

	-- output glitch detection variables
	VARIABLE CLROUT_GlitchData  : VitalGlitchDataType;
	VARIABLE ENOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE CLKOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        CLROUT_zd :=TO_X01(CLR_ipd);
        ENOUT_zd :=TO_X01(EN_ipd);
        CLKOUT_zd :=TO_X01(CLK_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => CLROUT,
	   GlitchData => CLROUT_GlitchData,
	   OutSignalName => "CLROUT",
	   OutTemp => CLROUT_zd,
	   Paths => (
	             0 => (CLR_ipd'last_event,tpd_CLR_CLROUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => ENOUT,
	   GlitchData => ENOUT_GlitchData,
	   OutSignalName => "ENOUT",
	   OutTemp => ENOUT_zd,
	   Paths => (
	             0 => (EN_ipd'last_event,tpd_EN_ENOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CLKOUT,
	   GlitchData => CLKOUT_GlitchData,
	   OutSignalName => "CLKOUT",
	   OutTemp => CLKOUT_zd,
	   Paths => (
	             0 => (CLK_ipd'last_event,tpd_CLK_CLKOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOOE_RCLK_CLR_EN_VITAL of IOOE_RCLK_CLR_EN is 
    for VITAL_ACT
    end for;
 end CFG_IOOE_RCLK_CLR_EN_VITAL;



 ---- CELL IOOE_RCLK_BUFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOOE_RCLK_BUFF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOOE_RCLK_BUFF :  entity is TRUE;
 end IOOE_RCLK_BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOOE_RCLK_BUFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, CLK_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS YOUT_zd : STD_LOGIC is Results(1);
	ALIAS CLKOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE YOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE CLKOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        YOUT_zd :=TO_X01(A_ipd);
        CLKOUT_zd :=TO_X01(CLK_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => YOUT,
	   GlitchData => YOUT_GlitchData,
	   OutSignalName => "YOUT",
	   OutTemp => YOUT_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_YOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CLKOUT,
	   GlitchData => CLKOUT_GlitchData,
	   OutSignalName => "CLKOUT",
	   OutTemp => CLKOUT_zd,
	   Paths => (
	             0 => (CLK_ipd'last_event,tpd_CLK_CLKOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOOE_RCLK_BUFF_VITAL of IOOE_RCLK_BUFF is 
    for VITAL_ACT
    end for;
 end CFG_IOOE_RCLK_BUFF_VITAL;



 ---- CELL IOOE_RCLK ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOOE_RCLK is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		: in    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOOE_RCLK :  entity is TRUE;
 end IOOE_RCLK;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOOE_RCLK is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL CLK_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (CLK_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS CLKOUT_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE CLKOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        CLKOUT_zd :=TO_X01(CLK_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => CLKOUT,
	   GlitchData => CLKOUT_GlitchData,
	   OutSignalName => "CLKOUT",
	   OutTemp => CLKOUT_zd,
	   Paths => (
	             0 => (CLK_ipd'last_event,tpd_CLK_CLKOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOOE_RCLK_VITAL of IOOE_RCLK is 
    for VITAL_ACT
    end for;
 end CFG_IOOE_RCLK_VITAL;



 ---- CELL PLLINT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity PLLINT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of PLLINT :  entity is TRUE;
 end PLLINT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of PLLINT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_PLLINT_VITAL of PLLINT is 
    for VITAL_ACT
    end for;
 end CFG_PLLINT_VITAL;



 ---- CELL PLLOUT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity PLLOUT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of PLLOUT :  entity is TRUE;
 end PLLOUT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of PLLOUT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_PLLOUT_VITAL of PLLOUT is 
    for VITAL_ACT
    end for;
 end CFG_PLLOUT_VITAL;



 ---- CELL BIBUF_HSTL_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_HSTL_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_HSTL_I :  entity is TRUE;
 end BIBUF_HSTL_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_HSTL_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_HSTL_I_VITAL of BIBUF_HSTL_I is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_HSTL_I_VITAL;



 ---- CELL BIBUF_SSTL3_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_SSTL3_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_SSTL3_I :  entity is TRUE;
 end BIBUF_SSTL3_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_SSTL3_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_SSTL3_I_VITAL of BIBUF_SSTL3_I is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_SSTL3_I_VITAL;



 ---- CELL BIBUF_SSTL3_II ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_SSTL3_II is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_SSTL3_II :  entity is TRUE;
 end BIBUF_SSTL3_II;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_SSTL3_II is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_SSTL3_II_VITAL of BIBUF_SSTL3_II is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_SSTL3_II_VITAL;



 ---- CELL BIBUF_SSTL2_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_SSTL2_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_SSTL2_I :  entity is TRUE;
 end BIBUF_SSTL2_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_SSTL2_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_SSTL2_I_VITAL of BIBUF_SSTL2_I is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_SSTL2_I_VITAL;



 ---- CELL BIBUF_SSTL2_II ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_SSTL2_II is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_SSTL2_II :  entity is TRUE;
 end BIBUF_SSTL2_II;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BIBUF_SSTL2_II is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_SSTL2_II_VITAL of BIBUF_SSTL2_II is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_SSTL2_II_VITAL;



 ---- CELL BUFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BUFF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BUFF :  entity is TRUE;
 end BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of BUFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BUFF_VITAL of BUFF is 
    for VITAL_ACT
    end for;
 end CFG_BUFF_VITAL;



 ---- CELL CLKINT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKINT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKINT :  entity is TRUE;
 end CLKINT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKINT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKINT_VITAL of CLKINT is 
    for VITAL_ACT
    end for;
 end CFG_CLKINT_VITAL;



 ---- CELL CLKINT_W ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKINT_W is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKINT_W :  entity is TRUE;
 end CLKINT_W;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKINT_W is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKINT_W_VITAL of CLKINT_W is 
    for VITAL_ACT
    end for;
 end CFG_CLKINT_W_VITAL;



 ---- CELL CLKOUT_E ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKOUT_E is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKOUT_E :  entity is TRUE;
 end CLKOUT_E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKOUT_E is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKOUT_E_VITAL of CLKOUT_E is 
    for VITAL_ACT
    end for;
 end CFG_CLKOUT_E_VITAL;



 ---- CELL CLKOUT_W ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKOUT_W is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKOUT_W :  entity is TRUE;
 end CLKOUT_W;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of CLKOUT_W is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKOUT_W_VITAL of CLKOUT_W is 
    for VITAL_ACT
    end for;
 end CFG_CLKOUT_W_VITAL;



 ---- CELL DFM ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFM is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFM :  entity is TRUE;
 end DFM;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFM is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (S_ipd, S, tipd_S);
	  VitalWireDelay (A_ipd, A, tipd_A);
	  VitalWireDelay (B_ipd, B, tipd_B);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (S_ipd, A_ipd, B_ipd, CLK_ipd)

	-- timing check results
	VARIABLE Tviol_S_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_S_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_A_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_A_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_B_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_CLK_posedge,
	 TimingData		=> Tmkr_S_CLK_posedge,
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_CLK_posedge_posedge,
	 SetupLow		=> tsetup_S_CLK_negedge_posedge,
	 HoldHigh		=> thold_S_CLK_posedge_posedge,
	 HoldLow		=> thold_S_CLK_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFM",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_CLK_posedge,
	 TimingData		=> Tmkr_A_CLK_posedge,
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_CLK_posedge_posedge,
	 SetupLow		=> tsetup_A_CLK_negedge_posedge,
	 HoldHigh		=> thold_A_CLK_posedge_posedge,
	 HoldLow		=> thold_A_CLK_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFM",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_CLK_posedge,
	 TimingData		=> Tmkr_B_CLK_posedge,
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_CLK_posedge_posedge,
	 SetupLow		=> tsetup_B_CLK_negedge_posedge,
	 HoldHigh		=> thold_B_CLK_posedge_posedge,
	 HoldLow		=> thold_B_CLK_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFM",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFM",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S_CLK_posedge or 
	 Tviol_A_CLK_posedge or 
	 Tviol_B_CLK_posedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, NET_0_2, '0', '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
         --- now combinatorial logic input to the DFF 
   NET_0_2 :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFM_VITAL of DFM is
   for VITAL_ACT
   end for;
end CFG_DFM_VITAL;



 ---- CELL DFM3B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFM3B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFM3B :  entity is TRUE;
 end DFM3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFM3B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (S_ipd, S, tipd_S);
	  VitalWireDelay (A_ipd, A, tipd_A);
	  VitalWireDelay (B_ipd, B, tipd_B);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (S_ipd, A_ipd, B_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_S_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_S_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_A_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_A_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_B_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_CLK_negedge, 
	 TimingData		=> Tmkr_S_CLK_negedge, 
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_CLK_posedge_negedge,
	 SetupLow		=> tsetup_S_CLK_negedge_negedge,
	 HoldHigh		=> thold_S_CLK_posedge_negedge,
	 HoldLow		=> thold_S_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFM3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_CLK_negedge, 
	 TimingData		=> Tmkr_A_CLK_negedge, 
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_CLK_posedge_negedge,
	 SetupLow		=> tsetup_A_CLK_negedge_negedge,
	 HoldHigh		=> thold_A_CLK_posedge_negedge,
	 HoldLow		=> thold_A_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFM3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_CLK_negedge, 
	 TimingData		=> Tmkr_B_CLK_negedge, 
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_CLK_posedge_negedge,
	 SetupLow		=> tsetup_B_CLK_negedge_negedge,
	 HoldHigh		=> thold_B_CLK_posedge_negedge,
	 HoldLow		=> thold_B_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFM3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>    TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFM3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFM3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFM3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S_CLK_negedge or 
	 Tviol_A_CLK_negedge or 
	 Tviol_B_CLK_negedge or 
	 Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, Q_zd, NET_0_2, '0', '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
         --- now combinatorial logic input to the DFF 
   NET_0_2 :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFM3B_VITAL of DFM3B is
   for VITAL_ACT
   end for;
end CFG_DFM3B_VITAL;



 ---- CELL DFM4A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFM4A is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFM4A :  entity is TRUE;
 end DFM4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFM4A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (S_ipd, S, tipd_S);
	  VitalWireDelay (A_ipd, A, tipd_A);
	  VitalWireDelay (B_ipd, B, tipd_B);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (S_ipd, A_ipd, B_ipd, PRE_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_S_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_S_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_A_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_A_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_B_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_CLK_posedge,
	 TimingData		=> Tmkr_S_CLK_posedge,
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_CLK_posedge_posedge,
	 SetupLow		=> tsetup_S_CLK_negedge_posedge,
	 HoldHigh		=> thold_S_CLK_posedge_posedge,
	 HoldLow		=> thold_S_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFM4A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_CLK_posedge,
	 TimingData		=> Tmkr_A_CLK_posedge,
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_CLK_posedge_posedge,
	 SetupLow		=> tsetup_A_CLK_negedge_posedge,
	 HoldHigh		=> thold_A_CLK_posedge_posedge,
	 HoldLow		=> thold_A_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFM4A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_CLK_posedge,
	 TimingData		=> Tmkr_B_CLK_posedge,
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_CLK_posedge_posedge,
	 SetupLow		=> tsetup_B_CLK_negedge_posedge,
	 HoldHigh		=> thold_B_CLK_posedge_posedge,
	 HoldLow		=> thold_B_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFM4A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFM4A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFM4A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFM4A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S_CLK_posedge or 
	 Tviol_A_CLK_posedge or 
	 Tviol_B_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, NET_0_2, '0', PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;
         --- now combinatorial logic input to the DFF 
   NET_0_2 :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFM4A_VITAL of DFM4A is
   for VITAL_ACT
   end for;
end CFG_DFM4A_VITAL;



 ---- CELL DFM4B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFM4B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFM4B :  entity is TRUE;
 end DFM4B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFM4B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (S_ipd, S, tipd_S);
	  VitalWireDelay (A_ipd, A, tipd_A);
	  VitalWireDelay (B_ipd, B, tipd_B);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (S_ipd, A_ipd, B_ipd, PRE_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_S_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_S_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_A_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_A_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_B_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_CLK_negedge, 
	 TimingData		=> Tmkr_S_CLK_negedge, 
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_CLK_posedge_negedge,
	 SetupLow		=> tsetup_S_CLK_negedge_negedge,
	 HoldHigh		=> thold_S_CLK_posedge_negedge,
	 HoldLow		=> thold_S_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFM4B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_CLK_negedge, 
	 TimingData		=> Tmkr_A_CLK_negedge, 
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_CLK_posedge_negedge,
	 SetupLow		=> tsetup_A_CLK_negedge_negedge,
	 HoldHigh		=> thold_A_CLK_posedge_negedge,
	 HoldLow		=> thold_A_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFM4B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_CLK_negedge, 
	 TimingData		=> Tmkr_B_CLK_negedge, 
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_CLK_posedge_negedge,
	 SetupLow		=> tsetup_B_CLK_negedge_negedge,
	 HoldHigh		=> thold_B_CLK_posedge_negedge,
	 HoldLow		=> thold_B_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFM4B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFM4B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFM4B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFM4B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S_CLK_negedge or 
	 Tviol_A_CLK_negedge or 
	 Tviol_B_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, NET_0_2, '0', PRE_ipd, CLK_delayed));
   Q_zd := Violation XOR Q_zd;
         --- now combinatorial logic input to the DFF 
   NET_0_2 :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFM4B_VITAL of DFM4B is
   for VITAL_ACT
   end for;
end CFG_DFM4B_VITAL;



 ---- CELL DFMA ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFMA is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFMA :  entity is TRUE;
 end DFMA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFMA is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (S_ipd, S, tipd_S);
	  VitalWireDelay (A_ipd, A, tipd_A);
	  VitalWireDelay (B_ipd, B, tipd_B);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (S_ipd, A_ipd, B_ipd, CLK_ipd)

	-- timing check results
	VARIABLE Tviol_S_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_S_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_A_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_A_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_B_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_CLK_negedge, 
	 TimingData		=> Tmkr_S_CLK_negedge, 
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_CLK_posedge_negedge,
	 SetupLow		=> tsetup_S_CLK_negedge_negedge,
	 HoldHigh		=> thold_S_CLK_posedge_negedge,
	 HoldLow		=> thold_S_CLK_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFMA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_CLK_negedge, 
	 TimingData		=> Tmkr_A_CLK_negedge, 
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_CLK_posedge_negedge,
	 SetupLow		=> tsetup_A_CLK_negedge_negedge,
	 HoldHigh		=> thold_A_CLK_posedge_negedge,
	 HoldLow		=> thold_A_CLK_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFMA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_CLK_negedge, 
	 TimingData		=> Tmkr_B_CLK_negedge, 
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_CLK_posedge_negedge,
	 SetupLow		=> tsetup_B_CLK_negedge_negedge,
	 HoldHigh		=> thold_B_CLK_posedge_negedge,
	 HoldLow		=> thold_B_CLK_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFMA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFMA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S_CLK_negedge or 
	 Tviol_A_CLK_negedge or 
	 Tviol_B_CLK_negedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, NET_0_2, '0', '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
         --- now combinatorial logic input to the DFF 
   NET_0_2 :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFMA_VITAL of DFMA is
   for VITAL_ACT
   end for;
end CFG_DFMA_VITAL;



 ---- CELL DFMB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFMB is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFMB :  entity is TRUE;
 end DFMB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFMB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (S_ipd, S, tipd_S);
	  VitalWireDelay (A_ipd, A, tipd_A);
	  VitalWireDelay (B_ipd, B, tipd_B);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (S_ipd, A_ipd, B_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_S_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_S_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_A_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_A_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_B_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_CLK_posedge,
	 TimingData		=> Tmkr_S_CLK_posedge,
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_CLK_posedge_posedge,
	 SetupLow		=> tsetup_S_CLK_negedge_posedge,
	 HoldHigh		=> thold_S_CLK_posedge_posedge,
	 HoldLow		=> thold_S_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFMB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_CLK_posedge,
	 TimingData		=> Tmkr_A_CLK_posedge,
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_CLK_posedge_posedge,
	 SetupLow		=> tsetup_A_CLK_negedge_posedge,
	 HoldHigh		=> thold_A_CLK_posedge_posedge,
	 HoldLow		=> thold_A_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFMB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_CLK_posedge,
	 TimingData		=> Tmkr_B_CLK_posedge,
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_CLK_posedge_posedge,
	 SetupLow		=> tsetup_B_CLK_negedge_posedge,
	 HoldHigh		=> thold_B_CLK_posedge_posedge,
	 HoldLow		=> thold_B_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFMB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>    TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFMB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFMB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFMB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S_CLK_posedge or 
	 Tviol_A_CLK_posedge or 
	 Tviol_B_CLK_posedge or 
	 Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, NET_0_2, '0', '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
         --- now combinatorial logic input to the DFF 
   NET_0_2 :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFMB_VITAL of DFMB is
   for VITAL_ACT
   end for;
end CFG_DFMB_VITAL;



 ---- CELL DFME1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFME1A is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFME1A :  entity is TRUE;
 end DFME1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFME1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (S_ipd, S, tipd_S);
	  VitalWireDelay (A_ipd, A, tipd_A);
	  VitalWireDelay (B_ipd, B, tipd_B);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (S_ipd, A_ipd, B_ipd, E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_S_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_S_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_A_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_A_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_B_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_CLK_posedge,
	 TimingData		=> Tmkr_S_CLK_posedge,
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_CLK_posedge_posedge,
	 SetupLow		=> tsetup_S_CLK_negedge_posedge,
	 HoldHigh		=> thold_S_CLK_posedge_posedge,
	 HoldLow		=> thold_S_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFME1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_CLK_posedge,
	 TimingData		=> Tmkr_A_CLK_posedge,
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_CLK_posedge_posedge,
	 SetupLow		=> tsetup_A_CLK_negedge_posedge,
	 HoldHigh		=> thold_A_CLK_posedge_posedge,
	 HoldLow		=> thold_A_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFME1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_CLK_posedge,
	 TimingData		=> Tmkr_B_CLK_posedge,
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_CLK_posedge_posedge,
	 SetupLow		=> tsetup_B_CLK_negedge_posedge,
	 HoldHigh		=> thold_B_CLK_posedge_posedge,
	 HoldLow		=> thold_B_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFME1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TRUE,	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFME1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFME1A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S_CLK_posedge or 
	 Tviol_A_CLK_posedge or 
	 Tviol_B_CLK_posedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, NET_0_2, E_delayed, '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
         --- now combinatorial logic input to the DFF 
   NET_0_2 :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFME1A_VITAL of DFME1A is
   for VITAL_ACT
   end for;
end CFG_DFME1A_VITAL;



 ---- CELL DFME1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFME1B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFME1B :  entity is TRUE;
 end DFME1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFME1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (S_ipd, S, tipd_S);
	  VitalWireDelay (A_ipd, A, tipd_A);
	  VitalWireDelay (B_ipd, B, tipd_B);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (S_ipd, A_ipd, B_ipd, E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_S_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_S_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_A_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_A_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_B_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_CLK_negedge, 
	 TimingData		=> Tmkr_S_CLK_negedge, 
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_CLK_posedge_negedge,
	 SetupLow		=> tsetup_S_CLK_negedge_negedge,
	 HoldHigh		=> thold_S_CLK_posedge_negedge,
	 HoldLow		=> thold_S_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFME1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_CLK_negedge, 
	 TimingData		=> Tmkr_A_CLK_negedge, 
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_CLK_posedge_negedge,
	 SetupLow		=> tsetup_A_CLK_negedge_negedge,
	 HoldHigh		=> thold_A_CLK_posedge_negedge,
	 HoldLow		=> thold_A_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFME1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_CLK_negedge, 
	 TimingData		=> Tmkr_B_CLK_negedge, 
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_CLK_posedge_negedge,
	 SetupLow		=> tsetup_B_CLK_negedge_negedge,
	 HoldHigh		=> thold_B_CLK_posedge_negedge,
	 HoldLow		=> thold_B_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFME1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TRUE,	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFME1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFME1B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S_CLK_negedge or 
	 Tviol_A_CLK_negedge or 
	 Tviol_B_CLK_negedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, NET_0_2, E_delayed, '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
         --- now combinatorial logic input to the DFF 
   NET_0_2 :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFME1B_VITAL of DFME1B is
   for VITAL_ACT
   end for;
end CFG_DFME1B_VITAL;



 ---- CELL DFME2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFME2A is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFME2A :  entity is TRUE;
 end DFME2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFME2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (S_ipd, S, tipd_S);
	  VitalWireDelay (A_ipd, A, tipd_A);
	  VitalWireDelay (B_ipd, B, tipd_B);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (S_ipd, A_ipd, B_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_S_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_S_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_A_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_A_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_B_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_CLK_posedge,
	 TimingData		=> Tmkr_S_CLK_posedge,
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_CLK_posedge_posedge,
	 SetupLow		=> tsetup_S_CLK_negedge_posedge,
	 HoldHigh		=> thold_S_CLK_posedge_posedge,
	 HoldLow		=> thold_S_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFME2A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_CLK_posedge,
	 TimingData		=> Tmkr_A_CLK_posedge,
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_CLK_posedge_posedge,
	 SetupLow		=> tsetup_A_CLK_negedge_posedge,
	 HoldHigh		=> thold_A_CLK_posedge_posedge,
	 HoldLow		=> thold_A_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFME2A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_CLK_posedge,
	 TimingData		=> Tmkr_B_CLK_posedge,
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_CLK_posedge_posedge,
	 SetupLow		=> tsetup_B_CLK_negedge_posedge,
	 HoldHigh		=> thold_B_CLK_posedge_posedge,
	 HoldLow		=> thold_B_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFME2A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFME2A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFME2A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFME2A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFME2A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S_CLK_posedge or 
	 Tviol_A_CLK_posedge or 
	 Tviol_B_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, NET_0_2, E_delayed, PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;
         --- now combinatorial logic input to the DFF 
   NET_0_2 :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFME2A_VITAL of DFME2A is
   for VITAL_ACT
   end for;
end CFG_DFME2A_VITAL;



 ---- CELL DFME2B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFME2B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFME2B :  entity is TRUE;
 end DFME2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFME2B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (S_ipd, S, tipd_S);
	  VitalWireDelay (A_ipd, A, tipd_A);
	  VitalWireDelay (B_ipd, B, tipd_B);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (S_ipd, A_ipd, B_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_S_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_S_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_A_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_A_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_B_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_CLK_negedge, 
	 TimingData		=> Tmkr_S_CLK_negedge, 
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_CLK_posedge_negedge,
	 SetupLow		=> tsetup_S_CLK_negedge_negedge,
	 HoldHigh		=> thold_S_CLK_posedge_negedge,
	 HoldLow		=> thold_S_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFME2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_CLK_negedge, 
	 TimingData		=> Tmkr_A_CLK_negedge, 
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_CLK_posedge_negedge,
	 SetupLow		=> tsetup_A_CLK_negedge_negedge,
	 HoldHigh		=> thold_A_CLK_posedge_negedge,
	 HoldLow		=> thold_A_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFME2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_CLK_negedge, 
	 TimingData		=> Tmkr_B_CLK_negedge, 
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_CLK_posedge_negedge,
	 SetupLow		=> tsetup_B_CLK_negedge_negedge,
	 HoldHigh		=> thold_B_CLK_posedge_negedge,
	 HoldLow		=> thold_B_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFME2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFME2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFME2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFME2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFME2B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S_CLK_negedge or 
	 Tviol_A_CLK_negedge or 
	 Tviol_B_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, NET_0_2, E_delayed, PRE_ipd, CLK_delayed));
   Q_zd := Violation XOR Q_zd;
         --- now combinatorial logic input to the DFF 
   NET_0_2 :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFME2B_VITAL of DFME2B is
   for VITAL_ACT
   end for;
end CFG_DFME2B_VITAL;



 ---- CELL DFME3A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFME3A is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFME3A :  entity is TRUE;
 end DFME3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFME3A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (S_ipd, S, tipd_S);
	  VitalWireDelay (A_ipd, A, tipd_A);
	  VitalWireDelay (B_ipd, B, tipd_B);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (S_ipd, A_ipd, B_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_S_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_S_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_A_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_A_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_B_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_CLK_posedge,
	 TimingData		=> Tmkr_S_CLK_posedge,
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_CLK_posedge_posedge,
	 SetupLow		=> tsetup_S_CLK_negedge_posedge,
	 HoldHigh		=> thold_S_CLK_posedge_posedge,
	 HoldLow		=> thold_S_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFME3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_CLK_posedge,
	 TimingData		=> Tmkr_A_CLK_posedge,
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_CLK_posedge_posedge,
	 SetupLow		=> tsetup_A_CLK_negedge_posedge,
	 HoldHigh		=> thold_A_CLK_posedge_posedge,
	 HoldLow		=> thold_A_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFME3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_CLK_posedge,
	 TimingData		=> Tmkr_B_CLK_posedge,
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_CLK_posedge_posedge,
	 SetupLow		=> tsetup_B_CLK_negedge_posedge,
	 HoldHigh		=> thold_B_CLK_posedge_posedge,
	 HoldLow		=> thold_B_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFME3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFME3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFME3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFME3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFME3A",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S_CLK_posedge or 
	 Tviol_A_CLK_posedge or 
	 Tviol_B_CLK_posedge or 
	 Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, NET_0_2, E_delayed, '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
         --- now combinatorial logic input to the DFF 
   NET_0_2 :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFME3A_VITAL of DFME3A is
   for VITAL_ACT
   end for;
end CFG_DFME3A_VITAL;



 ---- CELL DFME3B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFME3B is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFME3B :  entity is TRUE;
 end DFME3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFME3B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (S_ipd, S, tipd_S);
	  VitalWireDelay (A_ipd, A, tipd_A);
	  VitalWireDelay (B_ipd, B, tipd_B);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (S_ipd, A_ipd, B_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_S_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_S_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_A_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_A_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_B_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_CLK_negedge, 
	 TimingData		=> Tmkr_S_CLK_negedge, 
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_CLK_posedge_negedge,
	 SetupLow		=> tsetup_S_CLK_negedge_negedge,
	 HoldHigh		=> thold_S_CLK_posedge_negedge,
	 HoldLow		=> thold_S_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFME3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_CLK_negedge, 
	 TimingData		=> Tmkr_A_CLK_negedge, 
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_CLK_posedge_negedge,
	 SetupLow		=> tsetup_A_CLK_negedge_negedge,
	 HoldHigh		=> thold_A_CLK_posedge_negedge,
	 HoldLow		=> thold_A_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFME3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_CLK_negedge, 
	 TimingData		=> Tmkr_B_CLK_negedge, 
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_CLK_posedge_negedge,
	 SetupLow		=> tsetup_B_CLK_negedge_negedge,
	 HoldHigh		=> thold_B_CLK_posedge_negedge,
	 HoldLow		=> thold_B_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFME3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFME3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFME3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFME3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFME3B",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S_CLK_negedge or 
	 Tviol_A_CLK_negedge or 
	 Tviol_B_CLK_negedge or 
	 Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, Q_zd, NET_0_2, E_delayed, '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
         --- now combinatorial logic input to the DFF 
   NET_0_2 :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFME3B_VITAL of DFME3B is
   for VITAL_ACT
   end for;
end CFG_DFME3B_VITAL;



 ---- CELL DFMEG ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFMEG is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFMEG :  entity is TRUE;
 end DFMEG;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFMEG is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (S_ipd, S, tipd_S);
	  VitalWireDelay (A_ipd, A, tipd_A);
	  VitalWireDelay (B_ipd, B, tipd_B);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (S_ipd, A_ipd, B_ipd, PRE_ipd,CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_S_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_S_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_A_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_A_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_B_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_CLK_posedge,
	 TimingData		=> Tmkr_S_CLK_posedge,
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_CLK_posedge_posedge,
	 SetupLow		=> tsetup_S_CLK_negedge_posedge,
	 HoldHigh		=> thold_S_CLK_posedge_posedge,
	 HoldLow		=> thold_S_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFMEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_CLK_posedge,
	 TimingData		=> Tmkr_A_CLK_posedge,
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_CLK_posedge_posedge,
	 SetupLow		=> tsetup_A_CLK_negedge_posedge,
	 HoldHigh		=> thold_A_CLK_posedge_posedge,
	 HoldLow		=> thold_A_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFMEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_CLK_posedge,
	 TimingData		=> Tmkr_B_CLK_posedge,
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_CLK_posedge_posedge,
	 SetupLow		=> tsetup_B_CLK_negedge_posedge,
	 HoldHigh		=> thold_B_CLK_posedge_posedge,
	 HoldLow		=> thold_B_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFMEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFMEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFMEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFMEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFMEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFMEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DFMEG",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S_CLK_posedge or 
	 Tviol_A_CLK_posedge or 
	 Tviol_B_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, NET_0_2, E_delayed, PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;
         --- now combinatorial logic input to the DFF 
   NET_0_2 :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFMEG_VITAL of DFMEG is
   for VITAL_ACT
   end for;
end CFG_DFMEG_VITAL;



 ---- CELL DFMEH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFMEH is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFMEH :  entity is TRUE;
 end DFMEH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFMEH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (S_ipd, S, tipd_S);
	  VitalWireDelay (A_ipd, A, tipd_A);
	  VitalWireDelay (B_ipd, B, tipd_B);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (S_ipd, A_ipd, B_ipd, PRE_ipd,CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_S_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_S_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_A_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_A_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_B_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_CLK_negedge, 
	 TimingData		=> Tmkr_S_CLK_negedge, 
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_CLK_posedge_negedge,
	 SetupLow		=> tsetup_S_CLK_negedge_negedge,
	 HoldHigh		=> thold_S_CLK_posedge_negedge,
	 HoldLow		=> thold_S_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFMEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_CLK_negedge, 
	 TimingData		=> Tmkr_A_CLK_negedge, 
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_CLK_posedge_negedge,
	 SetupLow		=> tsetup_A_CLK_negedge_negedge,
	 HoldHigh		=> thold_A_CLK_posedge_negedge,
	 HoldLow		=> thold_A_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFMEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_CLK_negedge, 
	 TimingData		=> Tmkr_B_CLK_negedge, 
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_CLK_posedge_negedge,
	 SetupLow		=> tsetup_B_CLK_negedge_negedge,
	 HoldHigh		=> thold_B_CLK_posedge_negedge,
	 HoldLow		=> thold_B_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFMEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (CLR_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFMEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFMEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd) AND (NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFMEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFMEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFMEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DFMEH",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S_CLK_negedge or 
	 Tviol_A_CLK_negedge or 
	 Tviol_B_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, Q_zd, NET_0_2, E_delayed, PRE_ipd, CLK_delayed));
   Q_zd := Violation XOR Q_zd;
         --- now combinatorial logic input to the DFF 
   NET_0_2 :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFMEH_VITAL of DFMEH is
   for VITAL_ACT
   end for;
end CFG_DFMEH_VITAL;



 ---- CELL DFMPCA ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFMPCA is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFMPCA :  entity is TRUE;
 end DFMPCA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFMPCA is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (S_ipd, S, tipd_S);
	  VitalWireDelay (A_ipd, A, tipd_A);
	  VitalWireDelay (B_ipd, B, tipd_B);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (S_ipd, A_ipd, B_ipd, PRE_ipd,CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_S_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_S_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_A_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_A_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_B_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_CLK_posedge,
	 TimingData		=> Tmkr_S_CLK_posedge,
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_CLK_posedge_posedge,
	 SetupLow		=> tsetup_S_CLK_negedge_posedge,
	 HoldHigh		=> thold_S_CLK_posedge_posedge,
	 HoldLow		=> thold_S_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFMPCA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_CLK_posedge,
	 TimingData		=> Tmkr_A_CLK_posedge,
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_CLK_posedge_posedge,
	 SetupLow		=> tsetup_A_CLK_negedge_posedge,
	 HoldHigh		=> thold_A_CLK_posedge_posedge,
	 HoldLow		=> thold_A_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFMPCA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_CLK_posedge,
	 TimingData		=> Tmkr_B_CLK_posedge,
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_CLK_posedge_posedge,
	 SetupLow		=> tsetup_B_CLK_negedge_posedge,
	 HoldHigh		=> thold_B_CLK_posedge_posedge,
	 HoldLow		=> thold_B_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFMPCA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFMPCA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFMPCA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFMPCA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFMPCA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DFMPCA",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S_CLK_posedge or 
	 Tviol_A_CLK_posedge or 
	 Tviol_B_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, NET_0_2, '0', PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;
         --- now combinatorial logic input to the DFF 
   NET_0_2 :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFMPCA_VITAL of DFMPCA is
   for VITAL_ACT
   end for;
end CFG_DFMPCA_VITAL;



 ---- CELL DFMPCB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFMPCB is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_S_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_A_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_B_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		S		:  in    STD_ULOGIC;
		A		:  in    STD_ULOGIC;
		B		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFMPCB :  entity is TRUE;
 end DFMPCB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of DFMPCB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (S_ipd, S, tipd_S);
	  VitalWireDelay (A_ipd, A, tipd_A);
	  VitalWireDelay (B_ipd, B, tipd_B);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (S_ipd, A_ipd, B_ipd, PRE_ipd,CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_S_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_S_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_A_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_A_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_B_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_B_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE NET_0_2	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_S_CLK_negedge, 
	 TimingData		=> Tmkr_S_CLK_negedge, 
	 TestSignal		=> S_ipd,
	 TestSignalName		=> "S",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_S_CLK_posedge_negedge,
	 SetupLow		=> tsetup_S_CLK_negedge_negedge,
	 HoldHigh		=> thold_S_CLK_posedge_negedge,
	 HoldLow		=> thold_S_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFMPCB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_A_CLK_negedge, 
	 TimingData		=> Tmkr_A_CLK_negedge, 
	 TestSignal		=> A_ipd,
	 TestSignalName		=> "A",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_A_CLK_posedge_negedge,
	 SetupLow		=> tsetup_A_CLK_negedge_negedge,
	 HoldHigh		=> thold_A_CLK_posedge_negedge,
	 HoldLow		=> thold_A_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFMPCB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_B_CLK_negedge, 
	 TimingData		=> Tmkr_B_CLK_negedge, 
	 TestSignal		=> B_ipd,
	 TestSignalName		=> "B",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_B_CLK_posedge_negedge,
	 SetupLow		=> tsetup_B_CLK_negedge_negedge,
	 HoldHigh		=> thold_B_CLK_posedge_negedge,
	 HoldLow		=> thold_B_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFMPCB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((CLR_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFMPCB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((PRE_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFMPCB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) AND (CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFMPCB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFMPCB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 		TO_X01(CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DFMPCB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_S_CLK_negedge or 
	 Tviol_A_CLK_negedge or 
	 Tviol_B_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, Q_zd, NET_0_2, '0', PRE_ipd, CLK_delayed));
   Q_zd := Violation XOR Q_zd;
         --- now combinatorial logic input to the DFF 
   NET_0_2 :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFMPCB_VITAL of DFMPCB is
   for VITAL_ACT
   end for;
end CFG_DFMPCB_VITAL;



 ---- CELL HCLKMUX ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity HCLKMUX is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		
                tpw_A_posedge   : VitalDelayType :=  0.000 ns;
                tpw_A_negedge   : VitalDelayType :=  0.000 ns;
                tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of HCLKMUX :  entity is TRUE;
 end HCLKMUX;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of HCLKMUX is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- timing check results
	VARIABLE Pviol_A       : STD_ULOGIC := '0';
	VARIABLE PeriodData_A  : VitalPeriodDataType := VitalPeriodDataInit;


	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_A,
              PeriodData     => PeriodData_A,
              TestSignal     => A_ipd,
              TestSignalName => "A",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_A_posedge,
              PulseWidthLow  => tpw_A_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/HCLKMUX",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_HCLKMUX_VITAL of HCLKMUX is 
    for VITAL_ACT
    end for;
 end CFG_HCLKMUX_VITAL;



 ---- CELL IOFIFO_INBUF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOFIFO_INBUF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOFIFO_INBUF :  entity is TRUE;
 end IOFIFO_INBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOFIFO_INBUF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOFIFO_INBUF_VITAL of IOFIFO_INBUF is 
    for VITAL_ACT
    end for;
 end CFG_IOFIFO_INBUF_VITAL;



 ---- CELL IOFIFO_OUTBUF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOFIFO_OUTBUF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOFIFO_OUTBUF :  entity is TRUE;
 end IOFIFO_OUTBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOFIFO_OUTBUF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOFIFO_OUTBUF_VITAL of IOFIFO_OUTBUF is 
    for VITAL_ACT
    end for;
 end CFG_IOFIFO_OUTBUF_VITAL;



 ---- CELL IOOE_FCLK_BUFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOOE_FCLK_BUFF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOOE_FCLK_BUFF :  entity is TRUE;
 end IOOE_FCLK_BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOOE_FCLK_BUFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, CLK_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS YOUT_zd : STD_LOGIC is Results(1);
	ALIAS CLKOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE YOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE CLKOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        YOUT_zd :=TO_X01(A_ipd);
        CLKOUT_zd :=TO_X01(CLK_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => YOUT,
	   GlitchData => YOUT_GlitchData,
	   OutSignalName => "YOUT",
	   OutTemp => YOUT_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_YOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CLKOUT,
	   GlitchData => CLKOUT_GlitchData,
	   OutSignalName => "CLKOUT",
	   OutTemp => CLKOUT_zd,
	   Paths => (
	             0 => (CLK_ipd'last_event,tpd_CLK_CLKOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOOE_FCLK_BUFF_VITAL of IOOE_FCLK_BUFF is 
    for VITAL_ACT
    end for;
 end CFG_IOOE_FCLK_BUFF_VITAL;



 ---- CELL IOOE_OUT_FCLK ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOOE_OUT_FCLK is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOOE_OUT_FCLK :  entity is TRUE;
 end IOOE_OUT_FCLK;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOOE_OUT_FCLK is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, CLK_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS YOUT_zd : STD_LOGIC is Results(1);
	ALIAS CLKOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE YOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE CLKOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        YOUT_zd :=TO_X01(A_ipd);
        CLKOUT_zd :=TO_X01(CLK_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => YOUT,
	   GlitchData => YOUT_GlitchData,
	   OutSignalName => "YOUT",
	   OutTemp => YOUT_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_YOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CLKOUT,
	   GlitchData => CLKOUT_GlitchData,
	   OutSignalName => "CLKOUT",
	   OutTemp => CLKOUT_zd,
	   Paths => (
	             0 => (CLK_ipd'last_event,tpd_CLK_CLKOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOOE_OUT_FCLK_VITAL of IOOE_OUT_FCLK is 
    for VITAL_ACT
    end for;
 end CFG_IOOE_OUT_FCLK_VITAL;



 ---- CELL IOOE_OUT_FCLK_CLR_EN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOOE_OUT_FCLK_CLR_EN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_ENOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_CLROUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		CLR		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC;
		ENOUT		: out    STD_ULOGIC;
		CLROUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOOE_OUT_FCLK_CLR_EN :  entity is TRUE;
 end IOOE_OUT_FCLK_CLR_EN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOOE_OUT_FCLK_CLR_EN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
	VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, CLR_ipd, CLK_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 4)  := (others => 'X');
	ALIAS YOUT_zd : STD_LOGIC is Results(1);
	ALIAS ENOUT_zd : STD_LOGIC is Results(2);
	ALIAS CLROUT_zd : STD_LOGIC is Results(3);
	ALIAS CLKOUT_zd : STD_LOGIC is Results(4);

	-- output glitch detection variables
	VARIABLE YOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE ENOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE CLROUT_GlitchData  : VitalGlitchDataType;
	VARIABLE CLKOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        YOUT_zd :=TO_X01(A_ipd);
        ENOUT_zd :=TO_X01(EN_ipd);
        CLROUT_zd :=TO_X01(CLR_ipd);
        CLKOUT_zd :=TO_X01(CLK_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => YOUT,
	   GlitchData => YOUT_GlitchData,
	   OutSignalName => "YOUT",
	   OutTemp => YOUT_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_YOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => ENOUT,
	   GlitchData => ENOUT_GlitchData,
	   OutSignalName => "ENOUT",
	   OutTemp => ENOUT_zd,
	   Paths => (
	             0 => (EN_ipd'last_event,tpd_EN_ENOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CLROUT,
	   GlitchData => CLROUT_GlitchData,
	   OutSignalName => "CLROUT",
	   OutTemp => CLROUT_zd,
	   Paths => (
	             0 => (CLR_ipd'last_event,tpd_CLR_CLROUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CLKOUT,
	   GlitchData => CLKOUT_GlitchData,
	   OutSignalName => "CLKOUT",
	   OutTemp => CLKOUT_zd,
	   Paths => (
	             0 => (CLK_ipd'last_event,tpd_CLK_CLKOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOOE_OUT_FCLK_CLR_EN_VITAL of IOOE_OUT_FCLK_CLR_EN is 
    for VITAL_ACT
    end for;
 end CFG_IOOE_OUT_FCLK_CLR_EN_VITAL;



 ---- CELL IOOE_OUT_RCLK ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOOE_OUT_RCLK is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOOE_OUT_RCLK :  entity is TRUE;
 end IOOE_OUT_RCLK;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOOE_OUT_RCLK is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, CLK_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS YOUT_zd : STD_LOGIC is Results(1);
	ALIAS CLKOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE YOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE CLKOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        YOUT_zd :=TO_X01(A_ipd);
        CLKOUT_zd :=TO_X01(CLK_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => YOUT,
	   GlitchData => YOUT_GlitchData,
	   OutSignalName => "YOUT",
	   OutTemp => YOUT_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_YOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CLKOUT,
	   GlitchData => CLKOUT_GlitchData,
	   OutSignalName => "CLKOUT",
	   OutTemp => CLKOUT_zd,
	   Paths => (
	             0 => (CLK_ipd'last_event,tpd_CLK_CLKOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOOE_OUT_RCLK_VITAL of IOOE_OUT_RCLK is 
    for VITAL_ACT
    end for;
 end CFG_IOOE_OUT_RCLK_VITAL;



 ---- CELL IOOE_OUT_RCLK_CLR_EN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOOE_OUT_RCLK_CLR_EN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_YOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_ENOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_CLROUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		CLR		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		YOUT		: out    STD_ULOGIC;
		ENOUT		: out    STD_ULOGIC;
		CLROUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOOE_OUT_RCLK_CLR_EN :  entity is TRUE;
 end IOOE_OUT_RCLK_CLR_EN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOOE_OUT_RCLK_CLR_EN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
	VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, CLR_ipd, CLK_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 4)  := (others => 'X');
	ALIAS YOUT_zd : STD_LOGIC is Results(1);
	ALIAS ENOUT_zd : STD_LOGIC is Results(2);
	ALIAS CLROUT_zd : STD_LOGIC is Results(3);
	ALIAS CLKOUT_zd : STD_LOGIC is Results(4);

	-- output glitch detection variables
	VARIABLE YOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE ENOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE CLROUT_GlitchData  : VitalGlitchDataType;
	VARIABLE CLKOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        YOUT_zd :=TO_X01(A_ipd);
        ENOUT_zd :=TO_X01(EN_ipd);
        CLROUT_zd :=TO_X01(CLR_ipd);
        CLKOUT_zd :=TO_X01(CLK_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => YOUT,
	   GlitchData => YOUT_GlitchData,
	   OutSignalName => "YOUT",
	   OutTemp => YOUT_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_YOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => ENOUT,
	   GlitchData => ENOUT_GlitchData,
	   OutSignalName => "ENOUT",
	   OutTemp => ENOUT_zd,
	   Paths => (
	             0 => (EN_ipd'last_event,tpd_EN_ENOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CLROUT,
	   GlitchData => CLROUT_GlitchData,
	   OutSignalName => "CLROUT",
	   OutTemp => CLROUT_zd,
	   Paths => (
	             0 => (CLR_ipd'last_event,tpd_CLR_CLROUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CLKOUT,
	   GlitchData => CLKOUT_GlitchData,
	   OutSignalName => "CLKOUT",
	   OutTemp => CLKOUT_zd,
	   Paths => (
	             0 => (CLK_ipd'last_event,tpd_CLK_CLKOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOOE_OUT_RCLK_CLR_EN_VITAL of IOOE_OUT_RCLK_CLR_EN is 
    for VITAL_ACT
    end for;
 end CFG_IOOE_OUT_RCLK_CLR_EN_VITAL;



 ---- CELL IOOE_FCLK_CLR_EN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOOE_FCLK_CLR_EN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_EN_ENOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_CLROUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_CLKOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		EN		: in    STD_ULOGIC;
		CLR		: in    STD_ULOGIC;
		CLK		: in    STD_ULOGIC;
		ENOUT		: out    STD_ULOGIC;
		CLROUT		: out    STD_ULOGIC;
		CLKOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOOE_FCLK_CLR_EN :  entity is TRUE;
 end IOOE_FCLK_CLR_EN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOOE_FCLK_CLR_EN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
	VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (EN_ipd, CLR_ipd, CLK_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
	ALIAS ENOUT_zd : STD_LOGIC is Results(1);
	ALIAS CLROUT_zd : STD_LOGIC is Results(2);
	ALIAS CLKOUT_zd : STD_LOGIC is Results(3);

	-- output glitch detection variables
	VARIABLE ENOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE CLROUT_GlitchData  : VitalGlitchDataType;
	VARIABLE CLKOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        ENOUT_zd :=TO_X01(EN_ipd);
        CLROUT_zd :=TO_X01(CLR_ipd);
        CLKOUT_zd :=TO_X01(CLK_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => ENOUT,
	   GlitchData => ENOUT_GlitchData,
	   OutSignalName => "ENOUT",
	   OutTemp => ENOUT_zd,
	   Paths => (
	             0 => (EN_ipd'last_event,tpd_EN_ENOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CLROUT,
	   GlitchData => CLROUT_GlitchData,
	   OutSignalName => "CLROUT",
	   OutTemp => CLROUT_zd,
	   Paths => (
	             0 => (CLR_ipd'last_event,tpd_CLR_CLROUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => CLKOUT,
	   GlitchData => CLKOUT_GlitchData,
	   OutSignalName => "CLKOUT",
	   OutTemp => CLKOUT_zd,
	   Paths => (
	             0 => (CLK_ipd'last_event,tpd_CLK_CLKOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOOE_FCLK_CLR_EN_VITAL of IOOE_FCLK_CLR_EN is 
    for VITAL_ACT
    end for;
 end CFG_IOOE_FCLK_CLR_EN_VITAL;



 ---- CELL IOPAD_IN_U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_IN_U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_PAD_posedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge           : VitalDelayType := 0.000 ns;
                tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPAD_IN_U :  entity is TRUE;
 end IOPAD_IN_U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOPAD_IN_U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- timing check results
	VARIABLE Pviol_PAD       : STD_ULOGIC := '0';
	VARIABLE PeriodData_PAD  : VitalPeriodDataType := VitalPeriodDataInit;

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_IN_U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOPAD_IN_U_VITAL of IOPAD_IN_U is 
    for VITAL_ACT
    end for;
 end CFG_IOPAD_IN_U_VITAL;



 ---- CELL IOPAD_IN_D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_IN_D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		
                tpw_PAD_posedge 		: VitalDelayType := 0.000 ns;
                tpw_PAD_negedge           : VitalDelayType := 0.000 ns;
                tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPAD_IN_D :  entity is TRUE;
 end IOPAD_IN_D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOPAD_IN_D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	
        -- timing check results
	VARIABLE Pviol_PAD       : STD_ULOGIC := '0';
	VARIABLE PeriodData_PAD  : VitalPeriodDataType := VitalPeriodDataInit;

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_IN_D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','L'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOPAD_IN_D_VITAL of IOPAD_IN_D is 
    for VITAL_ACT
    end for;
 end CFG_IOPAD_IN_D_VITAL;



 ---- CELL IOPAD_TRI_U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_TRI_U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge 	    : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                
                tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPAD_TRI_U :  entity is TRUE;
 end IOPAD_TRI_U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOPAD_TRI_U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- timing check results
	VARIABLE Pviol_D       : STD_ULOGIC := '0';
        VARIABLE PeriodData_D : VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_E       : STD_ULOGIC := '0';
	VARIABLE PeriodData_E  : VitalPeriodDataType := VitalPeriodDataInit;

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_TRI_U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );
           
           VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_TRI_U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_IOPAD_TRI_U_VITAL of IOPAD_TRI_U is 
    for VITAL_ACT
    end for;
 end CFG_IOPAD_TRI_U_VITAL;



 ---- CELL IOPAD_TRI_D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_TRI_D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		
                tpw_D_posedge   : VitalDelayType := 0.000 ns;
                tpw_D_negedge   : VitalDelayType := 0.000 ns;
                tpw_E_posedge   : VitalDelayType := 0.000 ns;
                tpw_E_negedge   : VitalDelayType := 0.000 ns; 

                tpd_D_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPAD_TRI_D :  entity is TRUE;
 end IOPAD_TRI_D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOPAD_TRI_D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- timing check results
	VARIABLE Pviol_E       : STD_ULOGIC := '0';
	VARIABLE PeriodData_E  : VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_D       : STD_ULOGIC := '0';
	VARIABLE PeriodData_D  : VitalPeriodDataType := VitalPeriodDataInit;

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_TRI_D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_TRI_D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_IOPAD_TRI_D_VITAL of IOPAD_TRI_D is 
    for VITAL_ACT
    end for;
 end CFG_IOPAD_TRI_D_VITAL;



 ---- CELL IOPAD_BI_U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_BI_U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
	
		tpw_E_posedge       : VitalDelayType := 0.000 ns;
                tpw_E_negedge 	    : VitalDelayType := 0.000 ns;
		tpw_D_posedge       : VitalDelayType := 0.000 ns;
                tpw_D_negedge 	    : VitalDelayType := 0.000 ns;
		tpw_PAD_posedge     : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge     : VitalDelayType := 0.000 ns;

             	tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		
                tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPAD_BI_U :  entity is TRUE;
 end IOPAD_BI_U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOPAD_BI_U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- timing check results
	VARIABLE Pviol_D       : STD_ULOGIC := '0';
	VARIABLE PeriodData_D  : VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_E       : STD_ULOGIC := '0';
	VARIABLE PeriodData_E  : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE PViol_PAD     : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD :VitalPeriodDataType := VitalPeriodDataInit;

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        if ( TimingChecksOn) then
        
        
            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI_U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );
            
             VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI_U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

             VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI_U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

           end if;
	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOPAD_BI_U_VITAL of IOPAD_BI_U is 
    for VITAL_ACT
    end for;
 end CFG_IOPAD_BI_U_VITAL;



 ---- CELL IOPAD_BI_D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_BI_D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_E_posedge   : VitalDelayType := 0.000 ns;
                tpw_E_negedge 	: VitalDelayType := 0.000 ns;
		tpw_D_posedge   : VitalDelayType := 0.000 ns;
                tpw_D_negedge 	: VitalDelayType := 0.000 ns;
		tpw_PAD_posedge : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge : VitalDelayType := 0.000 ns;		

                tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
	        tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
	        tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPAD_BI_D :  entity is TRUE;
 end IOPAD_BI_D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of IOPAD_BI_D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

        -- timing check results
	VARIABLE Pviol_D       : STD_ULOGIC := '0';
	VARIABLE PeriodData_D  : VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_E       : STD_ULOGIC := '0';
	VARIABLE PeriodData_E  : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE PViol_PAD     : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD :VitalPeriodDataType := VitalPeriodDataInit;


	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin
        
        if ( TimingChecksOn ) then
        
            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI_D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );
 
            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI_D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            ); 
         
            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI_D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );
           end if;
	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

end process;

end VITAL_ACT;

 configuration CFG_IOPAD_BI_D_VITAL of IOPAD_BI_D is 
    for VITAL_ACT
    end for;
 end CFG_IOPAD_BI_D_VITAL;



 ---- CELL RCLKMUX ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity RCLKMUX is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		
                tpw_A_posedge   : VitalDelayType := 0.000 ns;
                tpw_A_negedge   : VitalDelayType := 0.000 ns;   
                tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of RCLKMUX :  entity is TRUE;
 end RCLKMUX;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of RCLKMUX is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- timing check results
	VARIABLE Pviol_A       : STD_ULOGIC := '0';
	VARIABLE PeriodData_A  : VitalPeriodDataType := VitalPeriodDataInit;


	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_A,
              PeriodData     => PeriodData_A,
              TestSignal     => A_ipd,
              TestSignalName => "A",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_A_posedge,
              PulseWidthLow  => tpw_A_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/RCLKMUX",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_RCLKMUX_VITAL of RCLKMUX is 
    for VITAL_ACT
    end for;
 end CFG_RCLKMUX_VITAL;



 ---- CELL TRIBUFF_HSTL_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_HSTL_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_HSTL_I :  entity is TRUE;
 end TRIBUFF_HSTL_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_HSTL_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_HSTL_I_VITAL of TRIBUFF_HSTL_I is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_HSTL_I_VITAL;



 ---- CELL TRIBUFF_SSTL3_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_SSTL3_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_SSTL3_I :  entity is TRUE;
 end TRIBUFF_SSTL3_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_SSTL3_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_SSTL3_I_VITAL of TRIBUFF_SSTL3_I is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_SSTL3_I_VITAL;



 ---- CELL TRIBUFF_SSTL3_II ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_SSTL3_II is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_SSTL3_II :  entity is TRUE;
 end TRIBUFF_SSTL3_II;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_SSTL3_II is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_SSTL3_II_VITAL of TRIBUFF_SSTL3_II is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_SSTL3_II_VITAL;



 ---- CELL TRIBUFF_SSTL2_I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_SSTL2_I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_SSTL2_I :  entity is TRUE;
 end TRIBUFF_SSTL2_I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_SSTL2_I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_SSTL2_I_VITAL of TRIBUFF_SSTL2_I is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_SSTL2_I_VITAL;



 ---- CELL TRIBUFF_SSTL2_II ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_SSTL2_II is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_SSTL2_II :  entity is TRUE;
 end TRIBUFF_SSTL2_II;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_SSTL2_II is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event,VitalExtendToFillDelay(tpd_E_PAD), true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_SSTL2_II_VITAL of TRIBUFF_SSTL2_II is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_SSTL2_II_VITAL;

-----------------------------------------------------------------
--
--  Actel IOFIFO_INFIFO VHDL behavioral model
--  64 X 1 I/O FIFO with rising write clock, rising read clock,
--  and active low WENB, RENB, and CLRB.
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - 9/25/00 - Dale Walter - Prototype version.
-- 2.0 - 9/27/02 - Krupa Singampalli - New Timing Arcs
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity IOFIFO_INFIFO is
  GENERIC (
        tipd_D       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_CLRB      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_Q   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLRB_Q    : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tsetup_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_negedge_posedge     :   VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLRB_WCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLRB_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True

        );
  PORT (
        D     : IN STD_ULOGIC ;
        WENB     : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RENB     : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        CLRB    : IN STD_ULOGIC ;
        Q     : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of IOFIFO_INFIFO : entity is FALSE;
  
end IOFIFO_INFIFO;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of IOFIFO_INFIFO is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal D_ipd   : std_ulogic := 'X';
  signal WENB_ipd   : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  signal RENB_ipd   : std_ulogic := 'X';
  signal RCLK_ipd : std_ulogic := 'X';
  signal CLRB_ipd  : std_ulogic := 'X';
  type MEM is array(0 to 63) of std_ulogic;
  --signal DUAL_PORT_RAM : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (D_ipd, D, VitalExtendToFillDelay(tipd_D));
    VitalWireDelay (WENB_ipd, WENB, VitalExtendToFillDelay(tipd_WENB));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (RENB_ipd, RENB, VitalExtendToFillDelay(tipd_RENB));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
    VitalWireDelay (CLRB_ipd, CLRB, VitalExtendToFillDelay(tipd_CLRB));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (D_ipd, WENB_ipd, WCLK_ipd, RENB_ipd, RCLK_ipd, CLRB_ipd)

      --  Memory
     variable DUAL_PORT_RAM : MEM;

     --  Read Timing Check Results
     variable Tviol_RENB_RCLK_posedge : X01 := '0';
     variable TmDt_RENB_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_D_WCLK_posedge : X01 := '0';
     variable TmDt_D_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WENB_WCLK_posedge : X01 := '0';
     variable TmDt_WENB_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  CLRB Timing Check Results
     variable Tviol_CLRB_RCLK_posedge : X01 := '0';
     variable TmDt_CLRB_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_CLRB_WCLK_posedge : X01 := '0';
     variable TmDt_CLRB_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_CLRB : X01 := '0';
     variable PeriodData_CLRB : VitalPeriodDataType := VitalPeriodDataInit;

     --  Functional Results
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT : SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1; -- free running counter
     variable RADDR : integer := -1; -- free running counter
     variable Q_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable Q_GlitchData : VitalGlitchDataType;

     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable RENB_delayed : std_ulogic := 'X';
     variable RENB_previous : std_ulogic := 'X';
     variable WENB_delayed : std_ulogic := 'X';
     variable WENB_previous : std_ulogic := 'X';
     variable D_delayed : std_ulogic := 'X';

  begin  --  process VITALBehavior 

    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RENB before RCLK rising
      --   Hold  RENB after RCLK rising

      VitalSetupHoldCheck ( Tviol_RENB_RCLK_posedge,
                            TmDt_RENB_RCLK_posedge,
                            RENB_ipd, "RENB",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RENB_RCLK_posedge_posedge,
			    tsetup_RENB_RCLK_negedge_posedge,
                            thold_RENB_RCLK_posedge_posedge,
                            thold_RENB_RCLK_negedge_posedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            '/',
                            InstancePath & "/IOFIFO_INFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            InstancePath & "/IOFIFO_INFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup D high or low before WCLK rising
      --   Hold  D high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_D_WCLK_posedge,
                            TmDt_D_WCLK_posedge,
                            D_ipd, "D",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_D_WCLK_posedge_posedge,
                            tsetup_D_WCLK_negedge_posedge,
                            thold_D_WCLK_posedge_posedge,
                            thold_D_WCLK_negedge_posedge,
                            TO_X01((CLRB_ipd) AND (NOT WENB_ipd)) /= '0',
                            '/',
                            InstancePath & "/IOFIFO_INFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup WENB high before WCLK rising
      --   Hold  WENB high after WCLK rising

      VitalSetupHoldCheck ( Tviol_WENB_WCLK_posedge,
                            TmDt_WENB_WCLK_posedge,
                            WENB_ipd, "WENB",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WENB_WCLK_posedge_posedge,
                            tsetup_WENB_WCLK_negedge_posedge,
                            thold_WENB_WCLK_posedge_posedge,
                            thold_WENB_WCLK_negedge_posedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            '/',
                            InstancePath & "/IOFIFO_INFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            InstancePath & "/IOFIFO_INFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup CLRB high before WCLK rising
      --   Hold  CLRB high after WCLK rising

         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLRB_RCLK_posedge,
          TimingData              => TmDt_CLRB_RCLK_posedge,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          RefSignal               => RCLK_ipd,
          RefSignalName           => "RCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLRB_RCLK_posedge_posedge,
          Removal                 => thold_CLRB_RCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TO_X01(NOT RENB_ipd) /='0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IOFIFO_INFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLRB_WCLK_posedge,
          TimingData              => TmDt_CLRB_WCLK_posedge,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          RefSignal               => RCLK_ipd,
          RefSignalName           => "WCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLRB_WCLK_posedge_posedge,
          Removal                 => thold_CLRB_WCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TO_X01(NOT WENB_ipd) /='0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IOFIFO_INFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLRB,
          PeriodData              => PeriodData_CLRB,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLRB_negedge,
          CheckEnabled            => TRUE,
          HeaderMsg               => InstancePath &"/IOFIFO_INFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);


    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################

      


      if (TO_X01(CLRB_ipd)='X') then
        assert false
        report ": CLRB unknown"
        severity Error;
      elsif (TO_X01(CLRB_ipd)='0') then
        WADDR := 0;
      else
        if (TO_X01(WCLK_ipd)='X') then
          if ((TO_X01(WENB_delayed) /= '1')) then
            if (TO_X01(WCLK_previous) /= 'X') then
              assert false
              report ": WCLK went unknown"
              severity Error;
            end if;
          end if;
        elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='1')) then
          case (TO_X01(WENB_delayed)) is
            when '1' =>
              null;
            when '0' =>
              -- Write first, then increment WADDR
              if (WADDR < 64) then
                DUAL_PORT_RAM(WADDR) := D_delayed ;
                WADDR := WADDR + 1;
              else
                assert false
                report ": Write failed - FIFO full."
                severity Error;
              end if;
            when others =>
              if (TO_X01(WENB_previous) = 'X') then
                assert false
                report ": WENB went unknown"
                severity Error;
              end if;
          end case;
        end if;
      end if;



      -- #########################################################
      -- # Read Functional Section
      -- #########################################################
     
      if (TO_X01(CLRB_ipd)='1') then
        if (TO_X01(RCLK_ipd) = 'X') then
          if ((TO_X01(RENB_delayed) /= '1')) then
            Q_zd := 'X';
            if (TO_X01(RCLK_previous) /= 'X') then
              assert false
              report ": RCLK went unknown"
              severity Warning;
            end if;
          end if;
        elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '1')) then
          case (TO_X01(RENB_delayed)) is
            when '1' =>
              null;
            when '0' =>
              -- Always read from address 0, then shift memory contents down.
              if (WADDR > 0) then -- 0 means memory empty
                Q_zd := DUAL_PORT_RAM(0);
                WADDR := WADDR - 1;
                if (WADDR > 0) then -- move everything down one slot
                  for I in 0 to (WADDR - 1) loop
                    DUAL_PORT_RAM(I) := DUAL_PORT_RAM(I + 1);
                  end loop;
                end if;
              else
                Q_zd := 'X';
                assert false
                report ": Read failed - FIFO empty."
                severity Error;
              end if;
            when others =>
              Q_zd := 'X';
              if (TO_X01(RENB_delayed) = 'X') and (TO_X01(RENB_previous) /= 'X') then
                assert false
                report ": RENB went unknown"
                severity Warning;
                RENB_previous := RENB_delayed;
              end if;
          end case;
        end if;
      end if;

      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      if WENB_ipd'event then
        WENB_previous := WENB_delayed;
        WENB_delayed := WENB_ipd;
      end if;
      if RENB_ipd'event then
        RENB_previous := RENB_delayed;
        RENB_delayed := RENB_ipd;
      end if;
      D_delayed := D_ipd;


    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => Q,
	GlitchData => Q_GlitchData,
	OutSignalName => "Q",
	OutTemp => Q_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_Q), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => Xon,
	MsgOn => MsgOn,
	MsgSeverity => WARNING
	);

    
  end process VITALBehavior;

end VITAL_ACT;

-----------------------------------------------------------------
-----------------------------------------------------------------
--
--  Actel IOFIFO_OUTFIFO VHDL behavioral model
--  64 X 1 I/O FIFO with rising write clock, rising read clock,
--  and active low WENB, RENB, and CLRB.
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - 9/25/00 - Dale Walter - Prototype version.
-- 2.0 - 9/27/02 - Krupa Singampalli - New Timing Arcs
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity IOFIFO_OUTFIFO is
  GENERIC (
        tipd_D       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_CLRB      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_Q   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLRB_Q    : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tsetup_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_negedge_posedge     :   VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLRB_WCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLRB_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True

        );
  PORT (
        D     : IN STD_ULOGIC ;
        WENB     : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RENB     : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        CLRB    : IN STD_ULOGIC ;
        Q     : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of IOFIFO_OUTFIFO : entity is FALSE;
  
end IOFIFO_OUTFIFO;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of IOFIFO_OUTFIFO is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal D_ipd   : std_ulogic := 'X';
  signal WENB_ipd   : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  signal RENB_ipd   : std_ulogic := 'X';
  signal RCLK_ipd : std_ulogic := 'X';
  signal CLRB_ipd  : std_ulogic := 'X';
  type MEM is array(0 to 63) of std_ulogic;
  signal DUAL_PORT_RAM : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (D_ipd, D, VitalExtendToFillDelay(tipd_D));
    VitalWireDelay (WENB_ipd, WENB, VitalExtendToFillDelay(tipd_WENB));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (RENB_ipd, RENB, VitalExtendToFillDelay(tipd_RENB));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
    VitalWireDelay (CLRB_ipd, CLRB, VitalExtendToFillDelay(tipd_CLRB));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (D_ipd, WENB_ipd, WCLK_ipd, RENB_ipd, RCLK_ipd, CLRB_ipd)

     --  Read Timing Check Results
     variable Tviol_RENB_RCLK_posedge : X01 := '0';
     variable TmDt_RENB_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_D_WCLK_posedge : X01 := '0';
     variable TmDt_D_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WENB_WCLK_posedge : X01 := '0';
     variable TmDt_WENB_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  CLRB Timing Check Results
     variable Tviol_CLRB_RCLK_posedge : X01 := '0';
     variable TmDt_CLRB_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_CLRB_WCLK_posedge : X01 := '0';
     variable TmDt_CLRB_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_CLRB : X01 := '0';
     variable PeriodData_CLRB : VitalPeriodDataType := VitalPeriodDataInit;

     --  Functional Results
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT : SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1; -- free running counter
     variable RADDR : integer := -1; -- free running counter
     variable Q_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable Q_GlitchData : VitalGlitchDataType;

     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable RENB_delayed : std_ulogic := 'X';
     variable RENB_previous : std_ulogic := 'X';
     variable WENB_delayed : std_ulogic := 'X';
     variable WENB_previous : std_ulogic := 'X';
     variable D_delayed : std_ulogic := 'X';

  begin  --  process VITALBehavior 

    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RENB before RCLK rising
      --   Hold  RENB after RCLK rising

      VitalSetupHoldCheck ( Tviol_RENB_RCLK_posedge,
                            TmDt_RENB_RCLK_posedge,
                            RENB_ipd, "RENB",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RENB_RCLK_posedge_posedge,
			    tsetup_RENB_RCLK_negedge_posedge,
                            thold_RENB_RCLK_posedge_posedge,
                            thold_RENB_RCLK_negedge_posedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            '/',
                            InstancePath & "/IOFIFO_OUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            InstancePath & "/IOFIFO_OUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup D high or low before WCLK rising
      --   Hold  D high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_D_WCLK_posedge,
                            TmDt_D_WCLK_posedge,
                            D_ipd, "D",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_D_WCLK_posedge_posedge,
                            tsetup_D_WCLK_negedge_posedge,
                            thold_D_WCLK_posedge_posedge,
                            thold_D_WCLK_negedge_posedge,
                            TO_X01((CLRB_ipd) AND (NOT WENB_ipd)) /= '0',
                            '/',
                            InstancePath & "/IOFIFO_OUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup WENB high before WCLK rising
      --   Hold  WENB high after WCLK rising

      VitalSetupHoldCheck ( Tviol_WENB_WCLK_posedge,
                            TmDt_WENB_WCLK_posedge,
                            WENB_ipd, "WENB",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WENB_WCLK_posedge_posedge,
                            tsetup_WENB_WCLK_negedge_posedge,
                            thold_WENB_WCLK_posedge_posedge,
                            thold_WENB_WCLK_negedge_posedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            '/',
                            InstancePath & "/IOFIFO_OUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            InstancePath & "/IOFIFO_OUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup CLRB high before WCLK rising
      --   Hold  CLRB high after WCLK rising

         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLRB_RCLK_posedge,
          TimingData              => TmDt_CLRB_RCLK_posedge,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          RefSignal               => RCLK_ipd,
          RefSignalName           => "RCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLRB_RCLK_posedge_posedge,
          Removal                 => thold_CLRB_RCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TO_X01(NOT RENB_ipd) /='0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IOFIFO_OUTFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLRB_WCLK_posedge,
          TimingData              => TmDt_CLRB_WCLK_posedge,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          RefSignal               => RCLK_ipd,
          RefSignalName           => "WCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLRB_WCLK_posedge_posedge,
          Removal                 => thold_CLRB_WCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TO_X01(NOT WENB_ipd) /='0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IOFIFO_OUTFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLRB,
          PeriodData              => PeriodData_CLRB,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLRB_negedge,
          CheckEnabled            => TRUE,
          HeaderMsg               => InstancePath &"/IOFIFO_OUTFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);


    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################


      if (TO_X01(CLRB_ipd)='X') then
        assert false
        report ": CLRB unknown"
        severity Error;
      elsif (TO_X01(CLRB_ipd)='0') then
        WADDR := -1;
        RADDR := -1;
      else
        if (TO_X01(WCLK_ipd)='X') then
	  if ((TO_X01(WENB_delayed) /= '1')) then
            if (TO_X01(WCLK_previous) /= 'X') then
	      assert false
	      report ": WCLK went unknown"
	      severity Error;
	    end if;
	  end if;
        elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='1')) then
	  case (TO_X01(WENB_delayed)) is
	    when '1' =>
	      null;
	    when '0' =>
              -- Increment WADDR
              WADDR := WADDR + 1;
              if ((RADDR > WADDR) or (WADDR - RADDR > 63)) then
                assert false
                report ": Write failed - FIFO full."
                severity Error;
              else
	        DUAL_PORT_RAM(WADDR mod 64) <= D_delayed ;
              end if;
	    when others =>
              if (TO_X01(WENB_previous) = 'X') then
                assert false
                report ": WENB went unknown"
                severity Error;
              end if;
	  end case;
        end if;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      if (TO_X01(CLRB_ipd)='1') then
        if (TO_X01(RCLK_ipd) = 'X') then
          if ((TO_X01(RENB_delayed) /= '1')) then
	    Q_zd := 'X';
	    if (TO_X01(RCLK_previous) /= 'X') then
	      assert false
	      report ": RCLK went unknown"
	      severity Warning;
	    end if;
	  end if;
        elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '1')) then
	  case (TO_X01(RENB_delayed)) is
	    when '1' =>
	      null;
	    when '0' =>
              -- Increment RADDR
              RADDR := RADDR + 1;
              if ((RADDR > WADDR) or (WADDR - RADDR > 63)) then
                assert false
                report ": Read failed - FIFO empty."
                severity Error;
              else
	        Q_zd := DUAL_PORT_RAM(RADDR mod 64);
              end if;
	    when others =>
	      Q_zd := 'X';
              if (TO_X01(RENB_delayed) = 'X') and (TO_X01(RENB_previous) /= 'X') then
	        assert false
	        report ": RENB went unknown"
	        severity Warning;
                RENB_previous := RENB_delayed;
              end if;
	  end case;
        end if;
      end if;

      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      if WENB_ipd'event then
        WENB_previous := WENB_delayed;
        WENB_delayed := WENB_ipd;
      end if;
      if RENB_ipd'event then
        RENB_previous := RENB_delayed;
        RENB_delayed := RENB_ipd;
      end if;
      D_delayed := D_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => Q,
	GlitchData => Q_GlitchData,
	OutSignalName => "Q",
	OutTemp => Q_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_Q), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => Xon,
	MsgOn => MsgOn,
	MsgSeverity => WARNING
	);

    
  end process VITALBehavior;

end VITAL_ACT;
--
--  Actel BIOFIFO_BIDIRINFIFO VHDL behavioral model
--  64 X 1 I/O FIFO with rising write clock, rising read clock,
--  and active low WENB, RENB, and CLRB.
--  AFL macro containing feed-through.
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - 5/17/02 - Dale Walter - Clone of IOFIFO_INFIFO.
-- 2.0 - 9/27/02 - Krupa Singampalli - New Timing Arcs
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity BIOFIFO_BIDIRINFIFO is
  GENERIC (
        tipd_A       : VitalDelayType01 := (0.00 ns, 0.00 ns);
        tipd_D       : VitalDelayType01 := (0.00 ns, 0.00 ns);
        tipd_WENB       : VitalDelayType01 := (0.00 ns, 0.00 ns);
        tipd_WCLK     : VitalDelayType01 := (0.00 ns, 0.00 ns);
        tipd_RENB       : VitalDelayType01 := (0.00 ns, 0.00 ns);
        tipd_RCLK     : VitalDelayType01 := (0.00 ns, 0.00 ns);
        tipd_CLRB      : VitalDelayType01 := (0.00 ns, 0.00 ns);
        tpd_A_Y   : VitalDelayType01 := (0.1000 ns, 0.1000 ns);
        tpd_RCLK_Q   : VitalDelayType01 := (0.1000 ns, 0.1000 ns);
        tpd_CLRB_Q    : VitalDelayType01 := (0.1000 ns, 0.1000 ns);
        tsetup_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_D_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_negedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLRB_WCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLRB_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True

        );
  PORT (
        A     : IN STD_ULOGIC ;
        D     : IN STD_ULOGIC ;
        WENB     : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RENB     : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        CLRB    : IN STD_ULOGIC ;
        Q     : OUT STD_ULOGIC ;
        Y     : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of BIOFIFO_BIDIRINFIFO : entity is FALSE;
  
end BIOFIFO_BIDIRINFIFO;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of BIOFIFO_BIDIRINFIFO is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal A_ipd   : std_ulogic := 'X';
  signal D_ipd   : std_ulogic := 'X';
  signal WENB_ipd   : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  signal RENB_ipd   : std_ulogic := 'X';
  signal RCLK_ipd : std_ulogic := 'X';
  signal CLRB_ipd  : std_ulogic := 'X';
  type MEM is array(0 to 63) of std_ulogic;
  signal DUAL_PORT_RAM : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (A_ipd, A, VitalExtendToFillDelay(tipd_A));
    VitalWireDelay (D_ipd, D, VitalExtendToFillDelay(tipd_D));
    VitalWireDelay (WENB_ipd, WENB, VitalExtendToFillDelay(tipd_WENB));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (RENB_ipd, RENB, VitalExtendToFillDelay(tipd_RENB));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
    VitalWireDelay (CLRB_ipd, CLRB, VitalExtendToFillDelay(tipd_CLRB));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (A_ipd, D_ipd, WENB_ipd, WCLK_ipd, RENB_ipd, RCLK_ipd, CLRB_ipd)

     --  Read Timing Check Results
     variable Tviol_RENB_RCLK_posedge : X01 := '0';
     variable TmDt_RENB_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_D_WCLK_posedge : X01 := '0';
     variable TmDt_D_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WENB_WCLK_posedge : X01 := '0';
     variable TmDt_WENB_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  CLRB Timing Check Results
     variable Tviol_CLRB_RCLK_posedge : X01 := '0';
     variable TmDt_CLRB_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_CLRB_WCLK_posedge : X01 := '0';
     variable TmDt_CLRB_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_CLRB : X01 := '0';
     variable PeriodData_CLRB : VitalPeriodDataType := VitalPeriodDataInit;

     --  Functional Results
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT : SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1; -- free running counter
     variable RADDR : integer := -1; -- free running counter
     variable Q_zd : std_ulogic;
     variable Y_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable Q_GlitchData : VitalGlitchDataType;
     variable Y_GlitchData : VitalGlitchDataType;

     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable RENB_delayed : std_ulogic := 'X';
     variable RENB_previous : std_ulogic := 'X';
     variable WENB_delayed : std_ulogic := 'X';
     variable WENB_previous : std_ulogic := 'X';
     variable D_delayed : std_ulogic := 'X';

  begin  --  process VITALBehavior 

    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RENB before RCLK rising
      --   Hold  RENB after RCLK rising

      VitalSetupHoldCheck ( Tviol_RENB_RCLK_posedge,
                            TmDt_RENB_RCLK_posedge,
                            RENB_ipd, "RENB",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RENB_RCLK_negedge_posedge,
                            thold_RENB_RCLK_negedge_posedge,
                            tsetup_RENB_RCLK_posedge_posedge,
                            thold_RENB_RCLK_posedge_posedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            '/',
                            InstancePath & "/BIOFIFO_BIDIRINFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            InstancePath & "/BIOFIFO_BIDIRINFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup D high or low before WCLK rising
      --   Hold  D high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_D_WCLK_posedge,
                            TmDt_D_WCLK_posedge,
                            D_ipd, "D",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_D_WCLK_negedge_posedge,
                            thold_D_WCLK_negedge_posedge,
                            tsetup_D_WCLK_posedge_posedge,
                            thold_D_WCLK_posedge_posedge,
                            TO_X01((CLRB_ipd) AND (NOT WENB_ipd)) /= '0',
                            '/',
                            InstancePath & "/BIOFIFO_BIDIRINFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup WENB high before WCLK rising
      --   Hold  WENB high after WCLK rising

      VitalSetupHoldCheck ( Tviol_WENB_WCLK_posedge,
                            TmDt_WENB_WCLK_posedge,
                            WENB_ipd, "WENB",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WENB_WCLK_negedge_posedge,
                            thold_WENB_WCLK_negedge_posedge,
                            tsetup_WENB_WCLK_posedge_posedge,
                            thold_WENB_WCLK_posedge_posedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            '/',
                            InstancePath & "/BIOFIFO_BIDIRINFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            InstancePath & "/BIOFIFO_BIDIRINFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup CLRB high before WCLK rising
      --   Hold  CLRB high after WCLK rising

         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLRB_RCLK_posedge,
          TimingData              => TmDt_CLRB_RCLK_posedge,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          RefSignal               => RCLK_ipd,
          RefSignalName           => "RCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLRB_RCLK_posedge_posedge,
          Removal                 => thold_CLRB_RCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TO_X01((NOT RENB_ipd) ) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/BIOFIFO_BIDIRINFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLRB_WCLK_posedge,
          TimingData              => TmDt_CLRB_WCLK_posedge,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          RefSignal               => RCLK_ipd,
          RefSignalName           => "WCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLRB_WCLK_posedge_posedge,
          Removal                 => thold_CLRB_WCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TO_X01((NOT WENB_ipd) ) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/BIOFIFO_BIDIRINFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLRB,
          PeriodData              => PeriodData_CLRB,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLRB_negedge,
          CheckEnabled            => TRUE,
          HeaderMsg               => InstancePath &"/BIOFIFO_BIDIRINFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);


    end if;

      Y_zd := TO_X01(A_ipd);

    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################


      if (TO_X01(CLRB_ipd)='X') then
        assert false
        report ": CLRB unknown"
        severity Warning;
      elsif (TO_X01(CLRB_ipd)='0') then
        WADDR := -1;
        RADDR := -1;
      else
        if (TO_X01(WCLK_ipd)='X') then
	  if ((TO_X01(WENB_delayed) /= '1')) then
            if (TO_X01(WCLK_previous) /= 'X') then
	      assert false
	      report ": WCLK went unknown"
	      severity Warning;
	    end if;
	  end if;
        elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='1')) then
	  case (TO_X01(WENB_delayed)) is
	    when '1' =>
	      null;
	    when '0' =>
              -- Increment WADDR
              WADDR := WADDR + 1;
              if ((RADDR > WADDR) or (WADDR - RADDR > 63)) then
                assert false
                report ": Write failed - FIFO full."
                severity Warning;
              else
	        DUAL_PORT_RAM(WADDR mod 64) <= D_delayed ;
              end if;
	    when others =>
              if (TO_X01(WENB_previous) = 'X') then
                assert false
                report ": WENB went unknown"
                severity Warning;
              end if;
	  end case;
        end if;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      if (TO_X01(CLRB_ipd)='1') then
        if (TO_X01(RCLK_ipd) = 'X') then
          if ((TO_X01(RENB_delayed) /= '1')) then
	    Q_zd := 'X';
	    if (TO_X01(RCLK_previous) /= 'X') then
	      assert false
	      report ": RCLK went unknown"
	      severity Warning;
	    end if;
	  end if;
        elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '1')) then
	  case (TO_X01(RENB_delayed)) is
	    when '1' =>
	      null;
	    when '0' =>
              -- Increment RADDR
              RADDR := RADDR + 1;
              if ((RADDR > WADDR) or (WADDR - RADDR > 63)) then
                assert false
                report ": Read failed - FIFO empty."
                severity Warning;
              else
	        Q_zd := DUAL_PORT_RAM(RADDR mod 64);
              end if;
	    when others =>
	      Q_zd := 'X';
              if (TO_X01(RENB_delayed) = 'X') and (TO_X01(RENB_previous) /= 'X') then
	        assert false
	        report ": RENB went unknown"
	        severity Warning;
                RENB_previous := RENB_delayed;
              end if;
	  end case;
        end if;
      end if;

      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      if WENB_ipd'event then
        WENB_previous := WENB_delayed;
        WENB_delayed := WENB_ipd;
      end if;
      if RENB_ipd'event then
        RENB_previous := RENB_delayed;
        RENB_delayed := RENB_ipd;
      end if;
      D_delayed := D_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => Q,
	GlitchData => Q_GlitchData,
	OutSignalName => "Q",
	OutTemp => Q_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_Q), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => Xon,
	MsgOn => MsgOn,
	MsgSeverity => WARNING
	);

   VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);


  end process VITALBehavior;

end VITAL_ACT;


-----------------------------------------------------------------
--
--  Actel BIOFIFO_BIDIROUTFIFO VHDL behavioral model
--  64 X 1 I/O FIFO with rising write clock, rising read clock,
--  and active low WENB, RENB, and CLRB.
--  AFL macro containing feed-through.
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - 5/17/02 - Dale Walter - Clone of IOFIFO_INFIFO.
-- 2.0 - 9/27/02 - Krupa Singampalli - New Timing Arcs
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity BIOFIFO_BIDIROUTFIFO is
  GENERIC (
       tipd_A       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_D       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_CLRB      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_A_Y   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_Q   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLRB_Q    : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tsetup_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_D_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_negedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLRB_WCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLRB_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True

        );
  PORT (
        A     : IN STD_ULOGIC ;
        D     : IN STD_ULOGIC ;
        WENB     : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RENB     : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        CLRB    : IN STD_ULOGIC ;
        Q     : OUT STD_ULOGIC ;
        Y     : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of BIOFIFO_BIDIROUTFIFO : entity is FALSE;
  
end BIOFIFO_BIDIROUTFIFO;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of BIOFIFO_BIDIROUTFIFO is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE; 

  signal A_ipd   : std_ulogic := 'X';
  signal D_ipd   : std_ulogic := 'X';
  signal WENB_ipd   : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  signal RENB_ipd   : std_ulogic := 'X';
  signal RCLK_ipd : std_ulogic := 'X';
  signal CLRB_ipd  : std_ulogic := 'X';
  type MEM is array(0 to 63) of std_ulogic;
  signal DUAL_PORT_RAM : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (A_ipd, A, VitalExtendToFillDelay(tipd_A));
    VitalWireDelay (D_ipd, D, VitalExtendToFillDelay(tipd_D));
    VitalWireDelay (WENB_ipd, WENB, VitalExtendToFillDelay(tipd_WENB));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (RENB_ipd, RENB, VitalExtendToFillDelay(tipd_RENB));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
    VitalWireDelay (CLRB_ipd, CLRB, VitalExtendToFillDelay(tipd_CLRB));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (A_ipd, D_ipd, WENB_ipd, WCLK_ipd, RENB_ipd, RCLK_ipd, CLRB_ipd)

     --  Read Timing Check Results
     variable Tviol_RENB_RCLK_posedge : X01 := '0';
     variable TmDt_RENB_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_D_WCLK_posedge : X01 := '0';
     variable TmDt_D_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WENB_WCLK_posedge : X01 := '0';
     variable TmDt_WENB_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  CLRB Timing Check Results
     variable Tviol_CLRB_RCLK_posedge : X01 := '0';
     variable TmDt_CLRB_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_CLRB_WCLK_posedge : X01 := '0';
     variable TmDt_CLRB_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_CLRB : X01 := '0';
     variable PeriodData_CLRB : VitalPeriodDataType := VitalPeriodDataInit;

     --  Functional Results
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT : SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1; -- free running counter
     variable RADDR : integer := -1; -- free running counter
     variable Q_zd : std_ulogic;
     variable Y_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable Q_GlitchData : VitalGlitchDataType;
     variable Y_GlitchData : VitalGlitchDataType;

     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable RENB_delayed : std_ulogic := 'X';
     variable RENB_previous : std_ulogic := 'X';
     variable WENB_delayed : std_ulogic := 'X';
     variable WENB_previous : std_ulogic := 'X';
     variable D_delayed : std_ulogic := 'X';

  begin  --  process VITALBehavior 

    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RENB before RCLK rising
      --   Hold  RENB after RCLK rising

      VitalSetupHoldCheck ( Tviol_RENB_RCLK_posedge,
                            TmDt_RENB_RCLK_posedge,
                            RENB_ipd, "RENB",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RENB_RCLK_negedge_posedge,
			    tsetup_RENB_RCLK_posedge_posedge,
                            thold_RENB_RCLK_negedge_posedge,
                            thold_RENB_RCLK_posedge_posedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            '/',
                            InstancePath & "/BIOFIFO_BIDIROUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            InstancePath & "/BIOFIFO_BIDIROUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup D high or low before WCLK rising
      --   Hold  D high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_D_WCLK_posedge,
                            TmDt_D_WCLK_posedge,
                            D_ipd, "D",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_D_WCLK_negedge_posedge,
                            tsetup_D_WCLK_posedge_posedge,
                            thold_D_WCLK_negedge_posedge,
                            thold_D_WCLK_posedge_posedge,
                            TO_X01((CLRB_ipd) AND (NOT WENB_ipd)) /= '0',
                            '/',
                            InstancePath & "/BIOFIFO_BIDIROUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup WENB high before WCLK rising
      --   Hold  WENB high after WCLK rising

      VitalSetupHoldCheck ( Tviol_WENB_WCLK_posedge,
                            TmDt_WENB_WCLK_posedge,
                            WENB_ipd, "WENB",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WENB_WCLK_negedge_posedge,
                            tsetup_WENB_WCLK_posedge_posedge,
                            thold_WENB_WCLK_negedge_posedge,
                            thold_WENB_WCLK_posedge_posedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            '/',
                            InstancePath & "/BIOFIFO_BIDIROUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            InstancePath & "/BIOFIFO_BIDIROUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup CLRB high before WCLK rising
      --   Hold  CLRB high after WCLK rising

         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLRB_RCLK_posedge,
          TimingData              => TmDt_CLRB_RCLK_posedge,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          RefSignal               => RCLK_ipd,
          RefSignalName           => "RCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLRB_RCLK_posedge_posedge,
          Removal                 => thold_CLRB_RCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/BIOFIFO_BIDIROUTFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLRB_WCLK_posedge,
          TimingData              => TmDt_CLRB_WCLK_posedge,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          RefSignal               => RCLK_ipd,
          RefSignalName           => "WCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLRB_WCLK_posedge_posedge,
          Removal                 => thold_CLRB_WCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/BIOFIFO_BIDIROUTFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLRB,
          PeriodData              => PeriodData_CLRB,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLRB_negedge,
          CheckEnabled            => TRUE,
          HeaderMsg               => InstancePath &"/BIOFIFO_BIDIROUTFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);


    end if;

      Y_zd := TO_X01(A_ipd);

    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################


      if (TO_X01(CLRB_ipd)='X') then
        assert false
        report ": CLRB unknown"
        severity Warning;
      elsif (TO_X01(CLRB_ipd)='0') then
        WADDR := -1;
        RADDR := -1;
      else
        if (TO_X01(WCLK_ipd)='X') then
	  if ((TO_X01(WENB_delayed) /= '1')) then
            if (TO_X01(WCLK_previous) /= 'X') then
	      assert false
	      report ": WCLK went unknown"
	      severity Warning;
	    end if;
	  end if;
        elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='1')) then
	  case (TO_X01(WENB_delayed)) is
	    when '1' =>
	      null;
	    when '0' =>
              -- Increment WADDR
              WADDR := WADDR + 1;
              if ((RADDR > WADDR) or (WADDR - RADDR > 63)) then
                assert false
                report ": Write failed - FIFO full."
                severity warning;
              else
	        DUAL_PORT_RAM(WADDR mod 64) <= D_delayed ;
              end if;
	    when others =>
              if (TO_X01(WENB_previous) = 'X') then
                assert false
                report ": WENB went unknown"
                severity Warning;
              end if;
	  end case;
        end if;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      if (TO_X01(CLRB_ipd)='1') then
        if (TO_X01(RCLK_ipd) = 'X') then
          if ((TO_X01(RENB_delayed) /= '1')) then
	    Q_zd := 'X';
	    if (TO_X01(RCLK_previous) /= 'X') then
	      assert false
	      report ": RCLK went unknown"
	      severity Warning;
	    end if;
	  end if;
        elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '1')) then
	  case (TO_X01(RENB_delayed)) is
	    when '1' =>
	      null;
	    when '0' =>
              -- Increment RADDR
              RADDR := RADDR + 1;
              if ((RADDR > WADDR) or (WADDR - RADDR > 63)) then
                assert false
                report ": Read failed - FIFO empty."
                severity Warning;
              else
	        Q_zd := DUAL_PORT_RAM(RADDR mod 64);
              end if;
	    when others =>
	      Q_zd := 'X';
              if (TO_X01(RENB_delayed) = 'X') and (TO_X01(RENB_previous) /= 'X') then
	        assert false
	        report ": RENB went unknown"
	        severity Warning;
                RENB_previous := RENB_delayed;
              end if;
	  end case;
        end if;
      end if;

      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      if WENB_ipd'event then
        WENB_previous := WENB_delayed;
        WENB_delayed := WENB_ipd;
      end if;
      if RENB_ipd'event then
        RENB_previous := RENB_delayed;
        RENB_delayed := RENB_ipd;
      end if;
      D_delayed := D_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => Q,
	GlitchData => Q_GlitchData,
	OutSignalName => "Q",
	OutTemp => Q_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_Q), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => Xon,
	MsgOn => MsgOn,
	MsgSeverity => WARNING
	);

   VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
  end process VITALBehavior;

end VITAL_ACT;

-----------------------------------------------------------------
--
--  Actel BIOFIFO_INFIFO VHDL behavioral model
--  64 X 1 I/O FIFO with rising write clock, rising read clock,
--  and active low WENB, RENB, and CLRB.
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - 9/25/00 - Dale Walter - Prototype version.
-- 2.0 - 9/27/02 - Krupa Singampalli - New Timing Arcs
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity BIOFIFO_INFIFO is
  GENERIC (
        tipd_D       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_CLRB      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_Q   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLRB_Q    : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tsetup_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_negedge_posedge     :   VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLRB_WCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLRB_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True

        );
  PORT (
        D     : IN STD_ULOGIC ;
        WENB     : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RENB     : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        CLRB    : IN STD_ULOGIC ;
        Q     : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of BIOFIFO_INFIFO : entity is FALSE;
  
end BIOFIFO_INFIFO;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of BIOFIFO_INFIFO is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal D_ipd   : std_ulogic := 'X';
  signal WENB_ipd   : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  signal RENB_ipd   : std_ulogic := 'X';
  signal RCLK_ipd : std_ulogic := 'X';
  signal CLRB_ipd  : std_ulogic := 'X';
  type MEM is array(0 to 63) of std_ulogic;
  signal DUAL_PORT_RAM : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (D_ipd, D, VitalExtendToFillDelay(tipd_D));
    VitalWireDelay (WENB_ipd, WENB, VitalExtendToFillDelay(tipd_WENB));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (RENB_ipd, RENB, VitalExtendToFillDelay(tipd_RENB));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
    VitalWireDelay (CLRB_ipd, CLRB, VitalExtendToFillDelay(tipd_CLRB));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (D_ipd, WENB_ipd, WCLK_ipd, RENB_ipd, RCLK_ipd, CLRB_ipd)

     --  Read Timing Check Results
     variable Tviol_RENB_RCLK_posedge : X01 := '0';
     variable TmDt_RENB_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_D_WCLK_posedge : X01 := '0';
     variable TmDt_D_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WENB_WCLK_posedge : X01 := '0';
     variable TmDt_WENB_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  CLRB Timing Check Results
     variable Tviol_CLRB_RCLK_posedge : X01 := '0';
     variable TmDt_CLRB_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_CLRB_WCLK_posedge : X01 := '0';
     variable TmDt_CLRB_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_CLRB : X01 := '0';
     variable PeriodData_CLRB : VitalPeriodDataType := VitalPeriodDataInit;

     --  Functional Results
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT : SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1; -- free running counter
     variable RADDR : integer := -1; -- free running counter
     variable Q_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable Q_GlitchData : VitalGlitchDataType;

     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable RENB_delayed : std_ulogic := 'X';
     variable RENB_previous : std_ulogic := 'X';
     variable WENB_delayed : std_ulogic := 'X';
     variable WENB_previous : std_ulogic := 'X';
     variable D_delayed : std_ulogic := 'X';

  begin  --  process VITALBehavior 

    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RENB before RCLK rising
      --   Hold  RENB after RCLK rising

      VitalSetupHoldCheck ( Tviol_RENB_RCLK_posedge,
                            TmDt_RENB_RCLK_posedge,
                            RENB_ipd, "RENB",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RENB_RCLK_negedge_posedge,
			    tsetup_RENB_RCLK_posedge_posedge,
                            thold_RENB_RCLK_negedge_posedge,
                            thold_RENB_RCLK_posedge_posedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            '/',
                            InstancePath & "/BIOFIFO_INFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            InstancePath & "/BIOFIFO_INFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup D high or low before WCLK rising
      --   Hold  D high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_D_WCLK_posedge,
                            TmDt_D_WCLK_posedge,
                            D_ipd, "D",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_D_WCLK_negedge_posedge,
                            tsetup_D_WCLK_posedge_posedge,
                            thold_D_WCLK_negedge_posedge,
                            thold_D_WCLK_posedge_posedge,
                            TO_X01((CLRB_ipd) AND (NOT WENB_ipd)) /= '0',
                            '/',
                            InstancePath & "/BIOFIFO_INFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup WENB high before WCLK rising
      --   Hold  WENB high after WCLK rising

      VitalSetupHoldCheck ( Tviol_WENB_WCLK_posedge,
                            TmDt_WENB_WCLK_posedge,
                            WENB_ipd, "WENB",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WENB_WCLK_negedge_posedge,
                            tsetup_WENB_WCLK_posedge_posedge,
                            thold_WENB_WCLK_negedge_posedge,
                            thold_WENB_WCLK_posedge_posedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            '/',
                            InstancePath & "/BIOFIFO_INFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            InstancePath & "/BIOFIFO_INFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup CLRB high before WCLK rising
      --   Hold  CLRB high after WCLK rising

         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLRB_RCLK_posedge,
          TimingData              => TmDt_CLRB_RCLK_posedge,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          RefSignal               => RCLK_ipd,
          RefSignalName           => "RCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLRB_RCLK_posedge_posedge,
          Removal                 => thold_CLRB_RCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TO_X01( NOT RENB_ipd) /='0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/BIOFIFO_INFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLRB_WCLK_posedge,
          TimingData              => TmDt_CLRB_WCLK_posedge,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          RefSignal               => RCLK_ipd,
          RefSignalName           => "WCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLRB_WCLK_posedge_posedge,
          Removal                 => thold_CLRB_WCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TO_X01( NOT WENB_ipd) /='0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/BIOFIFO_INFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLRB,
          PeriodData              => PeriodData_CLRB,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLRB_negedge,
          CheckEnabled            => TRUE,
          HeaderMsg               => InstancePath &"/BIOFIFO_INFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);


    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################


      if (TO_X01(CLRB_ipd)='X') then
        assert false
        report ": CLRB unknown"
        severity Error;
      elsif (TO_X01(CLRB_ipd)='0') then
        WADDR := -1;
        RADDR := -1;
      else
        if (TO_X01(WCLK_ipd)='X') then
	  if ((TO_X01(WENB_delayed) /= '1')) then
            if (TO_X01(WCLK_previous) /= 'X') then
	      assert false
	      report ": WCLK went unknown"
	      severity Error;
	    end if;
	  end if;
        elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='1')) then
	  case (TO_X01(WENB_delayed)) is
	    when '1' =>
	      null;
	    when '0' =>
              -- Increment WADDR
              WADDR := WADDR + 1;
              if ((RADDR > WADDR) or (WADDR - RADDR > 63)) then
                assert false
                report ": Write failed - FIFO full."
                severity Error;
              else
	        DUAL_PORT_RAM(WADDR mod 64) <= D_delayed ;
              end if;
	    when others =>
              if (TO_X01(WENB_previous) = 'X') then
                assert false
                report ": WENB went unknown"
                severity Error;
              end if;
	  end case;
        end if;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      if (TO_X01(CLRB_ipd)='1') then
        if (TO_X01(RCLK_ipd) = 'X') then
          if ((TO_X01(RENB_delayed) /= '1')) then
	    Q_zd := 'X';
	    if (TO_X01(RCLK_previous) /= 'X') then
	      assert false
	      report ": RCLK went unknown"
	      severity Warning;
	    end if;
	  end if;
        elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '1')) then
	  case (TO_X01(RENB_delayed)) is
	    when '1' =>
	      null;
	    when '0' =>
              -- Increment RADDR
              RADDR := RADDR + 1;
              if ((RADDR > WADDR) or (WADDR - RADDR > 63)) then
                assert false
                report ": Read failed - FIFO empty."
                severity Error;
              else
	        Q_zd := DUAL_PORT_RAM(RADDR mod 64);
              end if;
	    when others =>
	      Q_zd := 'X';
              if (TO_X01(RENB_delayed) = 'X') and (TO_X01(RENB_previous) /= 'X') then
	        assert false
	        report ": RENB went unknown"
	        severity Warning;
                RENB_previous := RENB_delayed;
              end if;
	  end case;
        end if;
      end if;

      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      if WENB_ipd'event then
        WENB_previous := WENB_delayed;
        WENB_delayed := WENB_ipd;
      end if;
      if RENB_ipd'event then
        RENB_previous := RENB_delayed;
        RENB_delayed := RENB_ipd;
      end if;
      D_delayed := D_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => Q,
	GlitchData => Q_GlitchData,
	OutSignalName => "Q",
	OutTemp => Q_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_Q), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => Xon,
	MsgOn => MsgOn,
	MsgSeverity => WARNING
	);

    
  end process VITALBehavior;

end VITAL_ACT;

-----------------------------------------------------------------
--
--  Actel BIOFIFO_OUTFIFO VHDL behavioral model
--  64 X 1 I/O FIFO with rising write clock, rising read clock,
--  and active low WENB, RENB, and CLRB.
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - 9/25/00 - Dale Walter - Prototype version.
-- 2.0 - 9/27/02 - Krupa Singampalli - New Timing Arcs
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity BIOFIFO_OUTFIFO is
  GENERIC (
        tipd_D       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_CLRB      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_Q   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLRB_Q    : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tsetup_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_negedge_posedge     :   VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLRB_WCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLRB_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True

        );
  PORT (
        D     : IN STD_ULOGIC ;
        WENB     : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RENB     : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        CLRB    : IN STD_ULOGIC ;
        Q     : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of BIOFIFO_OUTFIFO : entity is FALSE;
  
end BIOFIFO_OUTFIFO;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of BIOFIFO_OUTFIFO is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal D_ipd   : std_ulogic := 'X';
  signal WENB_ipd   : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  signal RENB_ipd   : std_ulogic := 'X';
  signal RCLK_ipd : std_ulogic := 'X';
  signal CLRB_ipd  : std_ulogic := 'X';
  type MEM is array(0 to 63) of std_ulogic;
  signal DUAL_PORT_RAM : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (D_ipd, D, VitalExtendToFillDelay(tipd_D));
    VitalWireDelay (WENB_ipd, WENB, VitalExtendToFillDelay(tipd_WENB));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (RENB_ipd, RENB, VitalExtendToFillDelay(tipd_RENB));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
    VitalWireDelay (CLRB_ipd, CLRB, VitalExtendToFillDelay(tipd_CLRB));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (D_ipd, WENB_ipd, WCLK_ipd, RENB_ipd, RCLK_ipd, CLRB_ipd)

     --  Read Timing Check Results
     variable Tviol_RENB_RCLK_posedge : X01 := '0';
     variable TmDt_RENB_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_D_WCLK_posedge : X01 := '0';
     variable TmDt_D_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WENB_WCLK_posedge : X01 := '0';
     variable TmDt_WENB_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  CLRB Timing Check Results
     variable Tviol_CLRB_RCLK_posedge : X01 := '0';
     variable TmDt_CLRB_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_CLRB_WCLK_posedge : X01 := '0';
     variable TmDt_CLRB_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_CLRB : X01 := '0';
     variable PeriodData_CLRB : VitalPeriodDataType := VitalPeriodDataInit;

     --  Functional Results
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT : SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1; -- free running counter
     variable RADDR : integer := -1; -- free running counter
     variable Q_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable Q_GlitchData : VitalGlitchDataType;

     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable RENB_delayed : std_ulogic := 'X';
     variable RENB_previous : std_ulogic := 'X';
     variable WENB_delayed : std_ulogic := 'X';
     variable WENB_previous : std_ulogic := 'X';
     variable D_delayed : std_ulogic := 'X';

  begin  --  process VITALBehavior 

    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RENB before RCLK rising
      --   Hold  RENB after RCLK rising

      VitalSetupHoldCheck ( Tviol_RENB_RCLK_posedge,
                            TmDt_RENB_RCLK_posedge,
                            RENB_ipd, "RENB",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RENB_RCLK_posedge_posedge,
			    tsetup_RENB_RCLK_negedge_posedge,
                            thold_RENB_RCLK_posedge_posedge,
                            thold_RENB_RCLK_negedge_posedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            '/',
                            InstancePath & "/BIOFIFO_OUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            InstancePath & "/BIOFIFO_OUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup D high or low before WCLK rising
      --   Hold  D high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_D_WCLK_posedge,
                            TmDt_D_WCLK_posedge,
                            D_ipd, "D",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_D_WCLK_posedge_posedge,
                            tsetup_D_WCLK_negedge_posedge,
                            thold_D_WCLK_posedge_posedge,
                            thold_D_WCLK_posedge_posedge,
                            TO_X01((CLRB_ipd) AND (NOT WENB_ipd)) /= '0',
                            '/',
                            InstancePath & "/BIOFIFO_OUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup WENB high before WCLK rising
      --   Hold  WENB high after WCLK rising

      VitalSetupHoldCheck ( Tviol_WENB_WCLK_posedge,
                            TmDt_WENB_WCLK_posedge,
                            WENB_ipd, "WENB",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WENB_WCLK_posedge_posedge,
                            tsetup_WENB_WCLK_negedge_posedge,
                            thold_WENB_WCLK_posedge_posedge,
                            thold_WENB_WCLK_negedge_posedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            '/',
                            InstancePath & "/BIOFIFO_OUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            InstancePath & "/BIOFIFO_OUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup CLRB high before WCLK rising
      --   Hold  CLRB high after WCLK rising

         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLRB_RCLK_posedge,
          TimingData              => TmDt_CLRB_RCLK_posedge,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          RefSignal               => RCLK_ipd,
          RefSignalName           => "RCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLRB_RCLK_posedge_posedge,
          Removal                 => thold_CLRB_RCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TO_X01(NOT RENB_ipd ) /='0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/BIOFIFO_OUTFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLRB_WCLK_posedge,
          TimingData              => TmDt_CLRB_WCLK_posedge,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          RefSignal               => RCLK_ipd,
          RefSignalName           => "WCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLRB_WCLK_posedge_posedge,
          Removal                 => thold_CLRB_WCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TO_X01(NOT WENB_ipd ) /='0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/BIOFIFO_OUTFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLRB,
          PeriodData              => PeriodData_CLRB,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLRB_negedge,
          CheckEnabled            => TRUE,
          HeaderMsg               => InstancePath &"/BIOFIFO_OUTFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);


    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################


      if (TO_X01(CLRB_ipd)='X') then
        assert false
        report ": CLRB unknown"
        severity Error;
      elsif (TO_X01(CLRB_ipd)='0') then
        WADDR := -1;
        RADDR := -1;
      else
        if (TO_X01(WCLK_ipd)='X') then
	  if ((TO_X01(WENB_delayed) /= '1')) then
            if (TO_X01(WCLK_previous) /= 'X') then
	      assert false
	      report ": WCLK went unknown"
	      severity Error;
	    end if;
	  end if;
        elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='1')) then
	  case (TO_X01(WENB_delayed)) is
	    when '1' =>
	      null;
	    when '0' =>
              -- Increment WADDR
              WADDR := WADDR + 1;
              if ((RADDR > WADDR) or (WADDR - RADDR > 63)) then
                assert false
                report ": Write failed - FIFO full."
                severity Error;
              else
	        DUAL_PORT_RAM(WADDR mod 64) <= D_delayed ;
              end if;
	    when others =>
              if (TO_X01(WENB_previous) = 'X') then
                assert false
                report ": WENB went unknown"
                severity Error;
              end if;
	  end case;
        end if;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      if (TO_X01(CLRB_ipd)='1') then
        if (TO_X01(RCLK_ipd) = 'X') then
          if ((TO_X01(RENB_delayed) /= '1')) then
	    Q_zd := 'X';
	    if (TO_X01(RCLK_previous) /= 'X') then
	      assert false
	      report ": RCLK went unknown"
	      severity Warning;
	    end if;
	  end if;
        elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '1')) then
	  case (TO_X01(RENB_delayed)) is
	    when '1' =>
	      null;
	    when '0' =>
              -- Increment RADDR
              RADDR := RADDR + 1;
              if ((RADDR > WADDR) or (WADDR - RADDR > 63)) then
                assert false
                report ": Read failed - FIFO empty."
                severity Error;
              else
	        Q_zd := DUAL_PORT_RAM(RADDR mod 64);
              end if;
	    when others =>
	      Q_zd := 'X';
              if (TO_X01(RENB_delayed) = 'X') and (TO_X01(RENB_previous) /= 'X') then
	        assert false
	        report ": RENB went unknown"
	        severity Warning;
                RENB_previous := RENB_delayed;
              end if;
	  end case;
        end if;
      end if;

      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      if WENB_ipd'event then
        WENB_previous := WENB_delayed;
        WENB_delayed := WENB_ipd;
      end if;
      if RENB_ipd'event then
        RENB_previous := RENB_delayed;
        RENB_delayed := RENB_ipd;
      end if;
      D_delayed := D_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => Q,
	GlitchData => Q_GlitchData,
	OutSignalName => "Q",
	OutTemp => Q_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_Q), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => Xon,
	MsgOn => MsgOn,
	MsgSeverity => WARNING
	);

    
  end process VITALBehavior;

end VITAL_ACT;

-----------------------------------------------------------------
--
--  Actel IOFIFO_BIDIRINFIFO VHDL behavioral model
--  64 X 1 I/O FIFO with rising write clock, rising read clock,
--  and active low WENB, RENB, and CLRB.
--  AFL macro containing feed-through.
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - 5/17/02 - Dale Walter - Clone of IOFIFO_INFIFO.
-- 2.0 - 9/27/02 - Krupa Singampalli - New Timing Arcs
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity IOFIFO_BIDIRINFIFO is
  GENERIC (
        tipd_A       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_D       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_CLRB      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_A_Y   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_Q   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLRB_Q    : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tsetup_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_D_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_negedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLRB_WCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLRB_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True

        );
  PORT (
        A     : IN STD_ULOGIC ;
        D     : IN STD_ULOGIC ;
        WENB     : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RENB     : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        CLRB    : IN STD_ULOGIC ;
        Q     : OUT STD_ULOGIC ;
        Y     : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of IOFIFO_BIDIRINFIFO : entity is FALSE;
  
end IOFIFO_BIDIRINFIFO;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of IOFIFO_BIDIRINFIFO is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal A_ipd   : std_ulogic := 'X';
  signal D_ipd   : std_ulogic := 'X';
  signal WENB_ipd   : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  signal RENB_ipd   : std_ulogic := 'X';
  signal RCLK_ipd : std_ulogic := 'X';
  signal CLRB_ipd  : std_ulogic := 'X';
  type MEM is array(0 to 63) of std_ulogic;
  signal DUAL_PORT_RAM : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (A_ipd, A, VitalExtendToFillDelay(tipd_A));
    VitalWireDelay (D_ipd, D, VitalExtendToFillDelay(tipd_D));
    VitalWireDelay (WENB_ipd, WENB, VitalExtendToFillDelay(tipd_WENB));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (RENB_ipd, RENB, VitalExtendToFillDelay(tipd_RENB));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
    VitalWireDelay (CLRB_ipd, CLRB, VitalExtendToFillDelay(tipd_CLRB));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (A_ipd, D_ipd, WENB_ipd, WCLK_ipd, RENB_ipd, RCLK_ipd, CLRB_ipd)

     --  Read Timing Check Results
     variable Tviol_RENB_RCLK_posedge : X01 := '0';
     variable TmDt_RENB_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_D_WCLK_posedge : X01 := '0';
     variable TmDt_D_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WENB_WCLK_posedge : X01 := '0';
     variable TmDt_WENB_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  CLRB Timing Check Results
     variable Tviol_CLRB_RCLK_posedge : X01 := '0';
     variable TmDt_CLRB_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_CLRB_WCLK_posedge : X01 := '0';
     variable TmDt_CLRB_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_CLRB : X01 := '0';
     variable PeriodData_CLRB : VitalPeriodDataType := VitalPeriodDataInit;

     --  Functional Results
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT : SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1; -- free running counter
     variable RADDR : integer := -1; -- free running counter
     variable Q_zd : std_ulogic;
     variable Y_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable Q_GlitchData : VitalGlitchDataType;
     variable Y_GlitchData : VitalGlitchDataType;

     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable RENB_delayed : std_ulogic := 'X';
     variable RENB_previous : std_ulogic := 'X';
     variable WENB_delayed : std_ulogic := 'X';
     variable WENB_previous : std_ulogic := 'X';
     variable D_delayed : std_ulogic := 'X';

  begin  --  process VITALBehavior 

    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RENB before RCLK rising
      --   Hold  RENB after RCLK rising

      VitalSetupHoldCheck ( Tviol_RENB_RCLK_posedge,
                            TmDt_RENB_RCLK_posedge,
                            RENB_ipd, "RENB",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RENB_RCLK_posedge_posedge,
			    tsetup_RENB_RCLK_negedge_posedge,
                            thold_RENB_RCLK_posedge_posedge,
                            thold_RENB_RCLK_negedge_posedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            '/',
                            InstancePath & "/IOFIFO_BIDIRINFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            InstancePath & "/IOFIFO_BIDIRINFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup D high or low before WCLK rising
      --   Hold  D high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_D_WCLK_posedge,
                            TmDt_D_WCLK_posedge,
                            D_ipd, "D",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_D_WCLK_posedge_posedge,
                            tsetup_D_WCLK_negedge_posedge,
                            thold_D_WCLK_posedge_posedge,
                            thold_D_WCLK_negedge_posedge,
                            TO_X01((CLRB_ipd) AND (NOT WENB_ipd)) /= '0',
                            '/',
                            InstancePath & "/IOFIFO_BIDIRINFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup WENB high before WCLK rising
      --   Hold  WENB high after WCLK rising

      VitalSetupHoldCheck ( Tviol_WENB_WCLK_posedge,
                            TmDt_WENB_WCLK_posedge,
                            WENB_ipd, "WENB",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WENB_WCLK_posedge_posedge,
                            tsetup_WENB_WCLK_negedge_posedge,
                            thold_WENB_WCLK_posedge_posedge,
                            thold_WENB_WCLK_negedge_posedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            '/',
                            InstancePath & "/IOFIFO_BIDIRINFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            InstancePath & "/IOFIFO_BIDIRINFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup CLRB high before WCLK rising
      --   Hold  CLRB high after WCLK rising

         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLRB_RCLK_posedge,
          TimingData              => TmDt_CLRB_RCLK_posedge,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          RefSignal               => RCLK_ipd,
          RefSignalName           => "RCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLRB_RCLK_posedge_posedge,
          Removal                 => thold_CLRB_RCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IOFIFO_BIDIRINFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLRB_WCLK_posedge,
          TimingData              => TmDt_CLRB_WCLK_posedge,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          RefSignal               => RCLK_ipd,
          RefSignalName           => "WCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLRB_WCLK_posedge_posedge,
          Removal                 => thold_CLRB_WCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IOFIFO_BIDIRINFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLRB,
          PeriodData              => PeriodData_CLRB,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLRB_negedge,
          CheckEnabled            => TRUE,
          HeaderMsg               => InstancePath &"/IOFIFO_BIDIRINFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);


    end if;

      Y_zd := TO_X01(A_ipd);

    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################


      if (TO_X01(CLRB_ipd)='X') then
        assert false
        report ": CLRB unknown"
        severity Warning;
      elsif (TO_X01(CLRB_ipd)='0') then
        WADDR := -1;
        RADDR := -1;
      else
        if (TO_X01(WCLK_ipd)='X') then
	  if ((TO_X01(WENB_delayed) /= '1')) then
            if (TO_X01(WCLK_previous) /= 'X') then
	      assert false
	      report ": WCLK went unknown"
	      severity Warning;
	    end if;
	  end if;
        elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='1')) then
	  case (TO_X01(WENB_delayed)) is
	    when '1' =>
	      null;
	    when '0' =>
              -- Increment WADDR
              WADDR := WADDR + 1;
              if ((RADDR > WADDR) or (WADDR - RADDR > 63)) then
                assert false
                report ": Write failed - FIFO full."
                severity Warning;
              else
	        DUAL_PORT_RAM(WADDR mod 64) <= D_delayed ;
              end if;
	    when others =>
              if (TO_X01(WENB_previous) = 'X') then
                assert false
                report ": WENB went unknown"
                severity warning;
              end if;
	  end case;
        end if;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      if (TO_X01(CLRB_ipd)='1') then
        if (TO_X01(RCLK_ipd) = 'X') then
          if ((TO_X01(RENB_delayed) /= '1')) then
	    Q_zd := 'X';
	    if (TO_X01(RCLK_previous) /= 'X') then
	      assert false
	      report ": RCLK went unknown"
	      severity Warning;
	    end if;
	  end if;
        elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '1')) then
	  case (TO_X01(RENB_delayed)) is
	    when '1' =>
	      null;
	    when '0' =>
              -- Increment RADDR
              RADDR := RADDR + 1;
              if ((RADDR > WADDR) or (WADDR - RADDR > 63)) then
                assert false
                report ": Read failed - FIFO empty."
                severity Warning;
              else
	        Q_zd := DUAL_PORT_RAM(RADDR mod 64);
              end if;
	    when others =>
	      Q_zd := 'X';
              if (TO_X01(RENB_delayed) = 'X') and (TO_X01(RENB_previous) /= 'X') then
	        assert false
	        report ": RENB went unknown"
	        severity Warning;
                RENB_previous := RENB_delayed;
              end if;
	  end case;
        end if;
      end if;

      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      if WENB_ipd'event then
        WENB_previous := WENB_delayed;
        WENB_delayed := WENB_ipd;
      end if;
      if RENB_ipd'event then
        RENB_previous := RENB_delayed;
        RENB_delayed := RENB_ipd;
      end if;
      D_delayed := D_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => Q,
	GlitchData => Q_GlitchData,
	OutSignalName => "Q",
	OutTemp => Q_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_Q), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => Xon,
	MsgOn => MsgOn,
	MsgSeverity => WARNING
	);

   VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

  end process VITALBehavior;

end VITAL_ACT;

----- CELL IOPADP_IN -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IOPADP_IN is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpw_PAD_posedge 		: VitalDelayType := 0.000 ns;
      tpw_PAD_negedge           : VitalDelayType := 0.000 ns;
      tpw_N2PIN_posedge         : VitalDelayType := 0.000 ns;
      tpw_N2PIN_negedge         : VitalDelayType := 0.000 ns;
      tpd_PAD_Y                      :        VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_N2PIN_Y                    :        VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PAD                       :        VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_N2PIN                     :        VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :        in    STD_ULOGIC;
      N2PIN                         :        in    STD_ULOGIC;
      Y                              :        out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IOPADP_IN : entity is FALSE;
end IOPADP_IN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of IOPADP_IN is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL PAD_ipd      : STD_ULOGIC := 'X';
   SIGNAL N2PIN_ipd    : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   VitalWireDelay (N2PIN_ipd, N2PIN, tipd_N2PIN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PAD_ipd, N2PIN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);
   ALIAS X_zd : STD_LOGIC is Results(2);
  
   -- timing check results
  VARIABLE Pviol_PAD       : STD_ULOGIC := '0';
  VARIABLE PeriodData_PAD  : VitalPeriodDataType := VitalPeriodDataInit;
  VARIABLE Pviol_N2PIN       : STD_ULOGIC := '0'; 
  VARIABLE PeriodData_N2PIN  : VitalPeriodDataType := VitalPeriodDataInit;

   -- output glitch detection variables
   VARIABLE Y_GlitchData      : VitalGlitchDataType;

   begin
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADP_IN",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

            VitalPeriodPulseCheck (
              Violation      => Pviol_N2PIN,
              PeriodData     => PeriodData_N2PIN,
              TestSignal     => PAD_ipd,
              TestSignalName => "N2PIN",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_N2PIN_posedge,
              PulseWidthLow  => tpw_N2PIN_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADP_IN",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(PAD_ipd);
      X_zd := TO_X01(N2PIN_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => VitalTransport,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_IOPADP_IN_VITAL of IOPADP_IN is
   for VITAL_ACT
   end for;
end CFG_IOPADP_IN_VITAL;


----- CELL IOPADN_IN -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IOPADN_IN is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      
      tpw_PAD_posedge 		: VitalDelayType := 0.000 ns;
      tpw_PAD_negedge           : VitalDelayType := 0.000 ns;      
      tpd_PAD_N2POUT                 :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      N2POUT                         :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IOPADN_IN : entity is FALSE;
end IOPADN_IN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;
architecture VITAL_ACT of IOPADN_IN is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS N2POUT_zd : STD_LOGIC is Results(1);

   -- timing check results
   VARIABLE Pviol_PAD       : STD_ULOGIC := '0';
   VARIABLE PeriodData_PAD  : VitalPeriodDataType := VitalPeriodDataInit;

   -- output glitch detection variables
   VARIABLE N2POUT_GlitchData	: VitalGlitchDataType;

   begin
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADN_IN",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

      -------------------------
      --  Functionality Section
      -------------------------
      N2POUT_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => N2POUT,
       GlitchData => N2POUT_GlitchData,
       OutSignalName => "N2POUT",
       OutTemp => N2POUT_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_N2POUT, TRUE)),
       Mode => VitalTransport,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_IOPADN_IN_VITAL of IOPADN_IN is
   for VITAL_ACT
   end for;
end CFG_IOPADN_IN_VITAL;


----- CELL IOPADP_TRI -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IOPADP_TRI is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      
      tpw_E_posedge                  :  VitalDelayType := 0.000 ns;
      tpw_E_negedge		     :  VitalDelayType := 0.000 ns;
      tpw_D_posedge		     :  VitalDelayType := 0.000 ns;
      tpw_D_negedge		     :  VitalDelayType := 0.000 ns;

      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IOPADP_TRI : entity is FALSE;
end IOPADP_TRI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;
architecture VITAL_ACT of IOPADP_TRI is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);
   
   -- timing check results
   VARIABLE Pviol_D       : STD_ULOGIC := '0'; 
   VARIABLE PeriodData_D  : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_E      : STD_ULOGIC := '0'; 
   VARIABLE PeriodData_E  : VitalPeriodDataType := VitalPeriodDataInit;

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADP_TRI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );
           
            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADP_TRI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_PAD), TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => VitalTransport,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL_ACT;

configuration CFG_IOPADP_TRI_VITAL of IOPADP_TRI is
   for VITAL_ACT
   end for;
end CFG_IOPADP_TRI_VITAL;


----- CELL IOPADN_TRI -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IOPADN_TRI is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      
      tpw_E_posedge              : VitalDelayType := 0.000 ns;    
      tpw_E_negedge		     : VitalDelayType := 0.000 ns;
      tpw_DB_posedge	     : VitalDelayType := 0.000 ns;
      tpw_DB_negedge             : VitalDelayType := 0.000 ns;
	
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_DB_PAD                     :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_DB                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      DB                             :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IOPADN_TRI : entity is FALSE;
end IOPADN_TRI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;
architecture VITAL_ACT of IOPADN_TRI is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL DB_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (DB_ipd, DB, tipd_DB);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (DB_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);

   -- timing check results
   VARIABLE Pviol_DB      : STD_ULOGIC := '0';
   VARIABLE PeriodData_DB : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_E       : STD_ULOGIC := '0';
   VARIABLE PeriodData_E  : VitalPeriodDataType := VitalPeriodDataInit;

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_DB,
              PeriodData     => PeriodData_DB,
              TestSignal     => DB_ipd,
              TestSignalName => "DB",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_DB_posedge,
              PulseWidthLow  => tpw_DB_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADN_TRI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADN_TRI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => (NOT DB_ipd),
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_PAD), TRUE),
                 1 => (DB_ipd'last_event, VitalExtendToFillDelay(tpd_DB_PAD), TRUE)),
       Mode => VitalTransport,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL_ACT;

configuration CFG_IOPADN_TRI_VITAL of IOPADN_TRI is
   for VITAL_ACT
   end for;
end CFG_IOPADN_TRI_VITAL;


----- CELL CLKBUF_LVDS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKBUF_LVDS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                     :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                     :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKBUF_LVDS : entity is TRUE;
end CLKBUF_LVDS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of CLKBUF_LVDS is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL PADP_ipd      : STD_ULOGIC := 'X';
   SIGNAL PADN_ipd      : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PADP_ipd, PADP, tipd_PADP);
   VitalWireDelay (PADN_ipd, PADN, tipd_PADN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PADP_ipd, PADN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData        : VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      if ((TO_X01(PADP_ipd) = '1') AND (TO_X01(PADN_ipd) = '0')) then
        Y_zd := '1';
      elsif ((TO_X01(PADP_ipd) = '0') AND (TO_X01(PADN_ipd) = '1')) then
        Y_zd := '0';
      else
        Y_zd := 'X';
      end if;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PADP_ipd'last_event, tpd_PADP_Y, TRUE),
                 1 => (PADN_ipd'last_event, tpd_PADN_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CLKBUF_LVDS_VITAL of CLKBUF_LVDS is
   for VITAL_ACT
   end for;
end CFG_CLKBUF_LVDS_VITAL;
----- CELL CLKBUF_LVPECL -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKBUF_LVPECL is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                     :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                     :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKBUF_LVPECL : entity is TRUE;
end CLKBUF_LVPECL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of CLKBUF_LVPECL is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL PADP_ipd      : STD_ULOGIC := 'X';
   SIGNAL PADN_ipd      : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PADP_ipd, PADP, tipd_PADP);
   VitalWireDelay (PADN_ipd, PADN, tipd_PADN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PADP_ipd, PADN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData        : VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      if ((TO_X01(PADP_ipd) = '1') AND (TO_X01(PADN_ipd) = '0')) then
        Y_zd := '1';
      elsif ((TO_X01(PADP_ipd) = '0') AND (TO_X01(PADN_ipd) = '1')) then
        Y_zd := '0';
      else
        Y_zd := 'X';
      end if;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PADP_ipd'last_event, tpd_PADP_Y, TRUE),
                 1 => (PADN_ipd'last_event, tpd_PADN_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CLKBUF_LVPECL_VITAL of CLKBUF_LVPECL is
   for VITAL_ACT
   end for;
end CFG_CLKBUF_LVPECL_VITAL;

----- CELL HCLKBUF_LVDS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity HCLKBUF_LVDS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                     :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                     :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);
attribute VITAL_LEVEL0 of HCLKBUF_LVDS : entity is TRUE;
end HCLKBUF_LVDS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of HCLKBUF_LVDS is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL PADP_ipd      : STD_ULOGIC := 'X';
   SIGNAL PADN_ipd      : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PADP_ipd, PADP, tipd_PADP);
   VitalWireDelay (PADN_ipd, PADN, tipd_PADN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PADP_ipd, PADN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData        : VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      if ((TO_X01(PADP_ipd) = '1') AND (TO_X01(PADN_ipd) = '0')) then
        Y_zd := '1';
      elsif ((TO_X01(PADP_ipd) = '0') AND (TO_X01(PADN_ipd) = '1')) then
        Y_zd := '0';
      else
        Y_zd := 'X';
      end if;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PADP_ipd'last_event, tpd_PADP_Y, TRUE),
                 1 => (PADN_ipd'last_event, tpd_PADN_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_HCLKBUF_LVDS_VITAL of HCLKBUF_LVDS is
   for VITAL_ACT
   end for;
end CFG_HCLKBUF_LVDS_VITAL;
----- CELL HCLKBUF_LVPECL -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity HCLKBUF_LVPECL is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                     :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                     :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);
attribute VITAL_LEVEL0 of HCLKBUF_LVPECL : entity is TRUE;
end HCLKBUF_LVPECL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of HCLKBUF_LVPECL is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL PADP_ipd      : STD_ULOGIC := 'X';
   SIGNAL PADN_ipd      : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PADP_ipd, PADP, tipd_PADP);
   VitalWireDelay (PADN_ipd, PADN, tipd_PADN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PADP_ipd, PADN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData        : VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      if ((TO_X01(PADP_ipd) = '1') AND (TO_X01(PADN_ipd) = '0')) then
        Y_zd := '1';
      elsif ((TO_X01(PADP_ipd) = '0') AND (TO_X01(PADN_ipd) = '1')) then
        Y_zd := '0';
      else
        Y_zd := 'X';
      end if;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PADP_ipd'last_event, tpd_PADP_Y, TRUE),
                 1 => (PADN_ipd'last_event, tpd_PADN_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_HCLKBUF_LVPECL_VITAL of HCLKBUF_LVPECL is
   for VITAL_ACT
   end for;
end CFG_HCLKBUF_LVPECL_VITAL;

----- CELL INBUF_LVDS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INBUF_LVDS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                     :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                     :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INBUF_LVDS : entity is TRUE;
end INBUF_LVDS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of INBUF_LVDS is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL PADP_ipd      : STD_ULOGIC := 'X';
   SIGNAL PADN_ipd      : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PADP_ipd, PADP, tipd_PADP);
   VitalWireDelay (PADN_ipd, PADN, tipd_PADN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PADP_ipd, PADN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData        : VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      if ((TO_X01(PADP_ipd) = '1') AND (TO_X01(PADN_ipd) = '0')) then
        Y_zd := '1';
      elsif ((TO_X01(PADP_ipd) = '0') AND (TO_X01(PADN_ipd) = '1')) then
        Y_zd := '0';
      else
        Y_zd := 'X';
      end if;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PADP_ipd'last_event, tpd_PADP_Y, TRUE),
                 1 => (PADN_ipd'last_event, tpd_PADN_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_INBUF_LVDS_VITAL of INBUF_LVDS is
   for VITAL_ACT
   end for;
end CFG_INBUF_LVDS_VITAL;
----- CELL INBUF_LVPECL -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INBUF_LVPECL is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                     :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                     :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INBUF_LVPECL : entity is TRUE;
end INBUF_LVPECL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of INBUF_LVPECL is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL PADP_ipd      : STD_ULOGIC := 'X';
   SIGNAL PADN_ipd      : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PADP_ipd, PADP, tipd_PADP);
   VitalWireDelay (PADN_ipd, PADN, tipd_PADN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PADP_ipd, PADN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData        : VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      if ((TO_X01(PADP_ipd) = '1') AND (TO_X01(PADN_ipd) = '0')) then
        Y_zd := '1';
      elsif ((TO_X01(PADP_ipd) = '0') AND (TO_X01(PADN_ipd) = '1')) then
        Y_zd := '0';
      else
        Y_zd := 'X';
      end if;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PADP_ipd'last_event, tpd_PADP_Y, TRUE),
                 1 => (PADN_ipd'last_event, tpd_PADN_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_INBUF_LVPECL_VITAL of INBUF_LVPECL is
   for VITAL_ACT
   end for;
end CFG_INBUF_LVPECL_VITAL;

----- CELL OUTBUF_LVDS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OUTBUF_LVDS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_PADP                     :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D_PADN                     :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      PADP                           :	out   STD_ULOGIC;
      PADN                           :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OUTBUF_LVDS : entity is TRUE;
end OUTBUF_LVDS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of OUTBUF_LVDS is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS PADP_zd : STD_LOGIC is Results(1);
   ALIAS PADN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE PADP_GlitchData	: VitalGlitchDataType;
   VARIABLE PADN_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PADP_zd := TO_X01(D_ipd);
      PADN_zd := NOT(TO_X01(D_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => PADP,
       GlitchData => PADP_GlitchData,
       OutSignalName => "PADP",
       OutTemp => PADP_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_PADP, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

      VitalPathDelay01 (
       OutSignal => PADN,
       GlitchData => PADN_GlitchData,
       OutSignalName => "PADN",
       OutTemp => PADN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_PADN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OUTBUF_LVDS_VITAL of OUTBUF_LVDS is
   for VITAL_ACT
   end for;
end CFG_OUTBUF_LVDS_VITAL;


----- CELL OUTBUF_LVPECL -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OUTBUF_LVPECL is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_PADP                     :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D_PADN                     :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      PADP                           :	out   STD_ULOGIC;
      PADN                           :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OUTBUF_LVPECL : entity is TRUE;
end OUTBUF_LVPECL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of OUTBUF_LVPECL is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS PADP_zd : STD_LOGIC is Results(1);
   ALIAS PADN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE PADP_GlitchData	: VitalGlitchDataType;
   VARIABLE PADN_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PADP_zd := TO_X01(D_ipd);
      PADN_zd := NOT(TO_X01(D_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => PADP,
       GlitchData => PADP_GlitchData,
       OutSignalName => "PADP",
       OutTemp => PADP_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_PADP, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

      VitalPathDelay01 (
       OutSignal => PADN,
       GlitchData => PADN_GlitchData,
       OutSignalName => "PADN",
       OutTemp => PADN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_PADN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OUTBUF_LVPECL_VITAL of OUTBUF_LVPECL is
   for VITAL_ACT
   end for;
end CFG_OUTBUF_LVPECL_VITAL;


----- CELL CM8F -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CM8F is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S11_Y                      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_S10_Y                      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_S01_Y                      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_S00_Y                      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D3_Y                       :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D2_Y                       :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D1_Y                       :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D0_Y                       :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_S11_FY                     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_S10_FY                     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_S01_FY                     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_S00_FY                     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D3_FY                      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D2_FY                      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D1_FY                      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D0_FY                      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_D0                        :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S00                       :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S01                       :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S10                       :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S11                       :  VitalDelayType01 := (0.000 ns, 0.000 ns));


   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S00                            :	in    STD_ULOGIC;
      S01                            :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      FY                             :	out   STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CM8F : entity is TRUE;
end CM8F;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of CM8F is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S00_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S01_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S11_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S00_ipd, S00, tipd_S00);
   VitalWireDelay (S01_ipd, S01, tipd_S01);
   VitalWireDelay (S10_ipd, S10, tipd_S10);
   VitalWireDelay (S11_ipd, S11, tipd_S11);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S00_ipd, S01_ipd, S10_ipd, S11_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);
   VARIABLE AND_Out, OR_Out, MUX1_Out, MUX2_Out : std_ulogic;

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;
   VARIABLE FY_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      AND_Out := VitalAND2(S00_ipd, S01_ipd);
      OR_Out := VitalOR2(S10_ipd, S11_ipd);
      MUX1_Out := VitalMUX2(D1_ipd, D0_ipd, AND_Out);
      MUX2_Out := VitalMUX2(D3_ipd, D2_ipd, AND_Out);
      Y_zd := VitalMUX2(MUX2_Out, MUX1_Out, OR_Out);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S11_ipd'last_event, tpd_S11_Y, TRUE),
                 1 => (S10_ipd'last_event, tpd_S10_Y, TRUE),
                 2 => (S01_ipd'last_event, tpd_S01_Y, TRUE),
                 3 => (S00_ipd'last_event, tpd_S00_Y, TRUE),
                 4 => (D3_ipd'last_event, tpd_D3_Y, TRUE),
                 5 => (D2_ipd'last_event, tpd_D2_Y, TRUE),
                 6 => (D1_ipd'last_event, tpd_D1_Y, TRUE),
                 7 => (D0_ipd'last_event, tpd_D0_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

      VitalPathDelay01 (
       OutSignal => FY,
       GlitchData => FY_GlitchData,
       OutSignalName => "FY",
       OutTemp => Y_zd,
       Paths => (0 => (S11_ipd'last_event, tpd_S11_FY, TRUE),
                 1 => (S10_ipd'last_event, tpd_S10_FY, TRUE),
                 2 => (S01_ipd'last_event, tpd_S01_FY, TRUE),
                 3 => (S00_ipd'last_event, tpd_S00_FY, TRUE),
                 4 => (D3_ipd'last_event, tpd_D3_FY, TRUE),
                 5 => (D2_ipd'last_event, tpd_D2_FY, TRUE),
                 6 => (D1_ipd'last_event, tpd_D1_FY, TRUE),
                 7 => (D0_ipd'last_event, tpd_D0_FY, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CM8F_VITAL of CM8F is
   for VITAL_ACT
   end for;
end CFG_CM8F_VITAL;

-----------------------------------------------------------------
--
--  Actel AX FIFO64K36 VHDL VITAL model
--  64K X 36 FIFO with rising write clock and rising read clock.
--  Allowable word widths x heights:
--    4096 x 1
--    2048 x 2
--    1024 x 4
--     512 x 9
--     256 x 18
--     128 x 36
--  Allowable depths: 1 to 16.
--
--  Assumptions:  
--    1. WEN, REN, and CLR active high.
--    2. WIDTH, DEPTH, AEVAL, and AFVAL static.
--    3. AEVAL and AFVAL specify the number of words between the
--       Read and Write address pointers.
--
--  Uses VITAL95 package
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - 2/8/01 - Dale Walter - Initial Version.  Not sure about timing arcs.
--                              Included all imaginable - some may need to be
--                              removed later.  Lowest DEPTH bit ignored.
-- 1.1 - 05/10/01 - Dale Walter - Change memory to variable instead of signal.
-- 1.2 - 05/31/01 - BT          _ modify the read/write operation, so both 
--                                operations can take care of all four flags.
-- 1.3 - 06/07/01 - Dale Walter - Change the CLR recovery/removal generics to 
--                                match NGT timing arcs.  Only check against
--                                WCLK, so RCLK checks removed.
-- 1.4 - 9/27/02 - Krupa Singampalli - New Timing Arcs
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity FIFO64K36 is
  GENERIC (
        tipd_DEPTH3   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH2   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH1   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH0   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WIDTH2   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WIDTH1   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WIDTH0   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AEVAL7   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AEVAL6   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AEVAL5   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AEVAL4   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AEVAL3   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AEVAL2   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AEVAL1   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AEVAL0   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AFVAL7   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AFVAL6   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AFVAL5   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AFVAL4   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AFVAL3   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AFVAL2   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AFVAL1   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_AFVAL0   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_REN      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD35     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD34     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD33     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD32     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD31     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD30     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD29     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD28     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD27     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD26     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD25     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD24     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD23     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD22     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD21     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD20     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD19     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD18     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD17     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD16     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD15     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD14     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD13     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD12     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD11     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD10     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD9      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD8      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD7      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD6      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD5      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD4      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD3      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WEN      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_CLR      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD1  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD2  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD3  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD4  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD5  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD6  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD7  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD8  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD9  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD10 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD11 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD12 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD13 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD14 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD15 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD16 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD17 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD18 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD19 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD20 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD21 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD22 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD23 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD24 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD25 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD26 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD27 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD28 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD29 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD30 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD31 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD32 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD33 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD34 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD35 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_FULL   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_AFULL  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_EMPTY  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_AEMPTY : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD0  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD1  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD2  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD3  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD4  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD5  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD6  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD7  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD8  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD9  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD10 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD11 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD12 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD13 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD14 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD15 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD16 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD17 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD18 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD19 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD20 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD21 : VitalDelayType01 := (0.100 ns, 0.10 ns);
        tpd_CLR_RD22 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD23 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD24 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD25 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD26 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD27 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD28 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD29 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD30 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD31 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD32 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD33 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_RD34 : VitalDelayType01 := (0.1000 ns, 0.100 ns);
        tpd_CLR_RD35 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_FULL   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_AFULL  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_EMPTY  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLR_AEMPTY : VitalDelayType01 := (0.100 ns, 0.100 ns);


        tsetup_WD35_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD34_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD33_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD32_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD31_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD30_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD29_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD28_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD27_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD26_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD25_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD24_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD23_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD22_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD21_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD20_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD19_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD18_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD17_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD16_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD15_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD14_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD13_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD12_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD11_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD10_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD9_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD8_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD35_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD34_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD33_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD32_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD31_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD30_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD29_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD28_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD27_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD26_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD25_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD24_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD23_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD22_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD21_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD20_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD19_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD18_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD17_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD16_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD15_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD14_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD13_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD12_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD11_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD10_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD9_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD8_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;

        tsetup_WEN_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

        tsetup_DEPTH3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        tsetup_WIDTH2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_AEVAL7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_AFVAL7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_DEPTH3_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH3_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_DEPTH0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        tsetup_WIDTH2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WIDTH0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        tsetup_AEVAL7_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL6_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL5_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL4_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL3_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL7_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL6_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL5_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL4_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL3_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AEVAL0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_AFVAL7_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL6_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL5_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL4_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL3_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL7_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL6_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL5_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL4_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL3_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_AFVAL0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_REN_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

        thold_WD35_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD34_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD33_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD32_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD31_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD30_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD29_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD28_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD27_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD26_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD25_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD24_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD23_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD22_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD21_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD20_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD19_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD18_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD17_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD16_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD15_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD14_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD13_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD12_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD11_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD10_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD9_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD8_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD35_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD34_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD33_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD32_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD31_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD30_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD29_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD28_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD27_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD26_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD25_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD24_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD23_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD22_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD21_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD20_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD19_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD18_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD17_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD16_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD15_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD14_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD13_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD12_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD11_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD10_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD9_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD8_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;


        thold_WEN_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

        thold_DEPTH3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        thold_WIDTH2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        thold_AEVAL7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        thold_AFVAL7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;



        thold_DEPTH3_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH3_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        thold_WIDTH2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WIDTH0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        thold_AEVAL7_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL6_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL5_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL4_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL3_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL7_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL6_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL5_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL4_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL3_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AEVAL0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        thold_AFVAL7_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL6_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL5_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL4_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL3_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL7_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL6_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL5_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL4_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL3_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_AFVAL0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        thold_REN_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

         
        trecovery_CLR_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLR_RCLK_posedge_posedge      :  VitalDelayType := 0.000 ns;
        trecovery_CLR_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLR_WCLK_posedge_posedge      :  VitalDelayType := 0.000 ns;

        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLR_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True
        );
  PORT (
        DEPTH3 : IN STD_ULOGIC ;
        DEPTH2 : IN STD_ULOGIC ;
        DEPTH1 : IN STD_ULOGIC ;
        DEPTH0 : IN STD_ULOGIC ;
        WIDTH2 : IN STD_ULOGIC ;
        WIDTH1 : IN STD_ULOGIC ;
        WIDTH0 : IN STD_ULOGIC ;
        AEVAL7 : IN STD_ULOGIC ;
        AEVAL6 : IN STD_ULOGIC ;
        AEVAL5 : IN STD_ULOGIC ;
        AEVAL4 : IN STD_ULOGIC ;
        AEVAL3 : IN STD_ULOGIC ;
        AEVAL2 : IN STD_ULOGIC ;
        AEVAL1 : IN STD_ULOGIC ;
        AEVAL0 : IN STD_ULOGIC ;
        AFVAL7 : IN STD_ULOGIC ;
        AFVAL6 : IN STD_ULOGIC ;
        AFVAL5 : IN STD_ULOGIC ;
        AFVAL4 : IN STD_ULOGIC ;
        AFVAL3 : IN STD_ULOGIC ;
        AFVAL2 : IN STD_ULOGIC ;
        AFVAL1 : IN STD_ULOGIC ;
        AFVAL0 : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        WD35   : IN STD_ULOGIC ;
        WD34   : IN STD_ULOGIC ;
        WD33   : IN STD_ULOGIC ;
        WD32   : IN STD_ULOGIC ;
        WD31   : IN STD_ULOGIC ;
        WD30   : IN STD_ULOGIC ;
        WD29   : IN STD_ULOGIC ;
        WD28   : IN STD_ULOGIC ;
        WD27   : IN STD_ULOGIC ;
        WD26   : IN STD_ULOGIC ;
        WD25   : IN STD_ULOGIC ;
        WD24   : IN STD_ULOGIC ;
        WD23   : IN STD_ULOGIC ;
        WD22   : IN STD_ULOGIC ;
        WD21   : IN STD_ULOGIC ;
        WD20   : IN STD_ULOGIC ;
        WD19   : IN STD_ULOGIC ;
        WD18   : IN STD_ULOGIC ;
        WD17   : IN STD_ULOGIC ;
        WD16   : IN STD_ULOGIC ;
        WD15   : IN STD_ULOGIC ;
        WD14   : IN STD_ULOGIC ;
        WD13   : IN STD_ULOGIC ;
        WD12   : IN STD_ULOGIC ;
        WD11   : IN STD_ULOGIC ;
        WD10   : IN STD_ULOGIC ;
        WD9    : IN STD_ULOGIC ;
        WD8    : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        CLR    : IN STD_ULOGIC ;
        RD35   : OUT STD_ULOGIC ;
        RD34   : OUT STD_ULOGIC ;
        RD33   : OUT STD_ULOGIC ;
        RD32   : OUT STD_ULOGIC ;
        RD31   : OUT STD_ULOGIC ;
        RD30   : OUT STD_ULOGIC ;
        RD29   : OUT STD_ULOGIC ;
        RD28   : OUT STD_ULOGIC ;
        RD27   : OUT STD_ULOGIC ;
        RD26   : OUT STD_ULOGIC ;
        RD25   : OUT STD_ULOGIC ;
        RD24   : OUT STD_ULOGIC ;
        RD23   : OUT STD_ULOGIC ;
        RD22   : OUT STD_ULOGIC ;
        RD21   : OUT STD_ULOGIC ;
        RD20   : OUT STD_ULOGIC ;
        RD19   : OUT STD_ULOGIC ;
        RD18   : OUT STD_ULOGIC ;
        RD17   : OUT STD_ULOGIC ;
        RD16   : OUT STD_ULOGIC ;
        RD15   : OUT STD_ULOGIC ;
        RD14   : OUT STD_ULOGIC ;
        RD13   : OUT STD_ULOGIC ;
        RD12   : OUT STD_ULOGIC ;
        RD11   : OUT STD_ULOGIC ;
        RD10   : OUT STD_ULOGIC ;
        RD9    : OUT STD_ULOGIC ;
        RD8    : OUT STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC ;
        RD6    : OUT STD_ULOGIC ;
        RD5    : OUT STD_ULOGIC ;
        RD4    : OUT STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC ;
        RD2    : OUT STD_ULOGIC ;
        RD1    : OUT STD_ULOGIC ;
        RD0    : OUT STD_ULOGIC ;
        FULL   : OUT STD_ULOGIC ;
        AFULL  : OUT STD_ULOGIC ;
        EMPTY  : OUT STD_ULOGIC ;
        AEMPTY : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of FIFO64K36 : entity is TRUE;
  
end FIFO64K36;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of FIFO64K36 is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal DEPTH3_ipd : std_ulogic := 'X';
  signal DEPTH2_ipd : std_ulogic := 'X';
  signal DEPTH1_ipd : std_ulogic := 'X';
  signal DEPTH0_ipd : std_ulogic := 'X';
  signal WIDTH2_ipd : std_ulogic := 'X';
  signal WIDTH1_ipd : std_ulogic := 'X';
  signal WIDTH0_ipd : std_ulogic := 'X';
  signal AEVAL7_ipd : std_ulogic := 'X';
  signal AEVAL6_ipd : std_ulogic := 'X';
  signal AEVAL5_ipd : std_ulogic := 'X';
  signal AEVAL4_ipd : std_ulogic := 'X';
  signal AEVAL3_ipd : std_ulogic := 'X';
  signal AEVAL2_ipd : std_ulogic := 'X';
  signal AEVAL1_ipd : std_ulogic := 'X';
  signal AEVAL0_ipd : std_ulogic := 'X';
  signal AFVAL7_ipd : std_ulogic := 'X';
  signal AFVAL6_ipd : std_ulogic := 'X';
  signal AFVAL5_ipd : std_ulogic := 'X';
  signal AFVAL4_ipd : std_ulogic := 'X';
  signal AFVAL3_ipd : std_ulogic := 'X';
  signal AFVAL2_ipd : std_ulogic := 'X';
  signal AFVAL1_ipd : std_ulogic := 'X';
  signal AFVAL0_ipd : std_ulogic := 'X';
  signal REN_ipd    : std_ulogic := 'X';
  signal RCLK_ipd   : std_ulogic := 'X';
  signal WD35_ipd   : std_ulogic := 'X';
  signal WD34_ipd   : std_ulogic := 'X';
  signal WD33_ipd   : std_ulogic := 'X';
  signal WD32_ipd   : std_ulogic := 'X';
  signal WD31_ipd   : std_ulogic := 'X';
  signal WD30_ipd   : std_ulogic := 'X';
  signal WD29_ipd   : std_ulogic := 'X';
  signal WD28_ipd   : std_ulogic := 'X';
  signal WD27_ipd   : std_ulogic := 'X';
  signal WD26_ipd   : std_ulogic := 'X';
  signal WD25_ipd   : std_ulogic := 'X';
  signal WD24_ipd   : std_ulogic := 'X';
  signal WD23_ipd   : std_ulogic := 'X';
  signal WD22_ipd   : std_ulogic := 'X';
  signal WD21_ipd   : std_ulogic := 'X';
  signal WD20_ipd   : std_ulogic := 'X';
  signal WD19_ipd   : std_ulogic := 'X';
  signal WD18_ipd   : std_ulogic := 'X';
  signal WD17_ipd   : std_ulogic := 'X';
  signal WD16_ipd   : std_ulogic := 'X';
  signal WD15_ipd   : std_ulogic := 'X';
  signal WD14_ipd   : std_ulogic := 'X';
  signal WD13_ipd   : std_ulogic := 'X';
  signal WD12_ipd   : std_ulogic := 'X';
  signal WD11_ipd   : std_ulogic := 'X';
  signal WD10_ipd   : std_ulogic := 'X';
  signal WD9_ipd    : std_ulogic := 'X';
  signal WD8_ipd    : std_ulogic := 'X';
  signal WD7_ipd    : std_ulogic := 'X';
  signal WD6_ipd    : std_ulogic := 'X';
  signal WD5_ipd    : std_ulogic := 'X';
  signal WD4_ipd    : std_ulogic := 'X';
  signal WD3_ipd    : std_ulogic := 'X';
  signal WD2_ipd    : std_ulogic := 'X';
  signal WD1_ipd    : std_ulogic := 'X';
  signal WD0_ipd    : std_ulogic := 'X';
  signal WEN_ipd    : std_ulogic := 'X';
  signal WCLK_ipd   : std_ulogic := 'X';
  signal CLR_ipd    : std_ulogic := '1';
  type MEM is array(0 to 65535) of std_ulogic_vector(35 downto 0);
  --signal RAM_TMP : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (DEPTH3_ipd, DEPTH3, VitalExtendToFillDelay(tipd_DEPTH3));
    VitalWireDelay (DEPTH2_ipd, DEPTH2, VitalExtendToFillDelay(tipd_DEPTH2));
    VitalWireDelay (DEPTH1_ipd, DEPTH1, VitalExtendToFillDelay(tipd_DEPTH1));
    VitalWireDelay (DEPTH0_ipd, DEPTH0, VitalExtendToFillDelay(tipd_DEPTH0));
    VitalWireDelay (WIDTH2_ipd, WIDTH2, VitalExtendToFillDelay(tipd_WIDTH2));
    VitalWireDelay (WIDTH1_ipd, WIDTH1, VitalExtendToFillDelay(tipd_WIDTH1));
    VitalWireDelay (WIDTH0_ipd, WIDTH0, VitalExtendToFillDelay(tipd_WIDTH0));
    VitalWireDelay (AEVAL7_ipd, AEVAL7, VitalExtendToFillDelay(tipd_AEVAL7));
    VitalWireDelay (AEVAL6_ipd, AEVAL6, VitalExtendToFillDelay(tipd_AEVAL6));
    VitalWireDelay (AEVAL5_ipd, AEVAL5, VitalExtendToFillDelay(tipd_AEVAL5));
    VitalWireDelay (AEVAL4_ipd, AEVAL4, VitalExtendToFillDelay(tipd_AEVAL4));
    VitalWireDelay (AEVAL3_ipd, AEVAL3, VitalExtendToFillDelay(tipd_AEVAL3));
    VitalWireDelay (AEVAL2_ipd, AEVAL2, VitalExtendToFillDelay(tipd_AEVAL2));
    VitalWireDelay (AEVAL1_ipd, AEVAL1, VitalExtendToFillDelay(tipd_AEVAL1));
    VitalWireDelay (AEVAL0_ipd, AEVAL0, VitalExtendToFillDelay(tipd_AEVAL0));
    VitalWireDelay (AFVAL7_ipd, AFVAL7, VitalExtendToFillDelay(tipd_AFVAL7));
    VitalWireDelay (AFVAL6_ipd, AFVAL6, VitalExtendToFillDelay(tipd_AFVAL6));
    VitalWireDelay (AFVAL5_ipd, AFVAL5, VitalExtendToFillDelay(tipd_AFVAL5));
    VitalWireDelay (AFVAL4_ipd, AFVAL4, VitalExtendToFillDelay(tipd_AFVAL4));
    VitalWireDelay (AFVAL3_ipd, AFVAL3, VitalExtendToFillDelay(tipd_AFVAL3));
    VitalWireDelay (AFVAL2_ipd, AFVAL2, VitalExtendToFillDelay(tipd_AFVAL2));
    VitalWireDelay (AFVAL1_ipd, AFVAL1, VitalExtendToFillDelay(tipd_AFVAL1));
    VitalWireDelay (AFVAL0_ipd, AFVAL0, VitalExtendToFillDelay(tipd_AFVAL0));
    VitalWireDelay (REN_ipd, REN, VitalExtendToFillDelay(tipd_REN));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
    VitalWireDelay (WD35_ipd, WD35, VitalExtendToFillDelay(tipd_WD35));
    VitalWireDelay (WD34_ipd, WD34, VitalExtendToFillDelay(tipd_WD34));
    VitalWireDelay (WD33_ipd, WD33, VitalExtendToFillDelay(tipd_WD33));
    VitalWireDelay (WD32_ipd, WD32, VitalExtendToFillDelay(tipd_WD32));
    VitalWireDelay (WD31_ipd, WD31, VitalExtendToFillDelay(tipd_WD31));
    VitalWireDelay (WD30_ipd, WD30, VitalExtendToFillDelay(tipd_WD30));
    VitalWireDelay (WD29_ipd, WD29, VitalExtendToFillDelay(tipd_WD29));
    VitalWireDelay (WD28_ipd, WD28, VitalExtendToFillDelay(tipd_WD28));
    VitalWireDelay (WD27_ipd, WD27, VitalExtendToFillDelay(tipd_WD27));
    VitalWireDelay (WD26_ipd, WD26, VitalExtendToFillDelay(tipd_WD26));
    VitalWireDelay (WD25_ipd, WD25, VitalExtendToFillDelay(tipd_WD25));
    VitalWireDelay (WD24_ipd, WD24, VitalExtendToFillDelay(tipd_WD24));
    VitalWireDelay (WD23_ipd, WD23, VitalExtendToFillDelay(tipd_WD23));
    VitalWireDelay (WD22_ipd, WD22, VitalExtendToFillDelay(tipd_WD22));
    VitalWireDelay (WD21_ipd, WD21, VitalExtendToFillDelay(tipd_WD21));
    VitalWireDelay (WD20_ipd, WD20, VitalExtendToFillDelay(tipd_WD20));
    VitalWireDelay (WD19_ipd, WD19, VitalExtendToFillDelay(tipd_WD19));
    VitalWireDelay (WD18_ipd, WD18, VitalExtendToFillDelay(tipd_WD18));
    VitalWireDelay (WD17_ipd, WD17, VitalExtendToFillDelay(tipd_WD17));
    VitalWireDelay (WD16_ipd, WD16, VitalExtendToFillDelay(tipd_WD16));
    VitalWireDelay (WD15_ipd, WD15, VitalExtendToFillDelay(tipd_WD15));
    VitalWireDelay (WD14_ipd, WD14, VitalExtendToFillDelay(tipd_WD14));
    VitalWireDelay (WD13_ipd, WD13, VitalExtendToFillDelay(tipd_WD13));
    VitalWireDelay (WD12_ipd, WD12, VitalExtendToFillDelay(tipd_WD12));
    VitalWireDelay (WD11_ipd, WD11, VitalExtendToFillDelay(tipd_WD11));
    VitalWireDelay (WD10_ipd, WD10, VitalExtendToFillDelay(tipd_WD10));
    VitalWireDelay (WD9_ipd, WD9, VitalExtendToFillDelay(tipd_WD9));
    VitalWireDelay (WD8_ipd, WD8, VitalExtendToFillDelay(tipd_WD8));
    VitalWireDelay (WD7_ipd, WD7, VitalExtendToFillDelay(tipd_WD7));
    VitalWireDelay (WD6_ipd, WD6, VitalExtendToFillDelay(tipd_WD6));
    VitalWireDelay (WD5_ipd, WD5, VitalExtendToFillDelay(tipd_WD5));
    VitalWireDelay (WD4_ipd, WD4, VitalExtendToFillDelay(tipd_WD4));
    VitalWireDelay (WD3_ipd, WD3, VitalExtendToFillDelay(tipd_WD3));
    VitalWireDelay (WD2_ipd, WD2, VitalExtendToFillDelay(tipd_WD2));
    VitalWireDelay (WD1_ipd, WD1, VitalExtendToFillDelay(tipd_WD1));
    VitalWireDelay (WD0_ipd, WD0, VitalExtendToFillDelay(tipd_WD0));
    VitalWireDelay (WEN_ipd, WEN, VitalExtendToFillDelay(tipd_WEN));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (CLR_ipd, CLR, VitalExtendToFillDelay(tipd_CLR));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (
                DEPTH3_ipd, DEPTH2_ipd, DEPTH1_ipd, DEPTH0_ipd, 
                WIDTH2_ipd, WIDTH1_ipd, WIDTH0_ipd,
                AEVAL7_ipd, AEVAL6_ipd, AEVAL5_ipd, AEVAL4_ipd, AEVAL3_ipd, 
                AEVAL2_ipd, AEVAL1_ipd, AEVAL0_ipd,
                AFVAL7_ipd, AFVAL6_ipd, AFVAL5_ipd, AFVAL4_ipd, AFVAL3_ipd, 
                AFVAL2_ipd, AFVAL1_ipd, AFVAL0_ipd,
                REN_ipd, RCLK_ipd,
                WD35_ipd, WD34_ipd, WD33_ipd, WD32_ipd, WD31_ipd, WD30_ipd,
                WD29_ipd, WD28_ipd, WD27_ipd, WD26_ipd, WD25_ipd, WD24_ipd,
                WD23_ipd, WD22_ipd, WD21_ipd, WD20_ipd, WD19_ipd, WD18_ipd,
                WD17_ipd, WD16_ipd, WD15_ipd, WD14_ipd, WD13_ipd, WD12_ipd,
                WD11_ipd, WD10_ipd, WD9_ipd, WD8_ipd, WD7_ipd, WD6_ipd,
                WD5_ipd, WD4_ipd, WD3_ipd, WD2_ipd, WD1_ipd, WD0_ipd,
                WEN_ipd, WCLK_ipd, CLR_ipd
                )

     --  Memory
     variable RAM_TMP : MEM;
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     --constant INT : SL_TO_INT := (-257, -257, 0, 1, -257, -257, 0, 1, -257);
     constant INT : SL_TO_INT := (-65537, -65537, 0, 1, -65537, -65537, 0, 1, -65537);

     --  Read Timing Check Results
     variable Tviol_DEPTH3_RCLK_posedge : X01 := '0';
     variable TmDt_DEPTH3_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DEPTH2_RCLK_posedge : X01 := '0';
     variable TmDt_DEPTH2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DEPTH1_RCLK_posedge : X01 := '0';
     variable TmDt_DEPTH1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DEPTH0_RCLK_posedge : X01 := '0';
     variable TmDt_DEPTH0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WIDTH2_RCLK_posedge : X01 := '0';
     variable TmDt_WIDTH2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WIDTH1_RCLK_posedge : X01 := '0';
     variable TmDt_WIDTH1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WIDTH0_RCLK_posedge : X01 := '0';
     variable TmDt_WIDTH0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AEVAL7_RCLK_posedge : X01 := '0';
     variable TmDt_AEVAL7_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AEVAL6_RCLK_posedge : X01 := '0';
     variable TmDt_AEVAL6_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AEVAL5_RCLK_posedge : X01 := '0';
     variable TmDt_AEVAL5_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AEVAL4_RCLK_posedge : X01 := '0';
     variable TmDt_AEVAL4_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AEVAL3_RCLK_posedge : X01 := '0';
     variable TmDt_AEVAL3_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AEVAL2_RCLK_posedge : X01 := '0';
     variable TmDt_AEVAL2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AEVAL1_RCLK_posedge : X01 := '0';
     variable TmDt_AEVAL1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AEVAL0_RCLK_posedge : X01 := '0';
     variable TmDt_AEVAL0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AFVAL7_RCLK_posedge : X01 := '0';
     variable TmDt_AFVAL7_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AFVAL6_RCLK_posedge : X01 := '0';
     variable TmDt_AFVAL6_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AFVAL5_RCLK_posedge : X01 := '0';
     variable TmDt_AFVAL5_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AFVAL4_RCLK_posedge : X01 := '0';
     variable TmDt_AFVAL4_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AFVAL3_RCLK_posedge : X01 := '0';
     variable TmDt_AFVAL3_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AFVAL2_RCLK_posedge : X01 := '0';
     variable TmDt_AFVAL2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AFVAL1_RCLK_posedge : X01 := '0';
     variable TmDt_AFVAL1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AFVAL0_RCLK_posedge : X01 := '0';
     variable TmDt_AFVAL0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_REN_RCLK_posedge : X01 := '0';
     variable TmDt_REN_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_CLR_RCLK_posedge : X01 := '0';
     variable Tmkr_CLR_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_DEPTH3_WCLK_posedge : X01 := '0';
     variable TmDt_DEPTH3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DEPTH2_WCLK_posedge : X01 := '0';
     variable TmDt_DEPTH2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DEPTH1_WCLK_posedge : X01 := '0';
     variable TmDt_DEPTH1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DEPTH0_WCLK_posedge : X01 := '0';
     variable TmDt_DEPTH0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WIDTH2_WCLK_posedge : X01 := '0';
     variable TmDt_WIDTH2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WIDTH1_WCLK_posedge : X01 := '0';
     variable TmDt_WIDTH1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WIDTH0_WCLK_posedge : X01 := '0';
     variable TmDt_WIDTH0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AEVAL7_WCLK_posedge : X01 := '0';
     variable TmDt_AEVAL7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AEVAL6_WCLK_posedge : X01 := '0';
     variable TmDt_AEVAL6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AEVAL5_WCLK_posedge : X01 := '0';
     variable TmDt_AEVAL5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AEVAL4_WCLK_posedge : X01 := '0';
     variable TmDt_AEVAL4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AEVAL3_WCLK_posedge : X01 := '0';
     variable TmDt_AEVAL3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AEVAL2_WCLK_posedge : X01 := '0';
     variable TmDt_AEVAL2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AEVAL1_WCLK_posedge : X01 := '0';
     variable TmDt_AEVAL1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AEVAL0_WCLK_posedge : X01 := '0';
     variable TmDt_AEVAL0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AFVAL7_WCLK_posedge : X01 := '0';
     variable TmDt_AFVAL7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AFVAL6_WCLK_posedge : X01 := '0';
     variable TmDt_AFVAL6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AFVAL5_WCLK_posedge : X01 := '0';
     variable TmDt_AFVAL5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AFVAL4_WCLK_posedge : X01 := '0';
     variable TmDt_AFVAL4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AFVAL3_WCLK_posedge : X01 := '0';
     variable TmDt_AFVAL3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AFVAL2_WCLK_posedge : X01 := '0';
     variable TmDt_AFVAL2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AFVAL1_WCLK_posedge : X01 := '0';
     variable TmDt_AFVAL1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_AFVAL0_WCLK_posedge : X01 := '0';
     variable TmDt_AFVAL0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD35_WCLK_posedge : X01 := '0';
     variable TmDt_WD35_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD34_WCLK_posedge : X01 := '0';
     variable TmDt_WD34_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD33_WCLK_posedge : X01 := '0';
     variable TmDt_WD33_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD32_WCLK_posedge : X01 := '0';
     variable TmDt_WD32_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD31_WCLK_posedge : X01 := '0';
     variable TmDt_WD31_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD30_WCLK_posedge : X01 := '0';
     variable TmDt_WD30_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD29_WCLK_posedge : X01 := '0';
     variable TmDt_WD29_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD28_WCLK_posedge : X01 := '0';
     variable TmDt_WD28_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD27_WCLK_posedge : X01 := '0';
     variable TmDt_WD27_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD26_WCLK_posedge : X01 := '0';
     variable TmDt_WD26_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD25_WCLK_posedge : X01 := '0';
     variable TmDt_WD25_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD24_WCLK_posedge : X01 := '0';
     variable TmDt_WD24_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD23_WCLK_posedge : X01 := '0';
     variable TmDt_WD23_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD22_WCLK_posedge : X01 := '0';
     variable TmDt_WD22_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD21_WCLK_posedge : X01 := '0';
     variable TmDt_WD21_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD20_WCLK_posedge : X01 := '0';
     variable TmDt_WD20_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD19_WCLK_posedge : X01 := '0';
     variable TmDt_WD19_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD18_WCLK_posedge : X01 := '0';
     variable TmDt_WD18_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD17_WCLK_posedge : X01 := '0';
     variable TmDt_WD17_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD16_WCLK_posedge : X01 := '0';
     variable TmDt_WD16_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD15_WCLK_posedge : X01 := '0';
     variable TmDt_WD15_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD14_WCLK_posedge : X01 := '0';
     variable TmDt_WD14_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD13_WCLK_posedge : X01 := '0';
     variable TmDt_WD13_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD12_WCLK_posedge : X01 := '0';
     variable TmDt_WD12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD11_WCLK_posedge : X01 := '0';
     variable TmDt_WD11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD10_WCLK_posedge : X01 := '0';
     variable TmDt_WD10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD9_WCLK_posedge : X01 := '0';
     variable TmDt_WD9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD8_WCLK_posedge : X01 := '0';
     variable TmDt_WD8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD7_WCLK_posedge : X01 := '0';
     variable TmDt_WD7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD6_WCLK_posedge : X01 := '0';
     variable TmDt_WD6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD5_WCLK_posedge : X01 := '0';
     variable TmDt_WD5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD4_WCLK_posedge : X01 := '0';
     variable TmDt_WD4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD3_WCLK_posedge : X01 := '0';
     variable TmDt_WD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD2_WCLK_posedge : X01 := '0';
     variable TmDt_WD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD1_WCLK_posedge : X01 := '0';
     variable TmDt_WD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD0_WCLK_posedge : X01 := '0';
     variable TmDt_WD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WEN_WCLK_posedge : X01 := '0';
     variable TmDt_WEN_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_CLR_WCLK_posedge : X01 := '0';
     variable Tmkr_CLR_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_CLR : X01 := '0';
     variable PeriodData_CLR : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  Functional Results
     variable WADDR : integer :=0;
     variable WADDR_P1 : integer :=0;
     variable WADDR_P2 : integer :=0;
     variable WADDR_wrap : integer :=0;
     variable RADDR : integer :=0;
     variable RADDR_P1: integer :=0;
     variable RADDR_P2 : integer :=0;
     variable RADDR_wrap : integer :=0;
     variable AEVAL : integer := 0; -- Almost empty threshold value
     variable AFVAL : integer := 0; -- Almost full threshold value
     variable AEVAL_temp : integer := 0;
     variable AFVAL_temp : integer := 0;
     variable WWIDTH : integer := -1; -- Word width
     variable HEIGTH : integer := -1; -- Word heigth
     variable DIVID  : integer := 1;  -- used to calculate the Almost FULL/EMPTY value 
     variable WDEPTH : integer := -1; -- Word depth
     variable MAX_ADDR : integer := -1; -- Maximum memory address
     variable MEM_USED : integer := 0; -- Memory addresses used
    
     variable WEN_int : std_ulogic;
     variable REN_int : std_ulogic; 
     variable RD35_zd : std_ulogic;
     variable RD34_zd : std_ulogic;
     variable RD33_zd : std_ulogic;
     variable RD32_zd : std_ulogic;
     variable RD31_zd : std_ulogic;
     variable RD30_zd : std_ulogic;
     variable RD29_zd : std_ulogic;
     variable RD28_zd : std_ulogic;
     variable RD27_zd : std_ulogic;
     variable RD26_zd : std_ulogic;
     variable RD25_zd : std_ulogic;
     variable RD24_zd : std_ulogic;
     variable RD23_zd : std_ulogic;
     variable RD22_zd : std_ulogic;
     variable RD21_zd : std_ulogic;
     variable RD20_zd : std_ulogic;
     variable RD19_zd : std_ulogic;
     variable RD18_zd : std_ulogic;
     variable RD17_zd : std_ulogic;
     variable RD16_zd : std_ulogic;
     variable RD15_zd : std_ulogic;
     variable RD14_zd : std_ulogic;
     variable RD13_zd : std_ulogic;
     variable RD12_zd : std_ulogic;
     variable RD11_zd : std_ulogic;
     variable RD10_zd : std_ulogic;
     variable RD9_zd : std_ulogic;
     variable RD8_zd : std_ulogic;
     variable RD7_zd : std_ulogic;
     variable RD6_zd : std_ulogic;
     variable RD5_zd : std_ulogic;
     variable RD4_zd : std_ulogic;
     variable RD3_zd : std_ulogic;
     variable RD2_zd : std_ulogic;
     variable RD1_zd : std_ulogic;
     variable RD0_zd : std_ulogic;
     variable FULL_zd : std_ulogic;
     variable AFULL_zd : std_ulogic;
     variable EMPTY_zd : std_ulogic;
     variable AEMPTY_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable RD35_GlitchData : VitalGlitchDataType;
     variable RD34_GlitchData : VitalGlitchDataType;
     variable RD33_GlitchData : VitalGlitchDataType;
     variable RD32_GlitchData : VitalGlitchDataType;
     variable RD31_GlitchData : VitalGlitchDataType;
     variable RD30_GlitchData : VitalGlitchDataType;
     variable RD29_GlitchData : VitalGlitchDataType;
     variable RD28_GlitchData : VitalGlitchDataType;
     variable RD27_GlitchData : VitalGlitchDataType;
     variable RD26_GlitchData : VitalGlitchDataType;
     variable RD25_GlitchData : VitalGlitchDataType;
     variable RD24_GlitchData : VitalGlitchDataType;
     variable RD23_GlitchData : VitalGlitchDataType;
     variable RD22_GlitchData : VitalGlitchDataType;
     variable RD21_GlitchData : VitalGlitchDataType;
     variable RD20_GlitchData : VitalGlitchDataType;
     variable RD19_GlitchData : VitalGlitchDataType;
     variable RD18_GlitchData : VitalGlitchDataType;
     variable RD17_GlitchData : VitalGlitchDataType;
     variable RD16_GlitchData : VitalGlitchDataType;
     variable RD15_GlitchData : VitalGlitchDataType;
     variable RD14_GlitchData : VitalGlitchDataType;
     variable RD13_GlitchData : VitalGlitchDataType;
     variable RD12_GlitchData : VitalGlitchDataType;
     variable RD11_GlitchData : VitalGlitchDataType;
     variable RD10_GlitchData : VitalGlitchDataType;
     variable RD9_GlitchData : VitalGlitchDataType;
     variable RD8_GlitchData : VitalGlitchDataType;
     variable RD7_GlitchData : VitalGlitchDataType;
     variable RD6_GlitchData : VitalGlitchDataType;
     variable RD5_GlitchData : VitalGlitchDataType;
     variable RD4_GlitchData : VitalGlitchDataType;
     variable RD3_GlitchData : VitalGlitchDataType;
     variable RD2_GlitchData : VitalGlitchDataType;
     variable RD1_GlitchData : VitalGlitchDataType;
     variable RD0_GlitchData : VitalGlitchDataType;
     variable FULL_GlitchData : VitalGlitchDataType;
     variable AFULL_GlitchData : VitalGlitchDataType;
     variable EMPTY_GlitchData : VitalGlitchDataType;
     variable AEMPTY_GlitchData : VitalGlitchDataType;

     -- Last value variables
     variable DEPTH3_delayed : std_ulogic := 'X';
     variable DEPTH2_delayed : std_ulogic := 'X';
     variable DEPTH1_delayed : std_ulogic := 'X';
     variable DEPTH0_delayed : std_ulogic := 'X';
     variable WIDTH2_delayed : std_ulogic := 'X';
     variable WIDTH1_delayed : std_ulogic := 'X';
     variable WIDTH0_delayed : std_ulogic := 'X';
     variable AEVAL7_delayed : std_ulogic := 'X';
     variable AEVAL6_delayed : std_ulogic := 'X';
     variable AEVAL5_delayed : std_ulogic := 'X';
     variable AEVAL4_delayed : std_ulogic := 'X';
     variable AEVAL3_delayed : std_ulogic := 'X';
     variable AEVAL2_delayed : std_ulogic := 'X';
     variable AEVAL1_delayed : std_ulogic := 'X';
     variable AEVAL0_delayed : std_ulogic := 'X';
     variable AFVAL7_delayed : std_ulogic := 'X';
     variable AFVAL6_delayed : std_ulogic := 'X';
     variable AFVAL5_delayed : std_ulogic := 'X';
     variable AFVAL4_delayed : std_ulogic := 'X';
     variable AFVAL3_delayed : std_ulogic := 'X';
     variable AFVAL2_delayed : std_ulogic := 'X';
     variable AFVAL1_delayed : std_ulogic := 'X';
     variable AFVAL0_delayed : std_ulogic := 'X';
     variable REN_delayed   : std_ulogic := 'X';
     variable REN_previous  : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable WD35_delayed : std_ulogic := 'X';
     variable WD34_delayed : std_ulogic := 'X';
     variable WD33_delayed : std_ulogic := 'X';
     variable WD32_delayed : std_ulogic := 'X';
     variable WD31_delayed : std_ulogic := 'X';
     variable WD30_delayed : std_ulogic := 'X';
     variable WD29_delayed : std_ulogic := 'X';
     variable WD28_delayed : std_ulogic := 'X';
     variable WD27_delayed : std_ulogic := 'X';
     variable WD26_delayed : std_ulogic := 'X';
     variable WD25_delayed : std_ulogic := 'X';
     variable WD24_delayed : std_ulogic := 'X';
     variable WD23_delayed : std_ulogic := 'X';
     variable WD22_delayed : std_ulogic := 'X';
     variable WD21_delayed : std_ulogic := 'X';
     variable WD20_delayed : std_ulogic := 'X';
     variable WD19_delayed : std_ulogic := 'X';
     variable WD18_delayed : std_ulogic := 'X';
     variable WD17_delayed : std_ulogic := 'X';
     variable WD16_delayed : std_ulogic := 'X';
     variable WD15_delayed : std_ulogic := 'X';
     variable WD14_delayed : std_ulogic := 'X';
     variable WD13_delayed : std_ulogic := 'X';
     variable WD12_delayed : std_ulogic := 'X';
     variable WD11_delayed : std_ulogic := 'X';
     variable WD10_delayed : std_ulogic := 'X';
     variable WD9_delayed : std_ulogic := 'X';
     variable WD8_delayed : std_ulogic := 'X';
     variable WD7_delayed : std_ulogic := 'X';
     variable WD6_delayed : std_ulogic := 'X';
     variable WD5_delayed : std_ulogic := 'X';
     variable WD4_delayed : std_ulogic := 'X';
     variable WD3_delayed : std_ulogic := 'X';
     variable WD2_delayed : std_ulogic := 'X';
     variable WD1_delayed : std_ulogic := 'X';
     variable WD0_delayed : std_ulogic := 'X';
     variable WEN_delayed   : std_ulogic := 'X';
     variable WEN_previous  : std_ulogic := 'X';
     variable WCLK_previous : std_ulogic := 'X';

  begin  --  process VITALBehavior 
    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup DEPTH high or low before RCLK rising
      --   Hold  DEPTH high or low after RCLK rising

      VitalSetupHoldCheck ( Tviol_DEPTH3_RCLK_posedge,
                            TmDt_DEPTH3_RCLK_posedge,
                            DEPTH3_ipd, "DEPTH3",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_DEPTH3_RCLK_posedge_posedge,
                            tsetup_DEPTH3_RCLK_negedge_posedge,
                            thold_DEPTH3_RCLK_posedge_posedge,
                            thold_DEPTH3_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_DEPTH2_RCLK_posedge,
                            TmDt_DEPTH2_RCLK_posedge,
                            DEPTH2_ipd, "DEPTH2",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_DEPTH2_RCLK_posedge_posedge,
                            tsetup_DEPTH2_RCLK_negedge_posedge,
                            thold_DEPTH2_RCLK_posedge_posedge,
                            thold_DEPTH2_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_DEPTH1_RCLK_posedge,
                            TmDt_DEPTH1_RCLK_posedge,
                            DEPTH1_ipd, "DEPTH1",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_DEPTH1_RCLK_posedge_posedge,
                            tsetup_DEPTH1_RCLK_negedge_posedge,
                            thold_DEPTH1_RCLK_posedge_posedge,
                            thold_DEPTH1_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_DEPTH0_RCLK_posedge,
                            TmDt_DEPTH0_RCLK_posedge,
                            DEPTH0_ipd, "DEPTH0",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_DEPTH0_RCLK_posedge_posedge,
                            tsetup_DEPTH0_RCLK_negedge_posedge,
                            thold_DEPTH0_RCLK_posedge_posedge,
                            thold_DEPTH0_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup WIDTH high or low before RCLK rising
      --   Hold  WIDTH high or low after RCLK rising

      VitalSetupHoldCheck ( Tviol_WIDTH2_RCLK_posedge,
                            TmDt_WIDTH2_RCLK_posedge,
                            WIDTH2_ipd, "WIDTH2",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_WIDTH2_RCLK_posedge_posedge,
                            tsetup_WIDTH2_RCLK_negedge_posedge,
                            thold_WIDTH2_RCLK_posedge_posedge,
                            thold_WIDTH2_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WIDTH1_RCLK_posedge,
                            TmDt_WIDTH1_RCLK_posedge,
                            WIDTH1_ipd, "WIDTH1",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_WIDTH1_RCLK_posedge_posedge,
                            tsetup_WIDTH1_RCLK_negedge_posedge,
                            thold_WIDTH1_RCLK_posedge_posedge,
                            thold_WIDTH1_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WIDTH0_RCLK_posedge,
                            TmDt_WIDTH0_RCLK_posedge,
                            WIDTH0_ipd, "WIDTH0",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_WIDTH0_RCLK_posedge_posedge,
                            tsetup_WIDTH0_RCLK_negedge_posedge,
                            thold_WIDTH0_RCLK_posedge_posedge,
                            thold_WIDTH0_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup AEVAL high or low before RCLK rising
      --   Hold  AEVAL high or low after RCLK rising

      VitalSetupHoldCheck ( Tviol_AEVAL7_RCLK_posedge,
                            TmDt_AEVAL7_RCLK_posedge,
                            AEVAL7_ipd, "AEVAL7",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_AEVAL7_RCLK_posedge_posedge,
                            tsetup_AEVAL7_RCLK_negedge_posedge,
                            thold_AEVAL7_RCLK_posedge_posedge,
                            thold_AEVAL7_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AEVAL6_RCLK_posedge,
                            TmDt_AEVAL6_RCLK_posedge,
                            AEVAL6_ipd, "AEVAL6",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_AEVAL6_RCLK_posedge_posedge,
                            tsetup_AEVAL6_RCLK_negedge_posedge,
                            thold_AEVAL6_RCLK_posedge_posedge,
                            thold_AEVAL6_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AEVAL5_RCLK_posedge,
                            TmDt_AEVAL5_RCLK_posedge,
                            AEVAL5_ipd, "AEVAL5",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_AEVAL5_RCLK_posedge_posedge,
                            tsetup_AEVAL5_RCLK_negedge_posedge,
                            thold_AEVAL5_RCLK_posedge_posedge,
                            thold_AEVAL5_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AEVAL4_RCLK_posedge,
                            TmDt_AEVAL4_RCLK_posedge,
                            AEVAL4_ipd, "AEVAL4",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_AEVAL4_RCLK_posedge_posedge,
                            tsetup_AEVAL4_RCLK_negedge_posedge,
                            thold_AEVAL4_RCLK_posedge_posedge,
                            thold_AEVAL4_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AEVAL3_RCLK_posedge,
                            TmDt_AEVAL3_RCLK_posedge,
                            AEVAL3_ipd, "AEVAL3",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_AEVAL3_RCLK_posedge_posedge,
                            tsetup_AEVAL3_RCLK_negedge_posedge,
                            thold_AEVAL3_RCLK_posedge_posedge,
                            thold_AEVAL3_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AEVAL2_RCLK_posedge,
                            TmDt_AEVAL2_RCLK_posedge,
                            AEVAL2_ipd, "AEVAL2",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_AEVAL2_RCLK_posedge_posedge,
                            tsetup_AEVAL2_RCLK_negedge_posedge,
                            thold_AEVAL2_RCLK_posedge_posedge,
                            thold_AEVAL2_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AEVAL1_RCLK_posedge,
                            TmDt_AEVAL1_RCLK_posedge,
                            AEVAL1_ipd, "AEVAL1",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_AEVAL1_RCLK_posedge_posedge,
                            tsetup_AEVAL1_RCLK_negedge_posedge,
                            thold_AEVAL1_RCLK_posedge_posedge,
                            thold_AEVAL1_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AEVAL0_RCLK_posedge,
                            TmDt_AEVAL0_RCLK_posedge,
                            AEVAL0_ipd, "AEVAL0",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_AEVAL0_RCLK_posedge_posedge,
                            tsetup_AEVAL0_RCLK_negedge_posedge,
                            thold_AEVAL0_RCLK_posedge_posedge,
                            thold_AEVAL0_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup AFVAL high before RCLK rising
      --   Hold  AFVAL high after RCLK rising

      VitalSetupHoldCheck ( Tviol_AFVAL7_RCLK_posedge,
                            TmDt_AFVAL7_RCLK_posedge,
                            AFVAL7_ipd, "AFVAL7",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_AFVAL7_RCLK_posedge_posedge,
                            tsetup_AFVAL7_RCLK_negedge_posedge,
                            thold_AFVAL7_RCLK_posedge_posedge,
                            thold_AFVAL7_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AFVAL6_RCLK_posedge,
                            TmDt_AFVAL6_RCLK_posedge,
                            AFVAL6_ipd, "AFVAL6",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_AFVAL6_RCLK_posedge_posedge,
                            tsetup_AFVAL6_RCLK_negedge_posedge,
                            thold_AFVAL6_RCLK_posedge_posedge,
                            thold_AFVAL6_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AFVAL5_RCLK_posedge,
                            TmDt_AFVAL5_RCLK_posedge,
                            AFVAL5_ipd, "AFVAL5",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_AFVAL5_RCLK_posedge_posedge,
                            tsetup_AFVAL5_RCLK_negedge_posedge,
                            thold_AFVAL5_RCLK_posedge_posedge,
                            thold_AFVAL5_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AFVAL4_RCLK_posedge,
                            TmDt_AFVAL4_RCLK_posedge,
                            AFVAL4_ipd, "AFVAL4",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_AFVAL4_RCLK_posedge_posedge,
                            tsetup_AFVAL4_RCLK_negedge_posedge,
                            thold_AFVAL4_RCLK_posedge_posedge,
                            thold_AFVAL4_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AFVAL3_RCLK_posedge,
                            TmDt_AFVAL3_RCLK_posedge,
                            AFVAL3_ipd, "AFVAL3",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_AFVAL3_RCLK_posedge_posedge,
                            tsetup_AFVAL3_RCLK_negedge_posedge,
                            thold_AFVAL3_RCLK_posedge_posedge,
                            thold_AFVAL3_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AFVAL2_RCLK_posedge,
                            TmDt_AFVAL2_RCLK_posedge,
                            AFVAL2_ipd, "AFVAL2",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_AFVAL2_RCLK_posedge_posedge,
                            tsetup_AFVAL2_RCLK_negedge_posedge,
                            thold_AFVAL2_RCLK_posedge_posedge,
                            thold_AFVAL2_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AFVAL1_RCLK_posedge,
                            TmDt_AFVAL1_RCLK_posedge,
                            AFVAL1_ipd, "AFVAL1",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_AFVAL1_RCLK_posedge_posedge,
                            tsetup_AFVAL1_RCLK_negedge_posedge,
                            thold_AFVAL1_RCLK_posedge_posedge,
                            thold_AFVAL1_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AFVAL0_RCLK_posedge,
                            TmDt_AFVAL0_RCLK_posedge,
                            AFVAL0_ipd, "AFVAL0",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_AFVAL0_RCLK_posedge_posedge,
                            tsetup_AFVAL0_RCLK_negedge_posedge,
                            thold_AFVAL0_RCLK_posedge_posedge,
                            thold_AFVAL0_RCLK_negedge_posedge,
                            ((To_X01(REN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup REN high before RCLK rising
      --   Hold  REN high after RCLK rising

      VitalSetupHoldCheck ( Tviol_REN_RCLK_posedge,
                            TmDt_REN_RCLK_posedge,
                            REN_ipd, "REN",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_REN_RCLK_posedge_posedge,
			    tsetup_REN_RCLK_negedge_posedge,
                            thold_REN_RCLK_posedge_posedge,
                            thold_REN_RCLK_negedge_posedge,
                            ((To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            ((To_X01(CLR_ipd)='0')),
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

     
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_RCLK_posedge,
          TimingData              => Tmkr_CLR_RCLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => RCLK_ipd,
          RefSignalName          => "RCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_RCLK_posedge_posedge,
          Removal                 => thold_CLR_RCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TimingCheckOn,
          RefTransition           => '/',
          HeaderMsg               => InstancePath & "/FIFO64K36",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);


      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup DEPTH high or low before WCLK rising
      --   Hold  DEPTH high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_DEPTH3_WCLK_posedge,
                            TmDt_DEPTH3_WCLK_posedge,
                            DEPTH3_ipd, "DEPTH3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_DEPTH3_WCLK_posedge_posedge,
                            tsetup_DEPTH3_WCLK_negedge_posedge,
                            thold_DEPTH3_WCLK_posedge_posedge,
                            thold_DEPTH3_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_DEPTH2_WCLK_posedge,
                            TmDt_DEPTH2_WCLK_posedge,
                            DEPTH2_ipd, "DEPTH2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_DEPTH2_WCLK_posedge_posedge,
                            tsetup_DEPTH2_WCLK_negedge_posedge,
                            thold_DEPTH2_WCLK_posedge_posedge,
                            thold_DEPTH2_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_DEPTH1_WCLK_posedge,
                            TmDt_DEPTH1_WCLK_posedge,
                            DEPTH1_ipd, "DEPTH1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_DEPTH1_WCLK_posedge_posedge,
                            tsetup_DEPTH1_WCLK_negedge_posedge,
                            thold_DEPTH1_WCLK_posedge_posedge,
                            thold_DEPTH1_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_DEPTH0_WCLK_posedge,
                            TmDt_DEPTH0_WCLK_posedge,
                            DEPTH0_ipd, "DEPTH0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_DEPTH0_WCLK_posedge_posedge,
                            tsetup_DEPTH0_WCLK_negedge_posedge,
                            thold_DEPTH0_WCLK_posedge_posedge,
                            thold_DEPTH0_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      --   Setup WIDTH high or low before WCLK rising
      --   Hold  WIDTH high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WIDTH2_WCLK_posedge,
                            TmDt_WIDTH2_WCLK_posedge,
                            WIDTH2_ipd, "WIDTH2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WIDTH2_WCLK_posedge_posedge,
                            tsetup_WIDTH2_WCLK_negedge_posedge,
                            thold_WIDTH2_WCLK_posedge_posedge,
                            thold_WIDTH2_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WIDTH1_WCLK_posedge,
                            TmDt_WIDTH1_WCLK_posedge,
                            WIDTH1_ipd, "WIDTH1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WIDTH1_WCLK_posedge_posedge,
                            tsetup_WIDTH1_WCLK_negedge_posedge,
                            thold_WIDTH1_WCLK_posedge_posedge,
                            thold_WIDTH1_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WIDTH0_WCLK_posedge,
                            TmDt_WIDTH0_WCLK_posedge,
                            WIDTH0_ipd, "WIDTH0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WIDTH0_WCLK_posedge_posedge,
                            tsetup_WIDTH0_WCLK_negedge_posedge,
                            thold_WIDTH0_WCLK_posedge_posedge,
                            thold_WIDTH0_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup AEVAL high or low before WCLK rising
      --   Hold  AEVAL high or low after WCLK rising

      VitalSetupHoldCheck ( Tviol_AEVAL7_WCLK_posedge,
                            TmDt_AEVAL7_WCLK_posedge,
                            AEVAL7_ipd, "AEVAL7",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_AEVAL7_WCLK_posedge_posedge,
                            tsetup_AEVAL7_WCLK_negedge_posedge,
                            thold_AEVAL7_WCLK_posedge_posedge,
                            thold_AEVAL7_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AEVAL6_WCLK_posedge,
                            TmDt_AEVAL6_WCLK_posedge,
                            AEVAL6_ipd, "AEVAL6",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_AEVAL6_WCLK_posedge_posedge,
                            tsetup_AEVAL6_WCLK_negedge_posedge,
                            thold_AEVAL6_WCLK_posedge_posedge,
                            thold_AEVAL6_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AEVAL5_WCLK_posedge,
                            TmDt_AEVAL5_WCLK_posedge,
                            AEVAL5_ipd, "AEVAL5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_AEVAL5_WCLK_posedge_posedge,
                            tsetup_AEVAL5_WCLK_negedge_posedge,
                            thold_AEVAL5_WCLK_posedge_posedge,
                            thold_AEVAL5_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AEVAL4_WCLK_posedge,
                            TmDt_AEVAL4_WCLK_posedge,
                            AEVAL4_ipd, "AEVAL4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_AEVAL4_WCLK_posedge_posedge,
                            tsetup_AEVAL4_WCLK_negedge_posedge,
                            thold_AEVAL4_WCLK_posedge_posedge,
                            thold_AEVAL4_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AEVAL3_WCLK_posedge,
                            TmDt_AEVAL3_WCLK_posedge,
                            AEVAL3_ipd, "AEVAL3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_AEVAL3_WCLK_posedge_posedge,
                            tsetup_AEVAL3_WCLK_negedge_posedge,
                            thold_AEVAL3_WCLK_posedge_posedge,
                            thold_AEVAL3_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AEVAL2_WCLK_posedge,
                            TmDt_AEVAL2_WCLK_posedge,
                            AEVAL2_ipd, "AEVAL2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_AEVAL2_WCLK_posedge_posedge,
                            tsetup_AEVAL2_WCLK_negedge_posedge,
                            thold_AEVAL2_WCLK_posedge_posedge,
                            thold_AEVAL2_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AEVAL1_WCLK_posedge,
                            TmDt_AEVAL1_WCLK_posedge,
                            AEVAL1_ipd, "AEVAL1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_AEVAL1_WCLK_posedge_posedge,
                            tsetup_AEVAL1_WCLK_negedge_posedge,
                            thold_AEVAL1_WCLK_posedge_posedge,
                            thold_AEVAL1_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AEVAL0_WCLK_posedge,
                            TmDt_AEVAL0_WCLK_posedge,
                            AEVAL0_ipd, "AEVAL0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_AEVAL0_WCLK_posedge_posedge,
                            tsetup_AEVAL0_WCLK_negedge_posedge,
                            thold_AEVAL0_WCLK_posedge_posedge,
                            thold_AEVAL0_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup AFVAL high before WCLK rising
      --   Hold  AFVAL high after WCLK rising

      VitalSetupHoldCheck ( Tviol_AFVAL7_WCLK_posedge,
                            TmDt_AFVAL7_WCLK_posedge,
                            AFVAL7_ipd, "AFVAL7",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_AFVAL7_WCLK_posedge_posedge,
                            tsetup_AFVAL7_WCLK_negedge_posedge,
                            thold_AFVAL7_WCLK_posedge_posedge,
                            thold_AFVAL7_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AFVAL6_WCLK_posedge,
                            TmDt_AFVAL6_WCLK_posedge,
                            AFVAL6_ipd, "AFVAL6",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_AFVAL6_WCLK_posedge_posedge,
                            tsetup_AFVAL6_WCLK_negedge_posedge,
                            thold_AFVAL6_WCLK_posedge_posedge,
                            thold_AFVAL6_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AFVAL5_WCLK_posedge,
                            TmDt_AFVAL5_WCLK_posedge,
                            AFVAL5_ipd, "AFVAL5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_AFVAL5_WCLK_posedge_posedge,
                            tsetup_AFVAL5_WCLK_negedge_posedge,
                            thold_AFVAL5_WCLK_posedge_posedge,
                            thold_AFVAL5_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AFVAL4_WCLK_posedge,
                            TmDt_AFVAL4_WCLK_posedge,
                            AFVAL4_ipd, "AFVAL4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_AFVAL4_WCLK_posedge_posedge,
                            tsetup_AFVAL4_WCLK_negedge_posedge,
                            thold_AFVAL4_WCLK_posedge_posedge,
                            thold_AFVAL4_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AFVAL3_WCLK_posedge,
                            TmDt_AFVAL3_WCLK_posedge,
                            AFVAL3_ipd, "AFVAL3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_AFVAL3_WCLK_posedge_posedge,
                            tsetup_AFVAL3_WCLK_negedge_posedge,
                            thold_AFVAL3_WCLK_posedge_posedge,
                            thold_AFVAL3_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AFVAL2_WCLK_posedge,
                            TmDt_AFVAL2_WCLK_posedge,
                            AFVAL2_ipd, "AFVAL2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_AFVAL2_WCLK_posedge_posedge,
                            tsetup_AFVAL2_WCLK_negedge_posedge,
                            thold_AFVAL2_WCLK_posedge_posedge,
                            thold_AFVAL2_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AFVAL1_WCLK_posedge,
                            TmDt_AFVAL1_WCLK_posedge,
                            AFVAL1_ipd, "AFVAL1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_AFVAL1_WCLK_posedge_posedge,
                            tsetup_AFVAL1_WCLK_negedge_posedge,
                            thold_AFVAL1_WCLK_posedge_posedge,
                            thold_AFVAL1_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_AFVAL0_WCLK_posedge,
                            TmDt_AFVAL0_WCLK_posedge,
                            AFVAL0_ipd, "AFVAL0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_AFVAL0_WCLK_posedge_posedge,
                            tsetup_AFVAL0_WCLK_negedge_posedge,
                            thold_AFVAL0_WCLK_posedge_posedge,
                            thold_AFVAL0_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup WD high or low before WCLK rising
      --   Hold  WD high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WD35_WCLK_posedge,
                            TmDt_WD35_WCLK_posedge,
                            WD35_ipd, "WD35",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD35_WCLK_posedge_posedge,
                            tsetup_WD35_WCLK_negedge_posedge,
                            thold_WD35_WCLK_posedge_posedge,
                            thold_WD35_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD34_WCLK_posedge,
                            TmDt_WD34_WCLK_posedge,
                            WD34_ipd, "WD34",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD34_WCLK_posedge_posedge,
                            tsetup_WD34_WCLK_negedge_posedge,
                            thold_WD34_WCLK_posedge_posedge,
                            thold_WD34_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD33_WCLK_posedge,
                            TmDt_WD33_WCLK_posedge,
                            WD33_ipd, "WD33",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD33_WCLK_posedge_posedge,
                            tsetup_WD33_WCLK_negedge_posedge,
                            thold_WD33_WCLK_posedge_posedge,
                            thold_WD33_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD32_WCLK_posedge,
                            TmDt_WD32_WCLK_posedge,
                            WD32_ipd, "WD32",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD32_WCLK_posedge_posedge,
                            tsetup_WD32_WCLK_negedge_posedge,
                            thold_WD32_WCLK_posedge_posedge,
                            thold_WD32_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD31_WCLK_posedge,
                            TmDt_WD31_WCLK_posedge,
                            WD31_ipd, "WD31",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD31_WCLK_posedge_posedge,
                            tsetup_WD31_WCLK_negedge_posedge,
                            thold_WD31_WCLK_posedge_posedge,
                            thold_WD31_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD30_WCLK_posedge,
                            TmDt_WD30_WCLK_posedge,
                            WD30_ipd, "WD30",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD30_WCLK_posedge_posedge,
                            tsetup_WD30_WCLK_negedge_posedge,
                            thold_WD30_WCLK_posedge_posedge,
                            thold_WD30_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD29_WCLK_posedge,
                            TmDt_WD29_WCLK_posedge,
                            WD29_ipd, "WD29",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD29_WCLK_posedge_posedge,
                            tsetup_WD29_WCLK_negedge_posedge,
                            thold_WD29_WCLK_posedge_posedge,
                            thold_WD29_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD28_WCLK_posedge,
                            TmDt_WD28_WCLK_posedge,
                            WD28_ipd, "WD28",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD28_WCLK_posedge_posedge,
                            tsetup_WD28_WCLK_negedge_posedge,
                            thold_WD28_WCLK_posedge_posedge,
                            thold_WD28_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD27_WCLK_posedge,
                            TmDt_WD27_WCLK_posedge,
                            WD27_ipd, "WD27",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD27_WCLK_posedge_posedge,
                            tsetup_WD27_WCLK_negedge_posedge,
                            thold_WD27_WCLK_posedge_posedge,
                            thold_WD27_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD26_WCLK_posedge,
                            TmDt_WD26_WCLK_posedge,
                            WD26_ipd, "WD26",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD26_WCLK_posedge_posedge,
                            tsetup_WD26_WCLK_negedge_posedge,
                            thold_WD26_WCLK_posedge_posedge,
                            thold_WD26_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD25_WCLK_posedge,
                            TmDt_WD25_WCLK_posedge,
                            WD25_ipd, "WD25",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD25_WCLK_posedge_posedge,
                            tsetup_WD25_WCLK_negedge_posedge,
                            thold_WD25_WCLK_posedge_posedge,
                            thold_WD25_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD24_WCLK_posedge,
                            TmDt_WD24_WCLK_posedge,
                            WD24_ipd, "WD24",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD24_WCLK_posedge_posedge,
                            tsetup_WD24_WCLK_negedge_posedge,
                            thold_WD24_WCLK_posedge_posedge,
                            thold_WD24_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='1')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD23_WCLK_posedge,
                            TmDt_WD23_WCLK_posedge,
                            WD23_ipd, "WD23",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD23_WCLK_posedge_posedge,
                            tsetup_WD23_WCLK_negedge_posedge,
                            thold_WD23_WCLK_posedge_posedge,
                            thold_WD23_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD22_WCLK_posedge,
                            TmDt_WD22_WCLK_posedge,
                            WD22_ipd, "WD22",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD22_WCLK_posedge_posedge,
                            tsetup_WD22_WCLK_negedge_posedge,
                            thold_WD22_WCLK_posedge_posedge,
                            thold_WD22_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD21_WCLK_posedge,
                            TmDt_WD21_WCLK_posedge,
                            WD21_ipd, "WD21",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD21_WCLK_posedge_posedge,
                            tsetup_WD21_WCLK_negedge_posedge,
                            thold_WD21_WCLK_posedge_posedge,
                            thold_WD21_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD20_WCLK_posedge,
                            TmDt_WD20_WCLK_posedge,
                            WD20_ipd, "WD20",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD20_WCLK_posedge_posedge,
                            tsetup_WD20_WCLK_negedge_posedge,
                            thold_WD20_WCLK_posedge_posedge,
                            thold_WD20_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD19_WCLK_posedge,
                            TmDt_WD19_WCLK_posedge,
                            WD19_ipd, "WD19",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD19_WCLK_posedge_posedge,
                            tsetup_WD19_WCLK_negedge_posedge,
                            thold_WD19_WCLK_posedge_posedge,
                            thold_WD19_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD18_WCLK_posedge,
                            TmDt_WD18_WCLK_posedge,
                            WD18_ipd, "WD18",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD18_WCLK_posedge_posedge,
                            tsetup_WD18_WCLK_negedge_posedge,
                            thold_WD18_WCLK_posedge_posedge,
                            thold_WD18_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD17_WCLK_posedge,
                            TmDt_WD17_WCLK_posedge,
                            WD17_ipd, "WD17",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD17_WCLK_posedge_posedge,
                            tsetup_WD17_WCLK_negedge_posedge,
                            thold_WD17_WCLK_posedge_posedge,
                            thold_WD17_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD16_WCLK_posedge,
                            TmDt_WD16_WCLK_posedge,
                            WD16_ipd, "WD16",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD16_WCLK_posedge_posedge,
                            tsetup_WD16_WCLK_negedge_posedge,
                            thold_WD16_WCLK_posedge_posedge,
                            thold_WD16_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD15_WCLK_posedge,
                            TmDt_WD15_WCLK_posedge,
                            WD15_ipd, "WD15",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD15_WCLK_posedge_posedge,
                            tsetup_WD15_WCLK_negedge_posedge,
                            thold_WD15_WCLK_posedge_posedge,
                            thold_WD15_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD14_WCLK_posedge,
                            TmDt_WD14_WCLK_posedge,
                            WD14_ipd, "WD14",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD14_WCLK_posedge_posedge,
                            tsetup_WD14_WCLK_negedge_posedge,
                            thold_WD14_WCLK_posedge_posedge,
                            thold_WD14_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD13_WCLK_posedge,
                            TmDt_WD13_WCLK_posedge,
                            WD13_ipd, "WD13",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD13_WCLK_posedge_posedge,
                            tsetup_WD13_WCLK_negedge_posedge,
                            thold_WD13_WCLK_posedge_posedge,
                            thold_WD13_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD12_WCLK_posedge,
                            TmDt_WD12_WCLK_posedge,
                            WD12_ipd, "WD12",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD12_WCLK_posedge_posedge,
                            tsetup_WD12_WCLK_negedge_posedge,
                            thold_WD12_WCLK_posedge_posedge,
                            thold_WD12_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD11_WCLK_posedge,
                            TmDt_WD11_WCLK_posedge,
                            WD11_ipd, "WD11",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD11_WCLK_posedge_posedge,
                            tsetup_WD11_WCLK_negedge_posedge,
                            thold_WD11_WCLK_posedge_posedge,
                            thold_WD11_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD10_WCLK_posedge,
                            TmDt_WD10_WCLK_posedge,
                            WD10_ipd, "WD10",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD10_WCLK_posedge_posedge,
                            tsetup_WD10_WCLK_negedge_posedge,
                            thold_WD10_WCLK_posedge_posedge,
                            thold_WD10_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD9_WCLK_posedge,
                            TmDt_WD9_WCLK_posedge,
                            WD9_ipd, "WD9",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD9_WCLK_posedge_posedge,
                            tsetup_WD9_WCLK_negedge_posedge,
                            thold_WD9_WCLK_posedge_posedge,
                            thold_WD9_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD8_WCLK_posedge,
                            TmDt_WD8_WCLK_posedge,
                            WD8_ipd, "WD8",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD8_WCLK_posedge_posedge,
                            tsetup_WD8_WCLK_negedge_posedge,
                            thold_WD8_WCLK_posedge_posedge,
                            thold_WD8_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD7_WCLK_posedge,
                            TmDt_WD7_WCLK_posedge,
                            WD7_ipd, "WD7",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD7_WCLK_posedge_posedge,
                            tsetup_WD7_WCLK_negedge_posedge,
                            thold_WD7_WCLK_posedge_posedge,
                            thold_WD7_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD6_WCLK_posedge,
                            TmDt_WD6_WCLK_posedge,
                            WD6_ipd, "WD6",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD6_WCLK_posedge_posedge,
                            tsetup_WD6_WCLK_negedge_posedge,
                            thold_WD6_WCLK_posedge_posedge,
                            thold_WD6_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD5_WCLK_posedge,
                            TmDt_WD5_WCLK_posedge,
                            WD5_ipd, "WD5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD5_WCLK_posedge_posedge,
                            tsetup_WD5_WCLK_negedge_posedge,
                            thold_WD5_WCLK_posedge_posedge,
                            thold_WD5_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD4_WCLK_posedge,
                            TmDt_WD4_WCLK_posedge,
                            WD4_ipd, "WD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD4_WCLK_posedge_posedge,
                            tsetup_WD4_WCLK_negedge_posedge,
                            thold_WD4_WCLK_posedge_posedge,
                            thold_WD4_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD3_WCLK_posedge,
                            TmDt_WD3_WCLK_posedge,
                            WD3_ipd, "WD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD3_WCLK_posedge_posedge,
                            tsetup_WD3_WCLK_negedge_posedge,
                            thold_WD3_WCLK_posedge_posedge,
                            thold_WD3_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD2_WCLK_posedge,
                            TmDt_WD2_WCLK_posedge,
                            WD2_ipd, "WD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD2_WCLK_posedge_posedge,
                            tsetup_WD2_WCLK_negedge_posedge,
                            thold_WD2_WCLK_posedge_posedge,
                            thold_WD2_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD1_WCLK_posedge,
                            TmDt_WD1_WCLK_posedge,
                            WD1_ipd, "WD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD1_WCLK_posedge_posedge,
                            tsetup_WD1_WCLK_negedge_posedge,
                            thold_WD1_WCLK_posedge_posedge,
                            thold_WD1_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD0_WCLK_posedge,
                            TmDt_WD0_WCLK_posedge,
                            WD0_ipd, "WD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD0_WCLK_posedge_posedge,
                            tsetup_WD0_WCLK_negedge_posedge,
                            thold_WD0_WCLK_posedge_posedge,
                            thold_WD0_WCLK_negedge_posedge,
                            ((To_X01(WEN_ipd)='1') and (To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup WEN high before WCLK rising
      --   Hold  WEN high after WCLK rising

      VitalSetupHoldCheck ( Tviol_WEN_WCLK_posedge,
                            TmDt_WEN_WCLK_posedge,
                            WEN_ipd, "WEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WEN_WCLK_posedge_posedge,
                            tsetup_WEN_WCLK_negedge_posedge,
                            thold_WEN_WCLK_posedge_posedge,
                            thold_WEN_WCLK_negedge_posedge,
                            ((To_X01(CLR_ipd)='0')),
                            '/',
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            ((To_X01(CLR_ipd)='0')),
                            InstancePath & "/FIFO64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Recovery CLR high before WCLK rising
      --   Hold  CLR high or low before WCLK rising

         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_WCLK_posedge,
          TimingData              => Tmkr_CLR_WCLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => WCLK_ipd,
          RefSignalName          => "WCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_WCLK_posedge_posedge,
          Removal                 => thold_CLR_WCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TimingCheckOn,
          RefTransition           => '/',
          HeaderMsg               => InstancePath & "/FIFO64K36",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);

      --   Pulse Width of CLR
 
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PeriodData_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => TRUE,
          HeaderMsg               => InstancePath &"/FIFO64K36",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);

    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################

     if(EMPTY_zd = '1') then
        REN_int := '0';
     else
        REN_int := REN_ipd;
     end if;

     if(FULL_zd = '1') then
       WEN_int :='0';
     else
       WEN_int := WEN_ipd;
     end if;


    if (TO_X01(CLR_ipd)='X') then
      assert false
      report ": CLR unknown"
      severity Warning;
    elsif (TO_X01(CLR_ipd)='1') then -- Clear the FIFO
      WADDR := 0;
      RADDR := 0;
      WADDR_P1 :=0;
      WADDR_P2 :=0;
      RADDR_P1 :=0;
      RADDR_P2 :=0;
      WADDR_wrap :=0;
      RADDR_wrap :=0;
      FULL_zd := '0';
      AFULL_zd := '0';
      EMPTY_zd := '1';
      AEMPTY_zd := '1';
      RD35_zd := 'X';
      RD34_zd := 'X';
      RD33_zd := 'X';
      RD32_zd := 'X';
      RD31_zd := 'X';
      RD30_zd := 'X';
      RD29_zd := 'X';
      RD28_zd := 'X';
      RD27_zd := 'X';
      RD26_zd := 'X';
      RD25_zd := 'X';
      RD24_zd := 'X';
      RD23_zd := 'X';
      RD22_zd := 'X';
      RD21_zd := 'X';
      RD20_zd := 'X';
      RD19_zd := 'X';
      RD18_zd := 'X';
      RD17_zd := 'X';
      RD16_zd := 'X';
      RD15_zd := 'X';
      RD14_zd := 'X';
      RD13_zd := 'X';
      RD12_zd := 'X';
      RD11_zd := 'X';
      RD10_zd := 'X';
      RD9_zd := 'X';
      RD8_zd := 'X';
      RD7_zd := 'X';
      RD6_zd := 'X';
      RD5_zd := 'X';
      RD4_zd := 'X';
      RD3_zd := 'X';
      RD2_zd := 'X';
      RD1_zd := 'X';
      RD0_zd := 'X';
    else

      -- Decode Word Width

      if (TO_X01(WIDTH2_delayed)='0' and TO_X01(WIDTH1_delayed)='0' and TO_X01(WIDTH0_delayed)='0') then
        WWIDTH := 1;
        DIVID  := 1;
        HEIGTH := 4096;
      elsif (TO_X01(WIDTH2_delayed)='0' and TO_X01(WIDTH1_delayed)='0' and TO_X01(WIDTH0_delayed)='1') then
        WWIDTH := 2;
        DIVID  := 2;
        HEIGTH := 2048;
      elsif (TO_X01(WIDTH2_delayed)='0' and TO_X01(WIDTH1_delayed)='1' and TO_X01(WIDTH0_delayed)='0') then
        WWIDTH := 4;
        DIVID  := 4;
        HEIGTH := 1024;
      elsif (TO_X01(WIDTH2_delayed)='0' and TO_X01(WIDTH1_delayed)='1' and TO_X01(WIDTH0_delayed)='1') then
        WWIDTH := 9;
        DIVID  := 8;
        HEIGTH := 512;
      elsif (TO_X01(WIDTH2_delayed)='1' and TO_X01(WIDTH1_delayed)='0' and TO_X01(WIDTH0_delayed)='0') then
        WWIDTH := 18;
        DIVID  := 16;
        HEIGTH := 256;
      elsif (TO_X01(WIDTH2_delayed)='1' and TO_X01(WIDTH1_delayed)='0' and TO_X01(WIDTH0_delayed)='1') then
        WWIDTH := 36;
        DIVID  := 32;
        HEIGTH := 128;
      else
	assert false
	report ": WIDTH value invalid"
	severity Error;
      end if;

      -- Decode Word Depth

      if (TO_X01(DEPTH3_delayed)='0' and TO_X01(DEPTH2_delayed)='0' and TO_X01(DEPTH1_delayed)='0' and TO_X01(DEPTH0_delayed)='0') then
        WDEPTH := 1;
      elsif (TO_X01(DEPTH3_delayed)='0' and TO_X01(DEPTH2_delayed)='0' and TO_X01(DEPTH1_delayed)='0' and TO_X01(DEPTH0_delayed)='1') then
        WDEPTH := 2;
      elsif (TO_X01(DEPTH3_delayed)='0' and TO_X01(DEPTH2_delayed)='0' and TO_X01(DEPTH1_delayed)='1' and TO_X01(DEPTH0_delayed)='0') then
        WDEPTH := 3;
      elsif (TO_X01(DEPTH3_delayed)='0' and TO_X01(DEPTH2_delayed)='0' and TO_X01(DEPTH1_delayed)='1' and TO_X01(DEPTH0_delayed)='1') then
        WDEPTH := 4;
      elsif (TO_X01(DEPTH3_delayed)='0' and TO_X01(DEPTH2_delayed)='1' and TO_X01(DEPTH1_delayed)='0' and TO_X01(DEPTH0_delayed)='0') then
        WDEPTH := 5;
      elsif (TO_X01(DEPTH3_delayed)='0' and TO_X01(DEPTH2_delayed)='1' and TO_X01(DEPTH1_delayed)='0' and TO_X01(DEPTH0_delayed)='1') then
        WDEPTH := 6;
      elsif (TO_X01(DEPTH3_delayed)='0' and TO_X01(DEPTH2_delayed)='1' and TO_X01(DEPTH1_delayed)='1' and TO_X01(DEPTH0_delayed)='0') then
        WDEPTH := 7;
      elsif (TO_X01(DEPTH3_delayed)='0' and TO_X01(DEPTH2_delayed)='1' and TO_X01(DEPTH1_delayed)='1' and TO_X01(DEPTH0_delayed)='1') then
        WDEPTH := 8;
      elsif (TO_X01(DEPTH3_delayed)='1' and TO_X01(DEPTH2_delayed)='0' and TO_X01(DEPTH1_delayed)='0' and TO_X01(DEPTH0_delayed)='0') then
        WDEPTH := 9;
      elsif (TO_X01(DEPTH3_delayed)='1' and TO_X01(DEPTH2_delayed)='0' and TO_X01(DEPTH1_delayed)='0' and TO_X01(DEPTH0_delayed)='1') then
        WDEPTH := 10;
      elsif (TO_X01(DEPTH3_delayed)='1' and TO_X01(DEPTH2_delayed)='0' and TO_X01(DEPTH1_delayed)='1' and TO_X01(DEPTH0_delayed)='0') then
        WDEPTH := 11;
      elsif (TO_X01(DEPTH3_delayed)='1' and TO_X01(DEPTH2_delayed)='0' and TO_X01(DEPTH1_delayed)='1' and TO_X01(DEPTH0_delayed)='1') then
        WDEPTH := 12;
      elsif (TO_X01(DEPTH3_delayed)='1' and TO_X01(DEPTH2_delayed)='1' and TO_X01(DEPTH1_delayed)='0' and TO_X01(DEPTH0_delayed)='0') then
        WDEPTH := 13;
      elsif (TO_X01(DEPTH3_delayed)='1' and TO_X01(DEPTH2_delayed)='1' and TO_X01(DEPTH1_delayed)='0' and TO_X01(DEPTH0_delayed)='1') then
        WDEPTH := 14;
      elsif (TO_X01(DEPTH3_delayed)='1' and TO_X01(DEPTH2_delayed)='1' and TO_X01(DEPTH1_delayed)='1' and TO_X01(DEPTH0_delayed)='0') then
        WDEPTH := 15;
      elsif (TO_X01(DEPTH3_delayed)='1' and TO_X01(DEPTH2_delayed)='1' and TO_X01(DEPTH1_delayed)='1' and TO_X01(DEPTH0_delayed)='1') then
        WDEPTH := 16;
      else
	assert false
	report ": DEPTH value invalid"
	severity Error;
      end if;

      -- Decode Almost Empty Value

      AEVAL_temp := ((INT(AEVAL7_delayed)*128)+(INT(AEVAL6_delayed)*64)
                +(INT(AEVAL5_delayed)*32)+(INT(AEVAL4_delayed)*16)+(INT(AEVAL3_delayed)*8)
                +(INT(AEVAL2_delayed)*4)+(INT(AEVAL1_delayed)*2)+(INT(AEVAL0_delayed)));

      -- Decode Almost Full Value

      AFVAL_temp := ((INT(AFVAL7_delayed)*128)+(INT(AFVAL6_delayed)*64)
                +(INT(AFVAL5_delayed)*32)+(INT(AFVAL4_delayed)*16)+(INT(AFVAL3_delayed)*8)
                +(INT(AFVAL2_delayed)*4)+(INT(AFVAL1_delayed)*2)+(INT(AFVAL0_delayed)));

      AEVAL :=AEVAL_temp * (256/DIVID);
      AFVAL :=AFVAL_temp * (256/DIVID);

      MAX_ADDR := HEIGTH * WDEPTH;
      if (TO_X01(WCLK_ipd)='X') then
        if ((TO_X01(WEN_delayed) /= '1')) then
          if (TO_X01(WCLK_previous) /= 'X') then
            assert false
            report ": WCLK went unknown"
            severity Error;
          end if;
        end if;
      elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='1')) then

        RADDR_P2 := RADDR_P1;
        RADDR_P1 := RADDR;

        case (TO_X01(WEN_int)) is
          when '0' =>
            null;
          when '1' =>
              RAM_TMP(WADDR) := WD35_delayed & WD34_delayed & WD33_delayed & WD32_delayed &
                                WD31_delayed & WD30_delayed & WD29_delayed & WD28_delayed &
                                WD27_delayed & WD26_delayed & WD25_delayed & WD24_delayed &
                                WD23_delayed & WD22_delayed & WD21_delayed & WD20_delayed &
                                WD19_delayed & WD18_delayed & WD17_delayed & WD16_delayed &
                                WD15_delayed & WD14_delayed & WD13_delayed & WD12_delayed &
                                WD11_delayed & WD10_delayed & WD9_delayed & WD8_delayed &
                                WD7_delayed & WD6_delayed & WD5_delayed & WD4_delayed &
                                WD3_delayed & WD2_delayed & WD1_delayed & WD0_delayed ;

              if(WADDR <MAX_ADDR-1  ) then 
                WADDR := WADDR + 1;
                --WADDR_wrap :=0;
               else 
                WADDR :=(WADDR +1) mod  MAX_ADDR;
                WADDR_wrap :=1 - WADDR_wrap;
               end if;

          when others =>
            if (TO_X01(WEN_previous) = 'X') then
              assert false
              report ": WEN went unknown"
              severity Error;
            end if;
        end case;

       if(WADDR   = RADDR_P2 ) then 
          if(RADDR_wrap /= WADDR_wrap) then
           FULL_zd := '1';
           WEN_int := '0';
          end if;
       else
           FULL_zd := '0';
       end if;

        if(WADDR_wrap = RADDR_wrap ) then 
         if((WADDR - RADDR) >=AFVAL ) then
           AFULL_zd := '1';
         else
           AFULL_zd := '0';
         end if;

         if((WADDR - RADDR) <= AEVAL) then
          AEMPTY_zd := '1';
          else
          AEMPTY_zd := '0';
         end if;
        else 
         if((MAX_ADDR + WADDR - RADDR) >=AFVAL ) then
            AFULL_zd := '1';
          else
            AFULL_zd := '0';
         end if;

         if((MAX_ADDR + WADDR - RADDR) <= AEVAL) then
           AEMPTY_zd := '1';
         else
           AEMPTY_zd := '0';
         end if;
        end if;
     end if; -- rising WCLK edge
  -- end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      if (TO_X01(RCLK_ipd)='X') then
        if ((TO_X01(REN_delayed) /= '1')) then
          if (TO_X01(RCLK_previous) /= 'X') then
            assert false
              report ": RCLK went unknown"
              severity Error;
            RD35_zd := 'X';
            RD34_zd := 'X';
            RD33_zd := 'X';
            RD32_zd := 'X';
            RD31_zd := 'X';
            RD30_zd := 'X';
            RD29_zd := 'X';
            RD28_zd := 'X';
            RD27_zd := 'X';
            RD26_zd := 'X';
            RD25_zd := 'X';
            RD24_zd := 'X';
            RD23_zd := 'X';
            RD22_zd := 'X';
            RD21_zd := 'X';
            RD20_zd := 'X';
            RD19_zd := 'X';
            RD18_zd := 'X';
            RD17_zd := 'X';
            RD16_zd := 'X';
            RD15_zd := 'X';
            RD14_zd := 'X';
            RD13_zd := 'X';
            RD12_zd := 'X';
            RD11_zd := 'X';
            RD10_zd := 'X';
            RD9_zd := 'X';
            RD8_zd := 'X';
            RD7_zd := 'X';
            RD6_zd := 'X';
            RD5_zd := 'X';
            RD4_zd := 'X';
            RD3_zd := 'X';
            RD2_zd := 'X';
            RD1_zd := 'X';
            RD0_zd := 'X';
          end if;
        end if;
      elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd)='1')) then

         WADDR_P2 := WADDR_P1;
         WADDR_P1 := WADDR;

        case (TO_X01(REN_int)) is
          when '0' =>
              null;
          when '1' =>

              RD35_zd := RAM_TMP(RADDR)(35);
              RD34_zd := RAM_TMP(RADDR)(34);
              RD33_zd := RAM_TMP(RADDR)(33);
              RD32_zd := RAM_TMP(RADDR)(32);
              RD31_zd := RAM_TMP(RADDR)(31);
              RD30_zd := RAM_TMP(RADDR)(30);
              RD29_zd := RAM_TMP(RADDR)(29);
              RD28_zd := RAM_TMP(RADDR)(28);
              RD27_zd := RAM_TMP(RADDR)(27);
              RD26_zd := RAM_TMP(RADDR)(26);
              RD25_zd := RAM_TMP(RADDR)(25);
              RD24_zd := RAM_TMP(RADDR)(24);
              RD23_zd := RAM_TMP(RADDR)(23);
              RD22_zd := RAM_TMP(RADDR)(22);
              RD21_zd := RAM_TMP(RADDR)(21);
              RD20_zd := RAM_TMP(RADDR)(20);
              RD19_zd := RAM_TMP(RADDR)(19);
              RD18_zd := RAM_TMP(RADDR)(18);
              RD17_zd := RAM_TMP(RADDR)(17);
              RD16_zd := RAM_TMP(RADDR)(16);
              RD15_zd := RAM_TMP(RADDR)(15);
              RD14_zd := RAM_TMP(RADDR)(14);
              RD13_zd := RAM_TMP(RADDR)(13);
              RD12_zd := RAM_TMP(RADDR)(12);
              RD11_zd := RAM_TMP(RADDR)(11);
              RD10_zd := RAM_TMP(RADDR)(10);
              RD9_zd := RAM_TMP(RADDR)(9);
              RD8_zd := RAM_TMP(RADDR)(8);
              RD7_zd := RAM_TMP(RADDR)(7);
              RD6_zd := RAM_TMP(RADDR)(6);
              RD5_zd := RAM_TMP(RADDR)(5);
              RD4_zd := RAM_TMP(RADDR)(4);
              RD3_zd := RAM_TMP(RADDR)(3);
              RD2_zd := RAM_TMP(RADDR)(2);
              RD1_zd := RAM_TMP(RADDR)(1);
              RD0_zd := RAM_TMP(RADDR)(0);

              if(RADDR <MAX_ADDR-1  ) then
                RADDR := RADDR + 1;
                --RADDR_wrap :=0;
              else
                RADDR :=(RADDR +1) mod  MAX_ADDR;
                RADDR_wrap :=1 - RADDR_wrap;
              end if;

       when others =>
        if (TO_X01(REN_previous) = 'X') then
          assert false
          report ": REN went unknown"
          severity Error;
          end if;
        end case;

        if(RADDR = WADDR_P2 ) then 
         if(RADDR_wrap = WADDR_wrap) then
           EMPTY_zd := '1';
           REN_int := '0';
         else
          EMPTY_zd  :=  '0';
          end if;
         else
          EMPTY_zd := '0';
         end if;

        if(WADDR_wrap = RADDR_wrap ) then
         if((WADDR - RADDR) >=AFVAL ) then
           AFULL_zd := '1';
         else
           AFULL_zd := '0';
         end if;

         if((WADDR - RADDR) <= AEVAL) then
          AEMPTY_zd := '1';
          else
          AEMPTY_zd := '0';
         end if;
        else
         if((MAX_ADDR + WADDR - RADDR) >=AFVAL ) then
            AFULL_zd := '1';
          else
            AFULL_zd := '0';
         end if;

         if((MAX_ADDR + WADDR - RADDR) <= AEVAL) then
           AEMPTY_zd := '1';
         else
           AEMPTY_zd := '0';
         end if;
        end if;
      end if; -- rising RCLK edge
    end if; -- CLR active

    WCLK_previous := WCLK_ipd;
    RCLK_previous := RCLK_ipd;
    WIDTH2_delayed := WIDTH2_ipd;
    WIDTH1_delayed := WIDTH1_ipd;
    WIDTH0_delayed := WIDTH0_ipd;
    if WEN_ipd'event then
      WEN_previous := WEN_delayed;
      WEN_delayed := WEN_ipd;
    end if;
    AFVAL7_delayed := AFVAL7_ipd;
    AFVAL6_delayed := AFVAL6_ipd;
    AFVAL5_delayed := AFVAL5_ipd;
    AFVAL4_delayed := AFVAL4_ipd;
    AFVAL3_delayed := AFVAL3_ipd;
    AFVAL2_delayed := AFVAL2_ipd;
    AFVAL1_delayed := AFVAL1_ipd;
    AFVAL0_delayed := AFVAL0_ipd;
    AEVAL7_delayed := AEVAL7_ipd;
    AEVAL6_delayed := AEVAL6_ipd;
    AEVAL5_delayed := AEVAL5_ipd;
    AEVAL4_delayed := AEVAL4_ipd;
    AEVAL3_delayed := AEVAL3_ipd;
    AEVAL2_delayed := AEVAL2_ipd;
    AEVAL1_delayed := AEVAL1_ipd;
    AEVAL0_delayed := AEVAL0_ipd;
    if REN_ipd'event then
      REN_previous := REN_delayed;
      REN_delayed := REN_ipd;
    end if;
    WD35_delayed := WD35_ipd;
    WD34_delayed := WD34_ipd;
    WD33_delayed := WD33_ipd;
    WD32_delayed := WD32_ipd;
    WD31_delayed := WD31_ipd;
    WD30_delayed := WD30_ipd;
    WD29_delayed := WD29_ipd;
    WD28_delayed := WD28_ipd;
    WD27_delayed := WD27_ipd;
    WD26_delayed := WD26_ipd;
    WD25_delayed := WD25_ipd;
    WD24_delayed := WD24_ipd;
    WD23_delayed := WD23_ipd;
    WD22_delayed := WD22_ipd;
    WD21_delayed := WD21_ipd;
    WD20_delayed := WD20_ipd;
    WD19_delayed := WD19_ipd;
    WD18_delayed := WD18_ipd;
    WD17_delayed := WD17_ipd;
    WD16_delayed := WD16_ipd;
    WD15_delayed := WD15_ipd;
    WD14_delayed := WD14_ipd;
    WD13_delayed := WD13_ipd;
    WD12_delayed := WD12_ipd;
    WD11_delayed := WD11_ipd;
    WD10_delayed := WD10_ipd;
    WD9_delayed := WD9_ipd;
    WD8_delayed := WD8_ipd;
    WD7_delayed := WD7_ipd;
    WD6_delayed := WD6_ipd;
    WD5_delayed := WD5_ipd;
    WD4_delayed := WD4_ipd;
    WD3_delayed := WD3_ipd;
    WD2_delayed := WD2_ipd;
    WD1_delayed := WD1_ipd;
    WD0_delayed := WD0_ipd;
    DEPTH3_delayed := DEPTH3_ipd;
    DEPTH2_delayed := DEPTH2_ipd;
    DEPTH1_delayed := DEPTH1_ipd;
    DEPTH0_delayed := DEPTH0_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => RD35,
	GlitchData => RD35_GlitchData,
	OutSignalName => "RD35",
	OutTemp => RD35_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD35), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD35), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => Xon,
	MsgOn => MsgOn,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
        OutSignal => RD34,
        GlitchData => RD34_GlitchData,
        OutSignalName => "RD34",
        OutTemp => RD34_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD34), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD34), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD33,
        GlitchData => RD33_GlitchData,
        OutSignalName => "RD33",
        OutTemp => RD33_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD33), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD33), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD32,
        GlitchData => RD32_GlitchData,
        OutSignalName => "RD32",
        OutTemp => RD32_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD32), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD32), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD31,
        GlitchData => RD31_GlitchData,
        OutSignalName => "RD31",
        OutTemp => RD31_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD31), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD31), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD30,
        GlitchData => RD30_GlitchData,
        OutSignalName => "RD30",
        OutTemp => RD30_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD30), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD30), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD29,
        GlitchData => RD29_GlitchData,
        OutSignalName => "RD29",
        OutTemp => RD29_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD29), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD29), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD28,
        GlitchData => RD28_GlitchData,
        OutSignalName => "RD28",
        OutTemp => RD28_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD28), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD28), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD27,
        GlitchData => RD27_GlitchData,
        OutSignalName => "RD27",
        OutTemp => RD27_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD27), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD27), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD26,
        GlitchData => RD26_GlitchData,
        OutSignalName => "RD26",
        OutTemp => RD26_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD26), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD26), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD25,
        GlitchData => RD25_GlitchData,
        OutSignalName => "RD25",
        OutTemp => RD25_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD25), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD25), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD24,
        GlitchData => RD24_GlitchData,
        OutSignalName => "RD24",
        OutTemp => RD24_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD24), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD24), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD23,
        GlitchData => RD23_GlitchData,
        OutSignalName => "RD23",
        OutTemp => RD23_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD23), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD23), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD22,
        GlitchData => RD22_GlitchData,
        OutSignalName => "RD22",
        OutTemp => RD22_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD22), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD22), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD21,
        GlitchData => RD21_GlitchData,
        OutSignalName => "RD21",
        OutTemp => RD21_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD21), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD21), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD20,
        GlitchData => RD20_GlitchData,
        OutSignalName => "RD20",
        OutTemp => RD20_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD20), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD20), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD19,
        GlitchData => RD19_GlitchData,
        OutSignalName => "RD19",
        OutTemp => RD19_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD19), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD19), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD18,
        GlitchData => RD18_GlitchData,
        OutSignalName => "RD18",
        OutTemp => RD18_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD18), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD18), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD17,
        GlitchData => RD17_GlitchData,
        OutSignalName => "RD17",
        OutTemp => RD17_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD17), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD17), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD16,
        GlitchData => RD16_GlitchData,
        OutSignalName => "RD16",
        OutTemp => RD16_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD16), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD16), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD15,
        GlitchData => RD15_GlitchData,
        OutSignalName => "RD15",
        OutTemp => RD15_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD15), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD15), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD14,
        GlitchData => RD14_GlitchData,
        OutSignalName => "RD14",
        OutTemp => RD14_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD14), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD14), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD13,
        GlitchData => RD13_GlitchData,
        OutSignalName => "RD13",
        OutTemp => RD13_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD13), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD13), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD12,
        GlitchData => RD12_GlitchData,
        OutSignalName => "RD12",
        OutTemp => RD12_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD12), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD12), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD11,
        GlitchData => RD11_GlitchData,
        OutSignalName => "RD11",
        OutTemp => RD11_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD11), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD11), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD10,
        GlitchData => RD10_GlitchData,
        OutSignalName => "RD10",
        OutTemp => RD10_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD10), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD10), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD9,
        GlitchData => RD9_GlitchData,
        OutSignalName => "RD9",
        OutTemp => RD9_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD9), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD9), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD8,
        GlitchData => RD8_GlitchData,
        OutSignalName => "RD8",
        OutTemp => RD8_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD8), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD8), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD7,
        GlitchData => RD7_GlitchData,
        OutSignalName => "RD7",
        OutTemp => RD7_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD7), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD7), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD6,
        GlitchData => RD6_GlitchData,
        OutSignalName => "RD6",
        OutTemp => RD6_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD6), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD6), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD5,
        GlitchData => RD5_GlitchData,
        OutSignalName => "RD5",
        OutTemp => RD5_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD5), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD5), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD4,
        GlitchData => RD4_GlitchData,
        OutSignalName => "RD4",
        OutTemp => RD4_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD4), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD4), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD3,
        GlitchData => RD3_GlitchData,
        OutSignalName => "RD3",
        OutTemp => RD3_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD3), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD3), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD2,
        GlitchData => RD2_GlitchData,
        OutSignalName => "RD2",
        OutTemp => RD2_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD2), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD2), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD1,
        GlitchData => RD1_GlitchData,
        OutSignalName => "RD1",
        OutTemp => RD1_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD1), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD1), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD0,
        GlitchData => RD0_GlitchData,
        OutSignalName => "RD0",
        OutTemp => RD0_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD0), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_RD0), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );
    
    VitalPathDelay01Z (
        OutSignal => FULL,
        GlitchData => FULL_GlitchData,
        OutSignalName => "FULL",
        OutTemp => FULL_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_FULL), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_FULL), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );
    
    VitalPathDelay01Z (
        OutSignal => AFULL,
        GlitchData => AFULL_GlitchData,
        OutSignalName => "AFULL",
        OutTemp => AFULL_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_AFULL), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_AFULL), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );
    
    VitalPathDelay01Z (
        OutSignal => EMPTY,
        GlitchData => EMPTY_GlitchData,
        OutSignalName => "EMPTY",
        OutTemp => EMPTY_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_EMPTY), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_EMPTY), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );
    
    VitalPathDelay01Z (
        OutSignal => AEMPTY,
        GlitchData => AEMPTY_GlitchData,
        OutSignalName => "AEMPTY",
        OutTemp => AEMPTY_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_AEMPTY), TRUE),
                  1 => (CLR_ipd'last_event, 
                        VitalExtendToFillDelay(tpd_CLR_AEMPTY), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );
  end process VITALBehavior;

end VITAL_ACT;

configuration CFG_FIFO64K36_VITAL of FIFO64K36 is
   for VITAL_ACT
   end for;
end CFG_FIFO64K36_VITAL;

-----------------------------------------------------------------
--
--  Actel AX RAM64K36 VHDL behavioral model
--  64K X 1 RAM with rising write clock and rising read clock.
--  Allows variable and independent Write and Read widths of only
--  4Kx1, 2Kx2, 1Kx4, 512x9, 256x18, or 128x36.
--  Depth pins functionally inert.  In model just to make sure 
--  they are connected.  Used by combiner to calculate cascading.
--
--  Future changes:  Need to be able to initialize RAM from text file.
--
--  Uses VITAL95 package
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - 11/22/00 - Dale Walter - Initial Version.
-- 1.1 - 03/13/01 - Dale Walter - Cloned from RAM4K36.
-- 1.2 - 05/09/01 - Dale Walter - Change memory to variable instead of signal.
--                              - Change WRAD & RDAD calculation to be the same
--                                regardless of WW and RR (i.e. low-order bits 
--                                assumed to be tied-off to GND for widths > 1.
-- 1.3 - 9/27/02 - Krupa Singampalli - New Timing Arcs
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
entity RAM64K36 is
  GENERIC (
        tipd_DEPTH3   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH2   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH1   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH0   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD15   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD14   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD13   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD12   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD11   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD10   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD9    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD8    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD7    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD6    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD5    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD35     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD34     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD33     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD32     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD31     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD30     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD29     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD28     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD27     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD26     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD25     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD24     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD23     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD22     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD21     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD20     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD19     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD18     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD17     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD16     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD15     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD14     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD13     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD12     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD11     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD10     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD9      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD8      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD7      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD6      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD5      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD4      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD3      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WW2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WW1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WW0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WEN      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD15   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD14   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD13   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD12   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD11   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD10   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD9    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD8    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD7    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD6    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD5    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD4    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RW2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RW1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RW0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_REN      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        

        tpd_RCLK_RD0  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD1  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD2  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD3  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD4  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD5  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD6  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD7  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD8  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD9  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD10 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD11 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD12 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD13 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD14 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD15 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD16 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD17 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD18 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD19 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD20 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD21 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD22 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD23 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD24 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD25 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD26 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD27 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD28 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD29 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD30 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD31 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD32 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD33 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD34 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD35 : VitalDelayType01 := (0.100 ns, 0.100 ns);


        tsetup_RDAD15_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD14_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD13_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD12_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD11_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD10_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD9_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD8_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD7_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD6_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD5_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD4_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_RDAD15_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD14_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD13_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD12_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD11_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD10_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD9_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD8_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD7_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD6_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD5_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD4_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        tsetup_RW2_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW1_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW0_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW2_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW1_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW0_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;


        tsetup_DEPTH3_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH2_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH1_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH0_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH3_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH2_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH1_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH0_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;



        tsetup_WRAD15_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD14_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD13_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD12_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD11_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD10_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD9_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD8_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_WRAD15_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD14_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD13_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD12_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD11_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD10_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD9_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD8_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_WD35_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD34_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD33_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD32_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD31_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD30_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD29_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD28_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD27_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD26_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD25_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD24_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD23_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD22_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD21_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD20_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD19_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD18_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD17_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD16_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD15_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD14_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD13_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD12_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD11_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD10_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD9_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD8_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD35_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD34_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD33_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD32_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD31_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD30_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD29_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD28_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD27_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD26_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD25_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD24_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD23_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD22_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD21_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD20_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD19_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD18_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD17_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD16_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD15_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD14_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD13_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD12_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD11_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD10_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD9_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD8_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;


        tsetup_WW2_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW2_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;


        thold_RDAD15_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD14_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD13_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD12_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD11_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD10_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD9_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD8_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD7_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD6_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD5_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;

        thold_RDAD15_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD14_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD13_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD12_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD11_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD10_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD9_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD8_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD7_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD6_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD5_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;



        thold_RW2_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW1_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW0_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW2_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW1_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW0_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

        thold_DEPTH3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        thold_WRAD15_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD14_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD13_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD12_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD11_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD10_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD9_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD8_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;

        thold_WRAD15_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD14_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD13_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD12_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD11_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD10_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD9_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD8_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        thold_WD35_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD34_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD33_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD32_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD31_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD30_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD29_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD28_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD27_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD26_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD25_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD24_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD23_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD22_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD21_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD20_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD19_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD18_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD17_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD16_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD15_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD14_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD13_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD12_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD11_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD10_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD9_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD8_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD35_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD34_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD33_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD32_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD31_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD30_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD29_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD28_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD27_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD26_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD25_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD24_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD23_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD22_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD21_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD20_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD19_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD18_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD17_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD16_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD15_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD14_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD13_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD12_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD11_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD10_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD9_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD8_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;


        thold_WW2_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW1_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW0_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW2_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW1_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW0_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

        tsetup_REN_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True
        );
  PORT (
        DEPTH3 : IN STD_ULOGIC ;
        DEPTH2 : IN STD_ULOGIC ;
        DEPTH1 : IN STD_ULOGIC ;
        DEPTH0 : IN STD_ULOGIC ;
        WRAD15 : IN STD_ULOGIC ;
        WRAD14 : IN STD_ULOGIC ;
        WRAD13 : IN STD_ULOGIC ;
        WRAD12 : IN STD_ULOGIC ;
        WRAD11 : IN STD_ULOGIC ;
        WRAD10 : IN STD_ULOGIC ;
        WRAD9  : IN STD_ULOGIC ;
        WRAD8  : IN STD_ULOGIC ;
        WRAD7  : IN STD_ULOGIC ;
        WRAD6  : IN STD_ULOGIC ;
        WRAD5  : IN STD_ULOGIC ;
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD35   : IN STD_ULOGIC ;
        WD34   : IN STD_ULOGIC ;
        WD33   : IN STD_ULOGIC ;
        WD32   : IN STD_ULOGIC ;
        WD31   : IN STD_ULOGIC ;
        WD30   : IN STD_ULOGIC ;
        WD29   : IN STD_ULOGIC ;
        WD28   : IN STD_ULOGIC ;
        WD27   : IN STD_ULOGIC ;
        WD26   : IN STD_ULOGIC ;
        WD25   : IN STD_ULOGIC ;
        WD24   : IN STD_ULOGIC ;
        WD23   : IN STD_ULOGIC ;
        WD22   : IN STD_ULOGIC ;
        WD21   : IN STD_ULOGIC ;
        WD20   : IN STD_ULOGIC ;
        WD19   : IN STD_ULOGIC ;
        WD18   : IN STD_ULOGIC ;
        WD17   : IN STD_ULOGIC ;
        WD16   : IN STD_ULOGIC ;
        WD15   : IN STD_ULOGIC ;
        WD14   : IN STD_ULOGIC ;
        WD13   : IN STD_ULOGIC ;
        WD12   : IN STD_ULOGIC ;
        WD11   : IN STD_ULOGIC ;
        WD10   : IN STD_ULOGIC ;
        WD9    : IN STD_ULOGIC ;
        WD8    : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        WW2    : IN STD_ULOGIC ;
        WW1    : IN STD_ULOGIC ;
        WW0    : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RDAD15 : IN STD_ULOGIC ;
        RDAD14 : IN STD_ULOGIC ;
        RDAD13 : IN STD_ULOGIC ;
        RDAD12 : IN STD_ULOGIC ;
        RDAD11 : IN STD_ULOGIC ;
        RDAD10 : IN STD_ULOGIC ;
        RDAD9  : IN STD_ULOGIC ;
        RDAD8  : IN STD_ULOGIC ;
        RDAD7  : IN STD_ULOGIC ;
        RDAD6  : IN STD_ULOGIC ;
        RDAD5  : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        RW2    : IN STD_ULOGIC ;
        RW1    : IN STD_ULOGIC ;
        RW0    : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD35   : OUT STD_ULOGIC ;
        RD34   : OUT STD_ULOGIC ;
        RD33   : OUT STD_ULOGIC ;
        RD32   : OUT STD_ULOGIC ;
        RD31   : OUT STD_ULOGIC ;
        RD30   : OUT STD_ULOGIC ;
        RD29   : OUT STD_ULOGIC ;
        RD28   : OUT STD_ULOGIC ;
        RD27   : OUT STD_ULOGIC ;
        RD26   : OUT STD_ULOGIC ;
        RD25   : OUT STD_ULOGIC ;
        RD24   : OUT STD_ULOGIC ;
        RD23   : OUT STD_ULOGIC ;
        RD22   : OUT STD_ULOGIC ;
        RD21   : OUT STD_ULOGIC ;
        RD20   : OUT STD_ULOGIC ;
        RD19   : OUT STD_ULOGIC ;
        RD18   : OUT STD_ULOGIC ;
        RD17   : OUT STD_ULOGIC ;
        RD16   : OUT STD_ULOGIC ;
        RD15   : OUT STD_ULOGIC ;
        RD14   : OUT STD_ULOGIC ;
        RD13   : OUT STD_ULOGIC ;
        RD12   : OUT STD_ULOGIC ;
        RD11   : OUT STD_ULOGIC ;
        RD10   : OUT STD_ULOGIC ;
        RD9    : OUT STD_ULOGIC ;
        RD8    : OUT STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC ;
        RD6    : OUT STD_ULOGIC ;
        RD5    : OUT STD_ULOGIC ;
        RD4    : OUT STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC ;
        RD2    : OUT STD_ULOGIC ;
        RD1    : OUT STD_ULOGIC ;
        RD0    : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of RAM64K36 : entity is TRUE;
  
end RAM64K36;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of RAM64K36 is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal DEPTH3_ipd : std_ulogic := 'X';
  signal DEPTH2_ipd : std_ulogic := 'X';
  signal DEPTH1_ipd : std_ulogic := 'X';
  signal DEPTH0_ipd : std_ulogic := 'X';
  signal WRAD15_ipd : std_ulogic := 'X';
  signal WRAD14_ipd : std_ulogic := 'X';
  signal WRAD13_ipd : std_ulogic := 'X';
  signal WRAD12_ipd : std_ulogic := 'X';
  signal WRAD11_ipd : std_ulogic := 'X';
  signal WRAD10_ipd : std_ulogic := 'X';
  signal WRAD9_ipd  : std_ulogic := 'X';
  signal WRAD8_ipd  : std_ulogic := 'X';
  signal WRAD7_ipd  : std_ulogic := 'X';
  signal WRAD6_ipd  : std_ulogic := 'X';
  signal WRAD5_ipd  : std_ulogic := 'X';
  signal WRAD4_ipd  : std_ulogic := 'X';
  signal WRAD3_ipd  : std_ulogic := 'X';
  signal WRAD2_ipd  : std_ulogic := 'X';
  signal WRAD1_ipd  : std_ulogic := 'X';
  signal WRAD0_ipd  : std_ulogic := 'X';
  signal WD35_ipd   : std_ulogic := 'X';
  signal WD34_ipd   : std_ulogic := 'X';
  signal WD33_ipd   : std_ulogic := 'X';
  signal WD32_ipd   : std_ulogic := 'X';
  signal WD31_ipd   : std_ulogic := 'X';
  signal WD30_ipd   : std_ulogic := 'X';
  signal WD29_ipd   : std_ulogic := 'X';
  signal WD28_ipd   : std_ulogic := 'X';
  signal WD27_ipd   : std_ulogic := 'X';
  signal WD26_ipd   : std_ulogic := 'X';
  signal WD25_ipd   : std_ulogic := 'X';
  signal WD24_ipd   : std_ulogic := 'X';
  signal WD23_ipd   : std_ulogic := 'X';
  signal WD22_ipd   : std_ulogic := 'X';
  signal WD21_ipd   : std_ulogic := 'X';
  signal WD20_ipd   : std_ulogic := 'X';
  signal WD19_ipd   : std_ulogic := 'X';
  signal WD18_ipd   : std_ulogic := 'X';
  signal WD17_ipd   : std_ulogic := 'X';
  signal WD16_ipd   : std_ulogic := 'X';
  signal WD15_ipd   : std_ulogic := 'X';
  signal WD14_ipd   : std_ulogic := 'X';
  signal WD13_ipd   : std_ulogic := 'X';
  signal WD12_ipd   : std_ulogic := 'X';
  signal WD11_ipd   : std_ulogic := 'X';
  signal WD10_ipd   : std_ulogic := 'X';
  signal WD9_ipd    : std_ulogic := 'X';
  signal WD8_ipd    : std_ulogic := 'X';
  signal WD7_ipd    : std_ulogic := 'X';
  signal WD6_ipd    : std_ulogic := 'X';
  signal WD5_ipd    : std_ulogic := 'X';
  signal WD4_ipd    : std_ulogic := 'X';
  signal WD3_ipd    : std_ulogic := 'X';
  signal WD2_ipd    : std_ulogic := 'X';
  signal WD1_ipd    : std_ulogic := 'X';
  signal WD0_ipd    : std_ulogic := 'X';
  signal WW2_ipd    : std_ulogic := 'X';
  signal WW1_ipd    : std_ulogic := 'X';
  signal WW0_ipd    : std_ulogic := 'X';
  signal WEN_ipd    : std_ulogic := 'X';
  signal WCLK_ipd   : std_ulogic := 'X';
  signal RDAD15_ipd : std_ulogic := 'X';
  signal RDAD14_ipd : std_ulogic := 'X';
  signal RDAD13_ipd : std_ulogic := 'X';
  signal RDAD12_ipd : std_ulogic := 'X';
  signal RDAD11_ipd : std_ulogic := 'X';
  signal RDAD10_ipd : std_ulogic := 'X';
  signal RDAD9_ipd  : std_ulogic := 'X';
  signal RDAD8_ipd  : std_ulogic := 'X';
  signal RDAD7_ipd  : std_ulogic := 'X';
  signal RDAD6_ipd  : std_ulogic := 'X';
  signal RDAD5_ipd  : std_ulogic := 'X';
  signal RDAD4_ipd  : std_ulogic := 'X';
  signal RDAD3_ipd  : std_ulogic := 'X';
  signal RDAD2_ipd  : std_ulogic := 'X';
  signal RDAD1_ipd  : std_ulogic := 'X';
  signal RDAD0_ipd  : std_ulogic := 'X';
  signal RW2_ipd    : std_ulogic := 'X';
  signal RW1_ipd    : std_ulogic := 'X';
  signal RW0_ipd    : std_ulogic := 'X';
  signal REN_ipd    : std_ulogic := 'X';
  signal RCLK_ipd   : std_ulogic := 'X';
  type MEM is array(0 to 65535) of std_ulogic; -- Internal memory
  type MEM9 is array(0 to 8191) of std_ulogic; -- Internal memory
  --signal RAM_TMP    : MEM;
  --signal RAM_TMP9   : MEM9;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (DEPTH3_ipd, DEPTH3, VitalExtendToFillDelay(tipd_DEPTH3));
    VitalWireDelay (DEPTH2_ipd, DEPTH2, VitalExtendToFillDelay(tipd_DEPTH2));
    VitalWireDelay (DEPTH1_ipd, DEPTH1, VitalExtendToFillDelay(tipd_DEPTH1));
    VitalWireDelay (DEPTH0_ipd, DEPTH0, VitalExtendToFillDelay(tipd_DEPTH0));
    VitalWireDelay (WRAD15_ipd, WRAD15, VitalExtendToFillDelay(tipd_WRAD15));
    VitalWireDelay (WRAD14_ipd, WRAD14, VitalExtendToFillDelay(tipd_WRAD14));
    VitalWireDelay (WRAD13_ipd, WRAD13, VitalExtendToFillDelay(tipd_WRAD13));
    VitalWireDelay (WRAD12_ipd, WRAD12, VitalExtendToFillDelay(tipd_WRAD12));
    VitalWireDelay (WRAD11_ipd, WRAD11, VitalExtendToFillDelay(tipd_WRAD11));
    VitalWireDelay (WRAD10_ipd, WRAD10, VitalExtendToFillDelay(tipd_WRAD10));
    VitalWireDelay (WRAD9_ipd, WRAD9, VitalExtendToFillDelay(tipd_WRAD9));
    VitalWireDelay (WRAD8_ipd, WRAD8, VitalExtendToFillDelay(tipd_WRAD8));
    VitalWireDelay (WRAD7_ipd, WRAD7, VitalExtendToFillDelay(tipd_WRAD7));
    VitalWireDelay (WRAD6_ipd, WRAD6, VitalExtendToFillDelay(tipd_WRAD6));
    VitalWireDelay (WRAD5_ipd, WRAD5, VitalExtendToFillDelay(tipd_WRAD5));
    VitalWireDelay (WRAD4_ipd, WRAD4, VitalExtendToFillDelay(tipd_WRAD4));
    VitalWireDelay (WRAD3_ipd, WRAD3, VitalExtendToFillDelay(tipd_WRAD3));
    VitalWireDelay (WRAD2_ipd, WRAD2, VitalExtendToFillDelay(tipd_WRAD2));
    VitalWireDelay (WRAD1_ipd, WRAD1, VitalExtendToFillDelay(tipd_WRAD1));
    VitalWireDelay (WRAD0_ipd, WRAD0, VitalExtendToFillDelay(tipd_WRAD0));
    VitalWireDelay (WD35_ipd, WD35, VitalExtendToFillDelay(tipd_WD35));
    VitalWireDelay (WD34_ipd, WD34, VitalExtendToFillDelay(tipd_WD34));
    VitalWireDelay (WD33_ipd, WD33, VitalExtendToFillDelay(tipd_WD33));
    VitalWireDelay (WD32_ipd, WD32, VitalExtendToFillDelay(tipd_WD32));
    VitalWireDelay (WD31_ipd, WD31, VitalExtendToFillDelay(tipd_WD31));
    VitalWireDelay (WD30_ipd, WD30, VitalExtendToFillDelay(tipd_WD30));
    VitalWireDelay (WD29_ipd, WD29, VitalExtendToFillDelay(tipd_WD29));
    VitalWireDelay (WD28_ipd, WD28, VitalExtendToFillDelay(tipd_WD28));
    VitalWireDelay (WD27_ipd, WD27, VitalExtendToFillDelay(tipd_WD27));
    VitalWireDelay (WD26_ipd, WD26, VitalExtendToFillDelay(tipd_WD26));
    VitalWireDelay (WD25_ipd, WD25, VitalExtendToFillDelay(tipd_WD25));
    VitalWireDelay (WD24_ipd, WD24, VitalExtendToFillDelay(tipd_WD24));
    VitalWireDelay (WD23_ipd, WD23, VitalExtendToFillDelay(tipd_WD23));
    VitalWireDelay (WD22_ipd, WD22, VitalExtendToFillDelay(tipd_WD22));
    VitalWireDelay (WD21_ipd, WD21, VitalExtendToFillDelay(tipd_WD21));
    VitalWireDelay (WD20_ipd, WD20, VitalExtendToFillDelay(tipd_WD20));
    VitalWireDelay (WD19_ipd, WD19, VitalExtendToFillDelay(tipd_WD19));
    VitalWireDelay (WD18_ipd, WD18, VitalExtendToFillDelay(tipd_WD18));
    VitalWireDelay (WD17_ipd, WD17, VitalExtendToFillDelay(tipd_WD17));
    VitalWireDelay (WD16_ipd, WD16, VitalExtendToFillDelay(tipd_WD16));
    VitalWireDelay (WD15_ipd, WD15, VitalExtendToFillDelay(tipd_WD15));
    VitalWireDelay (WD14_ipd, WD14, VitalExtendToFillDelay(tipd_WD14));
    VitalWireDelay (WD13_ipd, WD13, VitalExtendToFillDelay(tipd_WD13));
    VitalWireDelay (WD12_ipd, WD12, VitalExtendToFillDelay(tipd_WD12));
    VitalWireDelay (WD11_ipd, WD11, VitalExtendToFillDelay(tipd_WD11));
    VitalWireDelay (WD10_ipd, WD10, VitalExtendToFillDelay(tipd_WD10));
    VitalWireDelay (WD9_ipd, WD9, VitalExtendToFillDelay(tipd_WD9));
    VitalWireDelay (WD8_ipd, WD8, VitalExtendToFillDelay(tipd_WD8));
    VitalWireDelay (WD7_ipd, WD7, VitalExtendToFillDelay(tipd_WD7));
    VitalWireDelay (WD6_ipd, WD6, VitalExtendToFillDelay(tipd_WD6));
    VitalWireDelay (WD5_ipd, WD5, VitalExtendToFillDelay(tipd_WD5));
    VitalWireDelay (WD4_ipd, WD4, VitalExtendToFillDelay(tipd_WD4));
    VitalWireDelay (WD3_ipd, WD3, VitalExtendToFillDelay(tipd_WD3));
    VitalWireDelay (WD2_ipd, WD2, VitalExtendToFillDelay(tipd_WD2));
    VitalWireDelay (WD1_ipd, WD1, VitalExtendToFillDelay(tipd_WD1));
    VitalWireDelay (WD0_ipd, WD0, VitalExtendToFillDelay(tipd_WD0));
    VitalWireDelay (WW2_ipd, WW2, VitalExtendToFillDelay(tipd_WW2));
    VitalWireDelay (WW1_ipd, WW1, VitalExtendToFillDelay(tipd_WW1));
    VitalWireDelay (WW0_ipd, WW0, VitalExtendToFillDelay(tipd_WW0));
    VitalWireDelay (WEN_ipd, WEN, VitalExtendToFillDelay(tipd_WEN));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (RDAD15_ipd, RDAD15, VitalExtendToFillDelay(tipd_RDAD15));
    VitalWireDelay (RDAD14_ipd, RDAD14, VitalExtendToFillDelay(tipd_RDAD14));
    VitalWireDelay (RDAD13_ipd, RDAD13, VitalExtendToFillDelay(tipd_RDAD13));
    VitalWireDelay (RDAD12_ipd, RDAD12, VitalExtendToFillDelay(tipd_RDAD12));
    VitalWireDelay (RDAD11_ipd, RDAD11, VitalExtendToFillDelay(tipd_RDAD11));
    VitalWireDelay (RDAD10_ipd, RDAD10, VitalExtendToFillDelay(tipd_RDAD10));
    VitalWireDelay (RDAD9_ipd, RDAD9, VitalExtendToFillDelay(tipd_RDAD9));
    VitalWireDelay (RDAD8_ipd, RDAD8, VitalExtendToFillDelay(tipd_RDAD8));
    VitalWireDelay (RDAD7_ipd, RDAD7, VitalExtendToFillDelay(tipd_RDAD7));
    VitalWireDelay (RDAD6_ipd, RDAD6, VitalExtendToFillDelay(tipd_RDAD6));
    VitalWireDelay (RDAD5_ipd, RDAD5, VitalExtendToFillDelay(tipd_RDAD5));
    VitalWireDelay (RDAD4_ipd, RDAD4, VitalExtendToFillDelay(tipd_RDAD4));
    VitalWireDelay (RDAD3_ipd, RDAD3, VitalExtendToFillDelay(tipd_RDAD3));
    VitalWireDelay (RDAD2_ipd, RDAD2, VitalExtendToFillDelay(tipd_RDAD2));
    VitalWireDelay (RDAD1_ipd, RDAD1, VitalExtendToFillDelay(tipd_RDAD1));
    VitalWireDelay (RDAD0_ipd, RDAD0, VitalExtendToFillDelay(tipd_RDAD0));
    VitalWireDelay (RW2_ipd, RW2, VitalExtendToFillDelay(tipd_RW2));
    VitalWireDelay (RW1_ipd, RW1, VitalExtendToFillDelay(tipd_RW1));
    VitalWireDelay (RW0_ipd, RW0, VitalExtendToFillDelay(tipd_RW0));
    VitalWireDelay (REN_ipd, REN, VitalExtendToFillDelay(tipd_REN));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (DEPTH3_ipd, DEPTH2_ipd, DEPTH1_ipd, DEPTH0_ipd,
                WRAD15_ipd, WRAD14_ipd, WRAD13_ipd,
                WRAD12_ipd, WRAD11_ipd, WRAD10_ipd, WRAD9_ipd, 
                WRAD8_ipd, WRAD7_ipd, WRAD6_ipd, WRAD5_ipd, 
                WRAD4_ipd, WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd, 
                WD35_ipd, WD34_ipd, WD33_ipd, WD32_ipd, WD31_ipd, WD30_ipd,
                WD29_ipd, WD28_ipd, WD27_ipd, WD26_ipd, WD25_ipd, WD24_ipd,
                WD23_ipd, WD22_ipd, WD21_ipd, WD20_ipd, WD19_ipd, WD18_ipd,
                WD17_ipd, WD16_ipd, WD15_ipd, WD14_ipd, WD13_ipd, WD12_ipd,
                WD11_ipd, WD10_ipd, WD9_ipd, WD8_ipd, WD7_ipd, WD6_ipd,
                WD5_ipd, WD4_ipd, WD3_ipd, WD2_ipd, WD1_ipd, WD0_ipd,
                WW2_ipd, WW1_ipd, WW0_ipd, WEN_ipd, WCLK_ipd, 
                RDAD15_ipd, RDAD14_ipd, RDAD13_ipd, RDAD12_ipd, RDAD11_ipd, 
                RDAD10_ipd, RDAD9_ipd, RDAD8_ipd, RDAD7_ipd,
                RDAD6_ipd, RDAD5_ipd, RDAD4_ipd, RDAD3_ipd, RDAD2_ipd, 
                RDAD1_ipd, RDAD0_ipd, RW2_ipd, RW1_ipd, RW0_ipd,
                REN_ipd, RCLK_ipd)

     --  Memory 
     variable RAM_TMP    : MEM;
     variable RAM_TMP9   : MEM9;
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT : SL_TO_INT := (-65537, -65537, 0, 1, -65537, -65537, 0, 1, -65537);

     --  Read Timing Check Results
     variable Tviol_RDAD15_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD15_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD14_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD14_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD13_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD13_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD12_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD12_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD11_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD11_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD10_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD10_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD9_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD9_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD8_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD8_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD7_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD7_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD6_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD6_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD5_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD5_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD4_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD4_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD3_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD3_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD2_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD1_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD0_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RW2_RCLK_posedge : X01 := '0';
     variable TmDt_RW2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RW1_RCLK_posedge : X01 := '0';
     variable TmDt_RW1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RW0_RCLK_posedge : X01 := '0';
     variable TmDt_RW0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_REN_RCLK_posedge : X01 := '0';
     variable TmDt_REN_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_WD35_WCLK_posedge : X01 := '0';
     variable TmDt_WD35_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD34_WCLK_posedge : X01 := '0';
     variable TmDt_WD34_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD33_WCLK_posedge : X01 := '0';
     variable TmDt_WD33_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD32_WCLK_posedge : X01 := '0';
     variable TmDt_WD32_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD31_WCLK_posedge : X01 := '0';
     variable TmDt_WD31_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD30_WCLK_posedge : X01 := '0';
     variable TmDt_WD30_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD29_WCLK_posedge : X01 := '0';
     variable TmDt_WD29_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD28_WCLK_posedge : X01 := '0';
     variable TmDt_WD28_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD27_WCLK_posedge : X01 := '0';
     variable TmDt_WD27_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD26_WCLK_posedge : X01 := '0';
     variable TmDt_WD26_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD25_WCLK_posedge : X01 := '0';
     variable TmDt_WD25_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD24_WCLK_posedge : X01 := '0';
     variable TmDt_WD24_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD23_WCLK_posedge : X01 := '0';
     variable TmDt_WD23_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD22_WCLK_posedge : X01 := '0';
     variable TmDt_WD22_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD21_WCLK_posedge : X01 := '0';
     variable TmDt_WD21_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD20_WCLK_posedge : X01 := '0';
     variable TmDt_WD20_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD19_WCLK_posedge : X01 := '0';
     variable TmDt_WD19_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD18_WCLK_posedge : X01 := '0';
     variable TmDt_WD18_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD17_WCLK_posedge : X01 := '0';
     variable TmDt_WD17_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD16_WCLK_posedge : X01 := '0';
     variable TmDt_WD16_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD15_WCLK_posedge : X01 := '0';
     variable TmDt_WD15_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD14_WCLK_posedge : X01 := '0';
     variable TmDt_WD14_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD13_WCLK_posedge : X01 := '0';
     variable TmDt_WD13_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD12_WCLK_posedge : X01 := '0';
     variable TmDt_WD12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD11_WCLK_posedge : X01 := '0';
     variable TmDt_WD11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD10_WCLK_posedge : X01 := '0';
     variable TmDt_WD10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD9_WCLK_posedge : X01 := '0';
     variable TmDt_WD9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD8_WCLK_posedge : X01 := '0';
     variable TmDt_WD8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD7_WCLK_posedge : X01 := '0';
     variable TmDt_WD7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD6_WCLK_posedge : X01 := '0';
     variable TmDt_WD6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD5_WCLK_posedge : X01 := '0';
     variable TmDt_WD5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD4_WCLK_posedge : X01 := '0';
     variable TmDt_WD4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD3_WCLK_posedge : X01 := '0';
     variable TmDt_WD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD2_WCLK_posedge : X01 := '0';
     variable TmDt_WD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD1_WCLK_posedge : X01 := '0';
     variable TmDt_WD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD0_WCLK_posedge : X01 := '0';
     variable TmDt_WD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WW2_WCLK_posedge : X01 := '0';
     variable TmDt_WW2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WW1_WCLK_posedge : X01 := '0';
     variable TmDt_WW1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WW0_WCLK_posedge : X01 := '0';
     variable TmDt_WW0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD15_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD15_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD14_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD14_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD13_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD13_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD12_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD11_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD10_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD9_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD8_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD7_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD6_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD5_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD4_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD3_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD2_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD1_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD0_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DEPTH3_WCLK_posedge : X01 := '0';
     variable TmDt_DEPTH3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DEPTH2_WCLK_posedge : X01 := '0';
     variable TmDt_DEPTH2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DEPTH1_WCLK_posedge : X01 := '0';
     variable TmDt_DEPTH1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DEPTH0_WCLK_posedge : X01 := '0';
     variable TmDt_DEPTH0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WEN_WCLK_posedge : X01 := '0';
     variable TmDt_WEN_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  Functional Results
     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     variable WWIDTH : integer := -1;
     variable RWIDTH : integer := -1;
     variable RD35_zd : std_ulogic;
     variable RD34_zd : std_ulogic;
     variable RD33_zd : std_ulogic;
     variable RD32_zd : std_ulogic;
     variable RD31_zd : std_ulogic;
     variable RD30_zd : std_ulogic;
     variable RD29_zd : std_ulogic;
     variable RD28_zd : std_ulogic;
     variable RD27_zd : std_ulogic;
     variable RD26_zd : std_ulogic;
     variable RD25_zd : std_ulogic;
     variable RD24_zd : std_ulogic;
     variable RD23_zd : std_ulogic;
     variable RD22_zd : std_ulogic;
     variable RD21_zd : std_ulogic;
     variable RD20_zd : std_ulogic;
     variable RD19_zd : std_ulogic;
     variable RD18_zd : std_ulogic;
     variable RD17_zd : std_ulogic;
     variable RD16_zd : std_ulogic;
     variable RD15_zd : std_ulogic;
     variable RD14_zd : std_ulogic;
     variable RD13_zd : std_ulogic;
     variable RD12_zd : std_ulogic;
     variable RD11_zd : std_ulogic;
     variable RD10_zd : std_ulogic;
     variable RD9_zd : std_ulogic;
     variable RD8_zd : std_ulogic;
     variable RD7_zd : std_ulogic;
     variable RD6_zd : std_ulogic;
     variable RD5_zd : std_ulogic;
     variable RD4_zd : std_ulogic;
     variable RD3_zd : std_ulogic;
     variable RD2_zd : std_ulogic;
     variable RD1_zd : std_ulogic;
     variable RD0_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable RD35_GlitchData : VitalGlitchDataType;
     variable RD34_GlitchData : VitalGlitchDataType;
     variable RD33_GlitchData : VitalGlitchDataType;
     variable RD32_GlitchData : VitalGlitchDataType;
     variable RD31_GlitchData : VitalGlitchDataType;
     variable RD30_GlitchData : VitalGlitchDataType;
     variable RD29_GlitchData : VitalGlitchDataType;
     variable RD28_GlitchData : VitalGlitchDataType;
     variable RD27_GlitchData : VitalGlitchDataType;
     variable RD26_GlitchData : VitalGlitchDataType;
     variable RD25_GlitchData : VitalGlitchDataType;
     variable RD24_GlitchData : VitalGlitchDataType;
     variable RD23_GlitchData : VitalGlitchDataType;
     variable RD22_GlitchData : VitalGlitchDataType;
     variable RD21_GlitchData : VitalGlitchDataType;
     variable RD20_GlitchData : VitalGlitchDataType;
     variable RD19_GlitchData : VitalGlitchDataType;
     variable RD18_GlitchData : VitalGlitchDataType;
     variable RD17_GlitchData : VitalGlitchDataType;
     variable RD16_GlitchData : VitalGlitchDataType;
     variable RD15_GlitchData : VitalGlitchDataType;
     variable RD14_GlitchData : VitalGlitchDataType;
     variable RD13_GlitchData : VitalGlitchDataType;
     variable RD12_GlitchData : VitalGlitchDataType;
     variable RD11_GlitchData : VitalGlitchDataType;
     variable RD10_GlitchData : VitalGlitchDataType;
     variable RD9_GlitchData : VitalGlitchDataType;
     variable RD8_GlitchData : VitalGlitchDataType;
     variable RD7_GlitchData : VitalGlitchDataType;
     variable RD6_GlitchData : VitalGlitchDataType;
     variable RD5_GlitchData : VitalGlitchDataType;
     variable RD4_GlitchData : VitalGlitchDataType;
     variable RD3_GlitchData : VitalGlitchDataType;
     variable RD2_GlitchData : VitalGlitchDataType;
     variable RD1_GlitchData : VitalGlitchDataType;
     variable RD0_GlitchData : VitalGlitchDataType;

     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable REN_delayed  : std_ulogic := 'X';
     variable REN_previous : std_ulogic := 'X';
     variable WEN_delayed  : std_ulogic := 'X';
     variable WD35_delayed : std_ulogic := 'X';
     variable WD34_delayed : std_ulogic := 'X';
     variable WD33_delayed : std_ulogic := 'X';
     variable WD32_delayed : std_ulogic := 'X';
     variable WD31_delayed : std_ulogic := 'X';
     variable WD30_delayed : std_ulogic := 'X';
     variable WD29_delayed : std_ulogic := 'X';
     variable WD28_delayed : std_ulogic := 'X';
     variable WD27_delayed : std_ulogic := 'X';
     variable WD26_delayed : std_ulogic := 'X';
     variable WD25_delayed : std_ulogic := 'X';
     variable WD24_delayed : std_ulogic := 'X';
     variable WD23_delayed : std_ulogic := 'X';
     variable WD22_delayed : std_ulogic := 'X';
     variable WD21_delayed : std_ulogic := 'X';
     variable WD20_delayed : std_ulogic := 'X';
     variable WD19_delayed : std_ulogic := 'X';
     variable WD18_delayed : std_ulogic := 'X';
     variable WD17_delayed : std_ulogic := 'X';
     variable WD16_delayed : std_ulogic := 'X';
     variable WD15_delayed : std_ulogic := 'X';
     variable WD14_delayed : std_ulogic := 'X';
     variable WD13_delayed : std_ulogic := 'X';
     variable WD12_delayed : std_ulogic := 'X';
     variable WD11_delayed : std_ulogic := 'X';
     variable WD10_delayed : std_ulogic := 'X';
     variable WD9_delayed : std_ulogic := 'X';
     variable WD8_delayed : std_ulogic := 'X';
     variable WD7_delayed : std_ulogic := 'X';
     variable WD6_delayed : std_ulogic := 'X';
     variable WD5_delayed : std_ulogic := 'X';
     variable WD4_delayed : std_ulogic := 'X';
     variable WD3_delayed : std_ulogic := 'X';
     variable WD2_delayed : std_ulogic := 'X';
     variable WD1_delayed : std_ulogic := 'X';
     variable WD0_delayed : std_ulogic := 'X';
     variable WW2_delayed : std_ulogic := 'X';
     variable WW1_delayed : std_ulogic := 'X';
     variable WW0_delayed : std_ulogic := 'X';
     variable DEPTH3_delayed : std_ulogic := 'X';
     variable DEPTH2_delayed : std_ulogic := 'X';
     variable DEPTH1_delayed : std_ulogic := 'X';
     variable DEPTH0_delayed : std_ulogic := 'X';
     variable WRAD15_delayed : std_ulogic := 'X';
     variable WRAD14_delayed : std_ulogic := 'X';
     variable WRAD13_delayed : std_ulogic := 'X';
     variable WRAD12_delayed : std_ulogic := 'X';
     variable WRAD11_delayed : std_ulogic := 'X';
     variable WRAD10_delayed : std_ulogic := 'X';
     variable WRAD9_delayed : std_ulogic := 'X';
     variable WRAD8_delayed : std_ulogic := 'X';
     variable WRAD7_delayed : std_ulogic := 'X';
     variable WRAD6_delayed : std_ulogic := 'X';
     variable WRAD5_delayed : std_ulogic := 'X';
     variable WRAD4_delayed : std_ulogic := 'X';
     variable WRAD3_delayed : std_ulogic := 'X';
     variable WRAD2_delayed : std_ulogic := 'X';
     variable WRAD1_delayed : std_ulogic := 'X';
     variable WRAD0_delayed : std_ulogic := 'X';
     variable RDAD15_delayed : std_ulogic := 'X';
     variable RDAD14_delayed : std_ulogic := 'X';
     variable RDAD13_delayed : std_ulogic := 'X';
     variable RDAD12_delayed : std_ulogic := 'X';
     variable RDAD11_delayed : std_ulogic := 'X';
     variable RDAD10_delayed : std_ulogic := 'X';
     variable RDAD9_delayed : std_ulogic := 'X';
     variable RDAD8_delayed : std_ulogic := 'X';
     variable RDAD7_delayed : std_ulogic := 'X';
     variable RDAD6_delayed : std_ulogic := 'X';
     variable RDAD5_delayed : std_ulogic := 'X';
     variable RDAD4_delayed : std_ulogic := 'X';
     variable RDAD3_delayed : std_ulogic := 'X';
     variable RDAD2_delayed : std_ulogic := 'X';
     variable RDAD1_delayed : std_ulogic := 'X';
     variable RDAD0_delayed : std_ulogic := 'X';
     variable RW2_delayed : std_ulogic := 'X';
     variable RW1_delayed : std_ulogic := 'X';
     variable RW0_delayed : std_ulogic := 'X';
     variable RDAD15_previous : std_ulogic := 'X';
     variable RDAD14_previous : std_ulogic := 'X';
     variable RDAD13_previous : std_ulogic := 'X';
     variable RDAD12_previous : std_ulogic := 'X';
     variable RDAD11_previous : std_ulogic := 'X';
     variable RDAD10_previous : std_ulogic := 'X';
     variable RDAD9_previous : std_ulogic := 'X';
     variable RDAD8_previous : std_ulogic := 'X';
     variable RDAD7_previous : std_ulogic := 'X';
     variable RDAD6_previous : std_ulogic := 'X';
     variable RDAD5_previous : std_ulogic := 'X';
     variable RDAD4_previous : std_ulogic := 'X';
     variable RDAD3_previous : std_ulogic := 'X';
     variable RDAD2_previous : std_ulogic := 'X';
     variable RDAD1_previous : std_ulogic := 'X';
     variable RDAD0_previous : std_ulogic := 'X';
     variable RW2_previous : std_ulogic := 'X';
     variable RW1_previous : std_ulogic := 'X';
     variable RW0_previous : std_ulogic := 'X';

  begin  --  process VITALBehavior 


    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RDAD high or low before RCLK rising
      --   Hold  RDAD high or low after RCLK rising

      VitalSetupHoldCheck ( Tviol_RDAD15_RCLK_posedge,
                            TmDt_RDAD15_RCLK_posedge,
                            RDAD15_ipd, "RDAD15",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD15_RCLK_posedge_posedge,
                            tsetup_RDAD15_RCLK_negedge_posedge,
                            thold_RDAD15_RCLK_posedge_posedge,
                            thold_RDAD15_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD14_RCLK_posedge,
                            TmDt_RDAD14_RCLK_posedge,
                            RDAD14_ipd, "RDAD14",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD14_RCLK_posedge_posedge,
                            tsetup_RDAD14_RCLK_negedge_posedge,
                            thold_RDAD14_RCLK_posedge_posedge,
                            thold_RDAD14_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD13_RCLK_posedge,
                            TmDt_RDAD13_RCLK_posedge,
                            RDAD13_ipd, "RDAD13",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD13_RCLK_posedge_posedge,
                            tsetup_RDAD13_RCLK_negedge_posedge,
                            thold_RDAD13_RCLK_posedge_posedge,
                            thold_RDAD13_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD12_RCLK_posedge,
                            TmDt_RDAD12_RCLK_posedge,
                            RDAD12_ipd, "RDAD12",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD12_RCLK_posedge_posedge,
                            tsetup_RDAD12_RCLK_negedge_posedge,
                            thold_RDAD12_RCLK_posedge_posedge,
                            thold_RDAD12_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD11_RCLK_posedge,
                            TmDt_RDAD11_RCLK_posedge,
                            RDAD11_ipd, "RDAD11",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD11_RCLK_posedge_posedge,
                            tsetup_RDAD11_RCLK_negedge_posedge,
                            thold_RDAD11_RCLK_posedge_posedge,
                            thold_RDAD11_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD10_RCLK_posedge,
                            TmDt_RDAD10_RCLK_posedge,
                            RDAD10_ipd, "RDAD10",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD10_RCLK_posedge_posedge,
                            tsetup_RDAD10_RCLK_negedge_posedge,
                            thold_RDAD10_RCLK_posedge_posedge,
                            thold_RDAD10_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD9_RCLK_posedge,
                            TmDt_RDAD9_RCLK_posedge,
                            RDAD9_ipd, "RDAD9",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD9_RCLK_posedge_posedge,
                            tsetup_RDAD9_RCLK_negedge_posedge,
                            thold_RDAD9_RCLK_posedge_posedge,
                            thold_RDAD9_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD8_RCLK_posedge,
                            TmDt_RDAD8_RCLK_posedge,
                            RDAD8_ipd, "RDAD8",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD8_RCLK_posedge_posedge,
                            tsetup_RDAD8_RCLK_negedge_posedge,
                            thold_RDAD8_RCLK_posedge_posedge,
                            thold_RDAD8_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD7_RCLK_posedge,
                            TmDt_RDAD7_RCLK_posedge,
                            RDAD7_ipd, "RDAD7",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD7_RCLK_posedge_posedge,
                            tsetup_RDAD7_RCLK_negedge_posedge,
                            thold_RDAD7_RCLK_posedge_posedge,
                            thold_RDAD7_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD6_RCLK_posedge,
                            TmDt_RDAD6_RCLK_posedge,
                            RDAD6_ipd, "RDAD6",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD6_RCLK_posedge_posedge,
                            tsetup_RDAD6_RCLK_negedge_posedge,
                            thold_RDAD6_RCLK_posedge_posedge,
                            thold_RDAD6_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD5_RCLK_posedge,
                            TmDt_RDAD5_RCLK_posedge,
                            RDAD5_ipd, "RDAD5",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD5_RCLK_posedge_posedge,
                            tsetup_RDAD5_RCLK_negedge_posedge,
                            thold_RDAD5_RCLK_posedge_posedge,
                            thold_RDAD5_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD4_RCLK_posedge,
                            TmDt_RDAD4_RCLK_posedge,
                            RDAD4_ipd, "RDAD4",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD4_RCLK_posedge_posedge,
                            tsetup_RDAD4_RCLK_negedge_posedge,
                            thold_RDAD4_RCLK_posedge_posedge,
                            thold_RDAD4_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD3_RCLK_posedge,
                            TmDt_RDAD3_RCLK_posedge,
                            RDAD3_ipd, "RDAD3",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD3_RCLK_posedge_posedge,
                            tsetup_RDAD3_RCLK_negedge_posedge,
                            thold_RDAD3_RCLK_posedge_posedge,
                            thold_RDAD3_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD2_RCLK_posedge,
                            TmDt_RDAD2_RCLK_posedge,
                            RDAD2_ipd, "RDAD2",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD2_RCLK_posedge_posedge,
                            tsetup_RDAD2_RCLK_negedge_posedge,
                            thold_RDAD2_RCLK_posedge_posedge,
                            thold_RDAD2_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD1_RCLK_posedge,
                            TmDt_RDAD1_RCLK_posedge,
                            RDAD1_ipd, "RDAD1",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD1_RCLK_posedge_posedge,
                            tsetup_RDAD1_RCLK_negedge_posedge,
                            thold_RDAD1_RCLK_posedge_posedge,
                            thold_RDAD1_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD0_RCLK_posedge,
                            TmDt_RDAD0_RCLK_posedge,
                            RDAD0_ipd, "RDAD0",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD0_RCLK_posedge_posedge,
                            tsetup_RDAD0_RCLK_negedge_posedge,
                            thold_RDAD0_RCLK_posedge_posedge,
                            thold_RDAD0_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup RW high before RCLK rising
      --   Hold  RW high after RCLK rising

      VitalSetupHoldCheck ( Tviol_RW2_RCLK_posedge,
                            TmDt_RW2_RCLK_posedge,
                            RW2_ipd, "RW2",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RW2_RCLK_posedge_posedge,
                            tsetup_RW2_RCLK_negedge_posedge,
                            thold_RW2_RCLK_posedge_posedge,
                            thold_RW2_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RW1_RCLK_posedge,
                            TmDt_RW1_RCLK_posedge,
                            RW1_ipd, "RW1",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RW1_RCLK_posedge_posedge,
                            tsetup_RW1_RCLK_negedge_posedge,
                            thold_RW1_RCLK_posedge_posedge,
                            thold_RW1_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RW0_RCLK_posedge,
                            TmDt_RW0_RCLK_posedge,
                            RW0_ipd, "RW0",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RW0_RCLK_posedge_posedge,
                            tsetup_RW0_RCLK_negedge_posedge,
                            thold_RW0_RCLK_posedge_posedge,
                            thold_RW0_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup REN high before RCLK rising
      --   Hold  REN high after RCLK rising

      VitalSetupHoldCheck ( Tviol_REN_RCLK_posedge,
                            TmDt_REN_RCLK_posedge,
                            REN_ipd, "REN",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_REN_RCLK_posedge_posedge,
			    tsetup_REN_RCLK_negedge_posedge,
                            thold_REN_RCLK_posedge_posedge,
                            thold_REN_RCLK_negedge_posedge,
                            TimingCheckOn,
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup DEPTH high or low before WCLK rising
      --   Hold  DEPTH high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_DEPTH3_WCLK_posedge,
                            TmDt_DEPTH3_WCLK_posedge,
                            DEPTH3_ipd, "DEPTH3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_DEPTH3_WCLK_posedge_posedge,
                            tsetup_DEPTH3_WCLK_negedge_posedge,
                            thold_DEPTH3_WCLK_posedge_posedge,
                            thold_DEPTH3_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_DEPTH2_WCLK_posedge,
                            TmDt_DEPTH2_WCLK_posedge,
                            DEPTH2_ipd, "DEPTH2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_DEPTH2_WCLK_posedge_posedge,
                            tsetup_DEPTH2_WCLK_negedge_posedge,
                            thold_DEPTH2_WCLK_posedge_posedge,
                            thold_DEPTH2_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_DEPTH1_WCLK_posedge,
                            TmDt_DEPTH1_WCLK_posedge,
                            DEPTH1_ipd, "DEPTH1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_DEPTH1_WCLK_posedge_posedge,
                            tsetup_DEPTH1_WCLK_negedge_posedge,
                            thold_DEPTH1_WCLK_posedge_posedge,
                            thold_DEPTH1_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_DEPTH0_WCLK_posedge,
                            TmDt_DEPTH0_WCLK_posedge,
                            DEPTH0_ipd, "DEPTH0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_DEPTH0_WCLK_posedge_posedge,
                            tsetup_DEPTH0_WCLK_negedge_posedge,
                            thold_DEPTH0_WCLK_posedge_posedge,
                            thold_DEPTH0_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      --   Setup WRAD high or low before WCLK rising
      --   Hold  WRAD high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WRAD15_WCLK_posedge,
                            TmDt_WRAD15_WCLK_posedge,
                            WRAD15_ipd, "WRAD15",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD15_WCLK_posedge_posedge,
                            tsetup_WRAD15_WCLK_negedge_posedge,
                            thold_WRAD15_WCLK_posedge_posedge,
                            thold_WRAD15_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD14_WCLK_posedge,
                            TmDt_WRAD14_WCLK_posedge,
                            WRAD14_ipd, "WRAD14",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD14_WCLK_posedge_posedge,
                            tsetup_WRAD14_WCLK_negedge_posedge,
                            thold_WRAD14_WCLK_posedge_posedge,
                            thold_WRAD14_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD13_WCLK_posedge,
                            TmDt_WRAD13_WCLK_posedge,
                            WRAD13_ipd, "WRAD13",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD13_WCLK_posedge_posedge,
                            tsetup_WRAD13_WCLK_negedge_posedge,
                            thold_WRAD13_WCLK_posedge_posedge,
                            thold_WRAD13_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD12_WCLK_posedge,
                            TmDt_WRAD12_WCLK_posedge,
                            WRAD12_ipd, "WRAD12",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD12_WCLK_posedge_posedge,
                            tsetup_WRAD12_WCLK_negedge_posedge,
                            thold_WRAD12_WCLK_posedge_posedge,
                            thold_WRAD12_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD11_WCLK_posedge,
                            TmDt_WRAD11_WCLK_posedge,
                            WRAD11_ipd, "WRAD11",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD11_WCLK_posedge_posedge,
                            tsetup_WRAD11_WCLK_negedge_posedge,
                            thold_WRAD11_WCLK_posedge_posedge,
                            thold_WRAD11_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD10_WCLK_posedge,
                            TmDt_WRAD10_WCLK_posedge,
                            WRAD10_ipd, "WRAD10",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD10_WCLK_posedge_posedge,
                            tsetup_WRAD10_WCLK_negedge_posedge,
                            thold_WRAD10_WCLK_posedge_posedge,
                            thold_WRAD10_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD9_WCLK_posedge,
                            TmDt_WRAD9_WCLK_posedge,
                            WRAD9_ipd, "WRAD9",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD9_WCLK_posedge_posedge,
                            tsetup_WRAD9_WCLK_negedge_posedge,
                            thold_WRAD9_WCLK_posedge_posedge,
                            thold_WRAD9_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD8_WCLK_posedge,
                            TmDt_WRAD8_WCLK_posedge,
                            WRAD8_ipd, "WRAD8",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD8_WCLK_posedge_posedge,
                            tsetup_WRAD8_WCLK_negedge_posedge,
                            thold_WRAD8_WCLK_posedge_posedge,
                            thold_WRAD8_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD7_WCLK_posedge,
                            TmDt_WRAD7_WCLK_posedge,
                            WRAD7_ipd, "WRAD7",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD7_WCLK_posedge_posedge,
                            tsetup_WRAD7_WCLK_negedge_posedge,
                            thold_WRAD7_WCLK_posedge_posedge,
                            thold_WRAD7_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD6_WCLK_posedge,
                            TmDt_WRAD6_WCLK_posedge,
                            WRAD6_ipd, "WRAD6",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD6_WCLK_posedge_posedge,
                            tsetup_WRAD6_WCLK_negedge_posedge,
                            thold_WRAD6_WCLK_posedge_posedge,
                            thold_WRAD6_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD5_WCLK_posedge,
                            TmDt_WRAD5_WCLK_posedge,
                            WRAD5_ipd, "WRAD5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD5_WCLK_posedge_posedge,
                            tsetup_WRAD5_WCLK_negedge_posedge,
                            thold_WRAD5_WCLK_posedge_posedge,
                            thold_WRAD5_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD4_WCLK_posedge,
                            TmDt_WRAD4_WCLK_posedge,
                            WRAD4_ipd, "WRAD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD4_WCLK_posedge_posedge,
                            tsetup_WRAD4_WCLK_negedge_posedge,
                            thold_WRAD4_WCLK_posedge_posedge,
                            thold_WRAD4_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD3_WCLK_posedge,
                            TmDt_WRAD3_WCLK_posedge,
                            WRAD3_ipd, "WRAD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD3_WCLK_posedge_posedge,
                            tsetup_WRAD3_WCLK_negedge_posedge,
                            thold_WRAD3_WCLK_posedge_posedge,
                            thold_WRAD3_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD2_WCLK_posedge,
                            TmDt_WRAD2_WCLK_posedge,
                            WRAD2_ipd, "WRAD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD2_WCLK_posedge_posedge,
                            tsetup_WRAD2_WCLK_negedge_posedge,
                            thold_WRAD2_WCLK_posedge_posedge,
                            thold_WRAD2_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD1_WCLK_posedge,
                            TmDt_WRAD1_WCLK_posedge,
                            WRAD1_ipd, "WRAD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD1_WCLK_posedge_posedge,
                            tsetup_WRAD1_WCLK_negedge_posedge,
                            thold_WRAD1_WCLK_posedge_posedge,
                            thold_WRAD1_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD0_WCLK_posedge,
                            TmDt_WRAD0_WCLK_posedge,
                            WRAD0_ipd, "WRAD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD0_WCLK_posedge_posedge,
                            tsetup_WRAD0_WCLK_negedge_posedge,
                            thold_WRAD0_WCLK_posedge_posedge,
                            thold_WRAD0_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      --   Setup WD high or low before WCLK rising
      --   Hold  WD high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WD35_WCLK_posedge,
                            TmDt_WD35_WCLK_posedge,
                            WD35_ipd, "WD35",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD35_WCLK_posedge_posedge,
                            tsetup_WD35_WCLK_negedge_posedge,
                            thold_WD35_WCLK_posedge_posedge,
                            thold_WD35_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD34_WCLK_posedge,
                            TmDt_WD34_WCLK_posedge,
                            WD34_ipd, "WD34",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD34_WCLK_posedge_posedge,
                            tsetup_WD34_WCLK_negedge_posedge,
                            thold_WD34_WCLK_posedge_posedge,
                            thold_WD34_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD33_WCLK_posedge,
                            TmDt_WD33_WCLK_posedge,
                            WD33_ipd, "WD33",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD33_WCLK_posedge_posedge,
                            tsetup_WD33_WCLK_negedge_posedge,
                            thold_WD33_WCLK_posedge_posedge,
                            thold_WD33_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD32_WCLK_posedge,
                            TmDt_WD32_WCLK_posedge,
                            WD32_ipd, "WD32",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD32_WCLK_posedge_posedge,
                            tsetup_WD32_WCLK_negedge_posedge,
                            thold_WD32_WCLK_posedge_posedge,
                            thold_WD32_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD31_WCLK_posedge,
                            TmDt_WD31_WCLK_posedge,
                            WD31_ipd, "WD31",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD31_WCLK_posedge_posedge,
                            tsetup_WD31_WCLK_negedge_posedge,
                            thold_WD31_WCLK_posedge_posedge,
                            thold_WD31_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD30_WCLK_posedge,
                            TmDt_WD30_WCLK_posedge,
                            WD30_ipd, "WD30",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD30_WCLK_posedge_posedge,
                            tsetup_WD30_WCLK_negedge_posedge,
                            thold_WD30_WCLK_posedge_posedge,
                            thold_WD30_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD29_WCLK_posedge,
                            TmDt_WD29_WCLK_posedge,
                            WD29_ipd, "WD29",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD29_WCLK_posedge_posedge,
                            tsetup_WD29_WCLK_negedge_posedge,
                            thold_WD29_WCLK_posedge_posedge,
                            thold_WD29_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD28_WCLK_posedge,
                            TmDt_WD28_WCLK_posedge,
                            WD28_ipd, "WD28",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD28_WCLK_posedge_posedge,
                            tsetup_WD28_WCLK_negedge_posedge,
                            thold_WD28_WCLK_posedge_posedge,
                            thold_WD28_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD27_WCLK_posedge,
                            TmDt_WD27_WCLK_posedge,
                            WD27_ipd, "WD27",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD27_WCLK_posedge_posedge,
                            tsetup_WD27_WCLK_negedge_posedge,
                            thold_WD27_WCLK_posedge_posedge,
                            thold_WD27_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD26_WCLK_posedge,
                            TmDt_WD26_WCLK_posedge,
                            WD26_ipd, "WD26",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD26_WCLK_posedge_posedge,
                            tsetup_WD26_WCLK_negedge_posedge,
                            thold_WD26_WCLK_posedge_posedge,
                            thold_WD26_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD25_WCLK_posedge,
                            TmDt_WD25_WCLK_posedge,
                            WD25_ipd, "WD25",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD25_WCLK_posedge_posedge,
                            tsetup_WD25_WCLK_negedge_posedge,
                            thold_WD25_WCLK_posedge_posedge,
                            thold_WD25_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD24_WCLK_posedge,
                            TmDt_WD24_WCLK_posedge,
                            WD24_ipd, "WD24",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD24_WCLK_posedge_posedge,
                            tsetup_WD24_WCLK_negedge_posedge,
                            thold_WD24_WCLK_posedge_posedge,
                            thold_WD24_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD23_WCLK_posedge,
                            TmDt_WD23_WCLK_posedge,
                            WD23_ipd, "WD23",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD23_WCLK_posedge_posedge,
                            tsetup_WD23_WCLK_negedge_posedge,
                            thold_WD23_WCLK_posedge_posedge,
                            thold_WD23_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD22_WCLK_posedge,
                            TmDt_WD22_WCLK_posedge,
                            WD22_ipd, "WD22",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD22_WCLK_posedge_posedge,
                            tsetup_WD22_WCLK_negedge_posedge,
                            thold_WD22_WCLK_posedge_posedge,
                            thold_WD22_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD21_WCLK_posedge,
                            TmDt_WD21_WCLK_posedge,
                            WD21_ipd, "WD21",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD21_WCLK_posedge_posedge,
                            tsetup_WD21_WCLK_negedge_posedge,
                            thold_WD21_WCLK_posedge_posedge,
                            thold_WD21_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD20_WCLK_posedge,
                            TmDt_WD20_WCLK_posedge,
                            WD20_ipd, "WD20",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD20_WCLK_posedge_posedge,
                            tsetup_WD20_WCLK_negedge_posedge,
                            thold_WD20_WCLK_posedge_posedge,
                            thold_WD20_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD19_WCLK_posedge,
                            TmDt_WD19_WCLK_posedge,
                            WD19_ipd, "WD19",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD19_WCLK_posedge_posedge,
                            tsetup_WD19_WCLK_negedge_posedge,
                            thold_WD19_WCLK_posedge_posedge,
                            thold_WD19_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD18_WCLK_posedge,
                            TmDt_WD18_WCLK_posedge,
                            WD18_ipd, "WD18",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD18_WCLK_posedge_posedge,
                            tsetup_WD18_WCLK_negedge_posedge,
                            thold_WD18_WCLK_posedge_posedge,
                            thold_WD18_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD17_WCLK_posedge,
                            TmDt_WD17_WCLK_posedge,
                            WD17_ipd, "WD17",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD17_WCLK_posedge_posedge,
                            tsetup_WD17_WCLK_negedge_posedge,
                            thold_WD17_WCLK_posedge_posedge,
                            thold_WD17_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD16_WCLK_posedge,
                            TmDt_WD16_WCLK_posedge,
                            WD16_ipd, "WD16",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD16_WCLK_posedge_posedge,
                            tsetup_WD16_WCLK_negedge_posedge,
                            thold_WD16_WCLK_posedge_posedge,
                            thold_WD16_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD15_WCLK_posedge,
                            TmDt_WD15_WCLK_posedge,
                            WD15_ipd, "WD15",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD15_WCLK_posedge_posedge,
                            tsetup_WD15_WCLK_negedge_posedge,
                            thold_WD15_WCLK_posedge_posedge,
                            thold_WD15_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD14_WCLK_posedge,
                            TmDt_WD14_WCLK_posedge,
                            WD14_ipd, "WD14",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD14_WCLK_posedge_posedge,
                            tsetup_WD14_WCLK_negedge_posedge,
                            thold_WD14_WCLK_posedge_posedge,
                            thold_WD14_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD13_WCLK_posedge,
                            TmDt_WD13_WCLK_posedge,
                            WD13_ipd, "WD13",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD13_WCLK_posedge_posedge,
                            tsetup_WD13_WCLK_negedge_posedge,
                            thold_WD13_WCLK_posedge_posedge,
                            thold_WD13_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD12_WCLK_posedge,
                            TmDt_WD12_WCLK_posedge,
                            WD12_ipd, "WD12",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD12_WCLK_posedge_posedge,
                            tsetup_WD12_WCLK_negedge_posedge,
                            thold_WD12_WCLK_posedge_posedge,
                            thold_WD12_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD11_WCLK_posedge,
                            TmDt_WD11_WCLK_posedge,
                            WD11_ipd, "WD11",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD11_WCLK_posedge_posedge,
                            tsetup_WD11_WCLK_negedge_posedge,
                            thold_WD11_WCLK_posedge_posedge,
                            thold_WD11_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD10_WCLK_posedge,
                            TmDt_WD10_WCLK_posedge,
                            WD10_ipd, "WD10",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD10_WCLK_posedge_posedge,
                            tsetup_WD10_WCLK_negedge_posedge,
                            thold_WD10_WCLK_posedge_posedge,
                            thold_WD10_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD9_WCLK_posedge,
                            TmDt_WD9_WCLK_posedge,
                            WD9_ipd, "WD9",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD9_WCLK_posedge_posedge,
                            tsetup_WD9_WCLK_negedge_posedge,
                            thold_WD9_WCLK_posedge_posedge,
                            thold_WD9_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD8_WCLK_posedge,
                            TmDt_WD8_WCLK_posedge,
                            WD8_ipd, "WD8",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD8_WCLK_posedge_posedge,
                            tsetup_WD8_WCLK_negedge_posedge,
                            thold_WD8_WCLK_posedge_posedge,
                            thold_WD8_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD7_WCLK_posedge,
                            TmDt_WD7_WCLK_posedge,
                            WD7_ipd, "WD7",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD7_WCLK_posedge_posedge,
                            tsetup_WD7_WCLK_negedge_posedge,
                            thold_WD7_WCLK_posedge_posedge,
                            thold_WD7_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD6_WCLK_posedge,
                            TmDt_WD6_WCLK_posedge,
                            WD6_ipd, "WD6",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD6_WCLK_posedge_posedge,
                            tsetup_WD6_WCLK_negedge_posedge,
                            thold_WD6_WCLK_posedge_posedge,
                            thold_WD6_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD5_WCLK_posedge,
                            TmDt_WD5_WCLK_posedge,
                            WD5_ipd, "WD5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD5_WCLK_posedge_posedge,
                            tsetup_WD5_WCLK_negedge_posedge,
                            thold_WD5_WCLK_posedge_posedge,
                            thold_WD5_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD4_WCLK_posedge,
                            TmDt_WD4_WCLK_posedge,
                            WD4_ipd, "WD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD4_WCLK_posedge_posedge,
                            tsetup_WD4_WCLK_negedge_posedge,
                            thold_WD4_WCLK_posedge_posedge,
                            thold_WD4_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD3_WCLK_posedge,
                            TmDt_WD3_WCLK_posedge,
                            WD3_ipd, "WD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD3_WCLK_posedge_posedge,
                            tsetup_WD3_WCLK_negedge_posedge,
                            thold_WD3_WCLK_posedge_posedge,
                            thold_WD3_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD2_WCLK_posedge,
                            TmDt_WD2_WCLK_posedge,
                            WD2_ipd, "WD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD2_WCLK_posedge_posedge,
                            tsetup_WD2_WCLK_negedge_posedge,
                            thold_WD2_WCLK_posedge_posedge,
                            thold_WD2_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD1_WCLK_posedge,
                            TmDt_WD1_WCLK_posedge,
                            WD1_ipd, "WD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD1_WCLK_posedge_posedge,
                            tsetup_WD1_WCLK_negedge_posedge,
                            thold_WD1_WCLK_posedge_posedge,
                            thold_WD1_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD0_WCLK_posedge,
                            TmDt_WD0_WCLK_posedge,
                            WD0_ipd, "WD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD0_WCLK_posedge_posedge,
                            tsetup_WD0_WCLK_negedge_posedge,
                            thold_WD0_WCLK_posedge_posedge,
                            thold_WD0_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup WW high or low before WCLK rising
      --   Hold  WW high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WW2_WCLK_posedge,
                            TmDt_WW2_WCLK_posedge,
                            WW2_ipd, "WW2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WW2_WCLK_posedge_posedge,
                            tsetup_WW2_WCLK_negedge_posedge,
                            thold_WW2_WCLK_posedge_posedge,
                            thold_WW2_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WW1_WCLK_posedge,
                            TmDt_WW1_WCLK_posedge,
                            WW1_ipd, "WW1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WW1_WCLK_posedge_posedge,
                            tsetup_WW1_WCLK_negedge_posedge,
                            thold_WW1_WCLK_posedge_posedge,
                            thold_WW1_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WW0_WCLK_posedge,
                            TmDt_WW0_WCLK_posedge,
                            WW0_ipd, "WW0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WW0_WCLK_posedge_posedge,
                            tsetup_WW0_WCLK_negedge_posedge,
                            thold_WW0_WCLK_posedge_posedge,
                            thold_WW0_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup WEN high before WCLK rising
      --   Hold  WEN high after WCLK rising

      VitalSetupHoldCheck ( Tviol_WEN_WCLK_posedge,
                            TmDt_WEN_WCLK_posedge,
                            WEN_ipd, "WEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WEN_WCLK_posedge_posedge,
                            tsetup_WEN_WCLK_negedge_posedge,
                            thold_WEN_WCLK_posedge_posedge,
                            thold_WEN_WCLK_negedge_posedge,
                            TimingCheckOn,
                            '/',
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM64K36",
                            Xon,
                            MsgOn,
                            WARNING
                            );
    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################

      -- Decode Write Word Width
      if (TO_X01(WW2_delayed)='0' and TO_X01(WW1_delayed)='0' and TO_X01(WW0_delayed)='0') then
        WWIDTH := 1;
      elsif (TO_X01(WW2_delayed)='0' and TO_X01(WW1_delayed)='0' and TO_X01(WW0_delayed)='1') then
        WWIDTH := 2;
      elsif (TO_X01(WW2_delayed)='0' and TO_X01(WW1_delayed)='1' and TO_X01(WW0_delayed)='0') then
        WWIDTH := 4;
      elsif (TO_X01(WW2_delayed)='0' and TO_X01(WW1_delayed)='1' and TO_X01(WW0_delayed)='1') then
        WWIDTH := 9;
      elsif (TO_X01(WW2_delayed)='1' and TO_X01(WW1_delayed)='0' and TO_X01(WW0_delayed)='0') then
        WWIDTH := 18;
      elsif (TO_X01(WW2_delayed)='1' and TO_X01(WW1_delayed)='0' and TO_X01(WW0_delayed)='1') then
        WWIDTH := 36;
      else
	assert false
	report ": WW value invalid"
	severity Warning;
      end if;


      if (TO_X01(WCLK_ipd)='X') then
	if (TO_X01(WEN_delayed) /= '0') then
          if (TO_X01(WCLK_previous) /= 'X') then
	    assert false
	    report ": WCLK went unknown"
	    severity Warning;
	  end if;
	end if;
      elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='1')) then
	case (TO_X01(WEN_delayed)) is
	  when '0' =>
	    null;
	  when '1' =>

            -- Convert Write Address Signal to Integer
            if( INT(WRAD15_delayed) = -65537 ) then
              WADDR := -1;
            elsif( INT(WRAD14_delayed) = -65537 ) then
              WADDR := -1;
            else
              WADDR := ((INT(WRAD15_delayed)*32768)
                        +(INT(WRAD14_delayed)*16384)+(INT(WRAD13_delayed)*8192)+(INT(WRAD12_delayed)*4096)
                        +(INT(WRAD11_delayed)*2048)+(INT(WRAD10_delayed)*1024)+(INT(WRAD9_delayed)*512)
                        +(INT(WRAD8_delayed)*256)+(INT(WRAD7_delayed)*128)+(INT(WRAD6_delayed)*64)
                        +(INT(WRAD5_delayed)*32)+(INT(WRAD4_delayed)*16)+(INT(WRAD3_delayed)*8)
                        +(INT(WRAD2_delayed)*4)+(INT(WRAD1_delayed)*2)+(INT(WRAD0_delayed)));
            end if;

	    if (WADDR < 0) then
              if (TO_X01(WRAD15_delayed) = 'X' and WWIDTH = 1) then
                assert false
                report ": WRAD15 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD14_delayed) = 'X' and WWIDTH = 1) then
                assert false
                report ": WRAD14 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD13_delayed) = 'X' and WWIDTH = 1) then
                assert false
                report ": WRAD13 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD12_delayed) = 'X' and WWIDTH = 1) then
                assert false
                report ": WRAD12 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD11_delayed) = 'X' and WWIDTH = 1) then
                assert false
                report ": WRAD11 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD10_delayed) = 'X' and WWIDTH <= 2) then
                assert false
                report ": WRAD10 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD9_delayed) = 'X' and WWIDTH <= 4) then
                assert false
                report ": WRAD9 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD8_delayed) = 'X' and WWIDTH <= 9) then
                assert false
                report ": WRAD8 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD7_delayed) = 'X' and WWIDTH <= 18) then
                assert false
                report ": WRAD7 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD6_delayed) = 'X') then
                assert false
                report ": WRAD6 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD5_delayed) = 'X') then
                assert false
                report ": WRAD5 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD4_delayed) = 'X') then
                assert false
                report ": WRAD4 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD3_delayed) = 'X') then
                assert false
                report ": WRAD3 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD2_delayed) = 'X') then
                assert false
                report ": WRAD2 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD1_delayed) = 'X') then
                assert false
                report ": WRAD1 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD0_delayed) = 'X') then
                assert false
                report ": WRAD0 went unknown"
                severity Warning;
              end if;
	    else 
              case WWIDTH is
                when 1 => RAM_TMP(WADDR) := WD0_delayed ;
                when 2 => RAM_TMP(2*WADDR + 0) := WD0_delayed ;
                          RAM_TMP(2*WADDR + 1) := WD1_delayed ;
                when 4 => RAM_TMP(4*WADDR + 0) := WD0_delayed ;
                          RAM_TMP(4*WADDR + 1) := WD1_delayed ;
                          RAM_TMP(4*WADDR + 2) := WD2_delayed ;
                          RAM_TMP(4*WADDR + 3) := WD3_delayed ;
                when 9 => RAM_TMP(8*WADDR + 0) := WD0_delayed ;
                          RAM_TMP(8*WADDR + 1) := WD1_delayed ;
                          RAM_TMP(8*WADDR + 2) := WD2_delayed ;
                          RAM_TMP(8*WADDR + 3) := WD3_delayed ;
                          RAM_TMP(8*WADDR + 4) := WD4_delayed ;
                          RAM_TMP(8*WADDR + 5) := WD5_delayed ;
                          RAM_TMP(8*WADDR + 6) := WD6_delayed ;
                          RAM_TMP(8*WADDR + 7) := WD7_delayed ;
                          RAM_TMP9(WADDR) := WD8_delayed ;
                when 18 => RAM_TMP(16*WADDR + 0) := WD0_delayed ;
                           RAM_TMP(16*WADDR + 1) := WD1_delayed ;
                           RAM_TMP(16*WADDR + 2) := WD2_delayed ;
                           RAM_TMP(16*WADDR + 3) := WD3_delayed ;
                           RAM_TMP(16*WADDR + 4) := WD4_delayed ;
                           RAM_TMP(16*WADDR + 5) := WD5_delayed ;
                           RAM_TMP(16*WADDR + 6) := WD6_delayed ;
                           RAM_TMP(16*WADDR + 7) := WD7_delayed ;
                           RAM_TMP9((2*WADDR) + 0) := WD8_delayed ;
                           RAM_TMP(16*WADDR + 8) := WD9_delayed ;
                           RAM_TMP(16*WADDR + 9) := WD10_delayed ;
                           RAM_TMP(16*WADDR + 10) := WD11_delayed ;
                           RAM_TMP(16*WADDR + 11) := WD12_delayed ;
                           RAM_TMP(16*WADDR + 12) := WD13_delayed ;
                           RAM_TMP(16*WADDR + 13) := WD14_delayed ;
                           RAM_TMP(16*WADDR + 14) := WD15_delayed ;
                           RAM_TMP(16*WADDR + 15) := WD16_delayed ;
                           RAM_TMP9((2*WADDR) + 1) := WD17_delayed ;
                when 36 => RAM_TMP(32*WADDR + 0) := WD0_delayed ;
                           RAM_TMP(32*WADDR + 1) := WD1_delayed ;
                           RAM_TMP(32*WADDR + 2) := WD2_delayed ;
                           RAM_TMP(32*WADDR + 3) := WD3_delayed ;
                           RAM_TMP(32*WADDR + 4) := WD4_delayed ;
                           RAM_TMP(32*WADDR + 5) := WD5_delayed ;
                           RAM_TMP(32*WADDR + 6) := WD6_delayed ;
                           RAM_TMP(32*WADDR + 7) := WD7_delayed ;
                           RAM_TMP9((4*WADDR) + 0) := WD8_delayed ;
                           RAM_TMP(32*WADDR + 8) := WD9_delayed ;
                           RAM_TMP(32*WADDR + 9) := WD10_delayed ;
                           RAM_TMP(32*WADDR + 10) := WD11_delayed ;
                           RAM_TMP(32*WADDR + 11) := WD12_delayed ;
                           RAM_TMP(32*WADDR + 12) := WD13_delayed ;
                           RAM_TMP(32*WADDR + 13) := WD14_delayed ;
                           RAM_TMP(32*WADDR + 14) := WD15_delayed ;
                           RAM_TMP(32*WADDR + 15) := WD16_delayed ;
                           RAM_TMP9((4*WADDR) + 1) := WD17_delayed ;
                           RAM_TMP(32*WADDR + 16) := WD18_delayed ;
                           RAM_TMP(32*WADDR + 17) := WD19_delayed ;
                           RAM_TMP(32*WADDR + 18) := WD20_delayed ;
                           RAM_TMP(32*WADDR + 19) := WD21_delayed ;
                           RAM_TMP(32*WADDR + 20) := WD22_delayed ;
                           RAM_TMP(32*WADDR + 21) := WD23_delayed ;
                           RAM_TMP(32*WADDR + 22) := WD24_delayed ;
                           RAM_TMP(32*WADDR + 23) := WD25_delayed ;
                           RAM_TMP9((4*WADDR) + 2) := WD26_delayed ;
                           RAM_TMP(32*WADDR + 24) := WD27_delayed ;
                           RAM_TMP(32*WADDR + 25) := WD28_delayed ;
                           RAM_TMP(32*WADDR + 26) := WD29_delayed ;
                           RAM_TMP(32*WADDR + 27) := WD30_delayed ;
                           RAM_TMP(32*WADDR + 28) := WD31_delayed ;
                           RAM_TMP(32*WADDR + 29) := WD32_delayed ;
                           RAM_TMP(32*WADDR + 30) := WD33_delayed ;
                           RAM_TMP(32*WADDR + 31) := WD34_delayed ;
                           RAM_TMP9((4*WADDR) + 3) := WD35_delayed ;
                when others => 
	          assert false
	          report ": WWIDTH value invalid"
	          severity Warning;
              end case;
	    end if;
	  when others =>
            assert false
            report ": WEN went unknown"
            severity Warning;
	end case;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      -- Decode Read Word Width
      if (TO_X01(RW2_delayed)='0' and TO_X01(RW1_delayed)='0' and TO_X01(RW0_delayed)='0') then
        RWIDTH := 1;
      elsif (TO_X01(RW2_delayed)='0' and TO_X01(RW1_delayed)='0' and TO_X01(RW0_delayed)='1') then
        RWIDTH := 2;
      elsif (TO_X01(RW2_delayed)='0' and TO_X01(RW1_delayed)='1' and TO_X01(RW0_delayed)='0') then
        RWIDTH := 4;
      elsif (TO_X01(RW2_delayed)='0' and TO_X01(RW1_delayed)='1' and TO_X01(RW0_delayed)='1') then
        RWIDTH := 9;
      elsif (TO_X01(RW2_delayed)='1' and TO_X01(RW1_delayed)='0' and TO_X01(RW0_delayed)='0') then
        RWIDTH := 18;
      elsif (TO_X01(RW2_delayed)='1' and TO_X01(RW1_delayed)='0' and TO_X01(RW0_delayed)='1') then
        RWIDTH := 36;
      else
        assert false
        report ": RW value invalid"
        severity Warning;
      end if;

      -- Convert Read Address Signal to Integer
      if (INT(RDAD15_delayed) = -65537) then
        RADDR := -1;
      elsif (INT(RDAD14_delayed) = -65537) then
        RADDR := -1;
      else
        RADDR := ((INT(RDAD15_delayed)*32768)
                 +(INT(RDAD14_delayed)*16384)+(INT(RDAD13_delayed)*8192)+(INT(RDAD12_delayed)*4096)
                 +(INT(RDAD11_delayed)*2048)+(INT(RDAD10_delayed)*1024)+(INT(RDAD9_delayed)*512)
                 +(INT(RDAD8_delayed)*256)+(INT(RDAD7_delayed)*128)+(INT(RDAD6_delayed)*64)
                 +(INT(RDAD5_delayed)*32)+(INT(RDAD4_delayed)*16)+(INT(RDAD3_delayed)*8)
                 +(INT(RDAD2_delayed)*4)+(INT(RDAD1_delayed)*2)+(INT(RDAD0_delayed)));
      end if;
      if (TO_X01(RCLK_ipd) = 'X') then
	case RWIDTH is
          when 1 => RD0_zd := 'X';
          when 2 => RD0_zd := 'X';
                    RD1_zd := 'X';
          when 4 => RD0_zd := 'X';
                    RD1_zd := 'X';
                    RD2_zd := 'X';
                    RD3_zd := 'X';
          when 9 => RD0_zd := 'X';
                    RD1_zd := 'X';
                    RD2_zd := 'X';
                    RD3_zd := 'X';
                    RD4_zd := 'X';
                    RD5_zd := 'X';
                    RD6_zd := 'X';
                    RD7_zd := 'X';
                    RD8_zd := 'X';
          when 18 => RD0_zd := 'X';
                     RD1_zd := 'X';
                     RD2_zd := 'X';
                     RD3_zd := 'X';
                     RD4_zd := 'X';
                     RD5_zd := 'X';
                     RD6_zd := 'X';
                     RD7_zd := 'X';
                     RD8_zd := 'X';
                     RD9_zd := 'X';
                     RD10_zd := 'X';
                     RD11_zd := 'X';
                     RD12_zd := 'X';
                     RD13_zd := 'X';
                     RD14_zd := 'X';
                     RD15_zd := 'X';
                     RD16_zd := 'X';
                     RD17_zd := 'X';
          when 36 => RD0_zd := 'X';
                     RD1_zd := 'X';
                     RD2_zd := 'X';
                     RD3_zd := 'X';
                     RD4_zd := 'X';
                     RD5_zd := 'X';
                     RD6_zd := 'X';
                     RD7_zd := 'X';
                     RD8_zd := 'X';
                     RD9_zd := 'X';
                     RD10_zd := 'X';
                     RD11_zd := 'X';
                     RD12_zd := 'X';
                     RD13_zd := 'X';
                     RD14_zd := 'X';
                     RD15_zd := 'X';
                     RD16_zd := 'X';
                     RD17_zd := 'X';
                     RD18_zd := 'X';
                     RD19_zd := 'X';
                     RD20_zd := 'X';
                     RD21_zd := 'X';
                     RD22_zd := 'X';
                     RD23_zd := 'X';
                     RD24_zd := 'X';
                     RD25_zd := 'X';
                     RD26_zd := 'X';
                     RD27_zd := 'X';
                     RD28_zd := 'X';
                     RD29_zd := 'X';
                     RD30_zd := 'X';
                     RD31_zd := 'X';
                     RD32_zd := 'X';
                     RD33_zd := 'X';
                     RD34_zd := 'X';
                     RD35_zd := 'X';
          when others => 
            assert false
            report ": RWIDTH value invalid"
            severity Warning;
        end case;
	if (TO_X01(RCLK_previous) /= 'X') then
	  assert false
	  report ": RCLK went unknown"
	  severity Warning;
	end if;
      elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '1')) then
	case (TO_X01(REN_delayed)) is
          when '0' =>
                    assert true
                    report ": REN low - hold old output"
                    severity Note;
	  when '1' =>
	    if (RADDR < 0) then -- address invalid
              case RWIDTH is
                when 1 => RD0_zd := 'X';
                when 2 => RD0_zd := 'X';
                          RD1_zd := 'X';
                when 4 => RD0_zd := 'X';
                          RD1_zd := 'X';
                          RD2_zd := 'X';
                          RD3_zd := 'X';
                when 9 => RD0_zd := 'X';
                          RD1_zd := 'X';
                          RD2_zd := 'X';
                          RD3_zd := 'X';
                          RD4_zd := 'X';
                          RD5_zd := 'X';
                          RD6_zd := 'X';
                          RD7_zd := 'X';
                          RD8_zd := 'X';
                when 18 => RD0_zd := 'X';
                           RD1_zd := 'X';
                           RD2_zd := 'X';
                           RD3_zd := 'X';
                           RD4_zd := 'X';
                           RD5_zd := 'X';
                           RD6_zd := 'X';
                           RD7_zd := 'X';
                           RD8_zd := 'X';
                           RD9_zd := 'X';
                           RD10_zd := 'X';
                           RD11_zd := 'X';
                           RD12_zd := 'X';
                           RD13_zd := 'X';
                           RD14_zd := 'X';
                           RD15_zd := 'X';
                           RD16_zd := 'X';
                           RD17_zd := 'X';
                when 36 => RD0_zd := 'X';
                           RD1_zd := 'X';
                           RD2_zd := 'X';
                           RD3_zd := 'X';
                           RD4_zd := 'X';
                           RD5_zd := 'X';
                           RD6_zd := 'X';
                           RD7_zd := 'X';
                           RD8_zd := 'X';
                           RD9_zd := 'X';
                           RD10_zd := 'X';
                           RD11_zd := 'X';
                           RD12_zd := 'X';
                           RD13_zd := 'X';
                           RD14_zd := 'X';
                           RD15_zd := 'X';
                           RD16_zd := 'X';
                           RD17_zd := 'X';
                           RD18_zd := 'X';
                           RD19_zd := 'X';
                           RD20_zd := 'X';
                           RD21_zd := 'X';
                           RD22_zd := 'X';
                           RD23_zd := 'X';
                           RD24_zd := 'X';
                           RD25_zd := 'X';
                           RD26_zd := 'X';
                           RD27_zd := 'X';
                           RD28_zd := 'X';
                           RD29_zd := 'X';
                           RD30_zd := 'X';
                           RD31_zd := 'X';
                           RD32_zd := 'X';
                           RD33_zd := 'X';
                           RD34_zd := 'X';
                           RD35_zd := 'X';
                when others => 
	          assert false
	          report ": RWIDTH value invalid"
	          severity Warning;
              end case;
	      if (TO_X01(RDAD15_delayed) = 'X') and (TO_X01(RDAD15_previous) /= 'X' and RWIDTH = 1) then
		assert false
		report ": RDAD15 went unknown"
		severity Warning;
                RDAD15_previous := RDAD15_delayed;
	      end if;
	      if (TO_X01(RDAD14_delayed) = 'X') and (TO_X01(RDAD14_previous) /= 'X' and RWIDTH = 1) then
		assert false
		report ": RDAD14 went unknown"
		severity Warning;
                RDAD14_previous := RDAD14_delayed;
	      end if;
	      if (TO_X01(RDAD13_delayed) = 'X') and (TO_X01(RDAD13_previous) /= 'X' and RWIDTH = 1) then
		assert false
		report ": RDAD13 went unknown"
		severity Warning;
                RDAD13_previous := RDAD13_delayed;
	      end if;
	      if (TO_X01(RDAD12_delayed) = 'X') and (TO_X01(RDAD12_previous) /= 'X' and RWIDTH = 1) then
		assert false
		report ": RDAD12 went unknown"
		severity Warning;
                RDAD12_previous := RDAD12_delayed;
	      end if;
	      if (TO_X01(RDAD11_delayed) = 'X') and (TO_X01(RDAD11_previous) /= 'X' and RWIDTH = 1) then
		assert false
		report ": RDAD11 went unknown"
		severity Warning;
                RDAD11_previous := RDAD11_delayed;
	      end if;
	      if (TO_X01(RDAD10_delayed) = 'X') and (TO_X01(RDAD10_previous) /= 'X' and RWIDTH <= 2) then
		assert false
		report ": RDAD10 went unknown"
		severity Warning;
                RDAD10_previous := RDAD10_delayed;
	      end if;
	      if (TO_X01(RDAD9_delayed) = 'X') and (TO_X01(RDAD9_previous) /= 'X' and RWIDTH <= 4) then
		assert false
		report ": RDAD9 went unknown"
		severity Warning;
                RDAD9_previous := RDAD9_delayed;
	      end if;
	      if (TO_X01(RDAD8_delayed) = 'X') and (TO_X01(RDAD8_previous) /= 'X' and RWIDTH <= 9) then
		assert false
		report ": RDAD8 went unknown"
		severity Warning;
                RDAD8_previous := RDAD8_delayed;
	      end if;
	      if (TO_X01(RDAD7_delayed) = 'X') and (TO_X01(RDAD7_previous) /= 'X' and RWIDTH <= 18) then
		assert false
		report ": RDAD7 went unknown"
		severity Warning;
                RDAD7_previous := RDAD7_delayed;
	      end if;
	      if (TO_X01(RDAD6_delayed) = 'X') and (TO_X01(RDAD6_previous) /= 'X') then
		assert false
		report ": RDAD6 went unknown"
		severity Warning;
                RDAD6_previous := RDAD6_delayed;
	      end if;
	      if (TO_X01(RDAD5_delayed) = 'X') and (TO_X01(RDAD5_previous) /= 'X') then
		assert false
		report ": RDAD5 went unknown"
		severity Warning;
                RDAD5_previous := RDAD5_delayed;
	      end if;
	      if (TO_X01(RDAD4_delayed) = 'X') and (TO_X01(RDAD4_previous) /= 'X') then
		assert false
		report ": RDAD4 went unknown"
		severity Warning;
                RDAD4_previous := RDAD4_delayed;
	      end if;
	      if (TO_X01(RDAD3_delayed) = 'X') and (TO_X01(RDAD3_previous) /= 'X') then
		assert false
		report ": RDAD3 went unknown"
		severity Warning;
                RDAD3_previous := RDAD3_delayed;
	      end if;
	      if (TO_X01(RDAD2_delayed) = 'X') and (TO_X01(RDAD2_previous) /= 'X') then
		assert false
		report ": RDAD2 went unknown"
		severity Warning;
                RDAD2_previous := RDAD2_delayed;
	      end if;
	      if (TO_X01(RDAD1_delayed) = 'X') and (TO_X01(RDAD1_previous) /= 'X') then
		assert false
		report ": RDAD1 went unknown"
		severity Warning;
                RDAD1_previous := RDAD1_delayed;
	      end if;
	      if (TO_X01(RDAD0_delayed) = 'X') and (TO_X01(RDAD0_previous) /= 'X') then
		assert false
		report ": RDAD0 went unknown"
		severity Warning;
                RDAD0_previous := RDAD0_delayed;
	      end if;
	    else -- address OK
              case RWIDTH is
                when 1 => RD0_zd := RAM_TMP(RADDR) ;
                when 2 => RD0_zd := RAM_TMP(2*RADDR + 0) ;
                          RD1_zd := RAM_TMP(2*RADDR + 1) ;
                when 4 => RD0_zd := RAM_TMP(4*RADDR + 0) ;
                          RD1_zd := RAM_TMP(4*RADDR + 1) ;
                          RD2_zd := RAM_TMP(4*RADDR + 2) ;
                          RD3_zd := RAM_TMP(4*RADDR + 3) ;
                when 9 => RD0_zd := RAM_TMP(8*RADDR + 0) ;
                          RD1_zd := RAM_TMP(8*RADDR + 1) ;
                          RD2_zd := RAM_TMP(8*RADDR + 2) ;
                          RD3_zd := RAM_TMP(8*RADDR + 3) ;
                          RD4_zd := RAM_TMP(8*RADDR + 4) ;
                          RD5_zd := RAM_TMP(8*RADDR + 5) ;
                          RD6_zd := RAM_TMP(8*RADDR + 6) ;
                          RD7_zd := RAM_TMP(8*RADDR + 7) ;
                          RD8_zd := RAM_TMP9(RADDR) ;
                when 18 => RD0_zd := RAM_TMP(16*RADDR + 0) ;
                           RD1_zd := RAM_TMP(16*RADDR + 1) ;
                           RD2_zd := RAM_TMP(16*RADDR + 2) ;
                           RD3_zd := RAM_TMP(16*RADDR + 3) ;
                           RD4_zd := RAM_TMP(16*RADDR + 4) ;
                           RD5_zd := RAM_TMP(16*RADDR + 5) ;
                           RD6_zd := RAM_TMP(16*RADDR + 6) ;
                           RD7_zd := RAM_TMP(16*RADDR + 7) ;
                           RD8_zd := RAM_TMP9((2*RADDR) + 0) ;
                           RD9_zd := RAM_TMP(16*RADDR + 8) ;
                           RD10_zd := RAM_TMP(16*RADDR + 9) ;
                           RD11_zd := RAM_TMP(16*RADDR + 10) ;
                           RD12_zd := RAM_TMP(16*RADDR + 11) ;
                           RD13_zd := RAM_TMP(16*RADDR + 12) ;
                           RD14_zd := RAM_TMP(16*RADDR + 13) ;
                           RD15_zd := RAM_TMP(16*RADDR + 14) ;
                           RD16_zd := RAM_TMP(16*RADDR + 15) ;
                           RD17_zd := RAM_TMP9((2*RADDR) + 1) ;
                when 36 => RD0_zd := RAM_TMP(32*RADDR + 0) ;
                           RD1_zd := RAM_TMP(32*RADDR + 1) ;
                           RD2_zd := RAM_TMP(32*RADDR + 2) ;
                           RD3_zd := RAM_TMP(32*RADDR + 3) ;
                           RD4_zd := RAM_TMP(32*RADDR + 4) ;
                           RD5_zd := RAM_TMP(32*RADDR + 5) ;
                           RD6_zd := RAM_TMP(32*RADDR + 6) ;
                           RD7_zd := RAM_TMP(32*RADDR + 7) ;
                           RD8_zd := RAM_TMP9((4*RADDR) + 0) ;
                           RD9_zd := RAM_TMP(32*RADDR + 8) ;
                           RD10_zd := RAM_TMP(32*RADDR + 9) ;
                           RD11_zd := RAM_TMP(32*RADDR + 10) ;
                           RD12_zd := RAM_TMP(32*RADDR + 11) ;
                           RD13_zd := RAM_TMP(32*RADDR + 12) ;
                           RD14_zd := RAM_TMP(32*RADDR + 13) ;
                           RD15_zd := RAM_TMP(32*RADDR + 14) ;
                           RD16_zd := RAM_TMP(32*RADDR + 15) ;
                           RD17_zd := RAM_TMP9((4*RADDR) + 1) ;
                           RD18_zd := RAM_TMP(32*RADDR + 16) ;
                           RD19_zd := RAM_TMP(32*RADDR + 17) ;
                           RD20_zd := RAM_TMP(32*RADDR + 18) ;
                           RD21_zd := RAM_TMP(32*RADDR + 19) ;
                           RD22_zd := RAM_TMP(32*RADDR + 20) ;
                           RD23_zd := RAM_TMP(32*RADDR + 21) ;
                           RD24_zd := RAM_TMP(32*RADDR + 22) ;
                           RD25_zd := RAM_TMP(32*RADDR + 23) ;
                           RD26_zd := RAM_TMP9((4*RADDR) + 2) ;
                           RD27_zd := RAM_TMP(32*RADDR + 24) ;
                           RD28_zd := RAM_TMP(32*RADDR + 25) ;
                           RD29_zd := RAM_TMP(32*RADDR + 26) ;
                           RD30_zd := RAM_TMP(32*RADDR + 27) ;
                           RD31_zd := RAM_TMP(32*RADDR + 28) ;
                           RD32_zd := RAM_TMP(32*RADDR + 29) ;
                           RD33_zd := RAM_TMP(32*RADDR + 30) ;
                           RD34_zd := RAM_TMP(32*RADDR + 31) ;
                           RD35_zd := RAM_TMP9((4*RADDR ) + 3) ;
                when others => 
	          assert false
	          report ": RWIDTH value invalid"
	          severity Warning;
              end case;
	    end if;
	  when others =>
            case RWIDTH is
              when 1 => RD0_zd := 'X';
              when 2 => RD0_zd := 'X';
                        RD1_zd := 'X';
              when 4 => RD0_zd := 'X';
                        RD1_zd := 'X';
                        RD2_zd := 'X';
                        RD3_zd := 'X';
              when 9 => RD0_zd := 'X';
                        RD1_zd := 'X';
                        RD2_zd := 'X';
                        RD3_zd := 'X';
                        RD4_zd := 'X';
                        RD5_zd := 'X';
                        RD6_zd := 'X';
                        RD7_zd := 'X';
                        RD8_zd := 'X';
              when 18 => RD0_zd := 'X';
                         RD1_zd := 'X';
                         RD2_zd := 'X';
                         RD3_zd := 'X';
                         RD4_zd := 'X';
                         RD5_zd := 'X';
                         RD6_zd := 'X';
                         RD7_zd := 'X';
                         RD8_zd := 'X';
                         RD9_zd := 'X';
                         RD10_zd := 'X';
                         RD11_zd := 'X';
                         RD12_zd := 'X';
                         RD13_zd := 'X';
                         RD14_zd := 'X';
                         RD15_zd := 'X';
                         RD16_zd := 'X';
                         RD17_zd := 'X';
              when 36 => RD0_zd := 'X';
                         RD1_zd := 'X';
                         RD2_zd := 'X';
                         RD3_zd := 'X';
                         RD4_zd := 'X';
                         RD5_zd := 'X';
                         RD6_zd := 'X';
                         RD7_zd := 'X';
                         RD8_zd := 'X';
                         RD9_zd := 'X';
                         RD10_zd := 'X';
                         RD11_zd := 'X';
                         RD12_zd := 'X';
                         RD13_zd := 'X';
                         RD14_zd := 'X';
                         RD15_zd := 'X';
                         RD16_zd := 'X';
                         RD17_zd := 'X';
                         RD18_zd := 'X';
                         RD19_zd := 'X';
                         RD20_zd := 'X';
                         RD21_zd := 'X';
                         RD22_zd := 'X';
                         RD23_zd := 'X';
                         RD24_zd := 'X';
                         RD25_zd := 'X';
                         RD26_zd := 'X';
                         RD27_zd := 'X';
                         RD28_zd := 'X';
                         RD29_zd := 'X';
                         RD30_zd := 'X';
                         RD31_zd := 'X';
                         RD32_zd := 'X';
                         RD33_zd := 'X';
                         RD34_zd := 'X';
                         RD35_zd := 'X';
              when others => 
	        assert false
	        report ": RWIDTH value invalid"
	        severity Warning;
            end case; -- RWIDTH
            if (TO_X01(REN_delayed) = 'X') and (TO_X01(REN_previous) /= 'X') then
	      assert false
	      report ": REN went unknown"
	      severity Warning;
              REN_previous := REN_delayed;
            end if;
	end case; -- REN
      end if; -- Rising RCLK edge

      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      WW2_delayed := WW2_ipd;
      WW1_delayed := WW1_ipd;
      WW0_delayed := WW0_ipd;
      WEN_delayed := WEN_ipd;
      if RW2_ipd'event then
        RW2_previous := RW2_delayed;
        RW2_delayed := RW2_ipd;
      end if;
      if RW1_ipd'event then
        RW1_previous := RW1_delayed;
        RW1_delayed := RW1_ipd;
      end if;
      if RW0_ipd'event then
        RW0_previous := RW0_delayed;
        RW0_delayed := RW0_ipd;
      end if;
      if REN_ipd'event then
        REN_previous := REN_delayed;
        REN_delayed := REN_ipd;
      end if;
      WD35_delayed := WD35_ipd;
      WD34_delayed := WD34_ipd;
      WD33_delayed := WD33_ipd;
      WD32_delayed := WD32_ipd;
      WD31_delayed := WD31_ipd;
      WD30_delayed := WD30_ipd;
      WD29_delayed := WD29_ipd;
      WD28_delayed := WD28_ipd;
      WD27_delayed := WD27_ipd;
      WD26_delayed := WD26_ipd;
      WD25_delayed := WD25_ipd;
      WD24_delayed := WD24_ipd;
      WD23_delayed := WD23_ipd;
      WD22_delayed := WD22_ipd;
      WD21_delayed := WD21_ipd;
      WD20_delayed := WD20_ipd;
      WD19_delayed := WD19_ipd;
      WD18_delayed := WD18_ipd;
      WD17_delayed := WD17_ipd;
      WD16_delayed := WD16_ipd;
      WD15_delayed := WD15_ipd;
      WD14_delayed := WD14_ipd;
      WD13_delayed := WD13_ipd;
      WD12_delayed := WD12_ipd;
      WD11_delayed := WD11_ipd;
      WD10_delayed := WD10_ipd;
      WD9_delayed := WD9_ipd;
      WD8_delayed := WD8_ipd;
      WD7_delayed := WD7_ipd;
      WD6_delayed := WD6_ipd;
      WD5_delayed := WD5_ipd;
      WD4_delayed := WD4_ipd;
      WD3_delayed := WD3_ipd;
      WD2_delayed := WD2_ipd;
      WD1_delayed := WD1_ipd;
      WD0_delayed := WD0_ipd;
      WRAD15_delayed := WRAD15_ipd;
      WRAD14_delayed := WRAD14_ipd;
      WRAD13_delayed := WRAD13_ipd;
      WRAD12_delayed := WRAD12_ipd;
      WRAD11_delayed := WRAD11_ipd;
      WRAD10_delayed := WRAD10_ipd;
      WRAD9_delayed := WRAD9_ipd;
      WRAD8_delayed := WRAD8_ipd;
      WRAD7_delayed := WRAD7_ipd;
      WRAD6_delayed := WRAD6_ipd;
      WRAD5_delayed := WRAD5_ipd;
      WRAD4_delayed := WRAD4_ipd;
      WRAD3_delayed := WRAD3_ipd;
      WRAD2_delayed := WRAD2_ipd;
      WRAD1_delayed := WRAD1_ipd;
      WRAD0_delayed := WRAD0_ipd;
      if RDAD15_ipd'event then
        RDAD15_previous := RDAD15_delayed;
        RDAD15_delayed := RDAD15_ipd;
      end if;
      if RDAD14_ipd'event then
        RDAD14_previous := RDAD14_delayed;
        RDAD14_delayed := RDAD14_ipd;
      end if;
      if RDAD13_ipd'event then
        RDAD13_previous := RDAD13_delayed;
        RDAD13_delayed := RDAD13_ipd;
      end if;
      if RDAD12_ipd'event then
        RDAD12_previous := RDAD12_delayed;
        RDAD12_delayed := RDAD12_ipd;
      end if;
      if RDAD11_ipd'event then
        RDAD11_previous := RDAD11_delayed;
        RDAD11_delayed := RDAD11_ipd;
      end if;
      if RDAD10_ipd'event then
        RDAD10_previous := RDAD10_delayed;
        RDAD10_delayed := RDAD10_ipd;
      end if;
      if RDAD9_ipd'event then
        RDAD9_previous := RDAD9_delayed;
        RDAD9_delayed := RDAD9_ipd;
      end if;
      if RDAD8_ipd'event then
        RDAD8_previous := RDAD8_delayed;
        RDAD8_delayed := RDAD8_ipd;
      end if;
      if RDAD7_ipd'event then
        RDAD7_previous := RDAD7_delayed;
        RDAD7_delayed := RDAD7_ipd;
      end if;
      if RDAD6_ipd'event then
        RDAD6_previous := RDAD6_delayed;
        RDAD6_delayed := RDAD6_ipd;
      end if;
      if RDAD5_ipd'event then
        RDAD5_previous := RDAD5_delayed;
        RDAD5_delayed := RDAD5_ipd;
      end if;
      if RDAD4_ipd'event then
        RDAD4_previous := RDAD4_delayed;
        RDAD4_delayed := RDAD4_ipd;
      end if;
      if RDAD3_ipd'event then
        RDAD3_previous := RDAD3_delayed;
        RDAD3_delayed := RDAD3_ipd;
      end if;
      if RDAD2_ipd'event then
        RDAD2_previous := RDAD2_delayed;
        RDAD2_delayed := RDAD2_ipd;
      end if;
      if RDAD1_ipd'event then
        RDAD1_previous := RDAD1_delayed;
      end if;
        RDAD1_delayed := RDAD1_ipd;
      if RDAD0_ipd'event then
        RDAD0_previous := RDAD0_delayed;
        RDAD0_delayed := RDAD0_ipd;
      end if;


    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => RD35,
	GlitchData => RD35_GlitchData,
	OutSignalName => "RD35",
	OutTemp => RD35_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD35), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => Xon,
	MsgOn => MsgOn,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
        OutSignal => RD34,
        GlitchData => RD34_GlitchData,
        OutSignalName => "RD34",
        OutTemp => RD34_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD34), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD33,
        GlitchData => RD33_GlitchData,
        OutSignalName => "RD33",
        OutTemp => RD33_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD33), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD32,
        GlitchData => RD32_GlitchData,
        OutSignalName => "RD32",
        OutTemp => RD32_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD32), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD31,
        GlitchData => RD31_GlitchData,
        OutSignalName => "RD31",
        OutTemp => RD31_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD31), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD30,
        GlitchData => RD30_GlitchData,
        OutSignalName => "RD30",
        OutTemp => RD30_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD30), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD29,
        GlitchData => RD29_GlitchData,
        OutSignalName => "RD29",
        OutTemp => RD29_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD29), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD28,
        GlitchData => RD28_GlitchData,
        OutSignalName => "RD28",
        OutTemp => RD28_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD28), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD27,
        GlitchData => RD27_GlitchData,
        OutSignalName => "RD27",
        OutTemp => RD27_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD27), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD26,
        GlitchData => RD26_GlitchData,
        OutSignalName => "RD26",
        OutTemp => RD26_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD26), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD25,
        GlitchData => RD25_GlitchData,
        OutSignalName => "RD25",
        OutTemp => RD25_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD25), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD24,
        GlitchData => RD24_GlitchData,
        OutSignalName => "RD24",
        OutTemp => RD24_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD24), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD23,
        GlitchData => RD23_GlitchData,
        OutSignalName => "RD23",
        OutTemp => RD23_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD23), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD22,
        GlitchData => RD22_GlitchData,
        OutSignalName => "RD22",
        OutTemp => RD22_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD22), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD21,
        GlitchData => RD21_GlitchData,
        OutSignalName => "RD21",
        OutTemp => RD21_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD21), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD20,
        GlitchData => RD20_GlitchData,
        OutSignalName => "RD20",
        OutTemp => RD20_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD20), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD19,
        GlitchData => RD19_GlitchData,
        OutSignalName => "RD19",
        OutTemp => RD19_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD19), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD18,
        GlitchData => RD18_GlitchData,
        OutSignalName => "RD18",
        OutTemp => RD18_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD18), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD17,
        GlitchData => RD17_GlitchData,
        OutSignalName => "RD17",
        OutTemp => RD17_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD17), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD16,
        GlitchData => RD16_GlitchData,
        OutSignalName => "RD16",
        OutTemp => RD16_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD16), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD15,
        GlitchData => RD15_GlitchData,
        OutSignalName => "RD15",
        OutTemp => RD15_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD15), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD14,
        GlitchData => RD14_GlitchData,
        OutSignalName => "RD14",
        OutTemp => RD14_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD14), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD13,
        GlitchData => RD13_GlitchData,
        OutSignalName => "RD13",
        OutTemp => RD13_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD13), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD12,
        GlitchData => RD12_GlitchData,
        OutSignalName => "RD12",
        OutTemp => RD12_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD12), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD11,
        GlitchData => RD11_GlitchData,
        OutSignalName => "RD11",
        OutTemp => RD11_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD11), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD10,
        GlitchData => RD10_GlitchData,
        OutSignalName => "RD10",
        OutTemp => RD10_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD10), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD9,
        GlitchData => RD9_GlitchData,
        OutSignalName => "RD9",
        OutTemp => RD9_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD9), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD8,
        GlitchData => RD8_GlitchData,
        OutSignalName => "RD8",
        OutTemp => RD8_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD8), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD7,
        GlitchData => RD7_GlitchData,
        OutSignalName => "RD7",
        OutTemp => RD7_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD7), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD6,
        GlitchData => RD6_GlitchData,
        OutSignalName => "RD6",
        OutTemp => RD6_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD6), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD5,
        GlitchData => RD5_GlitchData,
        OutSignalName => "RD5",
        OutTemp => RD5_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD5), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD4,
        GlitchData => RD4_GlitchData,
        OutSignalName => "RD4",
        OutTemp => RD4_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD4), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD3,
        GlitchData => RD3_GlitchData,
        OutSignalName => "RD3",
        OutTemp => RD3_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD3), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD2,
        GlitchData => RD2_GlitchData,
        OutSignalName => "RD2",
        OutTemp => RD2_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD2), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD1,
        GlitchData => RD1_GlitchData,
        OutSignalName => "RD1",
        OutTemp => RD1_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD1), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD0,
        GlitchData => RD0_GlitchData,
        OutSignalName => "RD0",
        OutTemp => RD0_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD0), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );
    
  end process VITALBehavior;

end VITAL_ACT;

configuration CFG_RAM64K36_VITAL of RAM64K36 is
   for VITAL_ACT
   end for;
end CFG_RAM64K36_VITAL;

-----------------------------------------------------------------
--
--  Actel AX RAM64K36P VHDL behavioral model
--  64K X 1 pipelined RAM with rising write clock and rising read clock.
--  Allows variable and independent Write and Read widths of only
--  4Kx1, 2Kx2, 1Kx4, 512x9, 256x18, or 128x36.
--  Depth pins functionally inert.  In model just to make sure 
--  they are connected.  Used by combiner to calculate cascading.
--
--  Future changes:  Need to be able to initialize RAM from text file.
--
--  Uses VITAL95 package
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - 11/22/00 - Dale Walter - Initial Version.
-- 1.1 - 03/14/01 - Dale Walter - Cloned from RAM64K36.
-- 1.2 - 05/10/01 - Dale Walter - Change memory to variable instead of signal.
--                              - Change WRAD & RDAD calculation to be the same
--                                regardless of WW and RR (i.e. low-order bits
--                                assumed to be tied-off to GND for widths > 1.
-- 1.3 - 9/27/02 - Krupa Singampalli - New Timing Arcs
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
entity RAM64K36P is
  GENERIC (
        tipd_DEPTH3   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH2   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH1   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_DEPTH0   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD15   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD14   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD13   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD12   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD11   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD10   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD9    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD8    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD7    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD6    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD5    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD35     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD34     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD33     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD32     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD31     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD30     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD29     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD28     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD27     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD26     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD25     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD24     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD23     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD22     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD21     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD20     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD19     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD18     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD17     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD16     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD15     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD14     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD13     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD12     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD11     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD10     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD9      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD8      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD7      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD6      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD5      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD4      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD3      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WD0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WW2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WW1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WW0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WEN      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD15   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD14   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD13   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD12   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD11   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD10   : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD9    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD8    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD7    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD6    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD5    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD4    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RW2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RW1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RW0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_REN      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);

        
        tpd_RCLK_RD0  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD1  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD2  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD3  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD4  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD5  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD6  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD7  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD8  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD9  : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD10 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD11 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD12 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD13 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD14 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD15 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD16 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD17 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD18 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD19 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD20 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD21 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD22 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD23 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD24 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD25 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD26 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD27 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD28 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD29 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD30 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD31 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD32 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD33 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD34 : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_RD35 : VitalDelayType01 := (0.100 ns, 0.100 ns);



        tsetup_RDAD15_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD14_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD13_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD12_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD11_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD10_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD9_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD8_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD7_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD6_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD5_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD4_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_RDAD15_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD14_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD13_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD12_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD11_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD10_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_RDAD9_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD8_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD7_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD6_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD5_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD4_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;



        tsetup_RW2_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW1_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW0_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW2_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW1_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RW0_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;


        tsetup_DEPTH3_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH2_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH1_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH0_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH3_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH2_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH1_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_DEPTH0_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;



        tsetup_WRAD15_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD14_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD13_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD12_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD11_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD10_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD9_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD8_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_WRAD15_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD14_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD13_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD12_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD11_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD10_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_WRAD9_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD8_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        tsetup_WD35_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD34_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD33_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD32_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD31_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD30_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD29_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD28_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD27_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD26_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD25_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD24_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD23_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD22_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD21_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD20_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD19_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD18_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD17_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD16_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD15_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD14_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD13_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD12_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD11_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD10_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD9_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD8_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD35_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD34_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD33_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD32_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD31_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD30_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD29_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD28_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD27_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD26_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD25_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD24_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD23_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD22_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD21_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD20_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD19_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD18_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD17_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD16_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD15_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD14_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD13_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD12_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD11_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD10_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        tsetup_WD9_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD8_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;



        tsetup_WW2_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW2_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WW0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;


        thold_RDAD15_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD14_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD13_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD12_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD11_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD10_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD9_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD8_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD7_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD6_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD5_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;

        thold_RDAD15_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD14_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD13_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD12_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD11_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD10_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_RDAD9_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD8_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD7_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD6_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD5_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;

        thold_RW2_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW1_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW0_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW2_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW1_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RW0_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

        thold_DEPTH3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_DEPTH0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        thold_WRAD15_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD14_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD13_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD12_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD11_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD10_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD9_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD8_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;

        thold_WRAD15_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD14_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD13_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD12_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD11_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD10_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_WRAD9_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD8_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;


        thold_WD35_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD34_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD33_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD32_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD31_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD30_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD29_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD28_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD27_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD26_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD25_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD24_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD23_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD22_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD21_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD20_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD19_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD18_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD17_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD16_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD15_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD14_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD13_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD12_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD11_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD10_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD9_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD8_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD35_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD34_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD33_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD32_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD31_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD30_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD29_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD28_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD27_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD26_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD25_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD24_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD23_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD22_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD21_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD20_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD19_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD18_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD17_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD16_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD15_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD14_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD13_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD12_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD11_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD10_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD9_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD8_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;


        thold_WW2_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW1_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW0_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW2_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW1_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WW0_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

        tsetup_REN_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;



        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True
        );
  PORT (
        DEPTH3 : IN STD_ULOGIC ;
        DEPTH2 : IN STD_ULOGIC ;
        DEPTH1 : IN STD_ULOGIC ;
        DEPTH0 : IN STD_ULOGIC ;
        WRAD15 : IN STD_ULOGIC ;
        WRAD14 : IN STD_ULOGIC ;
        WRAD13 : IN STD_ULOGIC ;
        WRAD12 : IN STD_ULOGIC ;
        WRAD11 : IN STD_ULOGIC ;
        WRAD10 : IN STD_ULOGIC ;
        WRAD9  : IN STD_ULOGIC ;
        WRAD8  : IN STD_ULOGIC ;
        WRAD7  : IN STD_ULOGIC ;
        WRAD6  : IN STD_ULOGIC ;
        WRAD5  : IN STD_ULOGIC ;
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD35   : IN STD_ULOGIC ;
        WD34   : IN STD_ULOGIC ;
        WD33   : IN STD_ULOGIC ;
        WD32   : IN STD_ULOGIC ;
        WD31   : IN STD_ULOGIC ;
        WD30   : IN STD_ULOGIC ;
        WD29   : IN STD_ULOGIC ;
        WD28   : IN STD_ULOGIC ;
        WD27   : IN STD_ULOGIC ;
        WD26   : IN STD_ULOGIC ;
        WD25   : IN STD_ULOGIC ;
        WD24   : IN STD_ULOGIC ;
        WD23   : IN STD_ULOGIC ;
        WD22   : IN STD_ULOGIC ;
        WD21   : IN STD_ULOGIC ;
        WD20   : IN STD_ULOGIC ;
        WD19   : IN STD_ULOGIC ;
        WD18   : IN STD_ULOGIC ;
        WD17   : IN STD_ULOGIC ;
        WD16   : IN STD_ULOGIC ;
        WD15   : IN STD_ULOGIC ;
        WD14   : IN STD_ULOGIC ;
        WD13   : IN STD_ULOGIC ;
        WD12   : IN STD_ULOGIC ;
        WD11   : IN STD_ULOGIC ;
        WD10   : IN STD_ULOGIC ;
        WD9    : IN STD_ULOGIC ;
        WD8    : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        WW2    : IN STD_ULOGIC ;
        WW1    : IN STD_ULOGIC ;
        WW0    : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RDAD15 : IN STD_ULOGIC ;
        RDAD14 : IN STD_ULOGIC ;
        RDAD13 : IN STD_ULOGIC ;
        RDAD12 : IN STD_ULOGIC ;
        RDAD11 : IN STD_ULOGIC ;
        RDAD10 : IN STD_ULOGIC ;
        RDAD9  : IN STD_ULOGIC ;
        RDAD8  : IN STD_ULOGIC ;
        RDAD7  : IN STD_ULOGIC ;
        RDAD6  : IN STD_ULOGIC ;
        RDAD5  : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        RW2    : IN STD_ULOGIC ;
        RW1    : IN STD_ULOGIC ;
        RW0    : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD35   : OUT STD_ULOGIC ;
        RD34   : OUT STD_ULOGIC ;
        RD33   : OUT STD_ULOGIC ;
        RD32   : OUT STD_ULOGIC ;
        RD31   : OUT STD_ULOGIC ;
        RD30   : OUT STD_ULOGIC ;
        RD29   : OUT STD_ULOGIC ;
        RD28   : OUT STD_ULOGIC ;
        RD27   : OUT STD_ULOGIC ;
        RD26   : OUT STD_ULOGIC ;
        RD25   : OUT STD_ULOGIC ;
        RD24   : OUT STD_ULOGIC ;
        RD23   : OUT STD_ULOGIC ;
        RD22   : OUT STD_ULOGIC ;
        RD21   : OUT STD_ULOGIC ;
        RD20   : OUT STD_ULOGIC ;
        RD19   : OUT STD_ULOGIC ;
        RD18   : OUT STD_ULOGIC ;
        RD17   : OUT STD_ULOGIC ;
        RD16   : OUT STD_ULOGIC ;
        RD15   : OUT STD_ULOGIC ;
        RD14   : OUT STD_ULOGIC ;
        RD13   : OUT STD_ULOGIC ;
        RD12   : OUT STD_ULOGIC ;
        RD11   : OUT STD_ULOGIC ;
        RD10   : OUT STD_ULOGIC ;
        RD9    : OUT STD_ULOGIC ;
        RD8    : OUT STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC ;
        RD6    : OUT STD_ULOGIC ;
        RD5    : OUT STD_ULOGIC ;
        RD4    : OUT STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC ;
        RD2    : OUT STD_ULOGIC ;
        RD1    : OUT STD_ULOGIC ;
        RD0    : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of RAM64K36P : entity is TRUE;
  
end RAM64K36P;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of RAM64K36P is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal DEPTH3_ipd : std_ulogic := 'X';
  signal DEPTH2_ipd : std_ulogic := 'X';
  signal DEPTH1_ipd : std_ulogic := 'X';
  signal DEPTH0_ipd : std_ulogic := 'X';
  signal WRAD15_ipd : std_ulogic := 'X';
  signal WRAD14_ipd : std_ulogic := 'X';
  signal WRAD13_ipd : std_ulogic := 'X';
  signal WRAD12_ipd : std_ulogic := 'X';
  signal WRAD11_ipd : std_ulogic := 'X';
  signal WRAD10_ipd : std_ulogic := 'X';
  signal WRAD9_ipd  : std_ulogic := 'X';
  signal WRAD8_ipd  : std_ulogic := 'X';
  signal WRAD7_ipd  : std_ulogic := 'X';
  signal WRAD6_ipd  : std_ulogic := 'X';
  signal WRAD5_ipd  : std_ulogic := 'X';
  signal WRAD4_ipd  : std_ulogic := 'X';
  signal WRAD3_ipd  : std_ulogic := 'X';
  signal WRAD2_ipd  : std_ulogic := 'X';
  signal WRAD1_ipd  : std_ulogic := 'X';
  signal WRAD0_ipd  : std_ulogic := 'X';
  signal WD35_ipd   : std_ulogic := 'X';
  signal WD34_ipd   : std_ulogic := 'X';
  signal WD33_ipd   : std_ulogic := 'X';
  signal WD32_ipd   : std_ulogic := 'X';
  signal WD31_ipd   : std_ulogic := 'X';
  signal WD30_ipd   : std_ulogic := 'X';
  signal WD29_ipd   : std_ulogic := 'X';
  signal WD28_ipd   : std_ulogic := 'X';
  signal WD27_ipd   : std_ulogic := 'X';
  signal WD26_ipd   : std_ulogic := 'X';
  signal WD25_ipd   : std_ulogic := 'X';
  signal WD24_ipd   : std_ulogic := 'X';
  signal WD23_ipd   : std_ulogic := 'X';
  signal WD22_ipd   : std_ulogic := 'X';
  signal WD21_ipd   : std_ulogic := 'X';
  signal WD20_ipd   : std_ulogic := 'X';
  signal WD19_ipd   : std_ulogic := 'X';
  signal WD18_ipd   : std_ulogic := 'X';
  signal WD17_ipd   : std_ulogic := 'X';
  signal WD16_ipd   : std_ulogic := 'X';
  signal WD15_ipd   : std_ulogic := 'X';
  signal WD14_ipd   : std_ulogic := 'X';
  signal WD13_ipd   : std_ulogic := 'X';
  signal WD12_ipd   : std_ulogic := 'X';
  signal WD11_ipd   : std_ulogic := 'X';
  signal WD10_ipd   : std_ulogic := 'X';
  signal WD9_ipd    : std_ulogic := 'X';
  signal WD8_ipd    : std_ulogic := 'X';
  signal WD7_ipd    : std_ulogic := 'X';
  signal WD6_ipd    : std_ulogic := 'X';
  signal WD5_ipd    : std_ulogic := 'X';
  signal WD4_ipd    : std_ulogic := 'X';
  signal WD3_ipd    : std_ulogic := 'X';
  signal WD2_ipd    : std_ulogic := 'X';
  signal WD1_ipd    : std_ulogic := 'X';
  signal WD0_ipd    : std_ulogic := 'X';
  signal WW2_ipd    : std_ulogic := 'X';
  signal WW1_ipd    : std_ulogic := 'X';
  signal WW0_ipd    : std_ulogic := 'X';
  signal WEN_ipd    : std_ulogic := 'X';
  signal WCLK_ipd   : std_ulogic := 'X';
  signal RDAD15_ipd : std_ulogic := 'X';
  signal RDAD14_ipd : std_ulogic := 'X';
  signal RDAD13_ipd : std_ulogic := 'X';
  signal RDAD12_ipd : std_ulogic := 'X';
  signal RDAD11_ipd : std_ulogic := 'X';
  signal RDAD10_ipd : std_ulogic := 'X';
  signal RDAD9_ipd  : std_ulogic := 'X';
  signal RDAD8_ipd  : std_ulogic := 'X';
  signal RDAD7_ipd  : std_ulogic := 'X';
  signal RDAD6_ipd  : std_ulogic := 'X';
  signal RDAD5_ipd  : std_ulogic := 'X';
  signal RDAD4_ipd  : std_ulogic := 'X';
  signal RDAD3_ipd  : std_ulogic := 'X';
  signal RDAD2_ipd  : std_ulogic := 'X';
  signal RDAD1_ipd  : std_ulogic := 'X';
  signal RDAD0_ipd  : std_ulogic := 'X';
  signal RW2_ipd    : std_ulogic := 'X';
  signal RW1_ipd    : std_ulogic := 'X';
  signal RW0_ipd    : std_ulogic := 'X';
  signal REN_ipd    : std_ulogic := 'X';
  signal RCLK_ipd   : std_ulogic := 'X';
  type MEM is array(0 to 65535) of std_ulogic; -- Internal memory
  type MEM9 is array(0 to 8191) of std_ulogic; -- Internal memory
  --signal RAM_TMP    : MEM;
  --signal RAM_TMP9   : MEM9;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (DEPTH3_ipd, DEPTH3, VitalExtendToFillDelay(tipd_DEPTH3));
    VitalWireDelay (DEPTH2_ipd, DEPTH2, VitalExtendToFillDelay(tipd_DEPTH2));
    VitalWireDelay (DEPTH1_ipd, DEPTH1, VitalExtendToFillDelay(tipd_DEPTH1));
    VitalWireDelay (DEPTH0_ipd, DEPTH0, VitalExtendToFillDelay(tipd_DEPTH0));
    VitalWireDelay (WRAD15_ipd, WRAD15, VitalExtendToFillDelay(tipd_WRAD15));
    VitalWireDelay (WRAD14_ipd, WRAD14, VitalExtendToFillDelay(tipd_WRAD14));
    VitalWireDelay (WRAD13_ipd, WRAD13, VitalExtendToFillDelay(tipd_WRAD13));
    VitalWireDelay (WRAD12_ipd, WRAD12, VitalExtendToFillDelay(tipd_WRAD12));
    VitalWireDelay (WRAD11_ipd, WRAD11, VitalExtendToFillDelay(tipd_WRAD11));
    VitalWireDelay (WRAD10_ipd, WRAD10, VitalExtendToFillDelay(tipd_WRAD10));
    VitalWireDelay (WRAD9_ipd, WRAD9, VitalExtendToFillDelay(tipd_WRAD9));
    VitalWireDelay (WRAD8_ipd, WRAD8, VitalExtendToFillDelay(tipd_WRAD8));
    VitalWireDelay (WRAD7_ipd, WRAD7, VitalExtendToFillDelay(tipd_WRAD7));
    VitalWireDelay (WRAD6_ipd, WRAD6, VitalExtendToFillDelay(tipd_WRAD6));
    VitalWireDelay (WRAD5_ipd, WRAD5, VitalExtendToFillDelay(tipd_WRAD5));
    VitalWireDelay (WRAD4_ipd, WRAD4, VitalExtendToFillDelay(tipd_WRAD4));
    VitalWireDelay (WRAD3_ipd, WRAD3, VitalExtendToFillDelay(tipd_WRAD3));
    VitalWireDelay (WRAD2_ipd, WRAD2, VitalExtendToFillDelay(tipd_WRAD2));
    VitalWireDelay (WRAD1_ipd, WRAD1, VitalExtendToFillDelay(tipd_WRAD1));
    VitalWireDelay (WRAD0_ipd, WRAD0, VitalExtendToFillDelay(tipd_WRAD0));
    VitalWireDelay (WD35_ipd, WD35, VitalExtendToFillDelay(tipd_WD35));
    VitalWireDelay (WD34_ipd, WD34, VitalExtendToFillDelay(tipd_WD34));
    VitalWireDelay (WD33_ipd, WD33, VitalExtendToFillDelay(tipd_WD33));
    VitalWireDelay (WD32_ipd, WD32, VitalExtendToFillDelay(tipd_WD32));
    VitalWireDelay (WD31_ipd, WD31, VitalExtendToFillDelay(tipd_WD31));
    VitalWireDelay (WD30_ipd, WD30, VitalExtendToFillDelay(tipd_WD30));
    VitalWireDelay (WD29_ipd, WD29, VitalExtendToFillDelay(tipd_WD29));
    VitalWireDelay (WD28_ipd, WD28, VitalExtendToFillDelay(tipd_WD28));
    VitalWireDelay (WD27_ipd, WD27, VitalExtendToFillDelay(tipd_WD27));
    VitalWireDelay (WD26_ipd, WD26, VitalExtendToFillDelay(tipd_WD26));
    VitalWireDelay (WD25_ipd, WD25, VitalExtendToFillDelay(tipd_WD25));
    VitalWireDelay (WD24_ipd, WD24, VitalExtendToFillDelay(tipd_WD24));
    VitalWireDelay (WD23_ipd, WD23, VitalExtendToFillDelay(tipd_WD23));
    VitalWireDelay (WD22_ipd, WD22, VitalExtendToFillDelay(tipd_WD22));
    VitalWireDelay (WD21_ipd, WD21, VitalExtendToFillDelay(tipd_WD21));
    VitalWireDelay (WD20_ipd, WD20, VitalExtendToFillDelay(tipd_WD20));
    VitalWireDelay (WD19_ipd, WD19, VitalExtendToFillDelay(tipd_WD19));
    VitalWireDelay (WD18_ipd, WD18, VitalExtendToFillDelay(tipd_WD18));
    VitalWireDelay (WD17_ipd, WD17, VitalExtendToFillDelay(tipd_WD17));
    VitalWireDelay (WD16_ipd, WD16, VitalExtendToFillDelay(tipd_WD16));
    VitalWireDelay (WD15_ipd, WD15, VitalExtendToFillDelay(tipd_WD15));
    VitalWireDelay (WD14_ipd, WD14, VitalExtendToFillDelay(tipd_WD14));
    VitalWireDelay (WD13_ipd, WD13, VitalExtendToFillDelay(tipd_WD13));
    VitalWireDelay (WD12_ipd, WD12, VitalExtendToFillDelay(tipd_WD12));
    VitalWireDelay (WD11_ipd, WD11, VitalExtendToFillDelay(tipd_WD11));
    VitalWireDelay (WD10_ipd, WD10, VitalExtendToFillDelay(tipd_WD10));
    VitalWireDelay (WD9_ipd, WD9, VitalExtendToFillDelay(tipd_WD9));
    VitalWireDelay (WD8_ipd, WD8, VitalExtendToFillDelay(tipd_WD8));
    VitalWireDelay (WD7_ipd, WD7, VitalExtendToFillDelay(tipd_WD7));
    VitalWireDelay (WD6_ipd, WD6, VitalExtendToFillDelay(tipd_WD6));
    VitalWireDelay (WD5_ipd, WD5, VitalExtendToFillDelay(tipd_WD5));
    VitalWireDelay (WD4_ipd, WD4, VitalExtendToFillDelay(tipd_WD4));
    VitalWireDelay (WD3_ipd, WD3, VitalExtendToFillDelay(tipd_WD3));
    VitalWireDelay (WD2_ipd, WD2, VitalExtendToFillDelay(tipd_WD2));
    VitalWireDelay (WD1_ipd, WD1, VitalExtendToFillDelay(tipd_WD1));
    VitalWireDelay (WD0_ipd, WD0, VitalExtendToFillDelay(tipd_WD0));
    VitalWireDelay (WW2_ipd, WW2, VitalExtendToFillDelay(tipd_WW2));
    VitalWireDelay (WW1_ipd, WW1, VitalExtendToFillDelay(tipd_WW1));
    VitalWireDelay (WW0_ipd, WW0, VitalExtendToFillDelay(tipd_WW0));
    VitalWireDelay (WEN_ipd, WEN, VitalExtendToFillDelay(tipd_WEN));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (RDAD15_ipd, RDAD15, VitalExtendToFillDelay(tipd_RDAD15));
    VitalWireDelay (RDAD14_ipd, RDAD14, VitalExtendToFillDelay(tipd_RDAD14));
    VitalWireDelay (RDAD13_ipd, RDAD13, VitalExtendToFillDelay(tipd_RDAD13));
    VitalWireDelay (RDAD12_ipd, RDAD12, VitalExtendToFillDelay(tipd_RDAD12));
    VitalWireDelay (RDAD11_ipd, RDAD11, VitalExtendToFillDelay(tipd_RDAD11));
    VitalWireDelay (RDAD10_ipd, RDAD10, VitalExtendToFillDelay(tipd_RDAD10));
    VitalWireDelay (RDAD9_ipd, RDAD9, VitalExtendToFillDelay(tipd_RDAD9));
    VitalWireDelay (RDAD8_ipd, RDAD8, VitalExtendToFillDelay(tipd_RDAD8));
    VitalWireDelay (RDAD7_ipd, RDAD7, VitalExtendToFillDelay(tipd_RDAD7));
    VitalWireDelay (RDAD6_ipd, RDAD6, VitalExtendToFillDelay(tipd_RDAD6));
    VitalWireDelay (RDAD5_ipd, RDAD5, VitalExtendToFillDelay(tipd_RDAD5));
    VitalWireDelay (RDAD4_ipd, RDAD4, VitalExtendToFillDelay(tipd_RDAD4));
    VitalWireDelay (RDAD3_ipd, RDAD3, VitalExtendToFillDelay(tipd_RDAD3));
    VitalWireDelay (RDAD2_ipd, RDAD2, VitalExtendToFillDelay(tipd_RDAD2));
    VitalWireDelay (RDAD1_ipd, RDAD1, VitalExtendToFillDelay(tipd_RDAD1));
    VitalWireDelay (RDAD0_ipd, RDAD0, VitalExtendToFillDelay(tipd_RDAD0));
    VitalWireDelay (RW2_ipd, RW2, VitalExtendToFillDelay(tipd_RW2));
    VitalWireDelay (RW1_ipd, RW1, VitalExtendToFillDelay(tipd_RW1));
    VitalWireDelay (RW0_ipd, RW0, VitalExtendToFillDelay(tipd_RW0));
    VitalWireDelay (REN_ipd, REN, VitalExtendToFillDelay(tipd_REN));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (DEPTH3_ipd, DEPTH2_ipd, DEPTH1_ipd, DEPTH0_ipd,
                WRAD15_ipd, WRAD14_ipd, WRAD13_ipd,
                WRAD12_ipd, WRAD11_ipd, WRAD10_ipd, WRAD9_ipd, 
                WRAD8_ipd, WRAD7_ipd, WRAD6_ipd, WRAD5_ipd, 
                WRAD4_ipd, WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd, 
                WD35_ipd, WD34_ipd, WD33_ipd, WD32_ipd, WD31_ipd, WD30_ipd,
                WD29_ipd, WD28_ipd, WD27_ipd, WD26_ipd, WD25_ipd, WD24_ipd,
                WD23_ipd, WD22_ipd, WD21_ipd, WD20_ipd, WD19_ipd, WD18_ipd,
                WD17_ipd, WD16_ipd, WD15_ipd, WD14_ipd, WD13_ipd, WD12_ipd,
                WD11_ipd, WD10_ipd, WD9_ipd, WD8_ipd, WD7_ipd, WD6_ipd,
                WD5_ipd, WD4_ipd, WD3_ipd, WD2_ipd, WD1_ipd, WD0_ipd,
                WW2_ipd, WW1_ipd, WW0_ipd, WEN_ipd, WCLK_ipd, 
                RDAD15_ipd, RDAD14_ipd, RDAD13_ipd, RDAD12_ipd, RDAD11_ipd, 
                RDAD10_ipd, RDAD9_ipd, RDAD8_ipd, RDAD7_ipd,
                RDAD6_ipd, RDAD5_ipd, RDAD4_ipd, RDAD3_ipd, RDAD2_ipd, 
                RDAD1_ipd, RDAD0_ipd, RW2_ipd, RW1_ipd, RW0_ipd,
                REN_ipd, RCLK_ipd)

     --  Memory
     variable RAM_TMP    : MEM;
     variable RAM_TMP9   : MEM9;
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT : SL_TO_INT := (-65537, -65537, 0, 1, -65537, -65537, 0, 1, -65537);

     --  Read Timing Check Results
     variable Tviol_RDAD15_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD15_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD14_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD14_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD13_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD13_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD12_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD12_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD11_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD11_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD10_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD10_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD9_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD9_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD8_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD8_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD7_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD7_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD6_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD6_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD5_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD5_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD4_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD4_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD3_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD3_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD2_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD1_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD0_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RW2_RCLK_posedge : X01 := '0';
     variable TmDt_RW2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RW1_RCLK_posedge : X01 := '0';
     variable TmDt_RW1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RW0_RCLK_posedge : X01 := '0';
     variable TmDt_RW0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_REN_RCLK_posedge : X01 := '0';
     variable TmDt_REN_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_WD35_WCLK_posedge : X01 := '0';
     variable TmDt_WD35_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD34_WCLK_posedge : X01 := '0';
     variable TmDt_WD34_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD33_WCLK_posedge : X01 := '0';
     variable TmDt_WD33_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD32_WCLK_posedge : X01 := '0';
     variable TmDt_WD32_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD31_WCLK_posedge : X01 := '0';
     variable TmDt_WD31_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD30_WCLK_posedge : X01 := '0';
     variable TmDt_WD30_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD29_WCLK_posedge : X01 := '0';
     variable TmDt_WD29_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD28_WCLK_posedge : X01 := '0';
     variable TmDt_WD28_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD27_WCLK_posedge : X01 := '0';
     variable TmDt_WD27_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD26_WCLK_posedge : X01 := '0';
     variable TmDt_WD26_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD25_WCLK_posedge : X01 := '0';
     variable TmDt_WD25_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD24_WCLK_posedge : X01 := '0';
     variable TmDt_WD24_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD23_WCLK_posedge : X01 := '0';
     variable TmDt_WD23_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD22_WCLK_posedge : X01 := '0';
     variable TmDt_WD22_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD21_WCLK_posedge : X01 := '0';
     variable TmDt_WD21_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD20_WCLK_posedge : X01 := '0';
     variable TmDt_WD20_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD19_WCLK_posedge : X01 := '0';
     variable TmDt_WD19_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD18_WCLK_posedge : X01 := '0';
     variable TmDt_WD18_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD17_WCLK_posedge : X01 := '0';
     variable TmDt_WD17_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD16_WCLK_posedge : X01 := '0';
     variable TmDt_WD16_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD15_WCLK_posedge : X01 := '0';
     variable TmDt_WD15_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD14_WCLK_posedge : X01 := '0';
     variable TmDt_WD14_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD13_WCLK_posedge : X01 := '0';
     variable TmDt_WD13_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD12_WCLK_posedge : X01 := '0';
     variable TmDt_WD12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD11_WCLK_posedge : X01 := '0';
     variable TmDt_WD11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD10_WCLK_posedge : X01 := '0';
     variable TmDt_WD10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD9_WCLK_posedge : X01 := '0';
     variable TmDt_WD9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD8_WCLK_posedge : X01 := '0';
     variable TmDt_WD8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD7_WCLK_posedge : X01 := '0';
     variable TmDt_WD7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD6_WCLK_posedge : X01 := '0';
     variable TmDt_WD6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD5_WCLK_posedge : X01 := '0';
     variable TmDt_WD5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD4_WCLK_posedge : X01 := '0';
     variable TmDt_WD4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD3_WCLK_posedge : X01 := '0';
     variable TmDt_WD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD2_WCLK_posedge : X01 := '0';
     variable TmDt_WD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD1_WCLK_posedge : X01 := '0';
     variable TmDt_WD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD0_WCLK_posedge : X01 := '0';
     variable TmDt_WD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WW2_WCLK_posedge : X01 := '0';
     variable TmDt_WW2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WW1_WCLK_posedge : X01 := '0';
     variable TmDt_WW1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WW0_WCLK_posedge : X01 := '0';
     variable TmDt_WW0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD15_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD15_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD14_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD14_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD13_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD13_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD12_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD11_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD10_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD9_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD8_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD7_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD6_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD5_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD4_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD3_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD2_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD1_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD0_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DEPTH3_WCLK_posedge : X01 := '0';
     variable TmDt_DEPTH3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DEPTH2_WCLK_posedge : X01 := '0';
     variable TmDt_DEPTH2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DEPTH1_WCLK_posedge : X01 := '0';
     variable TmDt_DEPTH1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DEPTH0_WCLK_posedge : X01 := '0';
     variable TmDt_DEPTH0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WEN_WCLK_posedge : X01 := '0';
     variable TmDt_WEN_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  Functional Results
     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     variable WWIDTH : integer := -1;
     variable RWIDTH : integer := -1;
     variable RD35_zd : std_ulogic;
     variable RD34_zd : std_ulogic;
     variable RD33_zd : std_ulogic;
     variable RD32_zd : std_ulogic;
     variable RD31_zd : std_ulogic;
     variable RD30_zd : std_ulogic;
     variable RD29_zd : std_ulogic;
     variable RD28_zd : std_ulogic;
     variable RD27_zd : std_ulogic;
     variable RD26_zd : std_ulogic;
     variable RD25_zd : std_ulogic;
     variable RD24_zd : std_ulogic;
     variable RD23_zd : std_ulogic;
     variable RD22_zd : std_ulogic;
     variable RD21_zd : std_ulogic;
     variable RD20_zd : std_ulogic;
     variable RD19_zd : std_ulogic;
     variable RD18_zd : std_ulogic;
     variable RD17_zd : std_ulogic;
     variable RD16_zd : std_ulogic;
     variable RD15_zd : std_ulogic;
     variable RD14_zd : std_ulogic;
     variable RD13_zd : std_ulogic;
     variable RD12_zd : std_ulogic;
     variable RD11_zd : std_ulogic;
     variable RD10_zd : std_ulogic;
     variable RD9_zd : std_ulogic;
     variable RD8_zd : std_ulogic;
     variable RD7_zd : std_ulogic;
     variable RD6_zd : std_ulogic;
     variable RD5_zd : std_ulogic;
     variable RD4_zd : std_ulogic;
     variable RD3_zd : std_ulogic;
     variable RD2_zd : std_ulogic;
     variable RD1_zd : std_ulogic;
     variable RD0_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable RD35_GlitchData : VitalGlitchDataType;
     variable RD34_GlitchData : VitalGlitchDataType;
     variable RD33_GlitchData : VitalGlitchDataType;
     variable RD32_GlitchData : VitalGlitchDataType;
     variable RD31_GlitchData : VitalGlitchDataType;
     variable RD30_GlitchData : VitalGlitchDataType;
     variable RD29_GlitchData : VitalGlitchDataType;
     variable RD28_GlitchData : VitalGlitchDataType;
     variable RD27_GlitchData : VitalGlitchDataType;
     variable RD26_GlitchData : VitalGlitchDataType;
     variable RD25_GlitchData : VitalGlitchDataType;
     variable RD24_GlitchData : VitalGlitchDataType;
     variable RD23_GlitchData : VitalGlitchDataType;
     variable RD22_GlitchData : VitalGlitchDataType;
     variable RD21_GlitchData : VitalGlitchDataType;
     variable RD20_GlitchData : VitalGlitchDataType;
     variable RD19_GlitchData : VitalGlitchDataType;
     variable RD18_GlitchData : VitalGlitchDataType;
     variable RD17_GlitchData : VitalGlitchDataType;
     variable RD16_GlitchData : VitalGlitchDataType;
     variable RD15_GlitchData : VitalGlitchDataType;
     variable RD14_GlitchData : VitalGlitchDataType;
     variable RD13_GlitchData : VitalGlitchDataType;
     variable RD12_GlitchData : VitalGlitchDataType;
     variable RD11_GlitchData : VitalGlitchDataType;
     variable RD10_GlitchData : VitalGlitchDataType;
     variable RD9_GlitchData : VitalGlitchDataType;
     variable RD8_GlitchData : VitalGlitchDataType;
     variable RD7_GlitchData : VitalGlitchDataType;
     variable RD6_GlitchData : VitalGlitchDataType;
     variable RD5_GlitchData : VitalGlitchDataType;
     variable RD4_GlitchData : VitalGlitchDataType;
     variable RD3_GlitchData : VitalGlitchDataType;
     variable RD2_GlitchData : VitalGlitchDataType;
     variable RD1_GlitchData : VitalGlitchDataType;
     variable RD0_GlitchData : VitalGlitchDataType;

     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable REN_delayed  : std_ulogic := 'X';
     variable REN_previous : std_ulogic := 'X';
     variable WEN_delayed  : std_ulogic := 'X';
     variable WD35_delayed : std_ulogic := 'X';
     variable WD34_delayed : std_ulogic := 'X';
     variable WD33_delayed : std_ulogic := 'X';
     variable WD32_delayed : std_ulogic := 'X';
     variable WD31_delayed : std_ulogic := 'X';
     variable WD30_delayed : std_ulogic := 'X';
     variable WD29_delayed : std_ulogic := 'X';
     variable WD28_delayed : std_ulogic := 'X';
     variable WD27_delayed : std_ulogic := 'X';
     variable WD26_delayed : std_ulogic := 'X';
     variable WD25_delayed : std_ulogic := 'X';
     variable WD24_delayed : std_ulogic := 'X';
     variable WD23_delayed : std_ulogic := 'X';
     variable WD22_delayed : std_ulogic := 'X';
     variable WD21_delayed : std_ulogic := 'X';
     variable WD20_delayed : std_ulogic := 'X';
     variable WD19_delayed : std_ulogic := 'X';
     variable WD18_delayed : std_ulogic := 'X';
     variable WD17_delayed : std_ulogic := 'X';
     variable WD16_delayed : std_ulogic := 'X';
     variable WD15_delayed : std_ulogic := 'X';
     variable WD14_delayed : std_ulogic := 'X';
     variable WD13_delayed : std_ulogic := 'X';
     variable WD12_delayed : std_ulogic := 'X';
     variable WD11_delayed : std_ulogic := 'X';
     variable WD10_delayed : std_ulogic := 'X';
     variable WD9_delayed : std_ulogic := 'X';
     variable WD8_delayed : std_ulogic := 'X';
     variable WD7_delayed : std_ulogic := 'X';
     variable WD6_delayed : std_ulogic := 'X';
     variable WD5_delayed : std_ulogic := 'X';
     variable WD4_delayed : std_ulogic := 'X';
     variable WD3_delayed : std_ulogic := 'X';
     variable WD2_delayed : std_ulogic := 'X';
     variable WD1_delayed : std_ulogic := 'X';
     variable WD0_delayed : std_ulogic := 'X';
     variable WW2_delayed : std_ulogic := 'X';
     variable WW1_delayed : std_ulogic := 'X';
     variable WW0_delayed : std_ulogic := 'X';
     variable DEPTH3_delayed : std_ulogic := 'X';
     variable DEPTH2_delayed : std_ulogic := 'X';
     variable DEPTH1_delayed : std_ulogic := 'X';
     variable DEPTH0_delayed : std_ulogic := 'X';
     variable WRAD15_delayed : std_ulogic := 'X';
     variable WRAD14_delayed : std_ulogic := 'X';
     variable WRAD13_delayed : std_ulogic := 'X';
     variable WRAD12_delayed : std_ulogic := 'X';
     variable WRAD11_delayed : std_ulogic := 'X';
     variable WRAD10_delayed : std_ulogic := 'X';
     variable WRAD9_delayed : std_ulogic := 'X';
     variable WRAD8_delayed : std_ulogic := 'X';
     variable WRAD7_delayed : std_ulogic := 'X';
     variable WRAD6_delayed : std_ulogic := 'X';
     variable WRAD5_delayed : std_ulogic := 'X';
     variable WRAD4_delayed : std_ulogic := 'X';
     variable WRAD3_delayed : std_ulogic := 'X';
     variable WRAD2_delayed : std_ulogic := 'X';
     variable WRAD1_delayed : std_ulogic := 'X';
     variable WRAD0_delayed : std_ulogic := 'X';
     variable RDAD15_delayed : std_ulogic := 'X';
     variable RDAD14_delayed : std_ulogic := 'X';
     variable RDAD13_delayed : std_ulogic := 'X';
     variable RDAD12_delayed : std_ulogic := 'X';
     variable RDAD11_delayed : std_ulogic := 'X';
     variable RDAD10_delayed : std_ulogic := 'X';
     variable RDAD9_delayed : std_ulogic := 'X';
     variable RDAD8_delayed : std_ulogic := 'X';
     variable RDAD7_delayed : std_ulogic := 'X';
     variable RDAD6_delayed : std_ulogic := 'X';
     variable RDAD5_delayed : std_ulogic := 'X';
     variable RDAD4_delayed : std_ulogic := 'X';
     variable RDAD3_delayed : std_ulogic := 'X';
     variable RDAD2_delayed : std_ulogic := 'X';
     variable RDAD1_delayed : std_ulogic := 'X';
     variable RDAD0_delayed : std_ulogic := 'X';
     variable RW2_delayed : std_ulogic := 'X';
     variable RW1_delayed : std_ulogic := 'X';
     variable RW0_delayed : std_ulogic := 'X';
     variable RDAD15_previous : std_ulogic := 'X';
     variable RDAD14_previous : std_ulogic := 'X';
     variable RDAD13_previous : std_ulogic := 'X';
     variable RDAD12_previous : std_ulogic := 'X';
     variable RDAD11_previous : std_ulogic := 'X';
     variable RDAD10_previous : std_ulogic := 'X';
     variable RDAD9_previous : std_ulogic := 'X';
     variable RDAD8_previous : std_ulogic := 'X';
     variable RDAD7_previous : std_ulogic := 'X';
     variable RDAD6_previous : std_ulogic := 'X';
     variable RDAD5_previous : std_ulogic := 'X';
     variable RDAD4_previous : std_ulogic := 'X';
     variable RDAD3_previous : std_ulogic := 'X';
     variable RDAD2_previous : std_ulogic := 'X';
     variable RDAD1_previous : std_ulogic := 'X';
     variable RDAD0_previous : std_ulogic := 'X';
     variable RW2_previous : std_ulogic := 'X';
     variable RW1_previous : std_ulogic := 'X';
     variable RW0_previous : std_ulogic := 'X';

     --  Pipelined temporary results
     variable REN_stg1 : std_ulogic;
     
     variable RD35_stg1 : std_ulogic;
     variable RD34_stg1 : std_ulogic;
     variable RD33_stg1 : std_ulogic;
     variable RD32_stg1 : std_ulogic;
     variable RD31_stg1 : std_ulogic;
     variable RD30_stg1 : std_ulogic;
     variable RD29_stg1 : std_ulogic;
     variable RD28_stg1 : std_ulogic;
     variable RD27_stg1 : std_ulogic;
     variable RD26_stg1 : std_ulogic;
     variable RD25_stg1 : std_ulogic;
     variable RD24_stg1 : std_ulogic;
     variable RD23_stg1 : std_ulogic;
     variable RD22_stg1 : std_ulogic;
     variable RD21_stg1 : std_ulogic;
     variable RD20_stg1 : std_ulogic;
     variable RD19_stg1 : std_ulogic;
     variable RD18_stg1 : std_ulogic;
     variable RD17_stg1 : std_ulogic;
     variable RD16_stg1 : std_ulogic;
     variable RD15_stg1 : std_ulogic;
     variable RD14_stg1 : std_ulogic;
     variable RD13_stg1 : std_ulogic;
     variable RD12_stg1 : std_ulogic;
     variable RD11_stg1 : std_ulogic;
     variable RD10_stg1 : std_ulogic;
     variable RD9_stg1 : std_ulogic;
     variable RD8_stg1 : std_ulogic;
     variable RD7_stg1 : std_ulogic;
     variable RD6_stg1 : std_ulogic;
     variable RD5_stg1 : std_ulogic;
     variable RD4_stg1 : std_ulogic;
     variable RD3_stg1 : std_ulogic;
     variable RD2_stg1 : std_ulogic;
     variable RD1_stg1 : std_ulogic;
     variable RD0_stg1 : std_ulogic;

  begin  --  process VITALBehavior 

    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RDAD high or low before RCLK rising
      --   Hold  RDAD high or low after RCLK rising

      VitalSetupHoldCheck ( Tviol_RDAD15_RCLK_posedge,
                            TmDt_RDAD15_RCLK_posedge,
                            RDAD15_ipd, "RDAD15",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD15_RCLK_posedge_posedge,
                            tsetup_RDAD15_RCLK_negedge_posedge,
                            thold_RDAD15_RCLK_posedge_posedge,
                            thold_RDAD15_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD14_RCLK_posedge,
                            TmDt_RDAD14_RCLK_posedge,
                            RDAD14_ipd, "RDAD14",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD14_RCLK_posedge_posedge,
                            tsetup_RDAD14_RCLK_negedge_posedge,
                            thold_RDAD14_RCLK_posedge_posedge,
                            thold_RDAD14_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD13_RCLK_posedge,
                            TmDt_RDAD13_RCLK_posedge,
                            RDAD13_ipd, "RDAD13",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD13_RCLK_posedge_posedge,
                            tsetup_RDAD13_RCLK_negedge_posedge,
                            thold_RDAD13_RCLK_posedge_posedge,
                            thold_RDAD13_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD12_RCLK_posedge,
                            TmDt_RDAD12_RCLK_posedge,
                            RDAD12_ipd, "RDAD12",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD12_RCLK_posedge_posedge,
                            tsetup_RDAD12_RCLK_negedge_posedge,
                            thold_RDAD12_RCLK_posedge_posedge,
                            thold_RDAD12_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD11_RCLK_posedge,
                            TmDt_RDAD11_RCLK_posedge,
                            RDAD11_ipd, "RDAD11",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD11_RCLK_posedge_posedge,
                            tsetup_RDAD11_RCLK_negedge_posedge,
                            thold_RDAD11_RCLK_posedge_posedge,
                            thold_RDAD11_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD10_RCLK_posedge,
                            TmDt_RDAD10_RCLK_posedge,
                            RDAD10_ipd, "RDAD10",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD10_RCLK_posedge_posedge,
                            tsetup_RDAD10_RCLK_negedge_posedge,
                            thold_RDAD10_RCLK_posedge_posedge,
                            thold_RDAD10_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD9_RCLK_posedge,
                            TmDt_RDAD9_RCLK_posedge,
                            RDAD9_ipd, "RDAD9",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD9_RCLK_posedge_posedge,
                            tsetup_RDAD9_RCLK_negedge_posedge,
                            thold_RDAD9_RCLK_posedge_posedge,
                            thold_RDAD9_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD8_RCLK_posedge,
                            TmDt_RDAD8_RCLK_posedge,
                            RDAD8_ipd, "RDAD8",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD8_RCLK_posedge_posedge,
                            tsetup_RDAD8_RCLK_negedge_posedge,
                            thold_RDAD8_RCLK_posedge_posedge,
                            thold_RDAD8_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD7_RCLK_posedge,
                            TmDt_RDAD7_RCLK_posedge,
                            RDAD7_ipd, "RDAD7",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD7_RCLK_posedge_posedge,
                            tsetup_RDAD7_RCLK_negedge_posedge,
                            thold_RDAD7_RCLK_posedge_posedge,
                            thold_RDAD7_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD6_RCLK_posedge,
                            TmDt_RDAD6_RCLK_posedge,
                            RDAD6_ipd, "RDAD6",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD6_RCLK_posedge_posedge,
                            tsetup_RDAD6_RCLK_negedge_posedge,
                            thold_RDAD6_RCLK_posedge_posedge,
                            thold_RDAD6_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD5_RCLK_posedge,
                            TmDt_RDAD5_RCLK_posedge,
                            RDAD5_ipd, "RDAD5",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD5_RCLK_posedge_posedge,
                            tsetup_RDAD5_RCLK_negedge_posedge,
                            thold_RDAD5_RCLK_posedge_posedge,
                            thold_RDAD5_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD4_RCLK_posedge,
                            TmDt_RDAD4_RCLK_posedge,
                            RDAD4_ipd, "RDAD4",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD4_RCLK_posedge_posedge,
                            tsetup_RDAD4_RCLK_negedge_posedge,
                            thold_RDAD4_RCLK_posedge_posedge,
                            thold_RDAD4_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD3_RCLK_posedge,
                            TmDt_RDAD3_RCLK_posedge,
                            RDAD3_ipd, "RDAD3",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD3_RCLK_posedge_posedge,
                            tsetup_RDAD3_RCLK_negedge_posedge,
                            thold_RDAD3_RCLK_posedge_posedge,
                            thold_RDAD3_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD2_RCLK_posedge,
                            TmDt_RDAD2_RCLK_posedge,
                            RDAD2_ipd, "RDAD2",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD2_RCLK_posedge_posedge,
                            tsetup_RDAD2_RCLK_negedge_posedge,
                            thold_RDAD2_RCLK_posedge_posedge,
                            thold_RDAD2_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD1_RCLK_posedge,
                            TmDt_RDAD1_RCLK_posedge,
                            RDAD1_ipd, "RDAD1",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD1_RCLK_posedge_posedge,
                            tsetup_RDAD1_RCLK_negedge_posedge,
                            thold_RDAD1_RCLK_posedge_posedge,
                            thold_RDAD1_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RDAD0_RCLK_posedge,
                            TmDt_RDAD0_RCLK_posedge,
                            RDAD0_ipd, "RDAD0",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD0_RCLK_posedge_posedge,
                            tsetup_RDAD0_RCLK_negedge_posedge,
                            thold_RDAD0_RCLK_posedge_posedge,
                            thold_RDAD0_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup RW high before RCLK rising
      --   Hold  RW high after RCLK rising

      VitalSetupHoldCheck ( Tviol_RW2_RCLK_posedge,
                            TmDt_RW2_RCLK_posedge,
                            RW2_ipd, "RW2",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RW2_RCLK_posedge_posedge,
                            tsetup_RW2_RCLK_negedge_posedge,
                            thold_RW2_RCLK_posedge_posedge,
                            thold_RW2_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RW1_RCLK_posedge,
                            TmDt_RW1_RCLK_posedge,
                            RW1_ipd, "RW1",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RW1_RCLK_posedge_posedge,
                            tsetup_RW1_RCLK_negedge_posedge,
                            thold_RW1_RCLK_posedge_posedge,
                            thold_RW1_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_RW0_RCLK_posedge,
                            TmDt_RW0_RCLK_posedge,
                            RW0_ipd, "RW0",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RW0_RCLK_posedge_posedge,
                            tsetup_RW0_RCLK_negedge_posedge,
                            thold_RW0_RCLK_posedge_posedge,
                            thold_RW0_RCLK_negedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup REN high before RCLK rising
      --   Hold  REN high after RCLK rising

      VitalSetupHoldCheck ( Tviol_REN_RCLK_posedge,
                            TmDt_REN_RCLK_posedge,
                            REN_ipd, "REN",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_REN_RCLK_posedge_posedge,
			    tsetup_REN_RCLK_negedge_posedge,
                            thold_REN_RCLK_posedge_posedge,
                            thold_REN_RCLK_negedge_posedge,
                            TimingCheckOn,
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup DEPTH high or low before WCLK rising
      --   Hold  DEPTH high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_DEPTH3_WCLK_posedge,
                            TmDt_DEPTH3_WCLK_posedge,
                            DEPTH3_ipd, "DEPTH3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_DEPTH3_WCLK_posedge_posedge,
                            tsetup_DEPTH3_WCLK_negedge_posedge,
                            thold_DEPTH3_WCLK_posedge_posedge,
                            thold_DEPTH3_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_DEPTH2_WCLK_posedge,
                            TmDt_DEPTH2_WCLK_posedge,
                            DEPTH2_ipd, "DEPTH2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_DEPTH2_WCLK_posedge_posedge,
                            tsetup_DEPTH2_WCLK_negedge_posedge,
                            thold_DEPTH2_WCLK_posedge_posedge,
                            thold_DEPTH2_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_DEPTH1_WCLK_posedge,
                            TmDt_DEPTH1_WCLK_posedge,
                            DEPTH1_ipd, "DEPTH1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_DEPTH1_WCLK_posedge_posedge,
                            tsetup_DEPTH1_WCLK_negedge_posedge,
                            thold_DEPTH1_WCLK_posedge_posedge,
                            thold_DEPTH1_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_DEPTH0_WCLK_posedge,
                            TmDt_DEPTH0_WCLK_posedge,
                            DEPTH0_ipd, "DEPTH0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_DEPTH0_WCLK_posedge_posedge,
                            tsetup_DEPTH0_WCLK_negedge_posedge,
                            thold_DEPTH0_WCLK_posedge_posedge,
                            thold_DEPTH0_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      --   Setup WRAD high or low before WCLK rising
      --   Hold  WRAD high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WRAD15_WCLK_posedge,
                            TmDt_WRAD15_WCLK_posedge,
                            WRAD15_ipd, "WRAD15",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD15_WCLK_posedge_posedge,
                            tsetup_WRAD15_WCLK_negedge_posedge,
                            thold_WRAD15_WCLK_posedge_posedge,
                            thold_WRAD15_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD14_WCLK_posedge,
                            TmDt_WRAD14_WCLK_posedge,
                            WRAD14_ipd, "WRAD14",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD14_WCLK_posedge_posedge,
                            tsetup_WRAD14_WCLK_negedge_posedge,
                            thold_WRAD14_WCLK_posedge_posedge,
                            thold_WRAD14_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD13_WCLK_posedge,
                            TmDt_WRAD13_WCLK_posedge,
                            WRAD13_ipd, "WRAD13",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD13_WCLK_posedge_posedge,
                            tsetup_WRAD13_WCLK_negedge_posedge,
                            thold_WRAD13_WCLK_posedge_posedge,
                            thold_WRAD13_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD12_WCLK_posedge,
                            TmDt_WRAD12_WCLK_posedge,
                            WRAD12_ipd, "WRAD12",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD12_WCLK_posedge_posedge,
                            tsetup_WRAD12_WCLK_negedge_posedge,
                            thold_WRAD12_WCLK_posedge_posedge,
                            thold_WRAD12_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD11_WCLK_posedge,
                            TmDt_WRAD11_WCLK_posedge,
                            WRAD11_ipd, "WRAD11",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD11_WCLK_posedge_posedge,
                            tsetup_WRAD11_WCLK_negedge_posedge,
                            thold_WRAD11_WCLK_posedge_posedge,
                            thold_WRAD11_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD10_WCLK_posedge,
                            TmDt_WRAD10_WCLK_posedge,
                            WRAD10_ipd, "WRAD10",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD10_WCLK_posedge_posedge,
                            tsetup_WRAD10_WCLK_negedge_posedge,
                            thold_WRAD10_WCLK_posedge_posedge,
                            thold_WRAD10_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD9_WCLK_posedge,
                            TmDt_WRAD9_WCLK_posedge,
                            WRAD9_ipd, "WRAD9",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD9_WCLK_posedge_posedge,
                            tsetup_WRAD9_WCLK_negedge_posedge,
                            thold_WRAD9_WCLK_posedge_posedge,
                            thold_WRAD9_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD8_WCLK_posedge,
                            TmDt_WRAD8_WCLK_posedge,
                            WRAD8_ipd, "WRAD8",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD8_WCLK_posedge_posedge,
                            tsetup_WRAD8_WCLK_negedge_posedge,
                            thold_WRAD8_WCLK_posedge_posedge,
                            thold_WRAD8_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD7_WCLK_posedge,
                            TmDt_WRAD7_WCLK_posedge,
                            WRAD7_ipd, "WRAD7",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD7_WCLK_posedge_posedge,
                            tsetup_WRAD7_WCLK_negedge_posedge,
                            thold_WRAD7_WCLK_posedge_posedge,
                            thold_WRAD7_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD6_WCLK_posedge,
                            TmDt_WRAD6_WCLK_posedge,
                            WRAD6_ipd, "WRAD6",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD6_WCLK_posedge_posedge,
                            tsetup_WRAD6_WCLK_negedge_posedge,
                            thold_WRAD6_WCLK_posedge_posedge,
                            thold_WRAD6_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD5_WCLK_posedge,
                            TmDt_WRAD5_WCLK_posedge,
                            WRAD5_ipd, "WRAD5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD5_WCLK_posedge_posedge,
                            tsetup_WRAD5_WCLK_negedge_posedge,
                            thold_WRAD5_WCLK_posedge_posedge,
                            thold_WRAD5_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD4_WCLK_posedge,
                            TmDt_WRAD4_WCLK_posedge,
                            WRAD4_ipd, "WRAD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD4_WCLK_posedge_posedge,
                            tsetup_WRAD4_WCLK_negedge_posedge,
                            thold_WRAD4_WCLK_posedge_posedge,
                            thold_WRAD4_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD3_WCLK_posedge,
                            TmDt_WRAD3_WCLK_posedge,
                            WRAD3_ipd, "WRAD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD3_WCLK_posedge_posedge,
                            tsetup_WRAD3_WCLK_negedge_posedge,
                            thold_WRAD3_WCLK_posedge_posedge,
                            thold_WRAD3_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD2_WCLK_posedge,
                            TmDt_WRAD2_WCLK_posedge,
                            WRAD2_ipd, "WRAD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD2_WCLK_posedge_posedge,
                            tsetup_WRAD2_WCLK_negedge_posedge,
                            thold_WRAD2_WCLK_posedge_posedge,
                            thold_WRAD2_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD1_WCLK_posedge,
                            TmDt_WRAD1_WCLK_posedge,
                            WRAD1_ipd, "WRAD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD1_WCLK_posedge_posedge,
                            tsetup_WRAD1_WCLK_negedge_posedge,
                            thold_WRAD1_WCLK_posedge_posedge,
                            thold_WRAD1_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD0_WCLK_posedge,
                            TmDt_WRAD0_WCLK_posedge,
                            WRAD0_ipd, "WRAD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD0_WCLK_posedge_posedge,
                            tsetup_WRAD0_WCLK_negedge_posedge,
                            thold_WRAD0_WCLK_posedge_posedge,
                            thold_WRAD0_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
                            
      --   Setup WD high or low before WCLK rising
      --   Hold  WD high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WD35_WCLK_posedge,
                            TmDt_WD35_WCLK_posedge,
                            WD35_ipd, "WD35",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD35_WCLK_posedge_posedge,
                            tsetup_WD35_WCLK_negedge_posedge,
                            thold_WD35_WCLK_posedge_posedge,
                            thold_WD35_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD34_WCLK_posedge,
                            TmDt_WD34_WCLK_posedge,
                            WD34_ipd, "WD34",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD34_WCLK_posedge_posedge,
                            tsetup_WD34_WCLK_negedge_posedge,
                            thold_WD34_WCLK_posedge_posedge,
                            thold_WD34_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD33_WCLK_posedge,
                            TmDt_WD33_WCLK_posedge,
                            WD33_ipd, "WD33",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD33_WCLK_posedge_posedge,
                            tsetup_WD33_WCLK_negedge_posedge,
                            thold_WD33_WCLK_posedge_posedge,
                            thold_WD33_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD32_WCLK_posedge,
                            TmDt_WD32_WCLK_posedge,
                            WD32_ipd, "WD32",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD32_WCLK_posedge_posedge,
                            tsetup_WD32_WCLK_negedge_posedge,
                            thold_WD32_WCLK_posedge_posedge,
                            thold_WD32_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD31_WCLK_posedge,
                            TmDt_WD31_WCLK_posedge,
                            WD31_ipd, "WD31",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD31_WCLK_posedge_posedge,
                            tsetup_WD31_WCLK_negedge_posedge,
                            thold_WD31_WCLK_posedge_posedge,
                            thold_WD31_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD30_WCLK_posedge,
                            TmDt_WD30_WCLK_posedge,
                            WD30_ipd, "WD30",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD30_WCLK_posedge_posedge,
                            tsetup_WD30_WCLK_negedge_posedge,
                            thold_WD30_WCLK_posedge_posedge,
                            thold_WD30_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD29_WCLK_posedge,
                            TmDt_WD29_WCLK_posedge,
                            WD29_ipd, "WD29",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD29_WCLK_posedge_posedge,
                            tsetup_WD29_WCLK_negedge_posedge,
                            thold_WD29_WCLK_posedge_posedge,
                            thold_WD29_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD28_WCLK_posedge,
                            TmDt_WD28_WCLK_posedge,
                            WD28_ipd, "WD28",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD28_WCLK_posedge_posedge,
                            tsetup_WD28_WCLK_negedge_posedge,
                            thold_WD28_WCLK_posedge_posedge,
                            thold_WD28_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD27_WCLK_posedge,
                            TmDt_WD27_WCLK_posedge,
                            WD27_ipd, "WD27",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD27_WCLK_posedge_posedge,
                            tsetup_WD27_WCLK_negedge_posedge,
                            thold_WD27_WCLK_posedge_posedge,
                            thold_WD27_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD26_WCLK_posedge,
                            TmDt_WD26_WCLK_posedge,
                            WD26_ipd, "WD26",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD26_WCLK_posedge_posedge,
                            tsetup_WD26_WCLK_negedge_posedge,
                            thold_WD26_WCLK_posedge_posedge,
                            thold_WD26_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD25_WCLK_posedge,
                            TmDt_WD25_WCLK_posedge,
                            WD25_ipd, "WD25",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD25_WCLK_posedge_posedge,
                            tsetup_WD25_WCLK_negedge_posedge,
                            thold_WD25_WCLK_posedge_posedge,
                            thold_WD25_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD24_WCLK_posedge,
                            TmDt_WD24_WCLK_posedge,
                            WD24_ipd, "WD24",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD24_WCLK_posedge_posedge,
                            tsetup_WD24_WCLK_negedge_posedge,
                            thold_WD24_WCLK_posedge_posedge,
                            thold_WD24_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD23_WCLK_posedge,
                            TmDt_WD23_WCLK_posedge,
                            WD23_ipd, "WD23",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD23_WCLK_posedge_posedge,
                            tsetup_WD23_WCLK_negedge_posedge,
                            thold_WD23_WCLK_posedge_posedge,
                            thold_WD23_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD22_WCLK_posedge,
                            TmDt_WD22_WCLK_posedge,
                            WD22_ipd, "WD22",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD22_WCLK_posedge_posedge,
                            tsetup_WD22_WCLK_negedge_posedge,
                            thold_WD22_WCLK_posedge_posedge,
                            thold_WD22_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD21_WCLK_posedge,
                            TmDt_WD21_WCLK_posedge,
                            WD21_ipd, "WD21",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD21_WCLK_posedge_posedge,
                            tsetup_WD21_WCLK_negedge_posedge,
                            thold_WD21_WCLK_posedge_posedge,
                            thold_WD21_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD20_WCLK_posedge,
                            TmDt_WD20_WCLK_posedge,
                            WD20_ipd, "WD20",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD20_WCLK_posedge_posedge,
                            tsetup_WD20_WCLK_negedge_posedge,
                            thold_WD20_WCLK_posedge_posedge,
                            thold_WD20_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD19_WCLK_posedge,
                            TmDt_WD19_WCLK_posedge,
                            WD19_ipd, "WD19",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD19_WCLK_posedge_posedge,
                            tsetup_WD19_WCLK_negedge_posedge,
                            thold_WD19_WCLK_posedge_posedge,
                            thold_WD19_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD18_WCLK_posedge,
                            TmDt_WD18_WCLK_posedge,
                            WD18_ipd, "WD18",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD18_WCLK_posedge_posedge,
                            tsetup_WD18_WCLK_negedge_posedge,
                            thold_WD18_WCLK_posedge_posedge,
                            thold_WD18_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD17_WCLK_posedge,
                            TmDt_WD17_WCLK_posedge,
                            WD17_ipd, "WD17",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD17_WCLK_posedge_posedge,
                            tsetup_WD17_WCLK_negedge_posedge,
                            thold_WD17_WCLK_posedge_posedge,
                            thold_WD17_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD16_WCLK_posedge,
                            TmDt_WD16_WCLK_posedge,
                            WD16_ipd, "WD16",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD16_WCLK_posedge_posedge,
                            tsetup_WD16_WCLK_negedge_posedge,
                            thold_WD16_WCLK_posedge_posedge,
                            thold_WD16_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD15_WCLK_posedge,
                            TmDt_WD15_WCLK_posedge,
                            WD15_ipd, "WD15",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD15_WCLK_posedge_posedge,
                            tsetup_WD15_WCLK_negedge_posedge,
                            thold_WD15_WCLK_posedge_posedge,
                            thold_WD15_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD14_WCLK_posedge,
                            TmDt_WD14_WCLK_posedge,
                            WD14_ipd, "WD14",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD14_WCLK_posedge_posedge,
                            tsetup_WD14_WCLK_negedge_posedge,
                            thold_WD14_WCLK_posedge_posedge,
                            thold_WD14_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD13_WCLK_posedge,
                            TmDt_WD13_WCLK_posedge,
                            WD13_ipd, "WD13",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD13_WCLK_posedge_posedge,
                            tsetup_WD13_WCLK_negedge_posedge,
                            thold_WD13_WCLK_posedge_posedge,
                            thold_WD13_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD12_WCLK_posedge,
                            TmDt_WD12_WCLK_posedge,
                            WD12_ipd, "WD12",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD12_WCLK_posedge_posedge,
                            tsetup_WD12_WCLK_negedge_posedge,
                            thold_WD12_WCLK_posedge_posedge,
                            thold_WD12_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD11_WCLK_posedge,
                            TmDt_WD11_WCLK_posedge,
                            WD11_ipd, "WD11",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD11_WCLK_posedge_posedge,
                            tsetup_WD11_WCLK_negedge_posedge,
                            thold_WD11_WCLK_posedge_posedge,
                            thold_WD11_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD10_WCLK_posedge,
                            TmDt_WD10_WCLK_posedge,
                            WD10_ipd, "WD10",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD10_WCLK_posedge_posedge,
                            tsetup_WD10_WCLK_negedge_posedge,
                            thold_WD10_WCLK_posedge_posedge,
                            thold_WD10_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD9_WCLK_posedge,
                            TmDt_WD9_WCLK_posedge,
                            WD9_ipd, "WD9",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD9_WCLK_posedge_posedge,
                            tsetup_WD9_WCLK_negedge_posedge,
                            thold_WD9_WCLK_posedge_posedge,
                            thold_WD9_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD8_WCLK_posedge,
                            TmDt_WD8_WCLK_posedge,
                            WD8_ipd, "WD8",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD8_WCLK_posedge_posedge,
                            tsetup_WD8_WCLK_negedge_posedge,
                            thold_WD8_WCLK_posedge_posedge,
                            thold_WD8_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD7_WCLK_posedge,
                            TmDt_WD7_WCLK_posedge,
                            WD7_ipd, "WD7",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD7_WCLK_posedge_posedge,
                            tsetup_WD7_WCLK_negedge_posedge,
                            thold_WD7_WCLK_posedge_posedge,
                            thold_WD7_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD6_WCLK_posedge,
                            TmDt_WD6_WCLK_posedge,
                            WD6_ipd, "WD6",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD6_WCLK_posedge_posedge,
                            tsetup_WD6_WCLK_negedge_posedge,
                            thold_WD6_WCLK_posedge_posedge,
                            thold_WD6_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD5_WCLK_posedge,
                            TmDt_WD5_WCLK_posedge,
                            WD5_ipd, "WD5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD5_WCLK_posedge_posedge,
                            tsetup_WD5_WCLK_negedge_posedge,
                            thold_WD5_WCLK_posedge_posedge,
                            thold_WD5_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD4_WCLK_posedge,
                            TmDt_WD4_WCLK_posedge,
                            WD4_ipd, "WD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD4_WCLK_posedge_posedge,
                            tsetup_WD4_WCLK_negedge_posedge,
                            thold_WD4_WCLK_posedge_posedge,
                            thold_WD4_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD3_WCLK_posedge,
                            TmDt_WD3_WCLK_posedge,
                            WD3_ipd, "WD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD3_WCLK_posedge_posedge,
                            tsetup_WD3_WCLK_negedge_posedge,
                            thold_WD3_WCLK_posedge_posedge,
                            thold_WD3_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD2_WCLK_posedge,
                            TmDt_WD2_WCLK_posedge,
                            WD2_ipd, "WD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD2_WCLK_posedge_posedge,
                            tsetup_WD2_WCLK_negedge_posedge,
                            thold_WD2_WCLK_posedge_posedge,
                            thold_WD2_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD1_WCLK_posedge,
                            TmDt_WD1_WCLK_posedge,
                            WD1_ipd, "WD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD1_WCLK_posedge_posedge,
                            tsetup_WD1_WCLK_negedge_posedge,
                            thold_WD1_WCLK_posedge_posedge,
                            thold_WD1_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WD0_WCLK_posedge,
                            TmDt_WD0_WCLK_posedge,
                            WD0_ipd, "WD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD0_WCLK_posedge_posedge,
                            tsetup_WD0_WCLK_negedge_posedge,
                            thold_WD0_WCLK_posedge_posedge,
                            thold_WD0_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup WW high or low before WCLK rising
      --   Hold  WW high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WW2_WCLK_posedge,
                            TmDt_WW2_WCLK_posedge,
                            WW2_ipd, "WW2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WW2_WCLK_posedge_posedge,
                            tsetup_WW2_WCLK_negedge_posedge,
                            thold_WW2_WCLK_posedge_posedge,
                            thold_WW2_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WW1_WCLK_posedge,
                            TmDt_WW1_WCLK_posedge,
                            WW1_ipd, "WW1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WW1_WCLK_posedge_posedge,
                            tsetup_WW1_WCLK_negedge_posedge,
                            thold_WW1_WCLK_posedge_posedge,
                            thold_WW1_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      VitalSetupHoldCheck ( Tviol_WW0_WCLK_posedge,
                            TmDt_WW0_WCLK_posedge,
                            WW0_ipd, "WW0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WW0_WCLK_posedge_posedge,
                            tsetup_WW0_WCLK_negedge_posedge,
                            thold_WW0_WCLK_posedge_posedge,
                            thold_WW0_WCLK_negedge_posedge,
                            (To_X01(WEN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup WEN high before WCLK rising
      --   Hold  WEN high after WCLK rising

      VitalSetupHoldCheck ( Tviol_WEN_WCLK_posedge,
                            TmDt_WEN_WCLK_posedge,
                            WEN_ipd, "WEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WEN_WCLK_posedge_posedge,
                            tsetup_WEN_WCLK_negedge_posedge,
                            thold_WEN_WCLK_posedge_posedge,
                            thold_WEN_WCLK_negedge_posedge,
                            TimingCheckOn,
                            '/',
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM64K36P",
                            Xon,
                            MsgOn,
                            WARNING
                            );
    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################

      -- Decode Write Word Width
      if (TO_X01(WW2_delayed)='0' and TO_X01(WW1_delayed)='0' and TO_X01(WW0_delayed)='0') then
        WWIDTH := 1;
      elsif (TO_X01(WW2_delayed)='0' and TO_X01(WW1_delayed)='0' and TO_X01(WW0_delayed)='1') then
        WWIDTH := 2;
      elsif (TO_X01(WW2_delayed)='0' and TO_X01(WW1_delayed)='1' and TO_X01(WW0_delayed)='0') then
        WWIDTH := 4;
      elsif (TO_X01(WW2_delayed)='0' and TO_X01(WW1_delayed)='1' and TO_X01(WW0_delayed)='1') then
        WWIDTH := 9;
      elsif (TO_X01(WW2_delayed)='1' and TO_X01(WW1_delayed)='0' and TO_X01(WW0_delayed)='0') then
        WWIDTH := 18;
      elsif (TO_X01(WW2_delayed)='1' and TO_X01(WW1_delayed)='0' and TO_X01(WW0_delayed)='1') then
        WWIDTH := 36;
      else
	assert false
	report ": WW value invalid"
	severity Warning;
      end if;

      if (TO_X01(WCLK_ipd)='X') then
	if (TO_X01(WEN_delayed) /= '0') then
          if (TO_X01(WCLK_previous) /= 'X') then
	    assert false
	    report ": WCLK went unknown"
	    severity Warning;
	  end if;
	end if;
      elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='1')) then
	case (TO_X01(WEN_delayed)) is
	  when '0' =>
	    null;
	  when '1' =>

            -- Convert Write Address Signal to Integer
            if( INT(WRAD15_delayed) = -65537 ) then
              WADDR := -1;
            elsif( INT(WRAD14_delayed) = -65537 ) then
              WADDR := -1;
            else
              WADDR := ((INT(WRAD15_delayed)*32768)
                        +(INT(WRAD14_delayed)*16384)+(INT(WRAD13_delayed)*8192)+(INT(WRAD12_delayed)*4096)
                        +(INT(WRAD11_delayed)*2048)+(INT(WRAD10_delayed)*1024)+(INT(WRAD9_delayed)*512)
                        +(INT(WRAD8_delayed)*256)+(INT(WRAD7_delayed)*128)+(INT(WRAD6_delayed)*64)
                        +(INT(WRAD5_delayed)*32)+(INT(WRAD4_delayed)*16)+(INT(WRAD3_delayed)*8)
                        +(INT(WRAD2_delayed)*4)+(INT(WRAD1_delayed)*2)+(INT(WRAD0_delayed)));
            end if;

	    if (WADDR < 0) then
              if (TO_X01(WRAD15_delayed) = 'X' and WWIDTH = 1) then
                assert false
                report ": WRAD15 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD14_delayed) = 'X' and WWIDTH = 1) then
                assert false
                report ": WRAD14 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD13_delayed) = 'X' and WWIDTH = 1) then
                assert false
                report ": WRAD13 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD12_delayed) = 'X' and WWIDTH = 1) then
                assert false
                report ": WRAD12 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD11_delayed) = 'X' and WWIDTH = 1) then
                assert false
                report ": WRAD11 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD10_delayed) = 'X' and WWIDTH <= 2) then
                assert false
                report ": WRAD10 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD9_delayed) = 'X' and WWIDTH <= 4) then
                assert false
                report ": WRAD9 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD8_delayed) = 'X' and WWIDTH <= 9) then
                assert false
                report ": WRAD8 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD7_delayed) = 'X' and WWIDTH <= 18) then
                assert false
                report ": WRAD7 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD6_delayed) = 'X') then
                assert false
                report ": WRAD6 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD5_delayed) = 'X') then
                assert false
                report ": WRAD5 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD4_delayed) = 'X') then
                assert false
                report ": WRAD4 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD3_delayed) = 'X') then
                assert false
                report ": WRAD3 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD2_delayed) = 'X') then
                assert false
                report ": WRAD2 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD1_delayed) = 'X') then
                assert false
                report ": WRAD1 went unknown"
                severity Warning;
              end if;
              if (TO_X01(WRAD0_delayed) = 'X') then
                assert false
                report ": WRAD0 went unknown"
                severity Warning;
              end if;
	    else 
              case WWIDTH is
                when 1 => RAM_TMP(WADDR) := WD0_delayed ;
                when 2 => RAM_TMP(2*WADDR + 0) := WD0_delayed ;
                          RAM_TMP(2*WADDR + 1) := WD1_delayed ;
                when 4 => RAM_TMP(4*WADDR + 0) := WD0_delayed ;
                          RAM_TMP(4*WADDR + 1) := WD1_delayed ;
                          RAM_TMP(4*WADDR + 2) := WD2_delayed ;
                          RAM_TMP(4*WADDR + 3) := WD3_delayed ;
                when 9 => RAM_TMP(8*WADDR + 0) := WD0_delayed ;
                          RAM_TMP(8*WADDR + 1) := WD1_delayed ;
                          RAM_TMP(8*WADDR + 2) := WD2_delayed ;
                          RAM_TMP(8*WADDR + 3) := WD3_delayed ;
                          RAM_TMP(8*WADDR + 4) := WD4_delayed ;
                          RAM_TMP(8*WADDR + 5) := WD5_delayed ;
                          RAM_TMP(8*WADDR + 6) := WD6_delayed ;
                          RAM_TMP(8*WADDR + 7) := WD7_delayed ;
                          RAM_TMP9(WADDR) := WD8_delayed ;
                when 18 => RAM_TMP(16*WADDR + 0) := WD0_delayed ;
                           RAM_TMP(16*WADDR + 1) := WD1_delayed ;
                           RAM_TMP(16*WADDR + 2) := WD2_delayed ;
                           RAM_TMP(16*WADDR + 3) := WD3_delayed ;
                           RAM_TMP(16*WADDR + 4) := WD4_delayed ;
                           RAM_TMP(16*WADDR + 5) := WD5_delayed ;
                           RAM_TMP(16*WADDR + 6) := WD6_delayed ;
                           RAM_TMP(16*WADDR + 7) := WD7_delayed ;
                           RAM_TMP9((2*WADDR) + 0) := WD8_delayed ;
                           RAM_TMP(16*WADDR + 8) := WD9_delayed ;
                           RAM_TMP(16*WADDR + 9) := WD10_delayed ;
                           RAM_TMP(16*WADDR + 10) := WD11_delayed ;
                           RAM_TMP(16*WADDR + 11) := WD12_delayed ;
                           RAM_TMP(16*WADDR + 12) := WD13_delayed ;
                           RAM_TMP(16*WADDR + 13) := WD14_delayed ;
                           RAM_TMP(16*WADDR + 14) := WD15_delayed ;
                           RAM_TMP(16*WADDR + 15) := WD16_delayed ;
                           RAM_TMP9((2*WADDR) + 1) := WD17_delayed ;
                when 36 => RAM_TMP(32*WADDR + 0) := WD0_delayed ;
                           RAM_TMP(32*WADDR + 1) := WD1_delayed ;
                           RAM_TMP(32*WADDR + 2) := WD2_delayed ;
                           RAM_TMP(32*WADDR + 3) := WD3_delayed ;
                           RAM_TMP(32*WADDR + 4) := WD4_delayed ;
                           RAM_TMP(32*WADDR + 5) := WD5_delayed ;
                           RAM_TMP(32*WADDR + 6) := WD6_delayed ;
                           RAM_TMP(32*WADDR + 7) := WD7_delayed ;
                           RAM_TMP9((4*WADDR) + 0) := WD8_delayed ;
                           RAM_TMP(32*WADDR + 8) := WD9_delayed ;
                           RAM_TMP(32*WADDR + 9) := WD10_delayed ;
                           RAM_TMP(32*WADDR + 10) := WD11_delayed ;
                           RAM_TMP(32*WADDR + 11) := WD12_delayed ;
                           RAM_TMP(32*WADDR + 12) := WD13_delayed ;
                           RAM_TMP(32*WADDR + 13) := WD14_delayed ;
                           RAM_TMP(32*WADDR + 14) := WD15_delayed ;
                           RAM_TMP(32*WADDR + 15) := WD16_delayed ;
                           RAM_TMP9((4*WADDR) + 1) := WD17_delayed ;
                           RAM_TMP(32*WADDR + 16) := WD18_delayed ;
                           RAM_TMP(32*WADDR + 17) := WD19_delayed ;
                           RAM_TMP(32*WADDR + 18) := WD20_delayed ;
                           RAM_TMP(32*WADDR + 19) := WD21_delayed ;
                           RAM_TMP(32*WADDR + 20) := WD22_delayed ;
                           RAM_TMP(32*WADDR + 21) := WD23_delayed ;
                           RAM_TMP(32*WADDR + 22) := WD24_delayed ;
                           RAM_TMP(32*WADDR + 23) := WD25_delayed ;
                           RAM_TMP9((4*WADDR) + 2) := WD26_delayed ;
                           RAM_TMP(32*WADDR + 24) := WD27_delayed ;
                           RAM_TMP(32*WADDR + 25) := WD28_delayed ;
                           RAM_TMP(32*WADDR + 26) := WD29_delayed ;
                           RAM_TMP(32*WADDR + 27) := WD30_delayed ;
                           RAM_TMP(32*WADDR + 28) := WD31_delayed ;
                           RAM_TMP(32*WADDR + 29) := WD32_delayed ;
                           RAM_TMP(32*WADDR + 30) := WD33_delayed ;
                           RAM_TMP(32*WADDR + 31) := WD34_delayed ;
                           RAM_TMP9((4*WADDR ) + 3) := WD35_delayed ;
                when others => 
	          assert false
	          report ": WWIDTH value invalid"
	          severity Warning;
              end case;
	    end if;
	  when others =>
            assert false
            report ": WEN went unknown"
            severity Warning;
	end case;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      -- Decode Read Word Width
      if (TO_X01(RW2_delayed)='0' and TO_X01(RW1_delayed)='0' and TO_X01(RW0_delayed)='0') then
        RWIDTH := 1;
      elsif (TO_X01(RW2_delayed)='0' and TO_X01(RW1_delayed)='0' and TO_X01(RW0_delayed)='1') then
        RWIDTH := 2;
      elsif (TO_X01(RW2_delayed)='0' and TO_X01(RW1_delayed)='1' and TO_X01(RW0_delayed)='0') then
        RWIDTH := 4;
      elsif (TO_X01(RW2_delayed)='0' and TO_X01(RW1_delayed)='1' and TO_X01(RW0_delayed)='1') then
        RWIDTH := 9;
      elsif (TO_X01(RW2_delayed)='1' and TO_X01(RW1_delayed)='0' and TO_X01(RW0_delayed)='0') then
        RWIDTH := 18;
      elsif (TO_X01(RW2_delayed)='1' and TO_X01(RW1_delayed)='0' and TO_X01(RW0_delayed)='1') then
        RWIDTH := 36;
      else
        assert false
        report ": RW value invalid"
        severity Warning;
      end if;

      -- Convert Read Address Signal to Integer
      if (INT(RDAD15_delayed) = -65537) then
        RADDR := -1;
      elsif (INT(RDAD14_delayed) = -65537) then
        RADDR := -1;
      else
        RADDR := ((INT(RDAD15_delayed)*32768)
                 +(INT(RDAD14_delayed)*16384)+(INT(RDAD13_delayed)*8192)+(INT(RDAD12_delayed)*4096)
                 +(INT(RDAD11_delayed)*2048)+(INT(RDAD10_delayed)*1024)+(INT(RDAD9_delayed)*512)
                 +(INT(RDAD8_delayed)*256)+(INT(RDAD7_delayed)*128)+(INT(RDAD6_delayed)*64)
                 +(INT(RDAD5_delayed)*32)+(INT(RDAD4_delayed)*16)+(INT(RDAD3_delayed)*8)
                 +(INT(RDAD2_delayed)*4)+(INT(RDAD1_delayed)*2)+(INT(RDAD0_delayed)));
      end if;

      if (TO_X01(RCLK_ipd) = 'X') then
	case RWIDTH is
          when 1 => RD0_stg1 := 'X';
          when 2 => RD0_stg1 := 'X';
                    RD1_stg1 := 'X';
          when 4 => RD0_stg1 := 'X';
                    RD1_stg1 := 'X';
                    RD2_stg1 := 'X';
                    RD3_stg1 := 'X';
          when 9 => RD0_stg1 := 'X';
                    RD1_stg1 := 'X';
                    RD2_stg1 := 'X';
                    RD3_stg1 := 'X';
                    RD4_stg1 := 'X';
                    RD5_stg1 := 'X';
                    RD6_stg1 := 'X';
                    RD7_stg1 := 'X';
                    RD8_stg1 := 'X';
          when 18 => RD0_stg1 := 'X';
                     RD1_stg1 := 'X';
                     RD2_stg1 := 'X';
                     RD3_stg1 := 'X';
                     RD4_stg1 := 'X';
                     RD5_stg1 := 'X';
                     RD6_stg1 := 'X';
                     RD7_stg1 := 'X';
                     RD8_stg1 := 'X';
                     RD9_stg1 := 'X';
                     RD10_stg1 := 'X';
                     RD11_stg1 := 'X';
                     RD12_stg1 := 'X';
                     RD13_stg1 := 'X';
                     RD14_stg1 := 'X';
                     RD15_stg1 := 'X';
                     RD16_stg1 := 'X';
                     RD17_stg1 := 'X';
          when 36 => RD0_stg1 := 'X';
                     RD1_stg1 := 'X';
                     RD2_stg1 := 'X';
                     RD3_stg1 := 'X';
                     RD4_stg1 := 'X';
                     RD5_stg1 := 'X';
                     RD6_stg1 := 'X';
                     RD7_stg1 := 'X';
                     RD8_stg1 := 'X';
                     RD9_stg1 := 'X';
                     RD10_stg1 := 'X';
                     RD11_stg1 := 'X';
                     RD12_stg1 := 'X';
                     RD13_stg1 := 'X';
                     RD14_stg1 := 'X';
                     RD15_stg1 := 'X';
                     RD16_stg1 := 'X';
                     RD17_stg1 := 'X';
                     RD18_stg1 := 'X';
                     RD19_stg1 := 'X';
                     RD20_stg1 := 'X';
                     RD21_stg1 := 'X';
                     RD22_stg1 := 'X';
                     RD23_stg1 := 'X';
                     RD24_stg1 := 'X';
                     RD25_stg1 := 'X';
                     RD26_stg1 := 'X';
                     RD27_stg1 := 'X';
                     RD28_stg1 := 'X';
                     RD29_stg1 := 'X';
                     RD30_stg1 := 'X';
                     RD31_stg1 := 'X';
                     RD32_stg1 := 'X';
                     RD33_stg1 := 'X';
                     RD34_stg1 := 'X';
                     RD35_stg1 := 'X';
          when others => 
            assert false
            report ": RWIDTH value invalid"
            severity Warning;
        end case;
	if (TO_X01(RCLK_previous) /= 'X') then
	  assert false
	  report ": RCLK went unknown"
	  severity Warning;
	end if;
      elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '1')) then
	case (TO_X01(REN_stg1)) is
	  when '0' =>
                       assert true
                       report ": REN_stg1 low"
                       severity Note;
	  when '1' =>
            case RWIDTH is
              when 1 => RD0_zd := RD0_stg1;
              when 2 => RD0_zd := RD0_stg1;
                        RD1_zd := RD1_stg1;
              when 4 => RD0_zd := RD0_stg1;
                        RD1_zd := RD1_stg1;
                        RD2_zd := RD2_stg1;
                        RD3_zd := RD3_stg1;
              when 9 => RD0_zd := RD0_stg1;
                        RD1_zd := RD1_stg1;
                        RD2_zd := RD2_stg1;
                        RD3_zd := RD3_stg1;
                        RD4_zd := RD4_stg1;
                        RD5_zd := RD5_stg1;
                        RD6_zd := RD6_stg1;
                        RD7_zd := RD7_stg1;
                        RD8_zd := RD8_stg1;
             when 18 => RD0_zd := RD0_stg1;
                        RD1_zd := RD1_stg1;
                        RD2_zd := RD2_stg1;
                        RD3_zd := RD3_stg1;
                        RD4_zd := RD4_stg1;
                        RD5_zd := RD5_stg1;
                        RD6_zd := RD6_stg1;
                        RD7_zd := RD7_stg1;
                        RD8_zd := RD8_stg1;
                        RD9_zd := RD9_stg1;
                        RD10_zd := RD10_stg1;
                        RD11_zd := RD11_stg1;
                        RD12_zd := RD12_stg1;
                        RD13_zd := RD13_stg1;
                        RD14_zd := RD14_stg1;
                        RD15_zd := RD15_stg1;
                        RD16_zd := RD16_stg1;
                        RD17_zd := RD17_stg1;
             when 36 => RD0_zd := RD0_stg1;
                        RD1_zd := RD1_stg1;
                        RD2_zd := RD2_stg1;
                        RD3_zd := RD3_stg1;
                        RD4_zd := RD4_stg1;
                        RD5_zd := RD5_stg1;
                        RD6_zd := RD6_stg1;
                        RD7_zd := RD7_stg1;
                        RD8_zd := RD8_stg1;
                        RD9_zd := RD9_stg1;
                        RD10_zd := RD10_stg1;
                        RD11_zd := RD11_stg1;
                        RD12_zd := RD12_stg1;
                        RD13_zd := RD13_stg1;
                        RD14_zd := RD14_stg1;
                        RD15_zd := RD15_stg1;
                        RD16_zd := RD16_stg1;
                        RD17_zd := RD17_stg1;
                        RD18_zd := RD18_stg1;
                        RD19_zd := RD19_stg1;
                        RD20_zd := RD20_stg1;
                        RD21_zd := RD21_stg1;
                        RD22_zd := RD22_stg1;
                        RD23_zd := RD23_stg1;
                        RD24_zd := RD24_stg1;
                        RD25_zd := RD25_stg1;
                        RD26_zd := RD26_stg1;
                        RD27_zd := RD27_stg1;
                        RD28_zd := RD28_stg1;
                        RD29_zd := RD29_stg1;
                        RD30_zd := RD30_stg1;
                        RD31_zd := RD31_stg1;
                        RD32_zd := RD32_stg1;
                        RD33_zd := RD33_stg1;
                        RD34_zd := RD34_stg1;
                        RD35_zd := RD35_stg1;
             when others => 
	        assert false
	        report ": RWIDTH value invalid"
	        severity Warning;
            end case;
	  when others =>
            case RWIDTH is
              when 1 => 
                        RD0_zd := 'X';
              when 2 => 
                        RD0_zd := 'X';
                        RD1_zd := 'X';
              when 4 => 
                        RD0_zd := 'X';
                        RD1_zd := 'X';
                        RD2_zd := 'X';
                        RD3_zd := 'X';
              when 9 => 
                        RD0_zd := 'X';
                        RD1_zd := 'X';
                        RD2_zd := 'X';
                        RD3_zd := 'X';
                        RD4_zd := 'X';
                        RD5_zd := 'X';
                        RD6_zd := 'X';
                        RD7_zd := 'X';
                        RD8_zd := 'X';
              when 18 => 
                         RD0_zd := 'X';
                         RD1_zd := 'X';
                         RD2_zd := 'X';
                         RD3_zd := 'X';
                         RD4_zd := 'X';
                         RD5_zd := 'X';
                         RD6_zd := 'X';
                         RD7_zd := 'X';
                         RD8_zd := 'X';
                         RD9_zd := 'X';
                         RD10_zd := 'X';
                         RD11_zd := 'X';
                         RD12_zd := 'X';
                         RD13_zd := 'X';
                         RD14_zd := 'X';
                         RD15_zd := 'X';
                         RD16_zd := 'X';
                         RD17_zd := 'X';
              when 36 => 
                         RD0_zd := 'X';
                         RD1_zd := 'X';
                         RD2_zd := 'X';
                         RD3_zd := 'X';
                         RD4_zd := 'X';
                         RD5_zd := 'X';
                         RD6_zd := 'X';
                         RD7_zd := 'X';
                         RD8_zd := 'X';
                         RD9_zd := 'X';
                         RD10_zd := 'X';
                         RD11_zd := 'X';
                         RD12_zd := 'X';
                         RD13_zd := 'X';
                         RD14_zd := 'X';
                         RD15_zd := 'X';
                         RD16_zd := 'X';
                         RD17_zd := 'X';
                         RD18_zd := 'X';
                         RD19_zd := 'X';
                         RD20_zd := 'X';
                         RD21_zd := 'X';
                         RD22_zd := 'X';
                         RD23_zd := 'X';
                         RD24_zd := 'X';
                         RD25_zd := 'X';
                         RD26_zd := 'X';
                         RD27_zd := 'X';
                         RD28_zd := 'X';
                         RD29_zd := 'X';
                         RD30_zd := 'X';
                         RD31_zd := 'X';
                         RD32_zd := 'X';
                         RD33_zd := 'X';
                         RD34_zd := 'X';
                         RD35_zd := 'X';
              when others => 
	        assert false
	        report ": RWIDTH value invalid"
	        severity Warning;
            end case;
	end case; --REN_stg1
	case (TO_X01(REN_delayed)) is
	  when '0' =>
                       assert true
                       report ": REN low"
                       severity Note;
	  when '1' =>
	    if (RADDR < 0) then
              case RWIDTH is
                when 1 => RD0_stg1 := 'X';
                when 2 => RD0_stg1 := 'X';
                          RD1_stg1 := 'X';
                when 4 => RD0_stg1 := 'X';
                          RD1_stg1 := 'X';
                          RD2_stg1 := 'X';
                          RD3_stg1 := 'X';
                when 9 => RD0_stg1 := 'X';
                          RD1_stg1 := 'X';
                          RD2_stg1 := 'X';
                          RD3_stg1 := 'X';
                          RD4_stg1 := 'X';
                          RD5_stg1 := 'X';
                          RD6_stg1 := 'X';
                          RD7_stg1 := 'X';
                          RD8_stg1 := 'X';
                when 18 => RD0_stg1 := 'X';
                           RD1_stg1 := 'X';
                           RD2_stg1 := 'X';
                           RD3_stg1 := 'X';
                           RD4_stg1 := 'X';
                           RD5_stg1 := 'X';
                           RD6_stg1 := 'X';
                           RD7_stg1 := 'X';
                           RD8_stg1 := 'X';
                           RD9_stg1 := 'X';
                           RD10_stg1 := 'X';
                           RD11_stg1 := 'X';
                           RD12_stg1 := 'X';
                           RD13_stg1 := 'X';
                           RD14_stg1 := 'X';
                           RD15_stg1 := 'X';
                           RD16_stg1 := 'X';
                           RD17_stg1 := 'X';
                when 36 => RD0_stg1 := 'X';
                           RD1_stg1 := 'X';
                           RD2_stg1 := 'X';
                           RD3_stg1 := 'X';
                           RD4_stg1 := 'X';
                           RD5_stg1 := 'X';
                           RD6_stg1 := 'X';
                           RD7_stg1 := 'X';
                           RD8_stg1 := 'X';
                           RD9_stg1 := 'X';
                           RD10_stg1 := 'X';
                           RD11_stg1 := 'X';
                           RD12_stg1 := 'X';
                           RD13_stg1 := 'X';
                           RD14_stg1 := 'X';
                           RD15_stg1 := 'X';
                           RD16_stg1 := 'X';
                           RD17_stg1 := 'X';
                           RD18_stg1 := 'X';
                           RD19_stg1 := 'X';
                           RD20_stg1 := 'X';
                           RD21_stg1 := 'X';
                           RD22_stg1 := 'X';
                           RD23_stg1 := 'X';
                           RD24_stg1 := 'X';
                           RD25_stg1 := 'X';
                           RD26_stg1 := 'X';
                           RD27_stg1 := 'X';
                           RD28_stg1 := 'X';
                           RD29_stg1 := 'X';
                           RD30_stg1 := 'X';
                           RD31_stg1 := 'X';
                           RD32_stg1 := 'X';
                           RD33_stg1 := 'X';
                           RD34_stg1 := 'X';
                           RD35_stg1 := 'X';
                when others => 
	          assert false
	          report ": RWIDTH value invalid"
	          severity Warning;
              end case;
	      if (TO_X01(RDAD15_delayed) = 'X') and (TO_X01(RDAD15_previous) /= 'X' and RWIDTH = 1) then
		assert false
		report ": RDAD15 went unknown"
		severity Warning;
                RDAD15_previous := RDAD15_delayed;
	      end if;
	      if (TO_X01(RDAD14_delayed) = 'X') and (TO_X01(RDAD14_previous) /= 'X' and RWIDTH = 1) then
		assert false
		report ": RDAD14 went unknown"
		severity Warning;
                RDAD14_previous := RDAD14_delayed;
	      end if;
	      if (TO_X01(RDAD13_delayed) = 'X') and (TO_X01(RDAD13_previous) /= 'X' and RWIDTH = 1) then
		assert false
		report ": RDAD13 went unknown"
		severity Warning;
                RDAD13_previous := RDAD13_delayed;
	      end if;
	      if (TO_X01(RDAD12_delayed) = 'X') and (TO_X01(RDAD12_previous) /= 'X' and RWIDTH = 1) then
		assert false
		report ": RDAD12 went unknown"
		severity Warning;
                RDAD12_previous := RDAD12_delayed;
	      end if;
	      if (TO_X01(RDAD11_delayed) = 'X') and (TO_X01(RDAD11_previous) /= 'X' and RWIDTH = 1) then
		assert false
		report ": RDAD11 went unknown"
		severity Warning;
                RDAD11_previous := RDAD11_delayed;
	      end if;
	      if (TO_X01(RDAD10_delayed) = 'X') and (TO_X01(RDAD10_previous) /= 'X' and RWIDTH <= 2) then
		assert false
		report ": RDAD10 went unknown"
		severity Warning;
                RDAD10_previous := RDAD10_delayed;
	      end if;
	      if (TO_X01(RDAD9_delayed) = 'X') and (TO_X01(RDAD9_previous) /= 'X' and RWIDTH <= 4) then
		assert false
		report ": RDAD9 went unknown"
		severity Warning;
                RDAD9_previous := RDAD9_delayed;
	      end if;
	      if (TO_X01(RDAD8_delayed) = 'X') and (TO_X01(RDAD8_previous) /= 'X' and RWIDTH <= 9) then
		assert false
		report ": RDAD8 went unknown"
		severity Warning;
                RDAD8_previous := RDAD8_delayed;
	      end if;
	      if (TO_X01(RDAD7_delayed) = 'X') and (TO_X01(RDAD7_previous) /= 'X' and RWIDTH <= 18) then
		assert false
		report ": RDAD7 went unknown"
		severity Warning;
                RDAD7_previous := RDAD7_delayed;
	      end if;
	      if (TO_X01(RDAD6_delayed) = 'X') and (TO_X01(RDAD6_previous) /= 'X') then
		assert false
		report ": RDAD6 went unknown"
		severity Warning;
                RDAD6_previous := RDAD6_delayed;
	      end if;
	      if (TO_X01(RDAD5_delayed) = 'X') and (TO_X01(RDAD5_previous) /= 'X') then
		assert false
		report ": RDAD5 went unknown"
		severity Warning;
                RDAD5_previous := RDAD5_delayed;
	      end if;
	      if (TO_X01(RDAD4_delayed) = 'X') and (TO_X01(RDAD4_previous) /= 'X') then
		assert false
		report ": RDAD4 went unknown"
		severity Warning;
                RDAD4_previous := RDAD4_delayed;
	      end if;
	      if (TO_X01(RDAD3_delayed) = 'X') and (TO_X01(RDAD3_previous) /= 'X') then
		assert false
		report ": RDAD3 went unknown"
		severity Warning;
                RDAD3_previous := RDAD3_delayed;
	      end if;
	      if (TO_X01(RDAD2_delayed) = 'X') and (TO_X01(RDAD2_previous) /= 'X') then
		assert false
		report ": RDAD2 went unknown"
		severity Warning;
                RDAD2_previous := RDAD2_delayed;
	      end if;
	      if (TO_X01(RDAD1_delayed) = 'X') and (TO_X01(RDAD1_previous) /= 'X') then
		assert false
		report ": RDAD1 went unknown"
		severity Warning;
                RDAD1_previous := RDAD1_delayed;
	      end if;
	      if (TO_X01(RDAD0_delayed) = 'X') and (TO_X01(RDAD0_previous) /= 'X') then
		assert false
		report ": RDAD0 went unknown"
		severity Warning;
                RDAD0_previous := RDAD0_delayed;
	      end if;
	    else
              case RWIDTH is
                when 1 => RD0_stg1 := RAM_TMP(RADDR) ;
                when 2 => RD0_stg1 := RAM_TMP(2*RADDR + 0) ;
                          RD1_stg1 := RAM_TMP(2*RADDR + 1) ;
                when 4 => RD0_stg1 := RAM_TMP(4*RADDR + 0) ;
                          RD1_stg1 := RAM_TMP(4*RADDR + 1) ;
                          RD2_stg1 := RAM_TMP(4*RADDR + 2) ;
                          RD3_stg1 := RAM_TMP(4*RADDR + 3) ;
                when 9 => RD0_stg1 := RAM_TMP(8*RADDR + 0) ;
                          RD1_stg1 := RAM_TMP(8*RADDR + 1) ;
                          RD2_stg1 := RAM_TMP(8*RADDR + 2) ;
                          RD3_stg1 := RAM_TMP(8*RADDR + 3) ;
                          RD4_stg1 := RAM_TMP(8*RADDR + 4) ;
                          RD5_stg1 := RAM_TMP(8*RADDR + 5) ;
                          RD6_stg1 := RAM_TMP(8*RADDR + 6) ;
                          RD7_stg1 := RAM_TMP(8*RADDR + 7) ;
                          RD8_stg1 := RAM_TMP9(RADDR) ;
                when 18 => RD0_stg1 := RAM_TMP(16*RADDR + 0) ;
                           RD1_stg1 := RAM_TMP(16*RADDR + 1) ;
                           RD2_stg1 := RAM_TMP(16*RADDR + 2) ;
                           RD3_stg1 := RAM_TMP(16*RADDR + 3) ;
                           RD4_stg1 := RAM_TMP(16*RADDR + 4) ;
                           RD5_stg1 := RAM_TMP(16*RADDR + 5) ;
                           RD6_stg1 := RAM_TMP(16*RADDR + 6) ;
                           RD7_stg1 := RAM_TMP(16*RADDR + 7) ;
                           RD8_stg1 := RAM_TMP9((2*RADDR) + 0) ;
                           RD9_stg1 := RAM_TMP(16*RADDR + 8) ;
                           RD10_stg1 := RAM_TMP(16*RADDR + 9) ;
                           RD11_stg1 := RAM_TMP(16*RADDR + 10) ;
                           RD12_stg1 := RAM_TMP(16*RADDR + 11) ;
                           RD13_stg1 := RAM_TMP(16*RADDR + 12) ;
                           RD14_stg1 := RAM_TMP(16*RADDR + 13) ;
                           RD15_stg1 := RAM_TMP(16*RADDR + 14) ;
                           RD16_stg1 := RAM_TMP(16*RADDR + 15) ;
                           RD17_stg1 := RAM_TMP9((2*RADDR) + 1) ;
                when 36 => RD0_stg1 := RAM_TMP(32*RADDR + 0) ;
                           RD1_stg1 := RAM_TMP(32*RADDR + 1) ;
                           RD2_stg1 := RAM_TMP(32*RADDR + 2) ;
                           RD3_stg1 := RAM_TMP(32*RADDR + 3) ;
                           RD4_stg1 := RAM_TMP(32*RADDR + 4) ;
                           RD5_stg1 := RAM_TMP(32*RADDR + 5) ;
                           RD6_stg1 := RAM_TMP(32*RADDR + 6) ;
                           RD7_stg1 := RAM_TMP(32*RADDR + 7) ;
                           RD8_stg1 := RAM_TMP9((4*RADDR) + 0) ;
                           RD9_stg1 := RAM_TMP(32*RADDR + 8) ;
                           RD10_stg1 := RAM_TMP(32*RADDR + 9) ;
                           RD11_stg1 := RAM_TMP(32*RADDR + 10) ;
                           RD12_stg1 := RAM_TMP(32*RADDR + 11) ;
                           RD13_stg1 := RAM_TMP(32*RADDR + 12) ;
                           RD14_stg1 := RAM_TMP(32*RADDR + 13) ;
                           RD15_stg1 := RAM_TMP(32*RADDR + 14) ;
                           RD16_stg1 := RAM_TMP(32*RADDR + 15) ;
                           RD17_stg1 := RAM_TMP9((4*RADDR) + 1) ;
                           RD18_stg1 := RAM_TMP(32*RADDR + 16) ;
                           RD19_stg1 := RAM_TMP(32*RADDR + 17) ;
                           RD20_stg1 := RAM_TMP(32*RADDR + 18) ;
                           RD21_stg1 := RAM_TMP(32*RADDR + 19) ;
                           RD22_stg1 := RAM_TMP(32*RADDR + 20) ;
                           RD23_stg1 := RAM_TMP(32*RADDR + 21) ;
                           RD24_stg1 := RAM_TMP(32*RADDR + 22) ;
                           RD25_stg1 := RAM_TMP(32*RADDR + 23) ;
                           RD26_stg1 := RAM_TMP9((4*RADDR ) + 2) ;
                           RD27_stg1 := RAM_TMP(32*RADDR + 24) ;
                           RD28_stg1 := RAM_TMP(32*RADDR + 25) ;
                           RD29_stg1 := RAM_TMP(32*RADDR + 26) ;
                           RD30_stg1 := RAM_TMP(32*RADDR + 27) ;
                           RD31_stg1 := RAM_TMP(32*RADDR + 28) ;
                           RD32_stg1 := RAM_TMP(32*RADDR + 29) ;
                           RD33_stg1 := RAM_TMP(32*RADDR + 30) ;
                           RD34_stg1 := RAM_TMP(32*RADDR + 31) ;
                           RD35_stg1 := RAM_TMP9((4*RADDR) + 3) ;
                when others => 
	          assert false
	          report ": RWIDTH value invalid"
	          severity Warning;
              end case;
	    end if;
	  when others =>
            case RWIDTH is
              when 1 => 
                        RD0_stg1 := 'X';
              when 2 => 
                        RD0_stg1 := 'X';
                        RD1_stg1 := 'X';
              when 4 => 
                        RD0_stg1 := 'X';
                        RD1_stg1 := 'X';
                        RD2_stg1 := 'X';
                        RD3_stg1 := 'X';
              when 9 => 
                        RD0_stg1 := 'X';
                        RD1_stg1 := 'X';
                        RD2_stg1 := 'X';
                        RD3_stg1 := 'X';
                        RD4_stg1 := 'X';
                        RD5_stg1 := 'X';
                        RD6_stg1 := 'X';
                        RD7_stg1 := 'X';
                        RD8_stg1 := 'X';
              when 18 => 
                         RD0_stg1 := 'X';
                         RD1_stg1 := 'X';
                         RD2_stg1 := 'X';
                         RD3_stg1 := 'X';
                         RD4_stg1 := 'X';
                         RD5_stg1 := 'X';
                         RD6_stg1 := 'X';
                         RD7_stg1 := 'X';
                         RD8_stg1 := 'X';
                         RD9_stg1 := 'X';
                         RD10_stg1 := 'X';
                         RD11_stg1 := 'X';
                         RD12_stg1 := 'X';
                         RD13_stg1 := 'X';
                         RD14_stg1 := 'X';
                         RD15_stg1 := 'X';
                         RD16_stg1 := 'X';
                         RD17_stg1 := 'X';
              when 36 => 
                         RD0_stg1 := 'X';
                         RD1_stg1 := 'X';
                         RD2_stg1 := 'X';
                         RD3_stg1 := 'X';
                         RD4_stg1 := 'X';
                         RD5_stg1 := 'X';
                         RD6_stg1 := 'X';
                         RD7_stg1 := 'X';
                         RD8_stg1 := 'X';
                         RD9_stg1 := 'X';
                         RD10_stg1 := 'X';
                         RD11_stg1 := 'X';
                         RD12_stg1 := 'X';
                         RD13_stg1 := 'X';
                         RD14_stg1 := 'X';
                         RD15_stg1 := 'X';
                         RD16_stg1 := 'X';
                         RD17_stg1 := 'X';
                         RD18_stg1 := 'X';
                         RD19_stg1 := 'X';
                         RD20_stg1 := 'X';
                         RD21_stg1 := 'X';
                         RD22_stg1 := 'X';
                         RD23_stg1 := 'X';
                         RD24_stg1 := 'X';
                         RD25_stg1 := 'X';
                         RD26_stg1 := 'X';
                         RD27_stg1 := 'X';
                         RD28_stg1 := 'X';
                         RD29_stg1 := 'X';
                         RD30_stg1 := 'X';
                         RD31_stg1 := 'X';
                         RD32_stg1 := 'X';
                         RD33_stg1 := 'X';
                         RD34_stg1 := 'X';
                         RD35_stg1 := 'X';
              when others => 
	        assert false
	        report ": RWIDTH value invalid"
	        severity Warning;
            end case;
            if (TO_X01(REN_delayed) = 'X') and (TO_X01(REN_previous) /= 'X') then
	      assert false
	      report ": REN went unknown"
	      severity Warning;
              REN_previous := REN_delayed;
            end if;
	end case; -- REN
        REN_stg1 := REN_delayed;
      end if; -- Rising RCLK edge

      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      WW2_delayed := WW2_ipd;
      WW1_delayed := WW1_ipd;
      WW0_delayed := WW0_ipd;
      WEN_delayed := WEN_ipd;
      if RW2_ipd'event then
        RW2_previous := RW2_delayed;
        RW2_delayed := RW2_ipd;
      end if;
      if RW1_ipd'event then
        RW1_previous := RW1_delayed;
        RW1_delayed := RW1_ipd;
      end if;
      if RW0_ipd'event then
        RW0_previous := RW0_delayed;
        RW0_delayed := RW0_ipd;
      end if;
      if REN_ipd'event then
        REN_previous := REN_delayed;
        REN_delayed := REN_ipd;
      end if;
      WD35_delayed := WD35_ipd;
      WD34_delayed := WD34_ipd;
      WD33_delayed := WD33_ipd;
      WD32_delayed := WD32_ipd;
      WD31_delayed := WD31_ipd;
      WD30_delayed := WD30_ipd;
      WD29_delayed := WD29_ipd;
      WD28_delayed := WD28_ipd;
      WD27_delayed := WD27_ipd;
      WD26_delayed := WD26_ipd;
      WD25_delayed := WD25_ipd;
      WD24_delayed := WD24_ipd;
      WD23_delayed := WD23_ipd;
      WD22_delayed := WD22_ipd;
      WD21_delayed := WD21_ipd;
      WD20_delayed := WD20_ipd;
      WD19_delayed := WD19_ipd;
      WD18_delayed := WD18_ipd;
      WD17_delayed := WD17_ipd;
      WD16_delayed := WD16_ipd;
      WD15_delayed := WD15_ipd;
      WD14_delayed := WD14_ipd;
      WD13_delayed := WD13_ipd;
      WD12_delayed := WD12_ipd;
      WD11_delayed := WD11_ipd;
      WD10_delayed := WD10_ipd;
      WD9_delayed := WD9_ipd;
      WD8_delayed := WD8_ipd;
      WD7_delayed := WD7_ipd;
      WD6_delayed := WD6_ipd;
      WD5_delayed := WD5_ipd;
      WD4_delayed := WD4_ipd;
      WD3_delayed := WD3_ipd;
      WD2_delayed := WD2_ipd;
      WD1_delayed := WD1_ipd;
      WD0_delayed := WD0_ipd;
      WRAD15_delayed := WRAD15_ipd;
      WRAD14_delayed := WRAD14_ipd;
      WRAD13_delayed := WRAD13_ipd;
      WRAD12_delayed := WRAD12_ipd;
      WRAD11_delayed := WRAD11_ipd;
      WRAD10_delayed := WRAD10_ipd;
      WRAD9_delayed := WRAD9_ipd;
      WRAD8_delayed := WRAD8_ipd;
      WRAD7_delayed := WRAD7_ipd;
      WRAD6_delayed := WRAD6_ipd;
      WRAD5_delayed := WRAD5_ipd;
      WRAD4_delayed := WRAD4_ipd;
      WRAD3_delayed := WRAD3_ipd;
      WRAD2_delayed := WRAD2_ipd;
      WRAD1_delayed := WRAD1_ipd;
      WRAD0_delayed := WRAD0_ipd;
      if RDAD15_ipd'event then
        RDAD15_previous := RDAD15_delayed;
        RDAD15_delayed := RDAD15_ipd;
      end if;
      if RDAD14_ipd'event then
        RDAD14_previous := RDAD14_delayed;
        RDAD14_delayed := RDAD14_ipd;
      end if;
      if RDAD13_ipd'event then
        RDAD13_previous := RDAD13_delayed;
        RDAD13_delayed := RDAD13_ipd;
      end if;
      if RDAD12_ipd'event then
        RDAD12_previous := RDAD12_delayed;
        RDAD12_delayed := RDAD12_ipd;
      end if;
      if RDAD11_ipd'event then
        RDAD11_previous := RDAD11_delayed;
        RDAD11_delayed := RDAD11_ipd;
      end if;
      if RDAD10_ipd'event then
        RDAD10_previous := RDAD10_delayed;
        RDAD10_delayed := RDAD10_ipd;
      end if;
      if RDAD9_ipd'event then
        RDAD9_previous := RDAD9_delayed;
        RDAD9_delayed := RDAD9_ipd;
      end if;
      if RDAD8_ipd'event then
        RDAD8_previous := RDAD8_delayed;
        RDAD8_delayed := RDAD8_ipd;
      end if;
      if RDAD7_ipd'event then
        RDAD7_previous := RDAD7_delayed;
        RDAD7_delayed := RDAD7_ipd;
      end if;
      if RDAD6_ipd'event then
        RDAD6_previous := RDAD6_delayed;
        RDAD6_delayed := RDAD6_ipd;
      end if;
      if RDAD5_ipd'event then
        RDAD5_previous := RDAD5_delayed;
        RDAD5_delayed := RDAD5_ipd;
      end if;
      if RDAD4_ipd'event then
        RDAD4_previous := RDAD4_delayed;
        RDAD4_delayed := RDAD4_ipd;
      end if;
      if RDAD3_ipd'event then
        RDAD3_previous := RDAD3_delayed;
        RDAD3_delayed := RDAD3_ipd;
      end if;
      if RDAD2_ipd'event then
        RDAD2_previous := RDAD2_delayed;
        RDAD2_delayed := RDAD2_ipd;
      end if;
      if RDAD1_ipd'event then
        RDAD1_previous := RDAD1_delayed;
      end if;
        RDAD1_delayed := RDAD1_ipd;
      if RDAD0_ipd'event then
        RDAD0_previous := RDAD0_delayed;
        RDAD0_delayed := RDAD0_ipd;
      end if;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => RD35,
	GlitchData => RD35_GlitchData,
	OutSignalName => "RD35",
	OutTemp => RD35_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD35), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => Xon,
	MsgOn => MsgOn,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
        OutSignal => RD34,
        GlitchData => RD34_GlitchData,
        OutSignalName => "RD34",
        OutTemp => RD34_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD34), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD33,
        GlitchData => RD33_GlitchData,
        OutSignalName => "RD33",
        OutTemp => RD33_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD33), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD32,
        GlitchData => RD32_GlitchData,
        OutSignalName => "RD32",
        OutTemp => RD32_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD32), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD31,
        GlitchData => RD31_GlitchData,
        OutSignalName => "RD31",
        OutTemp => RD31_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD31), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD30,
        GlitchData => RD30_GlitchData,
        OutSignalName => "RD30",
        OutTemp => RD30_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD30), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD29,
        GlitchData => RD29_GlitchData,
        OutSignalName => "RD29",
        OutTemp => RD29_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD29), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD28,
        GlitchData => RD28_GlitchData,
        OutSignalName => "RD28",
        OutTemp => RD28_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD28), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD27,
        GlitchData => RD27_GlitchData,
        OutSignalName => "RD27",
        OutTemp => RD27_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD27), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD26,
        GlitchData => RD26_GlitchData,
        OutSignalName => "RD26",
        OutTemp => RD26_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD26), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD25,
        GlitchData => RD25_GlitchData,
        OutSignalName => "RD25",
        OutTemp => RD25_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD25), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD24,
        GlitchData => RD24_GlitchData,
        OutSignalName => "RD24",
        OutTemp => RD24_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD24), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD23,
        GlitchData => RD23_GlitchData,
        OutSignalName => "RD23",
        OutTemp => RD23_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD23), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD22,
        GlitchData => RD22_GlitchData,
        OutSignalName => "RD22",
        OutTemp => RD22_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD22), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD21,
        GlitchData => RD21_GlitchData,
        OutSignalName => "RD21",
        OutTemp => RD21_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD21), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD20,
        GlitchData => RD20_GlitchData,
        OutSignalName => "RD20",
        OutTemp => RD20_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD20), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD19,
        GlitchData => RD19_GlitchData,
        OutSignalName => "RD19",
        OutTemp => RD19_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD19), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD18,
        GlitchData => RD18_GlitchData,
        OutSignalName => "RD18",
        OutTemp => RD18_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD18), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD17,
        GlitchData => RD17_GlitchData,
        OutSignalName => "RD17",
        OutTemp => RD17_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD17), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD16,
        GlitchData => RD16_GlitchData,
        OutSignalName => "RD16",
        OutTemp => RD16_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD16), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD15,
        GlitchData => RD15_GlitchData,
        OutSignalName => "RD15",
        OutTemp => RD15_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD15), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD14,
        GlitchData => RD14_GlitchData,
        OutSignalName => "RD14",
        OutTemp => RD14_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD14), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD13,
        GlitchData => RD13_GlitchData,
        OutSignalName => "RD13",
        OutTemp => RD13_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD13), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD12,
        GlitchData => RD12_GlitchData,
        OutSignalName => "RD12",
        OutTemp => RD12_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD12), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD11,
        GlitchData => RD11_GlitchData,
        OutSignalName => "RD11",
        OutTemp => RD11_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD11), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD10,
        GlitchData => RD10_GlitchData,
        OutSignalName => "RD10",
        OutTemp => RD10_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD10), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD9,
        GlitchData => RD9_GlitchData,
        OutSignalName => "RD9",
        OutTemp => RD9_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD9), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD8,
        GlitchData => RD8_GlitchData,
        OutSignalName => "RD8",
        OutTemp => RD8_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD8), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD7,
        GlitchData => RD7_GlitchData,
        OutSignalName => "RD7",
        OutTemp => RD7_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD7), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD6,
        GlitchData => RD6_GlitchData,
        OutSignalName => "RD6",
        OutTemp => RD6_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD6), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD5,
        GlitchData => RD5_GlitchData,
        OutSignalName => "RD5",
        OutTemp => RD5_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD5), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD4,
        GlitchData => RD4_GlitchData,
        OutSignalName => "RD4",
        OutTemp => RD4_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD4), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD3,
        GlitchData => RD3_GlitchData,
        OutSignalName => "RD3",
        OutTemp => RD3_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD3), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD2,
        GlitchData => RD2_GlitchData,
        OutSignalName => "RD2",
        OutTemp => RD2_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD2), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD1,
        GlitchData => RD1_GlitchData,
        OutSignalName => "RD1",
        OutTemp => RD1_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD1), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );

    VitalPathDelay01Z (
        OutSignal => RD0,
        GlitchData => RD0_GlitchData,
        OutSignalName => "RD0",
        OutTemp => RD0_zd,
        Paths => (0 => (RCLK_ipd'last_event,
                        VitalExtendToFillDelay(tpd_RCLK_RD0), TRUE)
                 ),
        DefaultDelay => VitalZeroDelay01Z,
        Mode => Onevent,
        XON => Xon,
        MsgOn => MsgOn,
        MsgSeverity => WARNING
        );
    
  end process VITALBehavior;

end VITAL_ACT;

configuration CFG_RAM64K36P_VITAL of RAM64K36P is
   for VITAL_ACT
   end for;
end CFG_RAM64K36P_VITAL;

----- CELL PLL -----
-- 
-- Actel AX family PLL VITAL simulation model.
--
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

-- entity declaration --
entity PLL is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;

      f_REFCLK_LOCK          :	Integer := 3; -- Number of REFCLK pulses after which LOCK is raised

      tipd_PWRDWN            :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_REFCLK            :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_LOWFREQ           :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OSC2              :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OSC1              :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OSC0              :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI5             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI4             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI3             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI2             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI1             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI0             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ5             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ4             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ3             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ2             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ1             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ0             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE4        :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE3        :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE2        :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE1        :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE0        :  VitalDelayType01 := (0.000 ns, 0.000 ns);

      tpd_REFCLK_CLK1        :  VitalDelayType01 := (0.000 ns, 0.000 ns); -- unused
      tpd_REFCLK_CLK2        :  VitalDelayType01 := (0.000 ns, 0.000 ns); -- unused
      tpd_REFCLK_LOCK        :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PWRDWN                  :	in    STD_ULOGIC; -- Active low
      REFCLK                  :	in    STD_ULOGIC;
      LOWFREQ                 : in    STD_ULOGIC; 
      OSC2                    : in    STD_ULOGIC; 
      OSC1                    : in    STD_ULOGIC; 
      OSC0                    : in    STD_ULOGIC; 
      DIVI5                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI4                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI3                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI2                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI1                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI0                   : in    STD_ULOGIC; -- Clock multiplier
      DIVJ5                   : in    STD_ULOGIC; -- Clock divider
      DIVJ4                   : in    STD_ULOGIC; -- Clock divider
      DIVJ3                   : in    STD_ULOGIC; -- Clock divider
      DIVJ2                   : in    STD_ULOGIC; -- Clock divider
      DIVJ1                   : in    STD_ULOGIC; -- Clock divider
      DIVJ0                   : in    STD_ULOGIC; -- Clock divider
      DELAYLINE4              : in    STD_ULOGIC; -- Delay Value
      DELAYLINE3              : in    STD_ULOGIC; -- Delay Value
      DELAYLINE2              : in    STD_ULOGIC; -- Delay Value
      DELAYLINE1              : in    STD_ULOGIC; -- Delay Value
      DELAYLINE0              : in    STD_ULOGIC; -- Delay Value
      LOCK                    :	out   STD_ULOGIC;
      CLK1                    :	out   STD_ULOGIC;
      CLK2                    :	out   STD_ULOGIC);

attribute VITAL_LEVEL0 of PLL : entity is TRUE;
end PLL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of PLL is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL PWRDWN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL REFCLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LOWFREQ_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OSC2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OSC1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OSC0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVI5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVI4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVI3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVI2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVI1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVI0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVJ5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVJ4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVJ3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVJ2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVJ1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVJ0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DELAYLINE4_ipd : STD_ULOGIC := 'X';
   SIGNAL DELAYLINE3_ipd : STD_ULOGIC := 'X';
   SIGNAL DELAYLINE2_ipd : STD_ULOGIC := 'X';
   SIGNAL DELAYLINE1_ipd : STD_ULOGIC := 'X';
   SIGNAL DELAYLINE0_ipd : STD_ULOGIC := 'X';

   SIGNAL start_CLK2	 : STD_LOGIC := '0';
   SIGNAL restart_CLK2	 : STD_LOGIC := '0';
   SIGNAL CLK2_pw        : Time := 0.000 ns; -- CLK2 pulse width
   SIGNAL start_CLK1	 : STD_LOGIC := '0';
   SIGNAL restart_CLK1	 : STD_LOGIC := '0';
   SIGNAL CLK1_pw        : Time := 0.000 ns; -- CLK1 pulse width
   SIGNAL DIV            : Integer := 0;
   SIGNAL MULT           : Integer := 0;
   SIGNAL DELAY          : Time := 0.000 ns;

   SIGNAL REFCLK_period          : Time :=  0.000 ns; -- Current REFCLK period
   SIGNAL REFCLK_period_stable   : Integer := 0;      -- 1 when REFCLK period stable
   SIGNAL REFCLK_re              : Time :=  0.000 ns; -- Current REFCLK rising edge
   
   CONSTANT MINPER       : Time := 71.429 ns; -- 14 MHz
   CONSTANT MAXPER       : Time := 5.000 ns; -- 200 MHz
   
   SIGNAL ICLK1  : STD_ULOGIC := 'X';
   SIGNAL ICLK2  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
     VitalWireDelay (PWRDWN_ipd, PWRDWN, tipd_PWRDWN);
     VitalWireDelay (REFCLK_ipd, REFCLK, tipd_REFCLK);
     VitalWireDelay (LOWFREQ_ipd, LOWFREQ, tipd_LOWFREQ);
     VitalWireDelay (OSC2_ipd, OSC2, tipd_OSC2);
     VitalWireDelay (OSC1_ipd, OSC1, tipd_OSC1);
     VitalWireDelay (OSC0_ipd, OSC0, tipd_OSC0);
     VitalWireDelay (DIVI5_ipd, DIVI5, tipd_DIVI5);
     VitalWireDelay (DIVI4_ipd, DIVI4, tipd_DIVI4);
     VitalWireDelay (DIVI3_ipd, DIVI3, tipd_DIVI3);
     VitalWireDelay (DIVI2_ipd, DIVI2, tipd_DIVI2);
     VitalWireDelay (DIVI1_ipd, DIVI1, tipd_DIVI1);
     VitalWireDelay (DIVI0_ipd, DIVI0, tipd_DIVI0);
     VitalWireDelay (DIVJ5_ipd, DIVJ5, tipd_DIVJ5);
     VitalWireDelay (DIVJ4_ipd, DIVJ4, tipd_DIVJ4);
     VitalWireDelay (DIVJ3_ipd, DIVJ3, tipd_DIVJ3);
     VitalWireDelay (DIVJ2_ipd, DIVJ2, tipd_DIVJ2);
     VitalWireDelay (DIVJ1_ipd, DIVJ1, tipd_DIVJ1);
     VitalWireDelay (DIVJ0_ipd, DIVJ0, tipd_DIVJ0);
     VitalWireDelay (DELAYLINE4_ipd, DELAYLINE4, tipd_DELAYLINE4);
     VitalWireDelay (DELAYLINE3_ipd, DELAYLINE3, tipd_DELAYLINE3);
     VitalWireDelay (DELAYLINE2_ipd, DELAYLINE2, tipd_DELAYLINE2);
     VitalWireDelay (DELAYLINE1_ipd, DELAYLINE1, tipd_DELAYLINE1);
     VitalWireDelay (DELAYLINE0_ipd, DELAYLINE0, tipd_DELAYLINE0);

   end block WireDelay;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  ---------------------
  --  Get DELAYLINE, DIVI, DIVJ values 
  ---------------------

  GetDelay : process ( DELAYLINE4_ipd, DELAYLINE3_ipd, DELAYLINE2_ipd, DELAYLINE1_ipd, DELAYLINE0_ipd )

    variable DelayVal : Integer := 0;

  begin

    DelayVal := 0;
    if (TO_X01(DELAYLINE0_ipd) = '1') then
        DelayVal := DelayVal + 1;
    end if;
    if (TO_X01(DELAYLINE1_ipd) = '1') then
        DelayVal := DelayVal + 2;
    end if;
    if (TO_X01(DELAYLINE2_ipd) = '1') then
        DelayVal := DelayVal + 4;
    end if;
    if (TO_X01(DELAYLINE3_ipd) = '1') then
        DelayVal := DelayVal + 8;
    end if;
    if (TO_X01(DELAYLINE4_ipd) = '1') then
      DelayVal := 0 - DelayVal;
    end if;

    DELAY <= (real(DelayVal)) * 0.250 ns;

  end process GetDelay;

  GetDiv : process ( DIVJ5_ipd, DIVJ4_ipd, DIVJ3_ipd, DIVJ2_ipd, DIVJ1_ipd, DIVJ0_ipd )

    variable DivVal : Integer := 0;

  begin

    DivVal := 0;
    if (TO_X01(DIVJ0_ipd) = '1') then
      DivVal := DivVal + 1;
    end if;
    if (TO_X01(DIVJ1_ipd) = '1') then
      DivVal := DivVal + 2;
    end if;
    if (TO_X01(DIVJ2_ipd) = '1') then
      DivVal := DivVal + 4;
    end if;
    if (TO_X01(DIVJ3_ipd) = '1') then
      DivVal := DivVal + 8;
    end if;
    if (TO_X01(DIVJ4_ipd) = '1') then
      DivVal := DivVal + 16;
    end if;
    if (TO_X01(DIVJ5_ipd) = '1') then
      DivVal := DivVal + 32;
    end if;

    DIV <= DivVal + 1; -- "000000" means 1 and "111111" means 64

  end process GetDiv;

  GetMult : process ( DIVI5_ipd, DIVI4_ipd, DIVI3_ipd, DIVI2_ipd, DIVI1_ipd, DIVI0_ipd )

    variable MultVal : Integer := 0;

  begin

    MultVal := 0;
    if (TO_X01(DIVI0_ipd) = '1') then
      MultVal := MultVal + 1;
    end if;
    if (TO_X01(DIVI1_ipd) = '1') then
      MultVal := MultVal + 2;
    end if;
    if (TO_X01(DIVI2_ipd) = '1') then
      MultVal := MultVal + 4;
    end if;
    if (TO_X01(DIVI3_ipd) = '1') then
      MultVal := MultVal + 8;
    end if;
    if (TO_X01(DIVI4_ipd) = '1') then
      MultVal := MultVal + 16;
    end if;
    if (TO_X01(DIVI5_ipd) = '1') then
      MultVal := MultVal + 32;
    end if;


    MULT <= MultVal + 1; -- "000000" means 1 and "111111" means 64

  end process GetMult;

  --
  -- Get REFCLK period
  --

  GetRefclkPeriod : process ( REFCLK_ipd, PWRDWN_ipd, ICLK1, ICLK2 )

   VARIABLE period          : Time :=  0.000 ns; -- Current REFCLK period
   VARIABLE previous_period : Time := -1.000 ns; -- Previous REFCLK period
   VARIABLE re              : Time :=  0.000 ns; -- Current REFCLK rising edge
   VARIABLE previous_re     : Time :=  0.000 ns; -- Previous REFCLK rising edge
   VARIABLE last_re         : Time :=  0.000 ns; -- Last REFCLK rising edge

  begin

    if (PWRDWN_ipd = '1') then
      if (REFCLK_ipd'event and (TO_X01(REFCLK_ipd) = '1')) then
        previous_re := re;
        re := now;
        REFCLK_re <= re;
        period := re - previous_re;
        REFCLK_period <= period;
        if (previous_period /= period) then
          previous_period := period;
          REFCLK_period_stable <= 0;
        else
          REFCLK_period_stable <= 1;
        end if;
      elsif (now > 100 ns) then
        if ((now - 100 ns) > REFCLK_re) then
          REFCLK_period_stable <= 0;
        end if;
      end if;
    else
      previous_period := -1.000 ns;
      REFCLK_period_stable <= 0;
    end if;

  end process GetRefclkPeriod;

  --
  -- Raise Lock
  --

  RaiseLock : process ( REFCLK_ipd, REFCLK_period_stable )

    variable REFCLK_num_re           : Integer := 0; -- Number of REFCLK rising edges

  begin

    --
    -- Raise LOCK after REFCLK stabilizes and number of rising edges exceeds
    -- f_REFCLK_LOCK
    --

    if (REFCLK_period_stable = 1) then
      if (REFCLK_ipd'event and (TO_X01(REFCLK_ipd)='1')) then
        REFCLK_num_re := REFCLK_num_re + 1;
      end if;
    else
      REFCLK_num_re := 0;
    end if;
    if (REFCLK_num_re > f_REFCLK_LOCK) then
      LOCK <= '1' after tpd_REFCLK_LOCK(tr01);
    else
      LOCK <= '0' after tpd_REFCLK_LOCK(tr10);
    end if;

  end process RaiseLock;

  --
  -- Check REFCLK Frequency
  --

--  CheckFreq : process ( REFCLK_period )

    -- variable minper : Time := 0.000 ns;
    -- variable maxper : Time := 0.000 ns;

 -- begin

 --   if (REFCLK_period_stable = 1 and PWRDWN_ipd = '1') then
 --     -- minper := (1.0 / real(fmin_REFCLK));
 --     assert (REFCLK_period >= MINPER)
 --       report "REFCLK frequency below allowed minimum"
 --       severity error;
 --     -- maxper := (1.0 / real(fmax_REFCLK));
 --     assert (REFCLK_period <= MAXPER)
 --       report "REFCLK frequency above allowed maximum"
 --       severity error;
 --   end if;
 --
 -- end process CheckFreq;

  --
  -- Set CLK2 pulse width
  --

  SetClk2PW : process (PWRDWN_ipd, REFCLK_period_stable,
                       MULT, DELAY, restart_CLK2)

  begin

    if (REFCLK_period_stable = 1 and PWRDWN_ipd = '1') then
      if (DELAY'event) then
        start_CLK2 <= '0';
        restart_CLK2 <= '1' after REFCLK_period;
      elsif (restart_CLK2'event) then
        start_CLK2 <= '1';
        restart_CLK2 <= '0' after REFCLK_period;
      elsif (MULT > 0) then
        CLK2_pw <=  (REFCLK_period / (real(MULT) * 2.0));
        start_CLK2 <= '1';
      else
        CLK2_pw <=  (REFCLK_period / 2.0);
        start_CLK2 <= '1';
      end if;
    else
      start_CLK2 <= '0';
      restart_CLK2 <= '0';
    end if;

  end process SetClk2PW;

  --
  -- Set CLK1 pulse width
  --

  SetClk1PW : process (PWRDWN_ipd, REFCLK_period_stable,
                       DIV, DELAY, CLK2_pw, restart_CLK1)

  begin

    if (REFCLK_period_stable = 1 and PWRDWN_ipd = '1') then
      if (DELAY'event) then
        start_CLK1 <= '0';
        restart_CLK1 <= '1' after REFCLK_period;
      elsif (restart_CLK1'event) then
        start_CLK1 <= '1';
        restart_CLK1 <= '0' after REFCLK_period;
      elsif (DIV > 0) then
        CLK1_pw <=  CLK2_pw * DIV;
        start_CLK1 <= '1';
      else
        CLK1_pw <=  (REFCLK_period / 2.0);
        start_CLK1 <= '1';
      end if;
    else
      start_CLK1 <= '0';
      restart_CLK1 <= '0';
    end if;

  end process SetClk1PW;


  --
  -- Ouptut CLK1
  --

  OutputCLK1 : process

  begin

    wait until (start_CLK1'event and (TO_X01(start_CLK1) = '1'));
    wait until (REFCLK_ipd'event and (TO_X01(REFCLK_ipd) = '1'));
    wait for ((4 * REFCLK_period) + DELAY);
    while (start_CLK1 = '1') LOOP
      CLK1 <= '1';
      ICLK1 <= '1';
      wait for CLK1_pw;
      CLK1 <= '0';
      ICLK1 <= '0';
      wait for CLK1_pw;
    end loop;

    CLK1 <= 'X';

  end process OutputCLK1;

  --
  -- Output CLK2
  --

  OutputCLK2 : process 

  begin

    wait until (start_CLK2'event and (TO_X01(start_CLK2) = '1'));
    wait until (REFCLK_ipd'event and (TO_X01(REFCLK_ipd) = '1'));
    wait for ((4 * REFCLK_period) + DELAY);
    while (start_CLK2 = '1') LOOP
      CLK2 <= '1';
      ICLK2 <= '1';
      wait for CLK2_pw;
      CLK2 <= '0';
      ICLK2 <= '0';
      wait for CLK2_pw;
    end loop;

    CLK2 <= 'X';

  end process OutputCLK2;

end VITAL_ACT;

configuration CFG_PLL_VITAL of PLL is
   for VITAL_ACT
   end for;
end CFG_PLL_VITAL;

-- 
-- Actel AX family PLLFB VITAL simulation model.
--
-- 5/14/03:   Modified to take FB delay into account.
-- 7/17/03:   Modified to output X when REFCLK stuck @ 1/0.
-- 2/10/04:   Fixed to not use internal clock to catch stuck REFCLK.
-- 2/26/04:   Fixed Clk2_pw & clk1_pw - updated now after FB delay determined.
--
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

-- entity declaration --
entity PLLFB is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;

      f_REFCLK_LOCK          :	Integer := 3; -- Number of REFCLK pulses after which LOCK is raised.

      tipd_PWRDWN            :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_REFCLK            :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_FB                :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_LOWFREQ           :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OSC2              :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OSC1              :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OSC0              :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI5             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI4             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI3             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI2             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI1             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVI0             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ5             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ4             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ3             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ2             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ1             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DIVJ0             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE4        :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE3        :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE2        :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE1        :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DELAYLINE0        :  VitalDelayType01 := (0.000 ns, 0.000 ns);

      tpd_REFCLK_CLK1        :  VitalDelayType01 := (0.000 ns, 0.000 ns); -- unused
      tpd_REFCLK_CLK2        :  VitalDelayType01 := (0.000 ns, 0.000 ns); -- unused
      tpd_REFCLK_LOCK        :  VitalDelayType01 := (0.000 ns, 0.000 ns));



   port(
      PWRDWN                  :	in    STD_ULOGIC; -- Active low
      REFCLK                  :	in    STD_ULOGIC;
      FB                      :	in    STD_ULOGIC;
      LOWFREQ                 : in    STD_ULOGIC; 
      OSC2                    : in    STD_ULOGIC; 
      OSC1                    : in    STD_ULOGIC; 
      OSC0                    : in    STD_ULOGIC; 
      DIVI5                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI4                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI3                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI2                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI1                   : in    STD_ULOGIC; -- Clock multiplier
      DIVI0                   : in    STD_ULOGIC; -- Clock multiplier
      DIVJ5                   : in    STD_ULOGIC; -- Clock divider
      DIVJ4                   : in    STD_ULOGIC; -- Clock divider
      DIVJ3                   : in    STD_ULOGIC; -- Clock divider
      DIVJ2                   : in    STD_ULOGIC; -- Clock divider
      DIVJ1                   : in    STD_ULOGIC; -- Clock divider
      DIVJ0                   : in    STD_ULOGIC; -- Clock divider
      DELAYLINE4              : in    STD_ULOGIC; -- Delay Value
      DELAYLINE3              : in    STD_ULOGIC; -- Delay Value
      DELAYLINE2              : in    STD_ULOGIC; -- Delay Value
      DELAYLINE1              : in    STD_ULOGIC; -- Delay Value
      DELAYLINE0              : in    STD_ULOGIC; -- Delay Value
      LOCK                    :	out   STD_ULOGIC;
      CLK1                    :	out   STD_ULOGIC;
      CLK2                    :	out   STD_ULOGIC);

attribute VITAL_LEVEL0 of PLLFB : entity is TRUE;
end PLLFB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of PLLFB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL PWRDWN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL REFCLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL FB_ipd	 : STD_ULOGIC := 'X';
   SIGNAL LOWFREQ_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OSC2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OSC1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OSC0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVI5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVI4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVI3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVI2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVI1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVI0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVJ5_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVJ4_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVJ3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVJ2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVJ1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DIVJ0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL DELAYLINE4_ipd : STD_ULOGIC := 'X';
   SIGNAL DELAYLINE3_ipd : STD_ULOGIC := 'X';
   SIGNAL DELAYLINE2_ipd : STD_ULOGIC := 'X';
   SIGNAL DELAYLINE1_ipd : STD_ULOGIC := 'X';
   SIGNAL DELAYLINE0_ipd : STD_ULOGIC := 'X';

   SIGNAL start_CLK2	 : STD_LOGIC := '0';
   SIGNAL restart_CLK2	 : STD_LOGIC := '0';
   SIGNAL CLK2_pw        : Time := 0.000 ns; -- CLK2 pulse width
   SIGNAL start_CLK1	 : STD_LOGIC := '0';
   SIGNAL restart_CLK1	 : STD_LOGIC := '0';
   SIGNAL CLK1_pw        : Time := 0.000 ns; -- CLK1 pulse width
   SIGNAL DIV            : Integer := 0;
   SIGNAL MULT           : Integer := 0;
   SIGNAL DELAY          : Time := 0.000 ns;

   SIGNAL REFCLK_period          : Time :=  0.000 ns; -- Current REFCLK period
   SIGNAL REFCLK_period_stable   : Integer := 0;      -- 1 when REFCLK period stable
   SIGNAL REFCLK_re              : Time :=  0.000 ns; -- Current REFCLK rising edge

   SIGNAL FB_period              : Time :=  0.000 ns; -- Current FB period
   SIGNAL FB_period_stable       : Integer := 0;      -- 1 when FB period stable
   SIGNAL FB_re                  : Time :=  0.000 ns; -- Current FB rising edge
   SIGNAL FB_delay               : Time := -1.000 ns; -- FB delay
   SIGNAL FB_delay_determined    : Boolean := FALSE;  -- True when FB_delay determined

   CONSTANT MINPER       : Time := 71.429 ns; -- 14 MHz
   CONSTANT MAXPER       : Time := 5.000 ns;  -- 200 MHz
   
   SIGNAL ICLK1  : STD_ULOGIC := 'X';
   SIGNAL ICLK2  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
     VitalWireDelay (PWRDWN_ipd, PWRDWN, tipd_PWRDWN);
     VitalWireDelay (REFCLK_ipd, REFCLK, tipd_REFCLK);
     VitalWireDelay (FB_ipd, FB, tipd_FB);
     VitalWireDelay (LOWFREQ_ipd, LOWFREQ, tipd_LOWFREQ);
     VitalWireDelay (OSC2_ipd, OSC2, tipd_OSC2);
     VitalWireDelay (OSC1_ipd, OSC1, tipd_OSC1);
     VitalWireDelay (OSC0_ipd, OSC0, tipd_OSC0);
     VitalWireDelay (DIVI5_ipd, DIVI5, tipd_DIVI5);
     VitalWireDelay (DIVI4_ipd, DIVI4, tipd_DIVI4);
     VitalWireDelay (DIVI3_ipd, DIVI3, tipd_DIVI3);
     VitalWireDelay (DIVI2_ipd, DIVI2, tipd_DIVI2);
     VitalWireDelay (DIVI1_ipd, DIVI1, tipd_DIVI1);
     VitalWireDelay (DIVI0_ipd, DIVI0, tipd_DIVI0);
     VitalWireDelay (DIVJ5_ipd, DIVJ5, tipd_DIVJ5);
     VitalWireDelay (DIVJ4_ipd, DIVJ4, tipd_DIVJ4);
     VitalWireDelay (DIVJ3_ipd, DIVJ3, tipd_DIVJ3);
     VitalWireDelay (DIVJ2_ipd, DIVJ2, tipd_DIVJ2);
     VitalWireDelay (DIVJ1_ipd, DIVJ1, tipd_DIVJ1);
     VitalWireDelay (DIVJ0_ipd, DIVJ0, tipd_DIVJ0);
     VitalWireDelay (DELAYLINE4_ipd, DELAYLINE4, tipd_DELAYLINE4);
     VitalWireDelay (DELAYLINE3_ipd, DELAYLINE3, tipd_DELAYLINE3);
     VitalWireDelay (DELAYLINE2_ipd, DELAYLINE2, tipd_DELAYLINE2);
     VitalWireDelay (DELAYLINE1_ipd, DELAYLINE1, tipd_DELAYLINE1);
     VitalWireDelay (DELAYLINE0_ipd, DELAYLINE0, tipd_DELAYLINE0);

   end block WireDelay;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  ---------------------
  --  Get DELAYLINE, DIVI, DIVJ values 
  ---------------------

  GetDelay : process ( DELAYLINE4_ipd, DELAYLINE3_ipd, DELAYLINE2_ipd, DELAYLINE1_ipd, DELAYLINE0_ipd )

    variable DelayVal : Integer := 0;

  begin

    DelayVal := 0;
    if (TO_X01(DELAYLINE0_ipd) = '1') then
        DelayVal := DelayVal + 1;
    end if;
    if (TO_X01(DELAYLINE1_ipd) = '1') then
        DelayVal := DelayVal + 2;
    end if;
    if (TO_X01(DELAYLINE2_ipd) = '1') then
        DelayVal := DelayVal + 4;
    end if;
    if (TO_X01(DELAYLINE3_ipd) = '1') then
        DelayVal := DelayVal + 8;
    end if;
    if (TO_X01(DELAYLINE4_ipd) = '1') then
      DelayVal := 0 - DelayVal;
    end if;

    DELAY <= (real(DelayVal)) * 0.250 ns;

  end process GetDelay;

  GetDiv : process ( DIVJ5_ipd, DIVJ4_ipd, DIVJ3_ipd, DIVJ2_ipd, DIVJ1_ipd, DIVJ0_ipd )

    variable DivVal : Integer := 0;

  begin

    DivVal := 0;
    if (TO_X01(DIVJ0_ipd) = '1') then
      DivVal := DivVal + 1;
    end if;
    if (TO_X01(DIVJ1_ipd) = '1') then
      DivVal := DivVal + 2;
    end if;
    if (TO_X01(DIVJ2_ipd) = '1') then
      DivVal := DivVal + 4;
    end if;
    if (TO_X01(DIVJ3_ipd) = '1') then
      DivVal := DivVal + 8;
    end if;
    if (TO_X01(DIVJ4_ipd) = '1') then
      DivVal := DivVal + 16;
    end if;
    if (TO_X01(DIVJ5_ipd) = '1') then
      DivVal := DivVal + 32;
    end if;

    DIV <= DivVal + 1; -- "000000" means 1 and "111111" means 64

  end process GetDiv;

  GetMult : process ( DIVI5_ipd, DIVI4_ipd, DIVI3_ipd, DIVI2_ipd, DIVI1_ipd, DIVI0_ipd )

    variable MultVal : Integer := 0;

  begin

    MultVal := 0;
    if (TO_X01(DIVI0_ipd) = '1') then
      MultVal := MultVal + 1;
    end if;
    if (TO_X01(DIVI1_ipd) = '1') then
      MultVal := MultVal + 2;
    end if;
    if (TO_X01(DIVI2_ipd) = '1') then
      MultVal := MultVal + 4;
    end if;
    if (TO_X01(DIVI3_ipd) = '1') then
      MultVal := MultVal + 8;
    end if;
    if (TO_X01(DIVI4_ipd) = '1') then
      MultVal := MultVal + 16;
    end if;
    if (TO_X01(DIVI5_ipd) = '1') then
      MultVal := MultVal + 32;
    end if;


    MULT <= MultVal + 1; -- "000000" means 1 and "111111" means 64

  end process GetMult;

  --
  -- Get REFCLK period
  --

  GetRefclkPeriod : process ( REFCLK_ipd, PWRDWN_ipd, ICLK1, ICLK2 )

   VARIABLE period          : Time :=  0.000 ns; -- Current REFCLK period
   VARIABLE previous_period : Time := -1.000 ns; -- Previous REFCLK period
   VARIABLE re              : Time :=  0.000 ns; -- Current REFCLK rising edge
   VARIABLE previous_re     : Time :=  0.000 ns; -- Previous REFCLK rising edge
   VARIABLE last_re         : Time :=  0.000 ns; -- Last REFCLK rising edge

  begin

    if (PWRDWN_ipd = '1') then
      if (REFCLK_ipd'event and (TO_X01(REFCLK_ipd) = '1')) then
        previous_re := re;
        re := now;
        REFCLK_re <= re;
        period := re - previous_re;
        REFCLK_period <= period;
        if (previous_period /= period) then
          previous_period := period;
          REFCLK_period_stable <= 0;
        else
          REFCLK_period_stable <= 1;
        end if;
      elsif (now > 100 ns) then
        if ((now - 100 ns) > REFCLK_re) then
          REFCLK_period_stable <= 0;
        end if;
      end if;
    else
      previous_period := -1.000 ns;
      REFCLK_period_stable <= 0;
    end if;

  end process GetRefclkPeriod;

  --
  -- Get FB period
  --

  GetFBPeriod : process ( FB_ipd, PWRDWN_ipd )

   VARIABLE period              : Time :=  0.000 ns; -- Current FB period
   VARIABLE previous_period     : Time := -1.000 ns; -- Previous FB period
   VARIABLE re                  : Time :=  0.000 ns; -- Current FB rising edge
   VARIABLE previous_re         : Time :=  0.000 ns; -- Previous FB rising edge

  begin

    if (PWRDWN_ipd = '1') then
      if (FB_ipd'event) then
        if (TO_X01(FB_ipd) = '1') then
          previous_re := re;
          re := now;
          FB_re <= re;
          period := re - previous_re;
          FB_period <= period;
          if (previous_period /= period) then
            previous_period := period;
            FB_period_stable <= 0;
          else
            FB_period_stable <= 1;
          end if;
        elsif (TO_X01(FB_ipd) = 'X') then
          previous_period := -1.000 ns;
          FB_period_stable <= 0;
        end if;
      end if;
    else
      previous_period := -1.000 ns;
      FB_period_stable <= 0;
    end if;

  end process GetFBPeriod;

  --
  -- Get FB delay
  --

  GetFBDelay : process ( FB_period_stable, REFCLK_period_stable, PWRDWN_ipd )

    VARIABLE delay      : Time := -1.000 ns;
    VARIABLE prev_delay : Time := -1.000 ns;

  begin

    if (PWRDWN_ipd = '1') then
      if (FB_period_stable = 1 and REFCLK_period_stable = 1 and 
          FB_delay_determined = FALSE) then
        if (FB_re > REFCLK_re) then
          delay := FB_re - REFCLK_re;
          if (delay /= prev_delay) then
            prev_delay := delay;
            FB_delay <= delay;
            FB_delay_determined <= TRUE;
          end if;
        end if;
      end if;
    end if;

  end process GetFBDelay;

  --
  -- Raise Lock
  --

  RaiseLock : process ( REFCLK_ipd, REFCLK_period_stable, FB_delay_determined )

    variable REFCLK_num_re           : Integer := 0; -- Number of REFCLK rising edges

  begin

    --
    -- Raise LOCK after FB_delay determined, REFCLK stabilizes, and the
    -- number of rising edges exceeds f_REFCLK_LOCK
    --

    if (FB_delay_determined) then
      if (FB_period_stable = 1 and REFCLK_period_stable = 1) then
        if (REFCLK_ipd'event and (TO_X01(REFCLK_ipd)='1')) then
          REFCLK_num_re := REFCLK_num_re + 1;
        end if;
      else
        REFCLK_num_re := 0;
      end if;
      if (REFCLK_num_re > f_REFCLK_LOCK) then
        LOCK <= '1' after tpd_REFCLK_LOCK(tr01);
      else
        LOCK <= '0' after tpd_REFCLK_LOCK(tr10);
      end if;
    end if;

  end process RaiseLock;

  --
  -- Set CLK2 pulse width
  --

  SetClk2PW : process (PWRDWN_ipd, REFCLK_period_stable, FB_delay_determined,
                       MULT, DELAY, restart_CLK2)

  begin

    if (REFCLK_period_stable = 1 and PWRDWN_ipd = '1') then
      if (FB_delay_determined) then
        if (FB_delay_determined'event) then
          start_CLK2 <= '0';
          restart_CLK2 <= '1' after REFCLK_period;
        end if;
      else 
        CLK2_pw <=  (REFCLK_period / 2.0);
        start_CLK2 <= '1';
      end if;
      if (DELAY'event) then
        start_CLK2 <= '0';
        restart_CLK2 <= '1' after REFCLK_period;
      end if;
      if (MULT > 0) then
        CLK2_pw <=  (REFCLK_period / (real(MULT) * 2.0));
        if (start_CLK2 = '0') then
          start_CLK2 <= '1' after REFCLK_period;
        end if;
      else
        CLK2_pw <=  (REFCLK_period / 2.0);
        if (start_CLK2 = '0') then
          start_CLK2 <= '1' after REFCLK_period;
        end if;
      end if;
      if (restart_CLK2'event and restart_CLK2 = '1') then
        start_CLK2 <= '1';
        restart_CLK2 <= '0' after REFCLK_period;
      end if;
    else
      start_CLK2 <= '0';
      restart_CLK2 <= '0';
    end if;

  end process SetClk2PW;

  --
  -- Set CLK1 pulse width
  --

  SetClk1PW : process (PWRDWN_ipd, REFCLK_period_stable, FB_delay_determined,
                       DIV, DELAY, CLK2_pw, restart_CLK1)

  begin

    if (REFCLK_period_stable = 1 and PWRDWN_ipd = '1') then
      if (FB_delay_determined) then
        if (FB_delay_determined'event) then
          start_CLK1 <= '0';
          restart_CLK1 <= '1' after REFCLK_period;
        end if;
      else
        CLK1_pw <=  (REFCLK_period / 2.0);
        start_CLK1 <= '1';
      end if;
      if (DELAY'event) then
        start_CLK1 <= '0';
        restart_CLK1 <= '1' after REFCLK_period;
      end if;
      if (DIV > 0) then
        CLK1_pw <=  CLK2_pw * DIV;
        if (start_CLK1 = '0') then
          start_CLK1 <= '1' after REFCLK_period;
        end if;
      else
        CLK1_pw <=  (REFCLK_period / 2.0);
        if (start_CLK1 = '0') then
          start_CLK1 <= '1' after REFCLK_period;
        end if;
      end if;
      if (restart_CLK1'event and restart_CLK1 = '1') then
        start_CLK1 <= '1';
        restart_CLK1 <= '0' after REFCLK_period;
      end if;
    else
      start_CLK1 <= '0';
      restart_CLK1 <= '0';
    end if;

  end process SetClk1PW;


  --
  -- Ouptut CLK1
  --

  OutputCLK1 : process

  begin

    wait until (start_CLK1'event and (TO_X01(start_CLK1) = '1'));
    wait until (REFCLK_ipd'event and (TO_X01(REFCLK_ipd) = '1'));
    if (FB_delay_determined) then
      wait for ((4 * REFCLK_period) + DELAY - FB_delay);
    end if;
    while (start_CLK1 = '1') LOOP
      CLK1 <= '1';
      ICLK1 <= '1';
      wait for CLK1_pw;
      CLK1 <= '0';
      ICLK1 <= '0';
      wait for CLK1_pw;
    end loop;

    CLK1 <= 'X';

  end process OutputCLK1;

  --
  -- Output CLK2
  --

  OutputCLK2 : process 

  begin

    wait until (start_CLK2'event and (TO_X01(start_CLK2) = '1'));
    wait until (REFCLK_ipd'event and (TO_X01(REFCLK_ipd) = '1'));
    if (FB_delay_determined) then
      wait for ((4 * REFCLK_period) + DELAY - FB_delay);
    end if;
    while (start_CLK2 = '1') LOOP
      CLK2 <= '1';
      ICLK2 <= '1';
      wait for CLK2_pw;
      CLK2 <= '0';
      ICLK2 <= '0';
      wait for CLK2_pw;
    end loop;

    CLK2 <= 'X';

  end process OutputCLK2;

end VITAL_ACT;

configuration CFG_PLLFB_VITAL of PLLFB is
   for VITAL_ACT
   end for;
end CFG_PLLFB_VITAL;

-----------------------------------------------------------------
--
--  Actel IOFIFO_BIDIROUTFIFO VHDL behavioral model
--  64 X 1 I/O FIFO with rising write clock, rising read clock,
--  and active low WENB, RENB, and CLRB.
--  AFL macro containing feed-through.
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - 5/17/02 - Dale Walter - Clone of IOFIFO_INFIFO.
-- 2.0 - 9/27/02 - Krupa Singampalli - New Timing Arcs
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity IOFIFO_BIDIROUTFIFO is
  GENERIC (
        tipd_A       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_D       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RENB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tipd_CLRB      : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_A_Y   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_RCLK_Q   : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tpd_CLRB_Q    : VitalDelayType01 := (0.100 ns, 0.100 ns);
        tsetup_D_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_D_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_D_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_D_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_RENB_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WENB_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_RENB_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WENB_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        thold_CLRB_RCLK_negedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_RCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        thold_CLRB_WCLK_posedge_posedge     :   VitalDelayType := 0.000 ns;
        trecovery_CLRB_WCLK_posedge_posedge :  VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_CLRB_negedge     : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True

        );
  PORT (
        A     : IN STD_ULOGIC ;
        D     : IN STD_ULOGIC ;
        WENB     : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RENB     : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        CLRB    : IN STD_ULOGIC ;
        Q     : OUT STD_ULOGIC ;
        Y     : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of IOFIFO_BIDIROUTFIFO : entity is TRUE;
  
end IOFIFO_BIDIROUTFIFO;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of IOFIFO_BIDIROUTFIFO is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal A_ipd   : std_ulogic := 'X';
  signal D_ipd   : std_ulogic := 'X';
  signal WENB_ipd   : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  signal RENB_ipd   : std_ulogic := 'X';
  signal RCLK_ipd : std_ulogic := 'X';
  signal CLRB_ipd  : std_ulogic := 'X';
  type MEM is array(0 to 63) of std_ulogic;
  signal DUAL_PORT_RAM : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (A_ipd, A, VitalExtendToFillDelay(tipd_A));
    VitalWireDelay (D_ipd, D, VitalExtendToFillDelay(tipd_D));
    VitalWireDelay (WENB_ipd, WENB, VitalExtendToFillDelay(tipd_WENB));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (RENB_ipd, RENB, VitalExtendToFillDelay(tipd_RENB));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
    VitalWireDelay (CLRB_ipd, CLRB, VitalExtendToFillDelay(tipd_CLRB));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (A_ipd, D_ipd, WENB_ipd, WCLK_ipd, RENB_ipd, RCLK_ipd, CLRB_ipd)

     --  Read Timing Check Results
     variable Tviol_RENB_RCLK_posedge : X01 := '0';
     variable TmDt_RENB_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_D_WCLK_posedge : X01 := '0';
     variable TmDt_D_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WENB_WCLK_posedge : X01 := '0';
     variable TmDt_WENB_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  CLRB Timing Check Results
     variable Tviol_CLRB_RCLK_posedge : X01 := '0';
     variable TmDt_CLRB_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_CLRB_WCLK_posedge : X01 := '0';
     variable TmDt_CLRB_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_CLRB : X01 := '0';
     variable PeriodData_CLRB : VitalPeriodDataType := VitalPeriodDataInit;

     --  Functional Results
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT : SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1; -- free running counter
     variable RADDR : integer := -1; -- free running counter
     variable Q_zd : std_ulogic;
     variable Y_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable Q_GlitchData : VitalGlitchDataType;
     variable Y_GlitchData : VitalGlitchDataType;

     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable RENB_delayed : std_ulogic := 'X';
     variable RENB_previous : std_ulogic := 'X';
     variable WENB_delayed : std_ulogic := 'X';
     variable WENB_previous : std_ulogic := 'X';
     variable D_delayed : std_ulogic := 'X';

  begin  --  process VITALBehavior 

    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RENB before RCLK rising
      --   Hold  RENB after RCLK rising

      VitalSetupHoldCheck ( Tviol_RENB_RCLK_posedge,
                            TmDt_RENB_RCLK_posedge,
                            RENB_ipd, "RENB",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RENB_RCLK_posedge_posedge,
			    tsetup_RENB_RCLK_negedge_posedge,
                            thold_RENB_RCLK_posedge_posedge,
                            thold_RENB_RCLK_negedge_posedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            '/',
                            InstancePath & "/IOFIFO_BIDIROUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            InstancePath & "/IOFIFO_BIDIROUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup D high or low before WCLK rising
      --   Hold  D high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_D_WCLK_posedge,
                            TmDt_D_WCLK_posedge,
                            D_ipd, "D",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_D_WCLK_posedge_posedge,
                            tsetup_D_WCLK_negedge_posedge,
                            thold_D_WCLK_posedge_posedge,
                            thold_D_WCLK_negedge_posedge,
                            TO_X01((CLRB_ipd) AND (NOT WENB_ipd)) /= '0',
                            '/',
                            InstancePath & "/IOFIFO_BIDIROUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup WENB high before WCLK rising
      --   Hold  WENB high after WCLK rising

      VitalSetupHoldCheck ( Tviol_WENB_WCLK_posedge,
                            TmDt_WENB_WCLK_posedge,
                            WENB_ipd, "WENB",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WENB_WCLK_posedge_posedge,
                            tsetup_WENB_WCLK_negedge_posedge,
                            thold_WENB_WCLK_posedge_posedge,
                            thold_WENB_WCLK_negedge_posedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            '/',
                            InstancePath & "/IOFIFO_BIDIROUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TO_X01((CLRB_ipd) ) /= '0',
                            InstancePath & "/IOFIFO_BIDIROUTFIFO",
                            Xon,
                            MsgOn,
                            WARNING
                            );

      --   Setup CLRB high before WCLK rising
      --   Hold  CLRB high after WCLK rising

         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLRB_RCLK_posedge,
          TimingData              => TmDt_CLRB_RCLK_posedge,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          RefSignal               => RCLK_ipd,
          RefSignalName           => "RCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLRB_RCLK_posedge_posedge,
          Removal                 => thold_CLRB_RCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TO_X01(NOT RENB_ipd) /='0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IOFIFO_BIDIROUTFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLRB_WCLK_posedge,
          TimingData              => TmDt_CLRB_WCLK_posedge,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          RefSignal               => RCLK_ipd,
          RefSignalName           => "WCLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLRB_WCLK_posedge_posedge,
          Removal                 => thold_CLRB_WCLK_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => TO_X01(NOT WENB_ipd) /='0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IOFIFO_BIDIROUTFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLRB,
          PeriodData              => PeriodData_CLRB,
          TestSignal              => CLRB_ipd,
          TestSignalName          => "CLRB",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLRB_negedge,
          CheckEnabled            => TRUE,
          HeaderMsg               => InstancePath &"/IOFIFO_BIDIROUTFIFO",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);


    end if;

      Y_zd := TO_X01(A_ipd);

    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################


      if (TO_X01(CLRB_ipd)='X') then
        assert false
        report ": CLRB unknown"
        severity Warning;
      elsif (TO_X01(CLRB_ipd)='0') then
        WADDR := -1;
        RADDR := -1;
      else
        if (TO_X01(WCLK_ipd)='X') then
	  if ((TO_X01(WENB_delayed) /= '1')) then
            if (TO_X01(WCLK_previous) /= 'X') then
	      assert false
	      report ": WCLK went unknown"
	      severity Warning;
	    end if;
	  end if;
        elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='1')) then
	  case (TO_X01(WENB_delayed)) is
	    when '1' =>
	      null;
	    when '0' =>
              -- Increment WADDR
              WADDR := WADDR + 1;
              if ((RADDR > WADDR) or (WADDR - RADDR > 63)) then
                assert false
                report ": Write failed - FIFO full."
                severity Warning;
              else
	        DUAL_PORT_RAM(WADDR mod 64) <= D_delayed ;
              end if;
	    when others =>
              if (TO_X01(WENB_previous) = 'X') then
                assert false
                report ": WENB went unknown"
                severity Warning;
              end if;
	  end case;
        end if;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      if (TO_X01(CLRB_ipd)='1') then
        if (TO_X01(RCLK_ipd) = 'X') then
          if ((TO_X01(RENB_delayed) /= '1')) then
	    Q_zd := 'X';
	    if (TO_X01(RCLK_previous) /= 'X') then
	      assert false
	      report ": RCLK went unknown"
	      severity Warning;
	    end if;
	  end if;
        elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '1')) then
	  case (TO_X01(RENB_delayed)) is
	    when '1' =>
	      null;
	    when '0' =>
              -- Increment RADDR
              RADDR := RADDR + 1;
              if ((RADDR > WADDR) or (WADDR - RADDR > 63)) then
                assert false
                report ": Read failed - FIFO empty."
                severity Warning;
              else
	        Q_zd := DUAL_PORT_RAM(RADDR mod 64);
              end if;
	    when others =>
	      Q_zd := 'X';
              if (TO_X01(RENB_delayed) = 'X') and (TO_X01(RENB_previous) /= 'X') then
	        assert false
	        report ": RENB went unknown"
	        severity Warning;
                RENB_previous := RENB_delayed;
              end if;
	  end case;
        end if;
      end if;

      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      if WENB_ipd'event then
        WENB_previous := WENB_delayed;
        WENB_delayed := WENB_ipd;
      end if;
      if RENB_ipd'event then
        RENB_previous := RENB_delayed;
        RENB_delayed := RENB_ipd;
      end if;
      D_delayed := D_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => Q,
	GlitchData => Q_GlitchData,
	OutSignalName => "Q",
	OutTemp => Q_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_Q), true)),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => Xon,
	MsgOn => MsgOn,
	MsgSeverity => WARNING
	);

   VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, true)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

  end process VITALBehavior;

end VITAL_ACT;

----- CELL DDR_OUT ----
library ieee;
use ieee.std_logic_1164.all;
library axcelerator;

entity DDR_OUT is
    port(DR, DF, E, CLK, PRE, CLR : in std_logic;  Q : out std_logic) ;
end DDR_OUT;


architecture DEF_ARCH of  DDR_OUT is

    component DFEG
        port(D, E, CLK, CLR, PRE : in std_logic := 'U'; Q : out std_logic) ;
    end component;

    component DFEH
        port(D, E, CLK, CLR, PRE : in std_logic := 'U'; Q : out std_logic) ;
    end component;

    component MX2
        port(A, S, B : in std_logic := 'U'; Y : out std_logic) ;
    end component;

    signal QR   : std_ulogic := 'X';
    signal QF   : std_ulogic := 'X';

    begin

    U0 : DFEH
         port map(D => DF, E => E, CLK => CLK, CLR => CLR, PRE => PRE, Q => QF);
    U1 : DFEG
         port map(D => DR, E => E, CLK => CLK, CLR => CLR, PRE => PRE, Q => QR);
    U2 : MX2
         port map(A => QF, B => QR, S => CLK, Y => Q);

end DEF_ARCH;


----- CELL DDR_REG ----
library ieee;
use ieee.std_logic_1164.all;
library axcelerator;

entity DDR_REG is
    port(D, E, CLK, CLR, PRE : in std_logic;  QR, QF : out std_logic) ;
end DDR_REG;


architecture DEF_ARCH of  DDR_REG is

    component DFEG
        port(D, E, CLK, CLR, PRE : in std_logic := 'U'; Q : out std_logic) ;
    end component;

    component DFEH
        port(D, E, CLK, CLR, PRE : in std_logic := 'U'; Q : out std_logic) ;
    end component;

    begin

    U0 : DFEG
         port map(D => D, E => E, CLK => CLK, CLR => CLR, PRE => PRE, Q => QR);
    U1 : DFEH
         port map(D => D, E => E, CLK => CLK, CLR => CLR, PRE => PRE, Q => QF);

end DEF_ARCH;


library ieee;
use ieee.std_logic_1164.all;
library axcelerator;

----- CELL NAND5D ----
library ieee;
use ieee.std_logic_1164.all;
library axcelerator;

-- entity declaration --
entity NAND5D is
   port(
          A     : in std_logic;
          B     : in std_logic;
          C     : in std_logic;
          D     : in std_logic;
          E     : in std_logic;
          Y             : out std_logic);
end NAND5D;

-- architecture body --
architecture DEF_ARCH of  NAND5D is

-- component declaration --
COMPONENT OR5A
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


begin

     U1 : OR5A
          port map( A  => E,  B  => D,  C  => C,  D  => B,  E  => A,  Y  => Y);

end DEF_ARCH;


----- CELL NOR5D ----
library ieee;
use ieee.std_logic_1164.all;
library axcelerator;

-- entity declaration --
entity NOR5D is
   port(
          A     : in std_logic;
          B     : in std_logic;
          C     : in std_logic;
          D     : in std_logic;
          E     : in std_logic;
          Y             : out std_logic);
end NOR5D;

-- architecture body --
architecture DEF_ARCH of  NOR5D is

-- component declaration --
COMPONENT AND5A
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


begin

     U1 : AND5A
          port map( A  => E,  B  => D,  C  => C,  D  => B,  E  => A,  Y  => Y);

end DEF_ARCH;




 ---- CELL ADDSUB1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity ADDSUB1 is
    generic(
                TimingChecksOn:Boolean :=True;
                Xon: Boolean :=False;
                InstancePath: STRING :="*";
                MsgOn: Boolean :=True;
                tpd_A_S         : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_FCI_S               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_B_S         : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_A_FCO               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_B_FCO               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_AS_FCO              : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_FCI_FCO             : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_A          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_FCI                : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_B          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_AS         : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                A               : in    STD_ULOGIC;
                FCI             : in    STD_ULOGIC;
                B               : in    STD_ULOGIC;
                AS              : in    STD_ULOGIC;
                S               : out    STD_ULOGIC;
                FCO             : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of ADDSUB1 :  entity is TRUE;
 end ADDSUB1;


-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of ADDSUB1 is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL A_ipd  : STD_ULOGIC := 'X';
        SIGNAL FCI_ipd  : STD_ULOGIC := 'X';
        SIGNAL B_ipd  : STD_ULOGIC := 'X';
        SIGNAL AS_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (A_ipd, A, tipd_A);
        VitalWireDelay (FCI_ipd, FCI, tipd_FCI);
        VitalWireDelay (B_ipd, B, tipd_B);
        VitalWireDelay (AS_ipd, AS, tipd_AS);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (A_ipd, FCI_ipd, B_ipd, AS_ipd)


        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
        ALIAS S_zd : STD_LOGIC is Results(1);
        ALIAS FCO_zd : STD_LOGIC is Results(2);

        -- output glitch detection variables
        VARIABLE S_GlitchData  : VitalGlitchDataType;
        VARIABLE FCO_GlitchData  : VitalGlitchDataType;

        begin


           -------------------------
           --  Functionality Section
           -------------------------
           S_zd := (FCI_ipd) XOR ( NOT((B_ipd) XOR (A_ipd) XOR (AS_ipd)) );
           FCO_zd := ((( A_ipd  AND  NOT VitalMUX2( AS_ipd , (NOT AS_ipd) , (NOT B_ipd) )) OR ( A_ipd  AND  FCI_ipd )) OR ( FCI_ipd  AND  NOT VitalMUX2( AS_ipd
 , (NOT AS_ipd) , (NOT B_ipd) )));


           ----------------------
           --  Path Delay Section
           ----------------------

     VitalPathDelay01 (
           OutSignal => S,
           GlitchData => S_GlitchData,
           OutSignalName => "S",
           OutTemp => S_zd,
           Paths => (
                     0 => (A_ipd'last_event,tpd_A_S, true),
                     1 => (FCI_ipd'last_event,tpd_FCI_S, true),
                     2 => (B_ipd'last_event,tpd_B_S, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING);

     VitalPathDelay01 (
           OutSignal => FCO,
           GlitchData => FCO_GlitchData,
           OutSignalName => "FCO",
           OutTemp => FCO_zd,
           Paths => (
                     0 => (A_ipd'last_event,tpd_A_FCO, true),
                     1 => (B_ipd'last_event,tpd_B_FCO, true),
                     2 => (AS_ipd'last_event,tpd_AS_FCO, true),
                     3 => (FCI_ipd'last_event,tpd_FCI_FCO, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_ADDSUB1_VITAL of ADDSUB1 is
    for VITAL_ACT
    end for;
 end CFG_ADDSUB1_VITAL;


 ---- CELL FA1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity FA1A is
    generic(
                TimingChecksOn:Boolean :=True;
                Xon: Boolean :=False;
                InstancePath: STRING :="*";
                MsgOn: Boolean :=True;
                tpd_CI_CO               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_B_CO                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_A_CO                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CI_S                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_A_S         : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_B_S         : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_CI         : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_B          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_A          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                CI              : in    STD_ULOGIC;
                B               : in    STD_ULOGIC;
                A               : in    STD_ULOGIC;
                CO              : out    STD_ULOGIC;
                S               : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of FA1A :  entity is TRUE;
 end FA1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of FA1A is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL CI_ipd  : STD_ULOGIC := 'X';
        SIGNAL B_ipd  : STD_ULOGIC := 'X';
        SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (CI_ipd, CI, tipd_CI);
        VitalWireDelay (B_ipd, B, tipd_B);
        VitalWireDelay (A_ipd, A, tipd_A);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (CI_ipd, B_ipd, A_ipd)


        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
        ALIAS CO_zd : STD_LOGIC is Results(1);
        ALIAS S_zd : STD_LOGIC is Results(2);

        -- output glitch detection variables
        VARIABLE CO_GlitchData  : VitalGlitchDataType;
        VARIABLE S_GlitchData  : VitalGlitchDataType;

        begin

           -------------------------
           --  Functionality Section
           -------------------------

         S_zd :=
       (((NOT A_ipd)) AND ((((NOT B_ipd)) AND (A_ipd)) OR (((NOT B_ipd)) AND
         (CI_ipd) AND ((NOT A_ipd))) OR ((CI_ipd) AND (B_ipd) AND (A_ipd)))
         AND (CI_ipd)) OR (((NOT A_ipd)) AND (B_ipd) AND ((NOT CI_ipd))) OR
         ((A_ipd) AND ((((NOT B_ipd)) AND (A_ipd)) OR (((NOT B_ipd)) AND
         (CI_ipd) AND ((NOT A_ipd))) OR ((CI_ipd) AND (B_ipd) AND (A_ipd)))
         AND ((NOT CI_ipd))) OR ((A_ipd) AND (B_ipd) AND (CI_ipd));
      CO_zd :=
       (((NOT B_ipd)) AND (A_ipd)) OR (((NOT B_ipd)) AND (CI_ipd)) OR
       ((CI_ipd) AND (A_ipd));


           ----------------------
           --  Path Delay Section
           ----------------------

     VitalPathDelay01 (
           OutSignal => CO,
           GlitchData => CO_GlitchData,
           OutSignalName => "CO",
           OutTemp => CO_zd,
           Paths => (
                     0 => (CI_ipd'last_event,tpd_CI_CO, true),
                     1 => (B_ipd'last_event,tpd_B_CO, true),
                     2 => (A_ipd'last_event,tpd_A_CO, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING);

     VitalPathDelay01 (
           OutSignal => S,
           GlitchData => S_GlitchData,
           OutSignalName => "S",
           OutTemp => S_zd,
           Paths => (
                     0 => (CI_ipd'last_event,tpd_CI_S, true),
                     1 => (A_ipd'last_event,tpd_A_S, true),
                     2 => (B_ipd'last_event,tpd_B_S, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_FA1A_VITAL of FA1A is
    for VITAL_ACT
    end for;
 end CFG_FA1A_VITAL;



 ---- CELL FA1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity FA1B is
    generic(
                TimingChecksOn:Boolean :=True;
                Xon: Boolean :=False;
                InstancePath: STRING :="*";
                MsgOn: Boolean :=True;
                tpd_A_CO                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_B_CO                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CI_CO               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CI_S                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_A_S         : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_B_S         : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_A          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_B          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CI         : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                A               : in    STD_ULOGIC;
                B               : in    STD_ULOGIC;
                CI              : in    STD_ULOGIC;
                CO              : out    STD_ULOGIC;
                S               : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of FA1B :  entity is TRUE;
 end FA1B;
-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of FA1B is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL A_ipd  : STD_ULOGIC := 'X';
        SIGNAL B_ipd  : STD_ULOGIC := 'X';
        SIGNAL CI_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (A_ipd, A, tipd_A);
        VitalWireDelay (B_ipd, B, tipd_B);
        VitalWireDelay (CI_ipd, CI, tipd_CI);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (A_ipd, B_ipd, CI_ipd)


        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
        ALIAS CO_zd : STD_LOGIC is Results(1);
        ALIAS S_zd : STD_LOGIC is Results(2);

        -- output glitch detection variables
        VARIABLE CO_GlitchData  : VitalGlitchDataType;
        VARIABLE S_GlitchData  : VitalGlitchDataType;

        begin

           -------------------------
           --  Functionality Section
           -------------------------
           S_zd :=
       ((((((CI_ipd) AND ((NOT B_ipd)) AND (A_ipd)) OR ((((CI_ipd) AND
         (B_ipd)) OR ((NOT B_ipd))) AND ((NOT A_ipd)))) AND (CI_ipd)) OR
         ((B_ipd) AND ((NOT CI_ipd)))) AND (A_ipd)) OR ((((B_ipd) AND
         (CI_ipd)) OR ((((CI_ipd) AND ((NOT B_ipd)) AND (A_ipd)) OR
         ((((CI_ipd) AND (B_ipd)) OR ((NOT B_ipd))) AND ((NOT A_ipd)))) AND
         ((NOT CI_ipd)))) AND ((NOT A_ipd)));
      CO_zd :=
       ((CI_ipd) AND ((NOT B_ipd))) OR ((CI_ipd) AND ((NOT A_ipd)))
         OR (((NOT B_ipd)) AND ((NOT A_ipd)));



           ----------------------
           --  Path Delay Section
           ----------------------

     VitalPathDelay01 (
           OutSignal => CO,
           GlitchData => CO_GlitchData,
           OutSignalName => "CO",
           OutTemp => CO_zd,
           Paths => (
                     0 => (A_ipd'last_event,tpd_A_CO, true),
                     1 => (B_ipd'last_event,tpd_B_CO, true),
                     2 => (CI_ipd'last_event,tpd_CI_CO, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING);

     VitalPathDelay01 (
           OutSignal => S,
           GlitchData => S_GlitchData,
           OutSignalName => "S",
           OutTemp => S_zd,
           Paths => (
                     0 => (CI_ipd'last_event,tpd_CI_S, true),
                     1 => (A_ipd'last_event,tpd_A_S, true),
                     2 => (B_ipd'last_event,tpd_B_S, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING);

 end process;

end VITAL_ACT;


 configuration CFG_FA1B_VITAL of FA1B is
    for VITAL_ACT
    end for;
 end CFG_FA1B_VITAL;



 ---- CELL FA2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity FA2A is
    generic(
                TimingChecksOn:Boolean :=True;
                Xon: Boolean :=False;
                InstancePath: STRING :="*";
                MsgOn: Boolean :=True;
                tpd_CI_CO               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_B_CO                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_A0_CO               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_A1_CO               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_A0_S                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_A1_S                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_B_S         : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CI_S                : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_CI         : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_B          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_A0         : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_A1         : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                CI              : in    STD_ULOGIC;
                B               : in    STD_ULOGIC;
                A0              : in    STD_ULOGIC;
                A1              : in    STD_ULOGIC;
                CO              : out    STD_ULOGIC;
                S               : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of FA2A :  entity is TRUE;
 end FA2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library axcelerator;
use axcelerator.VTABLES.all;

architecture VITAL_ACT of FA2A is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL CI_ipd  : STD_ULOGIC := 'X';
        SIGNAL B_ipd  : STD_ULOGIC := 'X';
        SIGNAL A0_ipd  : STD_ULOGIC := 'X';
        SIGNAL A1_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (CI_ipd, CI, tipd_CI);
        VitalWireDelay (B_ipd, B, tipd_B);
        VitalWireDelay (A0_ipd, A0, tipd_A0);
        VitalWireDelay (A1_ipd, A1, tipd_A1);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (CI_ipd, B_ipd, A0_ipd, A1_ipd)


        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
        ALIAS CO_zd : STD_LOGIC is Results(1);
        ALIAS S_zd : STD_LOGIC is Results(2);

        -- output glitch detection variables
        VARIABLE CO_GlitchData  : VitalGlitchDataType;
        VARIABLE S_GlitchData  : VitalGlitchDataType;

        begin

           -------------------------
           --  Functionality Section
           -------------------------

              S_zd :=
       (((NOT ((A1_ipd) OR (A0_ipd)))) AND ((((A1_ipd) OR (A0_ipd)) AND
         ((NOT B_ipd))) OR (((NOT B_ipd)) AND (CI_ipd) AND ((NOT ((A1_ipd) OR
         (A0_ipd))))) OR ((CI_ipd) AND (B_ipd) AND ((A1_ipd) OR (A0_ipd))))
         AND (CI_ipd)) OR (((NOT ((A1_ipd) OR (A0_ipd)))) AND (B_ipd) AND
         ((NOT CI_ipd))) OR (((A1_ipd) OR (A0_ipd)) AND ((((A1_ipd) OR
         (A0_ipd)) AND ((NOT B_ipd))) OR (((NOT B_ipd)) AND (CI_ipd) AND
         ((NOT ((A1_ipd) OR (A0_ipd))))) OR ((CI_ipd) AND (B_ipd) AND
         ((A1_ipd) OR (A0_ipd)))) AND ((NOT CI_ipd))) OR (((A1_ipd) OR
         (A0_ipd)) AND (B_ipd) AND (CI_ipd));
      --CO_zd :=
      -- (((A1_ipd) OR (A0_ipd)) AND ((NOT B_ipd))) OR (((NOT B_ipd)) AND
      --   (CI_ipd) AND ((NOT ((A1_ipd) OR (A0_ipd))))) OR ((CI_ipd) AND
      --   (B_ipd) AND ((A1_ipd) OR (A0_ipd)));
      CO_zd :=
        (((A1_ipd) AND (NOT B_ipd)) OR ((A0_ipd) AND (NOT B_ipd)) OR
         ((A0_ipd) AND (CI_ipd)) OR ((A1_ipd) AND (CI_ipd)) OR
         ((NOT B_ipd) AND (CI_ipd)));


           ----------------------
           --  Path Delay Section
           ----------------------

     VitalPathDelay01 (
           OutSignal => CO,
           GlitchData => CO_GlitchData,
           OutSignalName => "CO",
           OutTemp => CO_zd,
           Paths => (
                     0 => (CI_ipd'last_event,tpd_CI_CO, true),
                     1 => (B_ipd'last_event,tpd_B_CO, true),
                     2 => (A0_ipd'last_event,tpd_A0_CO, true),
                     3 => (A1_ipd'last_event,tpd_A1_CO, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING);

    VitalPathDelay01 (
           OutSignal => S,
           GlitchData => S_GlitchData,
           OutSignalName => "S",
           OutTemp => S_zd,
           Paths => (
                     0 => (A0_ipd'last_event,tpd_A0_S, true),
                     1 => (A1_ipd'last_event,tpd_A1_S, true),
                     2 => (B_ipd'last_event,tpd_B_S, true),
                     3 => (CI_ipd'last_event,tpd_CI_S, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_FA2A_VITAL of FA2A is
    for VITAL_ACT
    end for;
 end CFG_FA2A_VITAL;




